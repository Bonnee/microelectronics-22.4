LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_unsigned.ALL;

ENTITY RCA IS
  PORT (
    A : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    B : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    Ci : IN STD_LOGIC;
    S : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    Co : OUT STD_LOGIC);
END RCA;

ARCHITECTURE STRUCTURAL OF RCA IS

  SIGNAL STMP : STD_LOGIC_VECTOR(5 DOWNTO 0);
  SIGNAL CTMP : STD_LOGIC_VECTOR(6 DOWNTO 0);

  COMPONENT FA
    PORT (
      A : IN STD_LOGIC;
      B : IN STD_LOGIC;
      Ci : IN STD_LOGIC;
      S : OUT STD_LOGIC;
      Co : OUT STD_LOGIC);
  END COMPONENT;

BEGIN

  CTMP(0) <= Ci;
  S <= STMP;
  Co <= CTMP(6);

  ADDER1 : FOR I IN 1 TO 6 GENERATE
    FAI : FA
    PORT MAP(A(I - 1), B(I - 1), CTMP(I - 1), STMP(I - 1), CTMP(I));
  END GENERATE;

END STRUCTURAL;
ARCHITECTURE BEHAVIORAL OF RCA IS

BEGIN

  S <= (A + B);

END BEHAVIORAL;

CONFIGURATION CFG_RCA_STRUCTURAL OF RCA IS
  FOR STRUCTURAL
    FOR ADDER1
      FOR ALL : FA
        USE CONFIGURATION WORK.CFG_FA_BEHAVIORAL;
      END FOR;
    END FOR;
  END FOR;
END CFG_RCA_STRUCTURAL;

CONFIGURATION CFG_RCA_BEHAVIORAL OF RCA IS
  FOR BEHAVIORAL
  END FOR;
END CFG_RCA_BEHAVIORAL;