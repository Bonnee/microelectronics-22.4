
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_BOOTHMUL_NBIT32 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_BOOTHMUL_NBIT32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT64_DW01_add_0 is

   port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (63 downto 0);  CO : out std_logic);

end RCA_NBIT64_DW01_add_0;

architecture SYN_rpl of RCA_NBIT64_DW01_add_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_29_port, carry_28_port, carry_27_port, carry_26_port, 
      carry_25_port, carry_24_port, carry_23_port, carry_22_port, carry_21_port
      , carry_20_port, carry_19_port, carry_18_port, carry_17_port, 
      carry_16_port, carry_15_port, carry_14_port, carry_13_port, carry_12_port
      , carry_11_port, carry_10_port, carry_9_port, carry_8_port, carry_7_port,
      carry_6_port, carry_5_port, carry_4_port, carry_3_port, carry_2_port, n1,
      n702, n716, n718, n719, n721, n730, n733, n734, n737, n739, n740, n742, 
      n743, n746, n753, n757, n758, n761, n763, n764, n766, n767, n769, n770, 
      n772, n773, n775, n776, n778, n779, n781, n782, n783, n784, n785, n786, 
      n787, n788, n789, n790, n791, n792, n793, n794, n796, n797, n798, n799, 
      n800, n801, n802, n803, net264871, net264877, net269988, net269993, 
      net270003, net270005, net270008, net270011, net270334, net270544, 
      net271683, net271681, net272167, net272197, net273975, net274069, 
      net274079, net270004, net276070, net273714, n715, n713, n712, net277992, 
      net278050, net278049, net278046, n755, n754, n752, n751, n749, n748, n745
      , n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
      n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, 
      n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, 
      n693, n694, n695, n696, n697, n698, n699, n700, n701, n703, n704, n705, 
      n706, n707, n708, n709, n710, n711, n714, n717, n720, n722, n723, n724, 
      n725, n726, n727, n728, n729, n731, n732, n735, n736, n738, n741, n744, 
      n747, n750, n756, n759, n760, n762, n765, n768, n771, n774, n777, n780, 
      n795, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, 
      n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, 
      n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, 
      n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, 
      n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, 
      n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, 
      n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885 : 
      std_logic;

begin
   
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U116 : XOR2_X1 port map( A => B(63), B => A(63), Z => n702);
   U149 : XOR2_X1 port map( A => n700, B => n753, Z => SUM(46));
   U161 : XOR2_X1 port map( A => n836, B => n770, Z => SUM(40));
   U162 : XOR2_X1 port map( A => A(40), B => B(40), Z => n770);
   U169 : XOR2_X1 port map( A => n750, B => n783, Z => SUM(36));
   U170 : XOR2_X1 port map( A => B(36), B => A(36), Z => n783);
   U171 : XOR2_X1 port map( A => n664, B => n786, Z => SUM(35));
   U172 : XOR2_X1 port map( A => B(35), B => n663, Z => n786);
   U173 : XOR2_X1 port map( A => n707, B => n789, Z => SUM(34));
   U174 : XOR2_X1 port map( A => B(34), B => A(34), Z => n789);
   U175 : XOR2_X1 port map( A => n820, B => n792, Z => SUM(33));
   U176 : XOR2_X1 port map( A => B(33), B => n811, Z => n792);
   U178 : XOR2_X1 port map( A => n873, B => n797, Z => SUM(31));
   U179 : XOR2_X1 port map( A => B(31), B => A(31), Z => n797);
   U180 : XOR2_X1 port map( A => n799, B => n801, Z => SUM(30));
   U181 : XOR2_X1 port map( A => B(30), B => A(30), Z => n801);
   U182 : XOR2_X1 port map( A => A(29), B => n803, Z => SUM(29));
   U183 : XOR2_X1 port map( A => carry_29_port, B => B(29), Z => n803);
   U184 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U150 : XOR2_X1 port map( A => n701, B => B(46), Z => n753);
   U1 : CLKBUF_X1 port map( A => A(56), Z => n657);
   U2 : INV_X1 port map( A => A(55), ZN => n658);
   U3 : CLKBUF_X1 port map( A => n751, Z => n700);
   U4 : CLKBUF_X1 port map( A => n712, Z => n659);
   U5 : INV_X1 port map( A => B(54), ZN => n680);
   U6 : INV_X1 port map( A => B(55), ZN => n681);
   U7 : INV_X1 port map( A => A(53), ZN => n684);
   U8 : INV_X1 port map( A => B(53), ZN => n677);
   U9 : AND2_X1 port map( A1 => n868, A2 => n838, ZN => n836);
   U10 : XNOR2_X1 port map( A => n690, B => n683, ZN => SUM(53));
   U11 : XNOR2_X1 port map( A => A(53), B => B(53), ZN => n683);
   U12 : XNOR2_X1 port map( A => n693, B => n682, ZN => SUM(55));
   U13 : XNOR2_X1 port map( A => B(55), B => n670, ZN => n682);
   U14 : INV_X1 port map( A => n702, ZN => n759);
   U15 : XNOR2_X1 port map( A => n736, B => n725, ZN => SUM(60));
   U16 : CLKBUF_X1 port map( A => n824, Z => n660);
   U17 : CLKBUF_X1 port map( A => n778, Z => n661);
   U18 : CLKBUF_X1 port map( A => A(49), Z => n662);
   U19 : CLKBUF_X1 port map( A => A(35), Z => n663);
   U20 : CLKBUF_X1 port map( A => n784, Z => n664);
   U21 : CLKBUF_X1 port map( A => A(59), Z => net277992);
   U22 : CLKBUF_X1 port map( A => n678, Z => n665);
   U23 : AND2_X1 port map( A1 => n671, A2 => n687, ZN => n666);
   U24 : AND2_X1 port map( A1 => n674, A2 => n673, ZN => n667);
   U25 : AND2_X1 port map( A1 => n673, A2 => n674, ZN => n668);
   U26 : AND2_X1 port map( A1 => n675, A2 => n681, ZN => n669);
   U27 : NAND2_X1 port map( A1 => n675, A2 => n676, ZN => n670);
   U28 : XNOR2_X1 port map( A => A(60), B => B(60), ZN => n725);
   U29 : XNOR2_X1 port map( A => B(59), B => net273714, ZN => net270004);
   U30 : OAI211_X1 port map( C1 => n717, C2 => n714, A => n720, B => n722, ZN 
                           => n711);
   U31 : INV_X1 port map( A => A(60), ZN => n717);
   U32 : INV_X1 port map( A => B(60), ZN => n714);
   U33 : OAI21_X1 port map( B1 => n681, B2 => n692, A => n685, ZN => n671);
   U34 : NAND2_X1 port map( A1 => n678, A2 => n677, ZN => n673);
   U35 : BUF_X1 port map( A => n840, Z => n771);
   U36 : CLKBUF_X1 port map( A => net278046, Z => n672);
   U37 : NAND2_X1 port map( A1 => n669, A2 => n676, ZN => n687);
   U38 : NAND2_X1 port map( A1 => n688, A2 => n684, ZN => n674);
   U39 : NAND2_X1 port map( A1 => n730, A2 => B(53), ZN => n688);
   U40 : BUF_X1 port map( A => A(54), Z => n691);
   U41 : NAND2_X1 port map( A1 => B(54), A2 => n691, ZN => n675);
   U42 : XNOR2_X1 port map( A => n691, B => B(54), ZN => net270008);
   U43 : INV_X1 port map( A => A(54), ZN => n679);
   U44 : INV_X1 port map( A => n730, ZN => n678);
   U45 : INV_X1 port map( A => n665, ZN => n690);
   U46 : OAI21_X1 port map( B1 => n692, B2 => n681, A => n685, ZN => n686);
   U47 : INV_X1 port map( A => A(55), ZN => n685);
   U48 : INV_X1 port map( A => n658, ZN => n693);
   U49 : NAND2_X1 port map( A1 => n667, A2 => n689, ZN => n676);
   U50 : AND2_X1 port map( A1 => n694, A2 => n675, ZN => n692);
   U51 : AND2_X1 port map( A1 => n686, A2 => n687, ZN => net264877);
   U52 : NAND2_X1 port map( A1 => n680, A2 => n679, ZN => n689);
   U53 : NAND2_X1 port map( A1 => n668, A2 => n689, ZN => n694);
   U54 : AND2_X1 port map( A1 => n671, A2 => n687, ZN => n695);
   U55 : AOI21_X1 port map( B1 => n697, B2 => n699, A => n749, ZN => n745);
   U56 : AND2_X1 port map( A1 => n745, A2 => A(48), ZN => net270334);
   U57 : CLKBUF_X1 port map( A => n745, Z => net271683);
   U58 : OAI21_X1 port map( B1 => n745, B2 => A(48), A => B(48), ZN => n746);
   U59 : AOI21_X1 port map( B1 => n698, B2 => A(47), A => B(47), ZN => n749);
   U60 : INV_X1 port map( A => n748, ZN => n698);
   U61 : INV_X1 port map( A => n698, ZN => n699);
   U62 : AOI22_X1 port map( A1 => n700, A2 => n703, B1 => n752, B2 => B(46), ZN
                           => n748);
   U63 : OR2_X1 port map( A1 => n751, A2 => A(46), ZN => n752);
   U64 : CLKBUF_X1 port map( A => A(46), Z => n703);
   U65 : CLKBUF_X1 port map( A => n703, Z => n701);
   U66 : INV_X1 port map( A => n699, ZN => net270544);
   U67 : INV_X1 port map( A => A(47), ZN => n697);
   U68 : CLKBUF_X1 port map( A => A(47), Z => n705);
   U69 : XNOR2_X1 port map( A => B(47), B => n705, ZN => net269993);
   U70 : AOI21_X1 port map( B1 => n696, B2 => n754, A => n755, ZN => n751);
   U71 : AOI21_X1 port map( B1 => net272197, B2 => A(45), A => B(45), ZN => 
                           n755);
   U72 : INV_X1 port map( A => net272197, ZN => n754);
   U73 : INV_X1 port map( A => n754, ZN => net276070);
   U74 : INV_X1 port map( A => A(45), ZN => n696);
   U75 : INV_X1 port map( A => n696, ZN => n704);
   U76 : XNOR2_X1 port map( A => B(45), B => n704, ZN => net269988);
   U77 : OR2_X1 port map( A1 => n781, A2 => n876, ZN => n706);
   U78 : NAND2_X1 port map( A1 => n782, A2 => n706, ZN => n778);
   U79 : INV_X1 port map( A => n787, ZN => n707);
   U80 : NAND2_X1 port map( A1 => n713, A2 => B(59), ZN => n708);
   U81 : CLKBUF_X1 port map( A => n659, Z => n709);
   U82 : NAND2_X1 port map( A1 => net278046, A2 => n708, ZN => n710);
   U83 : CLKBUF_X1 port map( A => n720, Z => n732);
   U84 : XNOR2_X1 port map( A => n729, B => B(61), ZN => net270005);
   U85 : NAND2_X1 port map( A1 => n711, A2 => n728, ZN => n724);
   U86 : NAND2_X1 port map( A1 => n710, A2 => B(60), ZN => n722);
   U87 : OAI211_X1 port map( C1 => n714, C2 => n717, A => n732, B => n731, ZN 
                           => net272167);
   U88 : NAND2_X1 port map( A1 => n726, A2 => A(60), ZN => n720);
   U89 : NAND2_X1 port map( A1 => n724, A2 => n738, ZN => n723);
   U90 : AOI21_X1 port map( B1 => n723, B2 => A(62), A => B(62), ZN => 
                           net278049);
   U91 : NOR2_X1 port map( A1 => n735, A2 => A(62), ZN => net278050);
   U92 : CLKBUF_X1 port map( A => n735, Z => net274069);
   U93 : NAND2_X1 port map( A1 => n727, A2 => net278046, ZN => n726);
   U94 : NAND2_X1 port map( A1 => n724, A2 => n738, ZN => n735);
   U95 : NAND2_X1 port map( A1 => n713, A2 => B(59), ZN => n727);
   U96 : NAND2_X1 port map( A1 => n741, A2 => n672, ZN => n736);
   U97 : OR2_X1 port map( A1 => A(61), A2 => B(61), ZN => n728);
   U98 : NAND2_X1 port map( A1 => n729, A2 => B(61), ZN => n738);
   U99 : BUF_X1 port map( A => A(61), Z => n729);
   U100 : CLKBUF_X1 port map( A => n727, Z => n741);
   U101 : CLKBUF_X1 port map( A => n722, Z => n731);
   U102 : BUF_X1 port map( A => n844, Z => n744);
   U103 : BUF_X1 port map( A => n763, Z => n844);
   U104 : CLKBUF_X1 port map( A => n829, Z => n747);
   U105 : INV_X1 port map( A => n781, ZN => n750);
   U106 : NAND2_X1 port map( A1 => n659, A2 => net277992, ZN => net278046);
   U107 : NOR2_X1 port map( A1 => net278049, A2 => net278050, ZN => n756);
   U108 : XNOR2_X1 port map( A => n756, B => n759, ZN => SUM(63));
   U109 : XNOR2_X1 port map( A => A(62), B => B(62), ZN => net270011);
   U110 : OR2_X1 port map( A1 => A(59), A2 => n712, ZN => n713);
   U111 : CLKBUF_X1 port map( A => net277992, Z => net273714);
   U112 : OAI21_X1 port map( B1 => n762, B2 => n760, A => n715, ZN => n712);
   U113 : OAI21_X1 port map( B1 => n716, B2 => A(58), A => B(58), ZN => n715);
   U114 : INV_X1 port map( A => A(58), ZN => n760);
   U115 : INV_X1 port map( A => n716, ZN => n762);
   U117 : XNOR2_X1 port map( A => B(58), B => A(58), ZN => net270003);
   U118 : CLKBUF_X1 port map( A => A(42), Z => n765);
   U119 : BUF_X1 port map( A => n739, Z => n840);
   U120 : CLKBUF_X1 port map( A => A(51), Z => n768);
   U121 : CLKBUF_X1 port map( A => n815, Z => n774);
   U122 : CLKBUF_X1 port map( A => n771, Z => n777);
   U123 : INV_X1 port map( A => n775, ZN => n780);
   U124 : AND2_X1 port map( A1 => n817, A2 => n871, ZN => n795);
   U125 : OR2_X1 port map( A1 => n805, A2 => n865, ZN => n804);
   U126 : AND2_X1 port map( A1 => n840, A2 => n814, ZN => n805);
   U127 : BUF_X1 port map( A => A(50), Z => n814);
   U128 : AND2_X1 port map( A1 => n844, A2 => A(42), ZN => n806);
   U129 : AND2_X1 port map( A1 => n869, A2 => n826, ZN => n807);
   U130 : CLKBUF_X1 port map( A => A(57), Z => n813);
   U131 : OR2_X1 port map( A1 => n806, A2 => n866, ZN => n808);
   U132 : OR2_X1 port map( A1 => n806, A2 => n866, ZN => n809);
   U133 : XNOR2_X1 port map( A => net270004, B => n709, ZN => SUM(59));
   U134 : INV_X1 port map( A => n872, ZN => n810);
   U135 : CLKBUF_X1 port map( A => A(33), Z => n811);
   U136 : INV_X1 port map( A => n774, ZN => n812);
   U137 : CLKBUF_X1 port map( A => net264871, Z => net274079);
   U138 : AOI21_X1 port map( B1 => n771, B2 => n814, A => n865, ZN => n815);
   U139 : CLKBUF_X1 port map( A => A(48), Z => net273975);
   U140 : AOI21_X1 port map( B1 => n809, B2 => A(43), A => B(43), ZN => n816);
   U141 : OR2_X1 port map( A1 => n790, A2 => A(33), ZN => n817);
   U142 : NAND2_X1 port map( A1 => n817, A2 => n871, ZN => n787);
   U143 : CLKBUF_X1 port map( A => n809, Z => n818);
   U144 : CLKBUF_X1 port map( A => A(37), Z => n839);
   U145 : AND2_X1 port map( A1 => n870, A2 => n837, ZN => n819);
   U146 : CLKBUF_X1 port map( A => n790, Z => n820);
   U147 : CLKBUF_X1 port map( A => n765, Z => n821);
   U148 : OR2_X1 port map( A1 => n695, A2 => A(56), ZN => n822);
   U151 : OR2_X1 port map( A1 => net264877, A2 => A(56), ZN => n721);
   U152 : INV_X1 port map( A => n660, ZN => n823);
   U153 : AOI22_X1 port map( A1 => n666, A2 => A(56), B1 => n822, B2 => B(56), 
                           ZN => n824);
   U154 : INV_X1 port map( A => n841, ZN => n825);
   U155 : OR2_X1 port map( A1 => n778, A2 => A(37), ZN => n826);
   U156 : NAND2_X1 port map( A1 => n869, A2 => n826, ZN => n775);
   U157 : AOI21_X1 port map( B1 => n744, B2 => n765, A => n866, ZN => n827);
   U158 : NAND2_X1 port map( A1 => n758, A2 => n828, ZN => net272197);
   U159 : NAND2_X1 port map( A1 => n829, A2 => A(44), ZN => n828);
   U160 : NOR2_X1 port map( A1 => n816, A2 => n843, ZN => n829);
   U163 : CLKBUF_X1 port map( A => n772, Z => n830);
   U164 : CLKBUF_X1 port map( A => A(38), Z => n831);
   U165 : INV_X1 port map( A => n762, ZN => net271681);
   U166 : INV_X1 port map( A => n864, ZN => n832);
   U167 : OR2_X1 port map( A1 => net274079, A2 => net270334, ZN => n833);
   U168 : CLKBUF_X1 port map( A => A(39), Z => n834);
   U177 : AND2_X1 port map( A1 => n868, A2 => n838, ZN => n835);
   U185 : OR2_X1 port map( A1 => n784, A2 => A(35), ZN => n837);
   U186 : NAND2_X1 port map( A1 => n870, A2 => n837, ZN => n781);
   U187 : OR2_X1 port map( A1 => n772, A2 => A(39), ZN => n838);
   U188 : INV_X1 port map( A => n867, ZN => n841);
   U189 : OR2_X1 port map( A1 => net264871, A2 => net270334, ZN => n842);
   U190 : NOR2_X1 port map( A1 => net270334, A2 => net264871, ZN => n742);
   U191 : AND2_X1 port map( A1 => n882, A2 => n827, ZN => n843);
   U192 : NOR2_X1 port map( A1 => n843, A2 => n761, ZN => n757);
   U193 : AND2_X1 port map( A1 => n881, A2 => n742, ZN => n845);
   U194 : NOR2_X1 port map( A1 => n743, A2 => n845, ZN => n739);
   U195 : AND2_X1 port map( A1 => n878, A2 => n824, ZN => n846);
   U196 : NOR2_X1 port map( A1 => n846, A2 => n719, ZN => n716);
   U197 : AND2_X1 port map( A1 => n815, A2 => n880, ZN => n847);
   U198 : NOR2_X1 port map( A1 => n737, A2 => n847, ZN => n734);
   U199 : XOR2_X1 port map( A => n830, B => n848, Z => SUM(39));
   U200 : XOR2_X1 port map( A => B(39), B => n834, Z => n848);
   U201 : XOR2_X1 port map( A => n661, B => n849, Z => SUM(37));
   U202 : XOR2_X1 port map( A => B(37), B => n839, Z => n849);
   U203 : XOR2_X1 port map( A => n744, B => n850, Z => SUM(42));
   U204 : XOR2_X1 port map( A => B(42), B => n821, Z => n850);
   U205 : XOR2_X1 port map( A => n747, B => n851, Z => SUM(44));
   U206 : XOR2_X1 port map( A => B(44), B => A(44), Z => n851);
   U207 : INV_X1 port map( A => A(32), ZN => n874);
   U208 : INV_X1 port map( A => A(51), ZN => n880);
   U209 : INV_X1 port map( A => A(41), ZN => n877);
   U210 : INV_X1 port map( A => A(43), ZN => n882);
   U211 : INV_X1 port map( A => A(34), ZN => n875);
   U212 : OAI21_X1 port map( B1 => n872, B2 => A(32), A => B(32), ZN => n794);
   U213 : INV_X1 port map( A => A(49), ZN => n881);
   U214 : INV_X1 port map( A => A(57), ZN => n878);
   U215 : INV_X1 port map( A => A(38), ZN => n883);
   U216 : INV_X1 port map( A => A(52), ZN => n879);
   U217 : INV_X1 port map( A => n791, ZN => n871);
   U218 : XNOR2_X1 port map( A => net274069, B => net270011, ZN => SUM(62));
   U219 : XNOR2_X1 port map( A => n666, B => n852, ZN => SUM(56));
   U220 : XNOR2_X1 port map( A => n657, B => B(56), ZN => n852);
   U221 : XNOR2_X1 port map( A => n667, B => net270008, ZN => SUM(54));
   U222 : XNOR2_X1 port map( A => n823, B => n853, ZN => SUM(57));
   U223 : XNOR2_X1 port map( A => n813, B => B(57), ZN => n853);
   U224 : XNOR2_X1 port map( A => net272167, B => net270005, ZN => SUM(61));
   U225 : XNOR2_X1 port map( A => net271681, B => net270003, ZN => SUM(58));
   U226 : XNOR2_X1 port map( A => n833, B => n854, ZN => SUM(49));
   U227 : XNOR2_X1 port map( A => n662, B => B(49), ZN => n854);
   U228 : XNOR2_X1 port map( A => net270544, B => net269993, ZN => SUM(47));
   U229 : XNOR2_X1 port map( A => n812, B => n855, ZN => SUM(51));
   U230 : XNOR2_X1 port map( A => n768, B => B(51), ZN => n855);
   U231 : XNOR2_X1 port map( A => net276070, B => net269988, ZN => SUM(45));
   U232 : XNOR2_X1 port map( A => n832, B => n856, ZN => SUM(52));
   U233 : XNOR2_X1 port map( A => A(52), B => B(52), ZN => n856);
   U234 : XNOR2_X1 port map( A => n777, B => n857, ZN => SUM(50));
   U235 : XNOR2_X1 port map( A => n814, B => B(50), ZN => n857);
   U236 : XNOR2_X1 port map( A => net271683, B => n858, ZN => SUM(48));
   U237 : XNOR2_X1 port map( A => net273975, B => B(48), ZN => n858);
   U238 : XNOR2_X1 port map( A => n872, B => n859, ZN => SUM(32));
   U239 : XOR2_X1 port map( A => B(32), B => n874, Z => n859);
   U240 : XNOR2_X1 port map( A => n818, B => n860, ZN => SUM(43));
   U241 : XNOR2_X1 port map( A => A(43), B => B(43), ZN => n860);
   U242 : XNOR2_X1 port map( A => n825, B => n861, ZN => SUM(41));
   U243 : XNOR2_X1 port map( A => B(41), B => A(41), ZN => n861);
   U244 : XNOR2_X1 port map( A => n780, B => n862, ZN => SUM(38));
   U245 : XNOR2_X1 port map( A => B(38), B => n831, ZN => n862);
   U246 : INV_X1 port map( A => n798, ZN => n873);
   U247 : OAI22_X1 port map( A1 => A(30), A2 => n799, B1 => B(30), B2 => n800, 
                           ZN => n798);
   U248 : AND2_X1 port map( A1 => n799, A2 => A(30), ZN => n800);
   U249 : AOI21_X1 port map( B1 => n885, B2 => n884, A => n802, ZN => n799);
   U250 : INV_X1 port map( A => B(29), ZN => n885);
   U251 : INV_X1 port map( A => A(29), ZN => n884);
   U252 : AOI21_X1 port map( B1 => A(29), B2 => B(29), A => carry_29_port, ZN 
                           => n802);
   U253 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U254 : INV_X1 port map( A => A(36), ZN => n876);
   U255 : OR2_X1 port map( A1 => n835, A2 => A(40), ZN => n769);
   U256 : AOI22_X1 port map( A1 => n836, A2 => A(40), B1 => n769, B2 => B(40), 
                           ZN => n766);
   U257 : OAI21_X1 port map( B1 => n807, B2 => A(38), A => B(38), ZN => n776);
   U258 : INV_X1 port map( A => n785, ZN => n870);
   U259 : OAI21_X1 port map( B1 => n819, B2 => A(36), A => B(36), ZN => n782);
   U260 : OAI21_X1 port map( B1 => n795, B2 => A(34), A => B(34), ZN => n788);
   U261 : AOI21_X1 port map( B1 => n867, B2 => A(41), A => B(41), ZN => n767);
   U262 : AOI21_X1 port map( B1 => n808, B2 => A(43), A => B(43), ZN => n761);
   U263 : INV_X1 port map( A => n764, ZN => n866);
   U264 : INV_X1 port map( A => n773, ZN => n868);
   U265 : AOI21_X1 port map( B1 => n784, B2 => A(35), A => B(35), ZN => n785);
   U266 : OAI21_X1 port map( B1 => n787, B2 => n875, A => n788, ZN => n784);
   U267 : OAI22_X1 port map( A1 => A(31), A2 => n873, B1 => n796, B2 => B(31), 
                           ZN => n793);
   U268 : AND2_X1 port map( A1 => n873, A2 => A(31), ZN => n796);
   U269 : OAI21_X1 port map( B1 => n739, B2 => A(50), A => B(50), ZN => n740);
   U270 : INV_X1 port map( A => n734, ZN => n864);
   U271 : OAI21_X1 port map( B1 => n734, B2 => A(52), A => B(52), ZN => n733);
   U272 : AOI22_X1 port map( A1 => n666, A2 => A(56), B1 => n721, B2 => B(56), 
                           ZN => n718);
   U273 : INV_X1 port map( A => n740, ZN => n865);
   U274 : AOI21_X1 port map( B1 => n772, B2 => A(39), A => B(39), ZN => n773);
   U275 : INV_X1 port map( A => n779, ZN => n869);
   U276 : AOI21_X1 port map( B1 => n778, B2 => A(37), A => B(37), ZN => n779);
   U277 : AOI21_X1 port map( B1 => n790, B2 => A(33), A => B(33), ZN => n791);
   U278 : OAI21_X1 port map( B1 => n810, B2 => n874, A => n794, ZN => n790);
   U279 : INV_X1 port map( A => n793, ZN => n872);
   U280 : OAI21_X1 port map( B1 => n864, B2 => n879, A => n733, ZN => n730);
   U281 : INV_X1 port map( A => n746, ZN => net264871);
   U282 : OAI21_X1 port map( B1 => n757, B2 => A(44), A => B(44), ZN => n758);
   U283 : OAI21_X1 port map( B1 => n763, B2 => A(42), A => B(42), ZN => n764);
   U284 : AOI21_X1 port map( B1 => n877, B2 => n841, A => n767, ZN => n763);
   U285 : INV_X1 port map( A => n766, ZN => n867);
   U286 : OAI21_X1 port map( B1 => n775, B2 => n883, A => n776, ZN => n772);
   U287 : INV_X1 port map( A => n718, ZN => n863);
   U288 : AOI21_X1 port map( B1 => n842, B2 => A(49), A => B(49), ZN => n743);
   U289 : AOI21_X1 port map( B1 => n804, B2 => A(51), A => B(51), ZN => n737);
   U290 : AOI21_X1 port map( B1 => n863, B2 => A(57), A => B(57), ZN => n719);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT62_DW01_add_0 is

   port( A, B : in std_logic_vector (61 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (61 downto 0);  CO : out std_logic);

end RCA_NBIT62_DW01_add_0;

architecture SYN_rpl of RCA_NBIT62_DW01_add_0 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_28_port, carry_27_port, carry_26_port, carry_25_port, 
      carry_24_port, carry_23_port, carry_22_port, carry_21_port, carry_20_port
      , carry_19_port, carry_18_port, carry_17_port, carry_16_port, 
      carry_15_port, carry_14_port, carry_13_port, carry_12_port, carry_11_port
      , carry_10_port, carry_9_port, carry_8_port, carry_7_port, carry_6_port, 
      carry_5_port, carry_4_port, carry_3_port, carry_2_port, n1, carry_59_port
      , carry_58_port, n600, n601, n602, n603, n604, n605, n606, n607, n610, 
      n611, n612, n613, n615, n621, n622, n625, n626, n627, n628, n629, n631, 
      n632, n633, n634, n635, n637, n638, n639, n642, n645, n646, n649, n650, 
      n651, n652, n653, n655, n656, n657, n658, n659, n661, n662, n663, n664, 
      n665, n667, n668, n669, n670, n671, n673, n674, n675, n676, n677, n679, 
      n680, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, 
      net264804, net264822, net264823, net270409, net270476, net270966, 
      net271876, net273837, net274638, net297750, n647, n644, n643, n620, n619,
      n617, n616, n614, n556, n557, n558, n559, n560, n561, n562, n563, n564, 
      n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, 
      n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, 
      n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n608, 
      n609, n618, n623, n624, n630, n636, n640, n641, n648, n654, n660, n666, 
      n672, n678, n681, n693, n694, n695, n696, n697, n698, n699, n700, n701, 
      n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, 
      n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, 
      n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, 
      n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, 
      n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, 
      n762, n763, n764, n765 : std_logic;

begin
   
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U1_58 : FA_X1 port map( A => A(58), B => B(58), CI => carry_58_port, CO => 
                           carry_59_port, S => SUM(58));
   U141 : XOR2_X1 port map( A => B(61), B => A(61), Z => n603);
   U142 : XOR2_X1 port map( A => B(60), B => A(60), Z => n606);
   U156 : XOR2_X1 port map( A => n642, B => n577, Z => SUM(45));
   U167 : XOR2_X1 port map( A => A(30), B => B(30), Z => n687);
   U168 : XOR2_X1 port map( A => B(29), B => n733, Z => n690);
   U169 : XOR2_X1 port map( A => A(28), B => n692, Z => SUM(28));
   U170 : XOR2_X1 port map( A => carry_28_port, B => B(28), Z => n692);
   U171 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U149 : XOR2_X1 port map( A => n561, B => B(52), Z => n621);
   U1 : INV_X1 port map( A => A(45), ZN => n556);
   U2 : CLKBUF_X1 port map( A => net270966, Z => n557);
   U3 : OR2_X1 port map( A1 => n613, A2 => net264804, ZN => n558);
   U4 : AND2_X2 port map( A1 => n579, A2 => n644, ZN => n578);
   U5 : XNOR2_X1 port map( A => n605, B => n606, ZN => SUM(60));
   U6 : BUF_X1 port map( A => n699, Z => n559);
   U7 : CLKBUF_X1 port map( A => n646, Z => n623);
   U8 : OAI21_X1 port map( B1 => n624, B2 => n623, A => n618, ZN => n560);
   U9 : BUF_X1 port map( A => A(52), Z => n561);
   U10 : CLKBUF_X1 port map( A => net264822, Z => n562);
   U11 : XNOR2_X1 port map( A => n623, B => n563, ZN => SUM(43));
   U12 : XNOR2_X1 port map( A => A(43), B => B(43), ZN => n563);
   U13 : AOI21_X1 port map( B1 => n756, B2 => n559, A => n683, ZN => n564);
   U14 : BUF_X1 port map( A => n593, Z => n565);
   U15 : NAND2_X1 port map( A1 => n585, A2 => n584, ZN => n566);
   U16 : BUF_X2 port map( A => A(49), Z => n719);
   U17 : CLKBUF_X1 port map( A => A(55), Z => n567);
   U18 : INV_X1 port map( A => n750, ZN => n568);
   U19 : CLKBUF_X1 port map( A => n566, Z => n569);
   U20 : CLKBUF_X1 port map( A => n745, Z => n570);
   U21 : BUF_X1 port map( A => A(54), Z => n609);
   U22 : CLKBUF_X1 port map( A => n746, Z => n695);
   U23 : BUF_X1 port map( A => n628, Z => n726);
   U24 : BUF_X1 port map( A => A(30), Z => n681);
   U25 : CLKBUF_X1 port map( A => n752, Z => n571);
   U26 : BUF_X1 port map( A => n652, Z => n735);
   U27 : BUF_X1 port map( A => n706, Z => n572);
   U28 : CLKBUF_X1 port map( A => A(56), Z => n730);
   U29 : XNOR2_X1 port map( A => n569, B => n573, ZN => SUM(57));
   U30 : XNOR2_X1 port map( A => A(57), B => B(57), ZN => n573);
   U31 : NAND2_X1 port map( A1 => n566, A2 => A(57), ZN => n574);
   U32 : NAND2_X1 port map( A1 => n586, A2 => B(57), ZN => n575);
   U33 : NAND2_X1 port map( A1 => A(57), A2 => B(57), ZN => n576);
   U34 : NAND3_X1 port map( A1 => n574, A2 => n575, A3 => n576, ZN => 
                           carry_58_port);
   U35 : INV_X1 port map( A => B(31), ZN => n710);
   U36 : INV_X1 port map( A => B(45), ZN => n630);
   U37 : INV_X1 port map( A => n578, ZN => n577);
   U38 : NAND2_X1 port map( A1 => net264822, A2 => A(44), ZN => n579);
   U39 : AOI21_X1 port map( B1 => n758, B2 => n707, A => n610, ZN => n580);
   U40 : NAND2_X1 port map( A1 => n593, A2 => n599, ZN => n581);
   U41 : NAND2_X1 port map( A1 => n598, A2 => B(51), ZN => n582);
   U42 : NAND2_X1 port map( A1 => n582, A2 => n581, ZN => n583);
   U43 : BUF_X1 port map( A => n622, Z => n593);
   U44 : NAND2_X1 port map( A1 => n580, A2 => n730, ZN => n584);
   U45 : NAND2_X1 port map( A1 => n601, A2 => B(56), ZN => n585);
   U46 : NAND2_X1 port map( A1 => n585, A2 => n584, ZN => n586);
   U47 : INV_X1 port map( A => B(54), ZN => n594);
   U48 : NAND2_X1 port map( A1 => n578, A2 => n587, ZN => net270966);
   U49 : INV_X1 port map( A => A(45), ZN => n587);
   U50 : XOR2_X1 port map( A => A(55), B => B(55), Z => n612);
   U51 : OAI21_X1 port map( B1 => n578, B2 => n556, A => n630, ZN => net264823)
                           ;
   U52 : OAI21_X1 port map( B1 => n682, B2 => n588, A => n710, ZN => n589);
   U53 : INV_X1 port map( A => A(31), ZN => n588);
   U54 : INV_X1 port map( A => n589, ZN => n683);
   U55 : OAI21_X1 port map( B1 => n597, B2 => n609, A => B(54), ZN => n614);
   U56 : NAND2_X1 port map( A1 => n614, A2 => net271876, ZN => n611);
   U57 : AND2_X1 port map( A1 => n591, A2 => n596, ZN => n597);
   U58 : INV_X1 port map( A => n617, ZN => n591);
   U59 : AND2_X1 port map( A1 => n591, A2 => n596, ZN => n608);
   U60 : NAND2_X1 port map( A1 => n591, A2 => n596, ZN => n613);
   U61 : AOI21_X1 port map( B1 => n616, B2 => A(53), A => B(53), ZN => n617);
   U62 : INV_X1 port map( A => A(54), ZN => net264804);
   U63 : XNOR2_X1 port map( A => A(54), B => n594, ZN => n615);
   U64 : OAI21_X1 port map( B1 => n609, B2 => n608, A => B(54), ZN => net273837
                           );
   U65 : OR2_X1 port map( A1 => A(53), A2 => n616, ZN => n596);
   U66 : NAND2_X1 port map( A1 => n620, A2 => n595, ZN => n616);
   U67 : CLKBUF_X1 port map( A => n616, Z => net274638);
   U68 : OR2_X1 port map( A1 => n619, A2 => n590, ZN => n595);
   U69 : INV_X1 port map( A => A(52), ZN => n590);
   U70 : OAI21_X1 port map( B1 => n583, B2 => n561, A => B(52), ZN => n620);
   U71 : OR2_X1 port map( A1 => n622, A2 => A(51), ZN => n598);
   U72 : CLKBUF_X1 port map( A => A(51), Z => n599);
   U73 : AOI22_X1 port map( A1 => n593, A2 => n599, B1 => net297750, B2 => 
                           B(51), ZN => n619);
   U74 : XNOR2_X1 port map( A => n565, B => n592, ZN => SUM(51));
   U75 : XNOR2_X1 port map( A => A(53), B => B(53), ZN => net270409);
   U76 : CLKBUF_X1 port map( A => n619, Z => net270476);
   U77 : XNOR2_X1 port map( A => A(51), B => B(51), ZN => n592);
   U78 : OAI21_X1 port map( B1 => n636, B2 => A(44), A => B(44), ZN => n644);
   U79 : INV_X1 port map( A => n643, ZN => n636);
   U80 : OAI21_X1 port map( B1 => n624, B2 => n623, A => n618, ZN => n643);
   U81 : INV_X1 port map( A => n647, ZN => n618);
   U82 : AOI21_X1 port map( B1 => n646, B2 => A(43), A => B(43), ZN => n647);
   U83 : CLKBUF_X1 port map( A => A(43), Z => n624);
   U84 : XNOR2_X1 port map( A => A(45), B => n630, ZN => n642);
   U85 : XNOR2_X1 port map( A => A(44), B => B(44), ZN => n645);
   U86 : INV_X1 port map( A => n560, ZN => net264822);
   U87 : OR2_X1 port map( A1 => n622, A2 => A(51), ZN => net297750);
   U88 : CLKBUF_X1 port map( A => A(29), Z => n733);
   U89 : AND2_X1 port map( A1 => n672, A2 => A(60), ZN => n640);
   U90 : XNOR2_X1 port map( A => A(40), B => B(40), ZN => n657);
   U91 : NAND2_X1 port map( A1 => n680, A2 => n712, ZN => n641);
   U92 : AOI21_X1 port map( B1 => A(33), B2 => n641, A => B(33), ZN => n648);
   U93 : INV_X1 port map( A => n664, ZN => n654);
   U94 : OR2_X1 port map( A1 => n751, A2 => n713, ZN => n702);
   U95 : CLKBUF_X1 port map( A => A(39), Z => n701);
   U96 : AND2_X1 port map( A1 => n765, A2 => n670, ZN => n660);
   U97 : NOR2_X1 port map( A1 => n660, A2 => n671, ZN => n708);
   U98 : AND2_X1 port map( A1 => n743, A2 => n672, ZN => n666);
   U99 : OR2_X1 port map( A1 => A(59), A2 => B(59), ZN => n672);
   U100 : NAND2_X1 port map( A1 => n743, A2 => n672, ZN => n605);
   U101 : CLKBUF_X1 port map( A => n731, Z => n678);
   U102 : NOR2_X1 port map( A1 => n671, A2 => n660, ZN => n667);
   U103 : INV_X1 port map( A => n711, ZN => n676);
   U104 : XNOR2_X1 port map( A => n602, B => n603, ZN => SUM(61));
   U105 : OAI21_X1 port map( B1 => n719, B2 => n726, A => n570, ZN => n693);
   U106 : CLKBUF_X1 port map( A => A(41), Z => n714);
   U107 : XOR2_X1 port map( A => n753, B => n687, Z => SUM(30));
   U108 : CLKBUF_X1 port map( A => n747, Z => n694);
   U109 : INV_X1 port map( A => n625, ZN => n696);
   U110 : AND2_X1 port map( A1 => n764, A2 => n664, ZN => n697);
   U111 : NOR2_X1 port map( A1 => n665, A2 => n697, ZN => n662);
   U112 : XNOR2_X1 port map( A => n698, B => n735, ZN => SUM(41));
   U113 : XNOR2_X1 port map( A => n714, B => B(41), ZN => n698);
   U114 : OAI22_X1 port map( A1 => n681, A2 => n753, B1 => n685, B2 => B(30), 
                           ZN => n699);
   U115 : OAI22_X1 port map( A1 => n681, A2 => n753, B1 => n685, B2 => B(30), 
                           ZN => n682);
   U116 : XOR2_X1 port map( A => n564, B => n700, Z => SUM(32));
   U117 : XOR2_X1 port map( A => A(32), B => B(32), Z => n700);
   U118 : XNOR2_X1 port map( A => n694, B => n651, ZN => SUM(42));
   U119 : AOI21_X1 port map( B1 => n757, B2 => n676, A => n648, ZN => n703);
   U120 : AOI21_X1 port map( B1 => n757, B2 => n676, A => n677, ZN => n673);
   U121 : INV_X1 port map( A => n727, ZN => n704);
   U122 : BUF_X1 port map( A => n754, Z => n727);
   U123 : OAI22_X1 port map( A1 => n733, A2 => n727, B1 => B(29), B2 => n688, 
                           ZN => n705);
   U124 : OAI22_X1 port map( A1 => n701, A2 => n734, B1 => B(39), B2 => n659, 
                           ZN => n706);
   U125 : AND2_X1 port map( A1 => n558, A2 => net273837, ZN => n707);
   U126 : CLKBUF_X1 port map( A => n634, Z => n709);
   U127 : XNOR2_X1 port map( A => A(31), B => n710, ZN => n684);
   U128 : NAND2_X1 port map( A1 => n680, A2 => n712, ZN => n711);
   U129 : NAND2_X1 port map( A1 => n564, A2 => A(32), ZN => n712);
   U130 : AND2_X1 port map( A1 => A(36), A2 => n708, ZN => n713);
   U131 : NOR2_X1 port map( A1 => n713, A2 => n751, ZN => n664);
   U132 : AND2_X1 port map( A1 => n695, A2 => n731, ZN => n715);
   U133 : XNOR2_X1 port map( A => n709, B => n716, ZN => SUM(47));
   U134 : XNOR2_X1 port map( A => A(47), B => B(47), ZN => n716);
   U135 : INV_X1 port map( A => n686, ZN => n717);
   U136 : XOR2_X1 port map( A => n734, B => n718, Z => SUM(39));
   U137 : XOR2_X1 port map( A => A(39), B => B(39), Z => n718);
   U138 : INV_X1 port map( A => A(50), ZN => n720);
   U139 : INV_X1 port map( A => n637, ZN => n721);
   U140 : AND2_X1 port map( A1 => net264823, A2 => net270966, ZN => n722);
   U143 : BUF_X1 port map( A => A(31), Z => n723);
   U144 : OR2_X1 port map( A1 => n571, A2 => n736, ZN => n724);
   U145 : OR2_X1 port map( A1 => n752, A2 => n736, ZN => n732);
   U146 : OR2_X1 port map( A1 => n761, A2 => n649, ZN => n725);
   U147 : NAND2_X1 port map( A1 => n650, A2 => n725, ZN => n646);
   U148 : INV_X1 port map( A => n655, ZN => n728);
   U150 : OR2_X1 port map( A1 => n613, A2 => net264804, ZN => net271876);
   U151 : AND2_X1 port map( A1 => n746, A2 => n731, ZN => n729);
   U152 : OR2_X1 port map( A1 => n634, A2 => A(47), ZN => n731);
   U153 : NAND2_X1 port map( A1 => n695, A2 => n678, ZN => n631);
   U154 : BUF_X1 port map( A => n658, Z => n734);
   U155 : NAND2_X1 port map( A1 => net264823, A2 => n557, ZN => n637);
   U157 : AND2_X1 port map( A1 => A(34), A2 => n703, ZN => n736);
   U158 : NOR2_X1 port map( A1 => n736, A2 => n752, ZN => n670);
   U159 : XNOR2_X1 port map( A => n737, B => n580, ZN => SUM(56));
   U160 : XNOR2_X1 port map( A => A(56), B => B(56), ZN => n737);
   U161 : XNOR2_X1 port map( A => n738, B => n726, ZN => SUM(49));
   U162 : XNOR2_X1 port map( A => n719, B => B(49), ZN => n738);
   U163 : XNOR2_X1 port map( A => net270409, B => net274638, ZN => SUM(53));
   U164 : INV_X1 port map( A => A(40), ZN => n762);
   U165 : XNOR2_X1 port map( A => A(38), B => B(38), ZN => n663);
   U166 : XNOR2_X1 port map( A => n711, B => n739, ZN => SUM(33));
   U172 : XNOR2_X1 port map( A => A(33), B => B(33), ZN => n739);
   U173 : XNOR2_X1 port map( A => n724, B => n740, ZN => SUM(35));
   U174 : XNOR2_X1 port map( A => A(35), B => B(35), ZN => n740);
   U175 : XNOR2_X1 port map( A => n741, B => n654, ZN => SUM(37));
   U176 : XNOR2_X1 port map( A => A(37), B => B(37), ZN => n741);
   U177 : INV_X1 port map( A => A(37), ZN => n764);
   U178 : XNOR2_X1 port map( A => n742, B => A(59), ZN => SUM(59));
   U179 : XNOR2_X1 port map( A => carry_59_port, B => B(59), ZN => n742);
   U180 : XNOR2_X1 port map( A => A(36), B => B(36), ZN => n669);
   U181 : INV_X1 port map( A => A(38), ZN => n763);
   U182 : AOI21_X1 port map( B1 => n707, B2 => n758, A => n610, ZN => n600);
   U183 : XNOR2_X1 port map( A => n613, B => n615, ZN => SUM(54));
   U184 : INV_X1 port map( A => n653, ZN => n748);
   U185 : XNOR2_X1 port map( A => n633, B => n715, ZN => SUM(48));
   U186 : OR2_X1 port map( A1 => n600, A2 => A(56), ZN => n601);
   U187 : INV_X1 port map( A => A(35), ZN => n765);
   U188 : AOI21_X1 port map( B1 => n732, B2 => A(35), A => B(35), ZN => n671);
   U189 : OAI21_X1 port map( B1 => n728, B2 => A(40), A => B(40), ZN => n656);
   U190 : INV_X1 port map( A => n567, ZN => n758);
   U191 : AND2_X1 port map( A1 => n640, A2 => n743, ZN => n604);
   U192 : XNOR2_X1 port map( A => A(34), B => B(34), ZN => n675);
   U193 : AND2_X1 port map( A1 => n717, A2 => A(30), ZN => n685);
   U194 : OAI22_X1 port map( A1 => n733, A2 => n727, B1 => n688, B2 => B(29), 
                           ZN => n686);
   U195 : AND2_X1 port map( A1 => n754, A2 => A(29), ZN => n688);
   U196 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U197 : AOI21_X1 port map( B1 => A(33), B2 => n641, A => B(33), ZN => n677);
   U198 : INV_X1 port map( A => A(33), ZN => n757);
   U199 : AOI21_X1 port map( B1 => n702, B2 => A(37), A => B(37), ZN => n665);
   U200 : XNOR2_X1 port map( A => A(48), B => B(48), ZN => n633);
   U201 : INV_X1 port map( A => A(48), ZN => n759);
   U202 : OAI21_X1 port map( B1 => n729, B2 => A(48), A => B(48), ZN => n632);
   U203 : INV_X1 port map( A => A(46), ZN => n760);
   U204 : OAI21_X1 port map( B1 => n722, B2 => A(46), A => B(46), ZN => n638);
   U205 : INV_X1 port map( A => n691, ZN => n755);
   U206 : INV_X1 port map( A => n674, ZN => n752);
   U207 : INV_X1 port map( A => A(42), ZN => n761);
   U208 : OAI21_X1 port map( B1 => n747, B2 => A(42), A => B(42), ZN => n650);
   U209 : XNOR2_X1 port map( A => A(42), B => B(42), ZN => n651);
   U210 : AOI21_X1 port map( B1 => n763, B2 => n750, A => n661, ZN => n658);
   U211 : OAI21_X1 port map( B1 => B(28), B2 => A(28), A => n755, ZN => n689);
   U212 : AOI21_X1 port map( B1 => A(28), B2 => B(28), A => carry_28_port, ZN 
                           => n691);
   U213 : XNOR2_X1 port map( A => A(50), B => B(50), ZN => n627);
   U214 : XNOR2_X1 port map( A => n562, B => n645, ZN => SUM(44));
   U215 : XNOR2_X1 port map( A => n704, B => n690, ZN => SUM(29));
   U216 : OAI22_X1 port map( A1 => n701, A2 => n734, B1 => n659, B2 => B(39), 
                           ZN => n655);
   U217 : AND2_X1 port map( A1 => n658, A2 => A(39), ZN => n659);
   U218 : INV_X1 port map( A => n668, ZN => n751);
   U219 : INV_X1 port map( A => n689, ZN => n754);
   U220 : INV_X1 port map( A => n635, ZN => n746);
   U221 : INV_X1 port map( A => n649, ZN => n747);
   U222 : OAI21_X1 port map( B1 => n572, B2 => n762, A => n656, ZN => n652);
   U223 : INV_X1 port map( A => n706, ZN => n749);
   U224 : XNOR2_X1 port map( A => n627, B => n744, ZN => SUM(50));
   U225 : OAI21_X1 port map( B1 => n696, B2 => A(50), A => B(50), ZN => n626);
   U226 : OAI21_X1 port map( B1 => n719, B2 => n726, A => n745, ZN => n625);
   U227 : AOI21_X1 port map( B1 => n628, B2 => A(49), A => B(49), ZN => n629);
   U228 : INV_X1 port map( A => n723, ZN => n756);
   U229 : XNOR2_X1 port map( A => n749, B => n657, ZN => SUM(40));
   U230 : INV_X1 port map( A => n629, ZN => n745);
   U231 : OAI21_X1 port map( B1 => n631, B2 => n759, A => n632, ZN => n628);
   U232 : AOI21_X1 port map( B1 => n634, B2 => A(47), A => B(47), ZN => n635);
   U233 : XNOR2_X1 port map( A => n612, B => n707, ZN => SUM(55));
   U234 : AOI21_X1 port map( B1 => A(59), B2 => B(59), A => carry_59_port, ZN 
                           => n607);
   U235 : AOI21_X1 port map( B1 => n611, B2 => A(55), A => B(55), ZN => n610);
   U236 : OAI21_X1 port map( B1 => n693, B2 => n720, A => n626, ZN => n622);
   U237 : INV_X1 port map( A => n693, ZN => n744);
   U238 : OAI21_X1 port map( B1 => n760, B2 => n637, A => n638, ZN => n634);
   U239 : OAI21_X1 port map( B1 => n714, B2 => n735, A => n748, ZN => n649);
   U240 : AOI21_X1 port map( B1 => n652, B2 => A(41), A => B(41), ZN => n653);
   U241 : XNOR2_X1 port map( A => n568, B => n663, ZN => SUM(38));
   U242 : INV_X1 port map( A => n662, ZN => n750);
   U243 : AOI21_X1 port map( B1 => n662, B2 => A(38), A => B(38), ZN => n661);
   U244 : INV_X1 port map( A => n607, ZN => n743);
   U245 : OAI22_X1 port map( A1 => n604, A2 => B(60), B1 => n666, B2 => A(60), 
                           ZN => n602);
   U246 : XNOR2_X1 port map( A => n708, B => n669, ZN => SUM(36));
   U247 : OAI21_X1 port map( B1 => n667, B2 => A(36), A => B(36), ZN => n668);
   U248 : XNOR2_X1 port map( A => n703, B => n675, ZN => SUM(34));
   U249 : OAI21_X1 port map( B1 => n673, B2 => A(34), A => B(34), ZN => n674);
   U250 : OAI21_X1 port map( B1 => n679, B2 => A(32), A => B(32), ZN => n680);
   U251 : XNOR2_X1 port map( A => n699, B => n684, ZN => SUM(31));
   U252 : AOI21_X1 port map( B1 => n756, B2 => n559, A => n683, ZN => n679);
   U253 : INV_X1 port map( A => n705, ZN => n753);
   U254 : XNOR2_X1 port map( A => net270476, B => n621, ZN => SUM(52));
   U255 : XNOR2_X1 port map( A => n639, B => n721, ZN => SUM(46));
   U256 : XNOR2_X1 port map( A => A(46), B => B(46), ZN => n639);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT60_DW01_add_0 is

   port( A, B : in std_logic_vector (59 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (59 downto 0);  CO : out std_logic);

end RCA_NBIT60_DW01_add_0;

architecture SYN_rpl of RCA_NBIT60_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_30_port, carry_26_port, carry_25_port, carry_24_port, 
      carry_23_port, carry_22_port, carry_21_port, carry_20_port, carry_19_port
      , carry_18_port, carry_17_port, carry_16_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_10_port
      , carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, n1, n518, n519, n520, n521, 
      n523, n524, n526, n527, n529, n530, n531, n535, n536, n537, n539, n541, 
      n542, n544, n545, n547, n548, n550, n551, n553, n554, n562, n565, n566, 
      n568, n569, n571, n572, n575, n577, n586, n589, n590, n592, n593, n594, 
      n595, n596, n597, n598, n599, n601, n603, n604, n607, n609, n610, n611, 
      n612, n613, net264781, net270179, net271514, net276021, net276366, 
      net282860, net270168, n563, n559, net287631, net272173, n560, n557, n556,
      n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, 
      n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, 
      n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, 
      n513, n514, n515, n516, n517, n522, n525, n528, n532, n533, n534, n538, 
      n540, n543, n546, n549, n552, n555, n558, n561, n564, n567, n570, n573, 
      n574, n576, n578, n579, n580, n581, n582, n583, n584, n585, n587, n588, 
      n591, n600, n602, n605, n606, n608, n614, n615, n616, n617, n618, n619, 
      n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, 
      n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, 
      n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, 
      n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, 
      n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, 
      n680, n681, n682, n683, n684, n685, n686, n687, n688 : std_logic;

begin
   
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U167 : XOR2_X1 port map( A => n609, B => n584, Z => SUM(28));
   U169 : XOR2_X1 port map( A => n641, B => n612, Z => SUM(27));
   U170 : XOR2_X1 port map( A => carry_26_port, B => n613, Z => SUM(26));
   U171 : XOR2_X1 port map( A => A(26), B => B(26), Z => n613);
   U172 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : CLKBUF_X1 port map( A => A(33), Z => n477);
   U2 : CLKBUF_X1 port map( A => n649, Z => n478);
   U3 : CLKBUF_X1 port map( A => A(49), Z => n616);
   U4 : BUF_X1 port map( A => A(37), Z => n479);
   U5 : AOI21_X1 port map( B1 => n631, B2 => n588, A => B(50), ZN => n480);
   U6 : OAI21_X1 port map( B1 => n573, B2 => n481, A => n538, ZN => n577);
   U7 : AOI21_X1 port map( B1 => n631, B2 => n588, A => B(50), ZN => n548);
   U8 : BUF_X1 port map( A => n490, Z => net276021);
   U9 : INV_X1 port map( A => B(29), ZN => n585);
   U10 : INV_X1 port map( A => B(39), ZN => n546);
   U11 : AND2_X1 port map( A1 => A(39), A2 => B(39), ZN => n481);
   U12 : BUF_X1 port map( A => n568, Z => n606);
   U13 : AND2_X2 port map( A1 => n555, A2 => n558, ZN => n482);
   U14 : BUF_X1 port map( A => n675, Z => n483);
   U15 : BUF_X1 port map( A => A(52), Z => n649);
   U16 : BUF_X1 port map( A => A(53), Z => n488);
   U17 : CLKBUF_X1 port map( A => A(35), Z => n484);
   U18 : XNOR2_X1 port map( A => n485, B => n482, ZN => SUM(38));
   U19 : XNOR2_X1 port map( A => A(38), B => n570, ZN => n485);
   U20 : INV_X1 port map( A => n685, ZN => n486);
   U21 : INV_X1 port map( A => B(42), ZN => n489);
   U22 : CLKBUF_X1 port map( A => n565, Z => n487);
   U23 : BUF_X1 port map( A => A(47), Z => n507);
   U24 : XNOR2_X1 port map( A => A(42), B => n489, ZN => n661);
   U25 : BUF_X1 port map( A => A(54), Z => n644);
   U26 : AND2_X1 port map( A1 => n567, A2 => n564, ZN => n490);
   U27 : OR2_X1 port map( A1 => n519, A2 => A(28), ZN => n520);
   U28 : CLKBUF_X1 port map( A => n559, Z => net282860);
   U29 : CLKBUF_X1 port map( A => A(48), Z => n510);
   U30 : NOR2_X1 port map( A1 => n480, A2 => n579, ZN => n491);
   U31 : AOI22_X1 port map( A1 => n650, A2 => B(51), B1 => n544, B2 => n545, ZN
                           => n492);
   U32 : INV_X1 port map( A => B(55), ZN => n498);
   U33 : INV_X1 port map( A => B(28), ZN => n637);
   U34 : INV_X1 port map( A => B(52), ZN => n629);
   U35 : NOR2_X1 port map( A1 => n494, A2 => n495, ZN => n493);
   U36 : NOR2_X1 port map( A1 => n541, A2 => B(52), ZN => n494);
   U37 : NOR2_X1 port map( A1 => n478, A2 => n514, ZN => n495);
   U38 : BUF_X1 port map( A => n670, Z => n514);
   U39 : INV_X1 port map( A => B(48), ZN => n506);
   U40 : INV_X1 port map( A => B(38), ZN => n570);
   U41 : OAI21_X1 port map( B1 => n497, B2 => n486, A => B(55), ZN => n496);
   U42 : AND2_X1 port map( A1 => n591, A2 => n669, ZN => n497);
   U43 : INV_X1 port map( A => B(44), ZN => n653);
   U44 : INV_X1 port map( A => B(53), ZN => n605);
   U45 : INV_X1 port map( A => B(36), ZN => n623);
   U46 : INV_X1 port map( A => B(46), ZN => n508);
   U47 : OAI21_X1 port map( B1 => n627, B2 => A(44), A => B(44), ZN => n566);
   U48 : XNOR2_X1 port map( A => n651, B => n491, ZN => SUM(51));
   U49 : BUF_X1 port map( A => A(36), Z => n499);
   U50 : XNOR2_X1 port map( A => n504, B => n511, ZN => SUM(48));
   U51 : XNOR2_X1 port map( A => A(48), B => n506, ZN => n504);
   U52 : OAI21_X1 port map( B1 => n507, B2 => n512, A => n503, ZN => n511);
   U53 : OR2_X1 port map( A1 => n511, A2 => n501, ZN => net271514);
   U54 : INV_X1 port map( A => n557, ZN => n503);
   U55 : OAI21_X1 port map( B1 => n507, B2 => n512, A => n503, ZN => n553);
   U56 : AOI21_X1 port map( B1 => A(47), B2 => n556, A => B(47), ZN => n557);
   U57 : NAND2_X1 port map( A1 => net272173, A2 => n560, ZN => n556);
   U58 : OAI21_X1 port map( B1 => n502, B2 => n509, A => B(46), ZN => n560);
   U59 : CLKBUF_X1 port map( A => A(46), Z => n509);
   U60 : OAI21_X1 port map( B1 => n502, B2 => n509, A => B(46), ZN => net287631
                           );
   U61 : INV_X1 port map( A => n559, ZN => n502);
   U62 : INV_X1 port map( A => A(48), ZN => n501);
   U63 : OAI21_X1 port map( B1 => net264781, B2 => n510, A => B(48), ZN => 
                           net276366);
   U64 : OAI21_X1 port map( B1 => net264781, B2 => n510, A => B(48), ZN => n554
                           );
   U65 : XNOR2_X1 port map( A => A(47), B => B(47), ZN => n505);
   U66 : NAND2_X1 port map( A1 => net272173, A2 => net287631, ZN => n512);
   U67 : XNOR2_X1 port map( A => A(46), B => n508, ZN => net270168);
   U68 : INV_X1 port map( A => A(46), ZN => n500);
   U69 : OR2_X1 port map( A1 => n559, A2 => n500, ZN => net272173);
   U70 : XNOR2_X1 port map( A => n505, B => n512, ZN => SUM(47));
   U71 : NAND2_X1 port map( A1 => n591, A2 => n669, ZN => n513);
   U72 : BUF_X1 port map( A => n562, Z => n522);
   U73 : OR2_X1 port map( A1 => n513, A2 => n685, ZN => n515);
   U74 : NAND2_X1 port map( A1 => n515, A2 => n496, ZN => n529);
   U75 : XNOR2_X1 port map( A => net282860, B => net270168, ZN => SUM(46));
   U76 : OAI21_X1 port map( B1 => n525, B2 => n522, A => n516, ZN => n559);
   U77 : INV_X1 port map( A => n563, ZN => n516);
   U78 : AOI21_X1 port map( B1 => A(45), B2 => n562, A => B(45), ZN => n563);
   U79 : XNOR2_X1 port map( A => n517, B => n522, ZN => SUM(45));
   U80 : CLKBUF_X1 port map( A => A(45), Z => n525);
   U81 : XNOR2_X1 port map( A => A(45), B => B(45), ZN => n517);
   U82 : BUF_X1 port map( A => n676, Z => n581);
   U83 : OAI22_X1 port map( A1 => n624, A2 => net276021, B1 => n575, B2 => 
                           B(41), ZN => n528);
   U84 : BUF_X1 port map( A => n519, Z => n584);
   U85 : NAND2_X1 port map( A1 => A(38), A2 => B(38), ZN => n534);
   U86 : NOR2_X1 port map( A1 => A(38), A2 => B(38), ZN => n533);
   U87 : INV_X1 port map( A => A(39), ZN => n543);
   U88 : INV_X1 port map( A => A(40), ZN => n540);
   U89 : XNOR2_X1 port map( A => A(37), B => B(37), ZN => n552);
   U90 : OAI21_X1 port map( B1 => B(37), B2 => n479, A => n586, ZN => n555);
   U91 : NAND2_X1 port map( A1 => n479, A2 => B(37), ZN => n558);
   U92 : NAND2_X1 port map( A1 => n540, A2 => n577, ZN => n564);
   U93 : OAI21_X1 port map( B1 => n540, B2 => n577, A => n561, ZN => n567);
   U94 : XNOR2_X1 port map( A => n549, B => n543, ZN => SUM(39));
   U95 : XNOR2_X1 port map( A => n532, B => n546, ZN => n549);
   U96 : INV_X1 port map( A => B(40), ZN => n561);
   U97 : XNOR2_X1 port map( A => A(40), B => n561, ZN => net270179);
   U98 : XNOR2_X1 port map( A => n552, B => n586, ZN => SUM(37));
   U99 : OAI21_X1 port map( B1 => n533, B2 => n482, A => n534, ZN => n532);
   U100 : CLKBUF_X1 port map( A => n532, Z => n573);
   U101 : NAND2_X1 port map( A1 => n543, A2 => n546, ZN => n538);
   U102 : AOI22_X1 port map( A1 => n584, A2 => n630, B1 => n520, B2 => B(28), 
                           ZN => n574);
   U103 : XNOR2_X1 port map( A => n576, B => n587, ZN => SUM(29));
   U104 : XNOR2_X1 port map( A => A(29), B => B(29), ZN => n576);
   U105 : AND2_X1 port map( A1 => n632, A2 => n668, ZN => n578);
   U106 : AND2_X1 port map( A1 => n688, A2 => n547, ZN => n579);
   U107 : NOR2_X1 port map( A1 => n548, A2 => n579, ZN => n545);
   U108 : NOR2_X1 port map( A1 => n607, A2 => n580, ZN => n636);
   U109 : NOR2_X1 port map( A1 => B(30), A2 => A(30), ZN => n580);
   U110 : NAND3_X1 port map( A1 => n620, A2 => n621, A3 => n622, ZN => n582);
   U111 : INV_X1 port map( A => n679, ZN => n583);
   U112 : OR2_X1 port map( A1 => n574, A2 => n585, ZN => n621);
   U113 : CLKBUF_X1 port map( A => n678, Z => n587);
   U114 : INV_X1 port map( A => n688, ZN => n588);
   U115 : BUF_X1 port map( A => n595, Z => n615);
   U116 : OR2_X1 port map( A1 => n608, A2 => n644, ZN => n591);
   U117 : OAI21_X1 port map( B1 => n493, B2 => n488, A => B(53), ZN => n600);
   U118 : OAI22_X1 port map( A1 => n484, A2 => n483, B1 => B(35), B2 => n592, 
                           ZN => n602);
   U119 : XNOR2_X1 port map( A => A(53), B => n605, ZN => n658);
   U120 : NAND2_X1 port map( A1 => n619, A2 => n539, ZN => n608);
   U121 : XNOR2_X1 port map( A => n675, B => n594, ZN => SUM(35));
   U122 : XNOR2_X1 port map( A => n521, B => n614, ZN => SUM(59));
   U123 : XOR2_X1 port map( A => B(59), B => A(59), Z => n614);
   U124 : OAI22_X1 port map( A1 => n478, A2 => n514, B1 => n541, B2 => B(52), 
                           ZN => n617);
   U125 : CLKBUF_X1 port map( A => A(30), Z => n634);
   U126 : CLKBUF_X1 port map( A => A(34), Z => n618);
   U127 : OR2_X1 port map( A1 => n617, A2 => n687, ZN => n619);
   U128 : NAND2_X1 port map( A1 => n600, A2 => n619, ZN => n535);
   U129 : NAND2_X1 port map( A1 => A(29), A2 => n678, ZN => n620);
   U130 : NAND2_X1 port map( A1 => A(29), A2 => B(29), ZN => n622);
   U131 : NAND3_X1 port map( A1 => n620, A2 => n621, A3 => n622, ZN => 
                           carry_30_port);
   U132 : XNOR2_X1 port map( A => A(36), B => n623, ZN => n657);
   U133 : CLKBUF_X1 port map( A => A(41), Z => n624);
   U134 : CLKBUF_X1 port map( A => A(32), Z => n625);
   U135 : XNOR2_X1 port map( A => n542, B => n626, ZN => SUM(52));
   U136 : XNOR2_X1 port map( A => A(52), B => n629, ZN => n626);
   U137 : AND2_X1 port map( A1 => n672, A2 => n639, ZN => n627);
   U138 : NAND2_X1 port map( A1 => net276366, A2 => net271514, ZN => n628);
   U139 : CLKBUF_X1 port map( A => A(28), Z => n630);
   U140 : AND2_X1 port map( A1 => n671, A2 => n642, ZN => n631);
   U141 : OR2_X1 port map( A1 => n647, A2 => n529, ZN => n632);
   U142 : NAND2_X1 port map( A1 => n632, A2 => n668, ZN => n526);
   U143 : CLKBUF_X1 port map( A => A(56), Z => n647);
   U144 : INV_X1 port map( A => n676, ZN => n633);
   U145 : CLKBUF_X1 port map( A => A(31), Z => n635);
   U146 : XNOR2_X1 port map( A => A(28), B => n637, ZN => n609);
   U147 : BUF_X1 port map( A => A(57), Z => n648);
   U148 : XNOR2_X1 port map( A => n526, B => n638, ZN => SUM(57));
   U149 : XOR2_X1 port map( A => A(57), B => B(57), Z => n638);
   U150 : OAI22_X1 port map( A1 => n624, A2 => net276021, B1 => n575, B2 => 
                           B(41), ZN => n571);
   U151 : OR2_X1 port map( A1 => n568, A2 => A(43), ZN => n639);
   U152 : NAND2_X1 port map( A1 => n672, A2 => n639, ZN => n565);
   U153 : OAI22_X1 port map( A1 => n484, A2 => n483, B1 => n592, B2 => B(35), 
                           ZN => n589);
   U154 : OR2_X1 port map( A1 => A(58), A2 => n523, ZN => n640);
   U155 : NAND2_X1 port map( A1 => n667, A2 => n640, ZN => n521);
   U156 : CLKBUF_X1 port map( A => n679, Z => n641);
   U157 : NAND2_X1 port map( A1 => n554, A2 => net271514, ZN => n550);
   U158 : OR2_X1 port map( A1 => n550, A2 => n616, ZN => n642);
   U159 : NAND2_X1 port map( A1 => n671, A2 => n642, ZN => n547);
   U160 : XNOR2_X1 port map( A => n615, B => n597, ZN => SUM(34));
   U161 : XNOR2_X1 port map( A => n523, B => n643, ZN => SUM(58));
   U162 : XNOR2_X1 port map( A => B(58), B => A(58), ZN => n643);
   U163 : BUF_X1 port map( A => n677, Z => n645);
   U164 : XOR2_X1 port map( A => A(50), B => B(50), Z => n665);
   U165 : BUF_X1 port map( A => n636, Z => n646);
   U166 : CLKBUF_X1 port map( A => A(51), Z => n650);
   U168 : XNOR2_X1 port map( A => A(51), B => B(51), ZN => n651);
   U173 : OR2_X1 port map( A1 => n565, A2 => n684, ZN => n652);
   U174 : NAND2_X1 port map( A1 => n566, A2 => n652, ZN => n562);
   U175 : XNOR2_X1 port map( A => A(55), B => n498, ZN => n666);
   U176 : XNOR2_X1 port map( A => A(44), B => n653, ZN => n662);
   U177 : XNOR2_X1 port map( A => n654, B => n606, ZN => SUM(43));
   U178 : XNOR2_X1 port map( A => A(43), B => B(43), ZN => n654);
   U179 : XNOR2_X1 port map( A => net276021, B => n655, ZN => SUM(41));
   U180 : XNOR2_X1 port map( A => A(41), B => B(41), ZN => n655);
   U181 : INV_X1 port map( A => A(50), ZN => n688);
   U182 : XNOR2_X1 port map( A => A(35), B => B(35), ZN => n594);
   U183 : INV_X1 port map( A => n553, ZN => net264781);
   U184 : XNOR2_X1 port map( A => n656, B => n634, ZN => SUM(30));
   U185 : XNOR2_X1 port map( A => n582, B => B(30), ZN => n656);
   U186 : XNOR2_X1 port map( A => n657, B => n602, ZN => SUM(36));
   U187 : XNOR2_X1 port map( A => n658, B => n617, ZN => SUM(53));
   U188 : XNOR2_X1 port map( A => A(34), B => B(34), ZN => n597);
   U189 : XNOR2_X1 port map( A => net270179, B => n577, ZN => SUM(40));
   U190 : XNOR2_X1 port map( A => n659, B => n581, ZN => SUM(33));
   U191 : XNOR2_X1 port map( A => A(33), B => B(33), ZN => n659);
   U192 : XNOR2_X1 port map( A => n660, B => n628, ZN => SUM(49));
   U193 : XNOR2_X1 port map( A => A(49), B => B(49), ZN => n660);
   U194 : XNOR2_X1 port map( A => n661, B => n528, ZN => SUM(42));
   U195 : XNOR2_X1 port map( A => n662, B => n487, ZN => SUM(44));
   U196 : XNOR2_X1 port map( A => n645, B => n663, ZN => SUM(32));
   U197 : XNOR2_X1 port map( A => A(32), B => B(32), ZN => n663);
   U198 : INV_X1 port map( A => n569, ZN => n672);
   U199 : XNOR2_X1 port map( A => n646, B => n664, ZN => SUM(31));
   U200 : XNOR2_X1 port map( A => A(31), B => B(31), ZN => n664);
   U201 : OAI22_X1 port map( A1 => n645, A2 => n625, B1 => n601, B2 => B(32), 
                           ZN => n598);
   U202 : AND2_X1 port map( A1 => n677, A2 => A(32), ZN => n601);
   U203 : AOI22_X1 port map( A1 => n650, A2 => B(51), B1 => n544, B2 => n491, 
                           ZN => n542);
   U204 : OR2_X1 port map( A1 => A(51), A2 => B(51), ZN => n544);
   U205 : INV_X1 port map( A => n551, ZN => n671);
   U206 : AOI21_X1 port map( B1 => n550, B2 => n616, A => B(49), ZN => n551);
   U207 : XNOR2_X1 port map( A => n665, B => n547, ZN => SUM(50));
   U208 : AOI21_X1 port map( B1 => A(30), B2 => B(30), A => carry_30_port, ZN 
                           => n607);
   U209 : INV_X1 port map( A => A(53), ZN => n687);
   U210 : AND2_X1 port map( A1 => n675, A2 => A(35), ZN => n592);
   U211 : XNOR2_X1 port map( A => B(27), B => n680, ZN => n612);
   U212 : XNOR2_X1 port map( A => n666, B => n513, ZN => SUM(55));
   U213 : XNOR2_X1 port map( A => n529, B => n531, ZN => SUM(56));
   U214 : XNOR2_X1 port map( A => A(56), B => B(56), ZN => n531);
   U215 : INV_X1 port map( A => n530, ZN => n668);
   U216 : AOI21_X1 port map( B1 => n529, B2 => n647, A => B(56), ZN => n530);
   U217 : INV_X1 port map( A => n518, ZN => n678);
   U218 : INV_X1 port map( A => n610, ZN => n679);
   U219 : AOI22_X1 port map( A1 => n613, A2 => carry_26_port, B1 => A(26), B2 
                           => B(26), ZN => n610);
   U220 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U221 : INV_X1 port map( A => n477, ZN => n681);
   U222 : XNOR2_X1 port map( A => A(54), B => B(54), ZN => n537);
   U223 : INV_X1 port map( A => A(44), ZN => n684);
   U224 : INV_X1 port map( A => n593, ZN => n675);
   U225 : OAI21_X1 port map( B1 => n578, B2 => n648, A => B(57), ZN => n527);
   U226 : OAI21_X1 port map( B1 => n583, B2 => n680, A => n611, ZN => n519);
   U227 : INV_X1 port map( A => A(42), ZN => n683);
   U228 : OAI21_X1 port map( B1 => n673, B2 => A(42), A => B(42), ZN => n572);
   U229 : AOI21_X1 port map( B1 => n676, B2 => A(33), A => B(33), ZN => n599);
   U230 : INV_X1 port map( A => n648, ZN => n686);
   U231 : INV_X1 port map( A => A(55), ZN => n685);
   U232 : INV_X1 port map( A => n524, ZN => n667);
   U233 : INV_X1 port map( A => n492, ZN => n670);
   U234 : INV_X1 port map( A => n603, ZN => n677);
   U235 : INV_X1 port map( A => A(27), ZN => n680);
   U236 : OAI21_X1 port map( B1 => A(27), B2 => n679, A => B(27), ZN => n611);
   U237 : OAI22_X1 port map( A1 => n635, A2 => n646, B1 => n604, B2 => B(31), 
                           ZN => n603);
   U238 : AND2_X1 port map( A1 => A(31), A2 => n636, ZN => n604);
   U239 : XNOR2_X1 port map( A => n537, B => n608, ZN => SUM(54));
   U240 : AOI21_X1 port map( B1 => n535, B2 => n644, A => B(54), ZN => n536);
   U241 : AOI21_X1 port map( B1 => n568, B2 => A(43), A => B(43), ZN => n569);
   U242 : OAI21_X1 port map( B1 => n528, B2 => n683, A => n572, ZN => n568);
   U243 : INV_X1 port map( A => n571, ZN => n673);
   U244 : AND2_X1 port map( A1 => A(41), A2 => n490, ZN => n575);
   U245 : OAI21_X1 port map( B1 => n602, B2 => n682, A => n590, ZN => n586);
   U246 : INV_X1 port map( A => n589, ZN => n674);
   U247 : OAI22_X1 port map( A1 => n618, A2 => n615, B1 => n596, B2 => B(34), 
                           ZN => n593);
   U248 : AND2_X1 port map( A1 => n595, A2 => A(34), ZN => n596);
   U249 : AOI21_X1 port map( B1 => n681, B2 => n633, A => n599, ZN => n595);
   U250 : INV_X1 port map( A => n598, ZN => n676);
   U251 : AOI22_X1 port map( A1 => n584, A2 => n630, B1 => n520, B2 => B(28), 
                           ZN => n518);
   U252 : OAI21_X1 port map( B1 => n674, B2 => n499, A => B(36), ZN => n590);
   U253 : INV_X1 port map( A => n499, ZN => n682);
   U254 : AOI21_X1 port map( B1 => n523, B2 => A(58), A => B(58), ZN => n524);
   U255 : OAI21_X1 port map( B1 => n526, B2 => n686, A => n527, ZN => n523);
   U256 : INV_X1 port map( A => n536, ZN => n669);
   U257 : OAI21_X1 port map( B1 => n493, B2 => n488, A => B(53), ZN => n539);
   U258 : AND2_X1 port map( A1 => n670, A2 => n649, ZN => n541);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT58_DW01_add_0 is

   port( A, B : in std_logic_vector (57 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (57 downto 0);  CO : out std_logic);

end RCA_NBIT58_DW01_add_0;

architecture SYN_rpl of RCA_NBIT58_DW01_add_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_24_port, carry_23_port, carry_22_port, carry_21_port, 
      carry_20_port, carry_19_port, carry_18_port, carry_17_port, carry_16_port
      , carry_15_port, carry_14_port, carry_13_port, carry_12_port, 
      carry_11_port, carry_10_port, carry_9_port, carry_8_port, carry_7_port, 
      carry_6_port, carry_5_port, carry_4_port, carry_3_port, carry_2_port, n1,
      n634, n635, n636, n637, n640, n652, n655, n675, n680, n691, n694, n708, 
      n711, n712, n714, n715, n717, n718, n719, n720, n721, n723, n724, n726, 
      n728, n729, n730, n731, n732, n733, net264713, net264718, net264731, 
      net270178, net270359, net270357, net270356, net270380, net270418, 
      net270569, net270590, net270617, net270890, net270933, net271088, 
      net271108, net271730, net272145, net272205, net272493, net272567, 
      net272615, net272904, net273379, net274336, net275467, net276035, 
      net276072, net276358, net276651, net276658, n709, n706, n705, n702, 
      net274074, net272360, n703, n699, n697, n696, n693, net276422, net270155,
      net296107, net264735, n679, n678, n658, n657, net270765, n676, n673, n672
      , net270360, net264719, n669, n661, net296154, net296099, net273368, 
      net271767, net271520, net270891, net270889, net270413, net270410, 
      net264739, net264715, n670, n667, n666, n664, n663, n660, net271467, 
      net270892, net264712, n685, n684, n682, n681, n590, n591, n592, n593, 
      n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, 
      n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, 
      n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, 
      n630, n631, n632, n633, n638, n639, n641, n642, n643, n644, n645, n646, 
      n647, n648, n649, n650, n651, n653, n654, n656, n659, n662, n665, n668, 
      n671, n674, n677, n683, n686, n687, n688, n689, n690, n692, n695, n698, 
      n700, n701, n704, n707, n710, n713, n716, n722, n725, n727, n734, n735, 
      n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, 
      n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, 
      n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, 
      n772, n773 : std_logic;

begin
   
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U115 : XOR2_X1 port map( A => B(57), B => A(57), Z => n635);
   U176 : XOR2_X1 port map( A => n747, B => n731, Z => SUM(25));
   U177 : XOR2_X1 port map( A => B(25), B => n737, Z => n731);
   U178 : XOR2_X1 port map( A => n704, B => n733, Z => SUM(24));
   U179 : XOR2_X1 port map( A => carry_24_port, B => B(24), Z => n733);
   U180 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : OAI21_X1 port map( B1 => n609, B2 => n596, A => B(48), ZN => n590);
   U2 : CLKBUF_X1 port map( A => n675, Z => n597);
   U3 : CLKBUF_X1 port map( A => A(42), Z => n591);
   U4 : BUF_X1 port map( A => n681, Z => net271467);
   U5 : INV_X1 port map( A => B(55), ZN => n625);
   U6 : BUF_X1 port map( A => n702, Z => net272567);
   U7 : CLKBUF_X1 port map( A => n726, Z => n698);
   U8 : CLKBUF_X1 port map( A => net270889, Z => n592);
   U9 : XNOR2_X1 port map( A => n755, B => n593, ZN => SUM(39));
   U10 : XOR2_X1 port map( A => A(39), B => n700, Z => n593);
   U11 : CLKBUF_X1 port map( A => n714, Z => n746);
   U12 : CLKBUF_X1 port map( A => n668, Z => net272145);
   U13 : CLKBUF_X1 port map( A => A(35), Z => n683);
   U14 : OAI21_X1 port map( B1 => n746, B2 => n743, A => n765, ZN => n594);
   U15 : BUF_X1 port map( A => A(28), Z => n606);
   U16 : CLKBUF_X1 port map( A => n604, Z => net276358);
   U17 : INV_X1 port map( A => n711, ZN => n595);
   U18 : CLKBUF_X1 port map( A => A(48), Z => n596);
   U19 : AND2_X1 port map( A1 => n602, A2 => n651, ZN => n598);
   U20 : OR2_X1 port map( A1 => net276072, A2 => net264718, ZN => net270890);
   U21 : NAND2_X1 port map( A1 => n763, A2 => n599, ZN => n615);
   U22 : NOR2_X1 port map( A1 => n619, A2 => n618, ZN => n599);
   U23 : BUF_X1 port map( A => net296107, Z => n639);
   U24 : NAND2_X1 port map( A1 => n600, A2 => n601, ZN => n602);
   U25 : INV_X1 port map( A => n654, ZN => n600);
   U26 : INV_X1 port map( A => n611, ZN => n601);
   U27 : CLKBUF_X1 port map( A => A(49), Z => n654);
   U28 : BUF_X1 port map( A => n669, Z => net270889);
   U29 : CLKBUF_X1 port map( A => net272360, Z => net274074);
   U30 : BUF_X1 port map( A => A(51), Z => net270590);
   U31 : OR2_X1 port map( A1 => n660, A2 => net264715, ZN => net270359);
   U32 : OR2_X1 port map( A1 => net276658, A2 => net270590, ZN => net270356);
   U33 : OR2_X1 port map( A1 => n691, A2 => n757, ZN => n742);
   U34 : INV_X1 port map( A => B(43), ZN => net272493);
   U35 : INV_X1 port map( A => B(39), ZN => n700);
   U36 : INV_X1 port map( A => net270356, ZN => n618);
   U37 : INV_X1 port map( A => B(53), ZN => n620);
   U38 : INV_X1 port map( A => B(27), ZN => n756);
   U39 : INV_X1 port map( A => B(50), ZN => n653);
   U40 : INV_X1 port map( A => B(46), ZN => net270413);
   U41 : INV_X1 port map( A => B(48), ZN => net273368);
   U42 : INV_X1 port map( A => B(29), ZN => n758);
   U43 : INV_X1 port map( A => B(42), ZN => n659);
   U44 : NOR3_X1 port map( A1 => A(38), A2 => net272205, A3 => net264731, ZN =>
                           n757);
   U45 : NAND2_X1 port map( A1 => n706, A2 => n689, ZN => n702);
   U46 : NOR2_X1 port map( A1 => n673, A2 => net270765, ZN => n669);
   U47 : AOI21_X1 port map( B1 => n741, B2 => n610, A => B(38), ZN => n691);
   U48 : XNOR2_X1 port map( A => n603, B => net271467, ZN => SUM(41));
   U49 : AOI22_X1 port map( A1 => net271467, A2 => n605, B1 => n682, B2 => 
                           B(41), ZN => n678);
   U50 : XNOR2_X1 port map( A => A(41), B => B(41), ZN => n603);
   U51 : NOR2_X1 port map( A1 => n685, A2 => net270892, ZN => n681);
   U52 : OR2_X1 port map( A1 => n681, A2 => A(41), ZN => n682);
   U53 : AND2_X1 port map( A1 => net264712, A2 => n684, ZN => net270892);
   U54 : NOR2_X1 port map( A1 => net271108, A2 => net274336, ZN => n684);
   U55 : INV_X1 port map( A => A(40), ZN => net264712);
   U56 : AOI21_X1 port map( B1 => n604, B2 => A(40), A => B(40), ZN => n685);
   U57 : CLKBUF_X1 port map( A => A(41), Z => n605);
   U58 : OR2_X1 port map( A1 => net274336, A2 => net271108, ZN => n604);
   U59 : XNOR2_X1 port map( A => A(40), B => B(40), ZN => net273379);
   U60 : XNOR2_X1 port map( A => net271767, B => n660, ZN => SUM(48));
   U61 : XNOR2_X1 port map( A => A(48), B => net273368, ZN => net271767);
   U62 : NAND2_X1 port map( A1 => n608, A2 => net270891, ZN => n660);
   U63 : INV_X1 port map( A => n664, ZN => n608);
   U64 : AND2_X1 port map( A1 => n608, A2 => net270891, ZN => n609);
   U65 : AOI21_X1 port map( B1 => n663, B2 => A(47), A => B(47), ZN => n664);
   U66 : NAND2_X1 port map( A1 => n667, A2 => net270360, ZN => n663);
   U67 : OAI21_X1 port map( B1 => net264739, B2 => net296154, A => B(46), ZN =>
                           n667);
   U68 : CLKBUF_X1 port map( A => A(46), Z => net296154);
   U69 : OAI21_X1 port map( B1 => net264739, B2 => net296154, A => B(46), ZN =>
                           net296099);
   U70 : INV_X1 port map( A => n666, ZN => net264739);
   U71 : OAI21_X1 port map( B1 => net271520, B2 => net270889, A => n607, ZN => 
                           n666);
   U72 : INV_X1 port map( A => n670, ZN => n607);
   U73 : OAI21_X1 port map( B1 => net271520, B2 => n592, A => n607, ZN => 
                           net276422);
   U74 : AOI21_X1 port map( B1 => n669, B2 => A(45), A => B(45), ZN => n670);
   U75 : XNOR2_X1 port map( A => net270889, B => net270410, ZN => SUM(45));
   U76 : CLKBUF_X1 port map( A => A(45), Z => net271520);
   U77 : OAI21_X1 port map( B1 => n609, B2 => n596, A => B(48), ZN => n661);
   U78 : INV_X1 port map( A => A(48), ZN => net264715);
   U79 : XNOR2_X1 port map( A => B(47), B => A(47), ZN => net270617);
   U80 : OR2_X1 port map( A1 => net276651, A2 => A(47), ZN => net270891);
   U81 : NAND2_X1 port map( A1 => net296099, A2 => net270360, ZN => net276651);
   U82 : INV_X1 port map( A => A(46), ZN => net264719);
   U83 : XNOR2_X1 port map( A => A(46), B => net270413, ZN => net270155);
   U84 : XNOR2_X1 port map( A => A(45), B => B(45), ZN => net270410);
   U85 : BUF_X1 port map( A => A(38), Z => n610);
   U86 : NAND2_X1 port map( A1 => n590, A2 => net270359, ZN => n611);
   U87 : NAND2_X1 port map( A1 => n627, A2 => B(52), ZN => n616);
   U88 : AOI21_X1 port map( B1 => n644, B2 => A(55), A => B(55), ZN => n640);
   U89 : INV_X1 port map( A => A(55), ZN => n621);
   U90 : CLKBUF_X1 port map( A => A(53), Z => n612);
   U91 : XNOR2_X1 port map( A => n672, B => n613, ZN => SUM(44));
   U92 : XOR2_X1 port map( A => A(44), B => B(44), Z => n613);
   U93 : NOR2_X1 port map( A1 => B(54), A2 => A(54), ZN => n633);
   U94 : NAND2_X1 port map( A1 => A(54), A2 => B(54), ZN => n632);
   U95 : NAND2_X1 port map( A1 => n630, A2 => n629, ZN => n631);
   U96 : AOI21_X1 port map( B1 => n631, B2 => n632, A => n633, ZN => n638);
   U97 : XNOR2_X1 port map( A => n638, B => n625, ZN => n623);
   U98 : INV_X1 port map( A => n644, ZN => net275467);
   U99 : XNOR2_X1 port map( A => n624, B => n642, ZN => SUM(54));
   U100 : NAND2_X1 port map( A1 => n615, A2 => n616, ZN => n614);
   U101 : NAND2_X1 port map( A1 => n615, A2 => n616, ZN => n641);
   U102 : INV_X1 port map( A => A(52), ZN => n619);
   U103 : AOI21_X1 port map( B1 => n643, B2 => n639, A => B(51), ZN => n617);
   U104 : OAI21_X1 port map( B1 => n617, B2 => n618, A => n619, ZN => n627);
   U105 : XNOR2_X1 port map( A => A(54), B => B(54), ZN => n624);
   U106 : NAND2_X1 port map( A1 => n614, A2 => B(53), ZN => n628);
   U107 : NAND2_X1 port map( A1 => n628, A2 => n626, ZN => n629);
   U108 : NAND2_X1 port map( A1 => n620, A2 => n645, ZN => n630);
   U109 : AND2_X1 port map( A1 => n629, A2 => n630, ZN => n642);
   U110 : XNOR2_X1 port map( A => A(53), B => B(53), ZN => n622);
   U111 : INV_X1 port map( A => n612, ZN => n626);
   U112 : CLKBUF_X1 port map( A => net270590, Z => n643);
   U113 : AOI21_X1 port map( B1 => n631, B2 => n632, A => n633, ZN => n644);
   U114 : XNOR2_X1 port map( A => n622, B => n641, ZN => SUM(53));
   U116 : XNOR2_X1 port map( A => n623, B => n621, ZN => SUM(55));
   U117 : AND2_X1 port map( A1 => n615, A2 => n616, ZN => n645);
   U118 : NAND2_X1 port map( A1 => net270359, A2 => n661, ZN => n657);
   U119 : OR2_X1 port map( A1 => n666, A2 => net264719, ZN => net270360);
   U120 : AND2_X1 port map( A1 => n672, A2 => n646, ZN => net270765);
   U121 : INV_X1 port map( A => A(44), ZN => n646);
   U122 : INV_X1 port map( A => n646, ZN => n649);
   U123 : AOI21_X1 port map( B1 => n650, B2 => n649, A => B(44), ZN => n673);
   U124 : OR2_X1 port map( A1 => n647, A2 => n648, ZN => n650);
   U125 : INV_X1 port map( A => n676, ZN => n647);
   U126 : NOR2_X1 port map( A1 => n647, A2 => n648, ZN => n672);
   U127 : OAI21_X1 port map( B1 => n675, B2 => A(43), A => B(43), ZN => n676);
   U128 : XOR2_X1 port map( A => A(43), B => net272493, Z => net276035);
   U129 : AND2_X1 port map( A1 => n675, A2 => A(43), ZN => n648);
   U130 : OAI21_X1 port map( B1 => n598, B2 => A(50), A => B(50), ZN => n656);
   U131 : NAND2_X1 port map( A1 => net270890, A2 => n656, ZN => net276658);
   U132 : OAI21_X1 port map( B1 => n598, B2 => A(50), A => B(50), ZN => n655);
   U133 : INV_X1 port map( A => n658, ZN => n651);
   U134 : OAI21_X1 port map( B1 => n654, B2 => n611, A => n651, ZN => net276072
                           );
   U135 : AOI21_X1 port map( B1 => n657, B2 => A(49), A => B(49), ZN => n658);
   U136 : XNOR2_X1 port map( A => net270418, B => n611, ZN => SUM(49));
   U137 : XNOR2_X1 port map( A => A(50), B => n653, ZN => net270380);
   U138 : INV_X1 port map( A => A(50), ZN => net264718);
   U139 : AOI21_X1 port map( B1 => net264735, B2 => A(42), A => B(42), ZN => 
                           n679);
   U140 : AOI21_X1 port map( B1 => net270357, B2 => net264713, A => n679, ZN =>
                           n675);
   U141 : INV_X1 port map( A => n678, ZN => net264735);
   U142 : INV_X1 port map( A => net264735, ZN => net270357);
   U143 : XNOR2_X1 port map( A => A(42), B => n659, ZN => n680);
   U144 : NAND2_X1 port map( A1 => n655, A2 => net270890, ZN => net296107);
   U145 : XNOR2_X1 port map( A => net270155, B => net276422, ZN => SUM(46));
   U146 : CLKBUF_X1 port map( A => n708, Z => net272615);
   U147 : BUF_X1 port map( A => A(25), Z => n737);
   U148 : CLKBUF_X1 port map( A => n690, Z => net270569);
   U149 : XNOR2_X1 port map( A => A(51), B => B(51), ZN => n695);
   U150 : OR2_X1 port map( A1 => net264731, A2 => net272205, ZN => n662);
   U151 : OR2_X1 port map( A1 => net264731, A2 => net272205, ZN => n741);
   U152 : XNOR2_X1 port map( A => A(34), B => B(34), ZN => net271730);
   U153 : AOI21_X1 port map( B1 => n665, B2 => n674, A => n697, ZN => n693);
   U154 : CLKBUF_X1 port map( A => n693, Z => net272904);
   U155 : AND2_X1 port map( A1 => n693, A2 => B(37), ZN => net272205);
   U156 : OAI21_X1 port map( B1 => n693, B2 => B(37), A => A(37), ZN => n694);
   U157 : AOI21_X1 port map( B1 => n668, B2 => A(36), A => B(36), ZN => n697);
   U158 : INV_X1 port map( A => n696, ZN => n668);
   U159 : INV_X1 port map( A => n668, ZN => n674);
   U160 : AOI22_X1 port map( A1 => net274074, A2 => n683, B1 => n699, B2 => 
                           B(35), ZN => n696);
   U161 : OR2_X1 port map( A1 => net272360, A2 => A(35), ZN => n699);
   U162 : XNOR2_X1 port map( A => net274074, B => n671, ZN => SUM(35));
   U163 : INV_X1 port map( A => A(36), ZN => n665);
   U164 : XNOR2_X1 port map( A => A(36), B => B(36), ZN => net270933);
   U165 : XNOR2_X1 port map( A => A(35), B => B(35), ZN => n671);
   U166 : NOR2_X1 port map( A1 => n703, A2 => n677, ZN => net272360);
   U167 : NOR2_X1 port map( A1 => n702, A2 => A(34), ZN => n677);
   U168 : AOI21_X1 port map( B1 => n702, B2 => A(34), A => B(34), ZN => n703);
   U169 : OR2_X1 port map( A1 => n686, A2 => n705, ZN => n689);
   U170 : NAND2_X1 port map( A1 => n687, A2 => n688, ZN => n705);
   U171 : INV_X1 port map( A => n709, ZN => n687);
   U172 : AND2_X1 port map( A1 => n687, A2 => n688, ZN => n690);
   U173 : AOI21_X1 port map( B1 => n708, B2 => A(32), A => B(32), ZN => n709);
   U174 : INV_X1 port map( A => A(33), ZN => n686);
   U175 : OAI21_X1 port map( B1 => n690, B2 => A(33), A => B(33), ZN => n706);
   U181 : OR2_X1 port map( A1 => A(32), A2 => n708, ZN => n688);
   U182 : XNOR2_X1 port map( A => A(32), B => B(32), ZN => net271088);
   U183 : XNOR2_X1 port map( A => A(33), B => B(33), ZN => net270178);
   U184 : CLKBUF_X1 port map( A => A(31), Z => n725);
   U185 : OAI21_X1 port map( B1 => n767, B2 => n707, A => B(27), ZN => n692);
   U186 : XNOR2_X1 port map( A => n695, B => net276658, ZN => SUM(51));
   U187 : NAND2_X1 port map( A1 => n692, A2 => n752, ZN => n701);
   U188 : CLKBUF_X1 port map( A => A(24), Z => n704);
   U189 : INV_X1 port map( A => n771, ZN => n707);
   U190 : XNOR2_X1 port map( A => n597, B => net276035, ZN => SUM(43));
   U191 : AND2_X1 port map( A1 => n766, A2 => n748, ZN => n710);
   U192 : AOI21_X1 port map( B1 => n713, B2 => n754, A => n700, ZN => net274336
                           );
   U193 : OR2_X1 port map( A1 => n736, A2 => n757, ZN => n713);
   U194 : CLKBUF_X1 port map( A => n729, Z => n716);
   U195 : AND2_X1 port map( A1 => net270356, A2 => n763, ZN => n722);
   U196 : CLKBUF_X1 port map( A => n636, Z => n727);
   U197 : XNOR2_X1 port map( A => n722, B => n734, ZN => SUM(52));
   U198 : XNOR2_X1 port map( A => A(52), B => B(52), ZN => n734);
   U199 : CLKBUF_X1 port map( A => A(26), Z => n735);
   U200 : AOI21_X1 port map( B1 => n662, B2 => n610, A => B(38), ZN => n736);
   U201 : XNOR2_X1 port map( A => net276358, B => net273379, ZN => SUM(40));
   U202 : XNOR2_X1 port map( A => n767, B => n738, ZN => SUM(27));
   U203 : XOR2_X1 port map( A => A(27), B => n756, Z => n738);
   U204 : XNOR2_X1 port map( A => n739, B => net272904, ZN => SUM(37));
   U205 : XNOR2_X1 port map( A => A(37), B => B(37), ZN => n739);
   U206 : XNOR2_X1 port map( A => n662, B => n740, ZN => SUM(38));
   U207 : XNOR2_X1 port map( A => A(38), B => B(38), ZN => n740);
   U208 : CLKBUF_X1 port map( A => A(30), Z => n743);
   U209 : XNOR2_X1 port map( A => n717, B => n719, ZN => SUM(29));
   U210 : OR2_X1 port map( A1 => n717, A2 => n770, ZN => n744);
   U211 : NAND2_X1 port map( A1 => n718, A2 => n744, ZN => n714);
   U212 : OAI22_X1 port map( A1 => n735, A2 => n751, B1 => n698, B2 => B(26), 
                           ZN => n745);
   U213 : CLKBUF_X1 port map( A => n716, Z => n747);
   U214 : OR2_X1 port map( A1 => n701, A2 => n606, ZN => n748);
   U215 : NAND2_X1 port map( A1 => n748, A2 => n766, ZN => n717);
   U216 : XNOR2_X1 port map( A => n751, B => n749, ZN => SUM(26));
   U217 : XNOR2_X1 port map( A => A(26), B => B(26), ZN => n749);
   U218 : XNOR2_X1 port map( A => n636, B => n750, ZN => SUM(56));
   U219 : XNOR2_X1 port map( A => B(56), B => A(56), ZN => n750);
   U220 : XNOR2_X1 port map( A => net272567, B => net271730, ZN => SUM(34));
   U221 : BUF_X1 port map( A => n768, Z => n751);
   U222 : OR2_X1 port map( A1 => n745, A2 => n771, ZN => n752);
   U223 : NAND2_X1 port map( A1 => n752, A2 => n724, ZN => n720);
   U224 : XNOR2_X1 port map( A => net270357, B => n680, ZN => SUM(42));
   U225 : AND2_X1 port map( A1 => net275467, A2 => n621, ZN => n753);
   U226 : NOR2_X1 port map( A1 => n640, A2 => n753, ZN => n636);
   U227 : NOR2_X1 port map( A1 => n742, A2 => n754, ZN => net271108);
   U228 : INV_X1 port map( A => A(39), ZN => n754);
   U229 : INV_X1 port map( A => n742, ZN => n755);
   U230 : XNOR2_X1 port map( A => net271088, B => net272615, ZN => SUM(32));
   U231 : XNOR2_X1 port map( A => net272145, B => net270933, ZN => SUM(36));
   U232 : XNOR2_X1 port map( A => net276651, B => net270617, ZN => SUM(47));
   U233 : XNOR2_X1 port map( A => A(29), B => n758, ZN => n719);
   U234 : OR2_X1 port map( A1 => n594, A2 => n769, ZN => n759);
   U235 : NAND2_X1 port map( A1 => n712, A2 => n759, ZN => n708);
   U236 : XNOR2_X1 port map( A => A(49), B => B(49), ZN => net270418);
   U237 : XNOR2_X1 port map( A => net270380, B => net276072, ZN => SUM(50));
   U238 : INV_X1 port map( A => n591, ZN => net264713);
   U239 : XNOR2_X1 port map( A => n760, B => n746, ZN => SUM(30));
   U240 : XNOR2_X1 port map( A => A(30), B => B(30), ZN => n760);
   U241 : XNOR2_X1 port map( A => net270569, B => net270178, ZN => SUM(33));
   U242 : XNOR2_X1 port map( A => n761, B => n764, ZN => SUM(31));
   U243 : XNOR2_X1 port map( A => A(31), B => B(31), ZN => n761);
   U244 : XNOR2_X1 port map( A => n762, B => n701, ZN => SUM(28));
   U245 : XNOR2_X1 port map( A => A(28), B => B(28), ZN => n762);
   U246 : OAI21_X1 port map( B1 => n767, B2 => n707, A => B(27), ZN => n724);
   U247 : INV_X1 port map( A => A(29), ZN => n770);
   U248 : OAI21_X1 port map( B1 => n710, B2 => A(29), A => B(29), ZN => n718);
   U249 : INV_X1 port map( A => n721, ZN => n766);
   U250 : INV_X1 port map( A => n652, ZN => n763);
   U251 : INV_X1 port map( A => n723, ZN => n767);
   U252 : INV_X1 port map( A => A(27), ZN => n771);
   U253 : XNOR2_X1 port map( A => n634, B => n635, ZN => SUM(57));
   U254 : INV_X1 port map( A => n728, ZN => n768);
   U255 : AOI21_X1 port map( B1 => n773, B2 => n772, A => n732, ZN => n729);
   U256 : INV_X1 port map( A => B(24), ZN => n773);
   U257 : INV_X1 port map( A => A(24), ZN => n772);
   U258 : AOI21_X1 port map( B1 => A(24), B2 => B(24), A => carry_24_port, ZN 
                           => n732);
   U259 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U260 : AOI21_X1 port map( B1 => n714, B2 => A(30), A => B(30), ZN => n715);
   U261 : AOI22_X1 port map( A1 => n727, A2 => A(56), B1 => n637, B2 => B(56), 
                           ZN => n634);
   U262 : OR2_X1 port map( A1 => n636, A2 => A(56), ZN => n637);
   U263 : OAI22_X1 port map( A1 => n737, A2 => n716, B1 => n730, B2 => B(25), 
                           ZN => n728);
   U264 : AND2_X1 port map( A1 => A(25), A2 => n729, ZN => n730);
   U265 : OAI22_X1 port map( A1 => n751, A2 => n735, B1 => n726, B2 => B(26), 
                           ZN => n723);
   U266 : AND2_X1 port map( A1 => n768, A2 => A(26), ZN => n726);
   U267 : INV_X1 port map( A => n594, ZN => n764);
   U268 : INV_X1 port map( A => A(31), ZN => n769);
   U269 : OAI21_X1 port map( B1 => n595, B2 => n725, A => B(31), ZN => n712);
   U270 : AOI21_X1 port map( B1 => n720, B2 => n606, A => B(28), ZN => n721);
   U271 : OAI21_X1 port map( B1 => n746, B2 => n743, A => n765, ZN => n711);
   U272 : INV_X1 port map( A => n715, ZN => n765);
   U273 : INV_X1 port map( A => n694, ZN => net264731);
   U274 : AOI21_X1 port map( B1 => net296107, B2 => net270590, A => B(51), ZN 
                           => n652);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT56_DW01_add_0 is

   port( A, B : in std_logic_vector (55 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (55 downto 0);  CO : out std_logic);

end RCA_NBIT56_DW01_add_0;

architecture SYN_rpl of RCA_NBIT56_DW01_add_0 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_25_port, carry_22_port, carry_21_port, carry_20_port, 
      carry_19_port, carry_18_port, carry_17_port, carry_16_port, carry_15_port
      , carry_14_port, carry_13_port, carry_12_port, carry_11_port, 
      carry_10_port, carry_9_port, carry_8_port, carry_7_port, carry_6_port, 
      carry_5_port, carry_4_port, carry_3_port, carry_2_port, n1, n567, n568, 
      n569, n571, n572, n573, n576, n577, n579, n580, n581, n582, n583, n584, 
      n585, n586, n587, n595, n619, n621, n622, n624, n625, n627, n628, n629, 
      n630, n631, n633, n634, n635, n636, n637, n638, n639, n640, n642, n643, 
      n644, n645, n646, n648, n649, n650, n651, n652, n654, n655, n656, n657, 
      n658, n659, n660, n662, n663, net264690, net264697, net270039, net270279,
      net270391, net271098, net272696, net273386, net276216, net276209, 
      net276208, net276206, net276201, net276197, net276542, net278453, 
      net278447, net278444, net278437, net272487, net278458, net272159, 
      net270453, n601, n600, n599, net271700, net264670, n598, n597, n596, n593
      , net273856, net272775, net271092, net264695, n594, n592, n591, n590, 
      n589, net273589, net273387, net271782, n523, n524, n525, n526, n527, n528
      , n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
      n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, 
      n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, 
      n565, n566, n570, n574, n575, n578, n588, n602, n603, n604, n605, n606, 
      n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, 
      n620, n623, n626, n632, n641, n647, n653, n661, n664, n665, n666, n667, 
      n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, 
      n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, 
      n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, 
      n704, n705, n706, n707, n708, n709, n710, n711, n712 : std_logic;

begin
   
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => n663, CO => 
                           carry_25_port, S => SUM(24));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U150 : XOR2_X1 port map( A => n703, B => B(53), Z => n576);
   U173 : XOR2_X1 port map( A => n653, B => n567, Z => SUM(23));
   U174 : XOR2_X1 port map( A => carry_22_port, B => n662, Z => SUM(22));
   U175 : XOR2_X1 port map( A => A(22), B => B(22), Z => n662);
   U176 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : BUF_X1 port map( A => A(31), Z => n523);
   U2 : NOR2_X1 port map( A1 => n622, A2 => n612, ZN => n524);
   U3 : CLKBUF_X1 port map( A => A(23), Z => n525);
   U4 : NOR2_X1 port map( A1 => net276201, A2 => net276208, ZN => n560);
   U5 : BUF_X1 port map( A => n695, Z => n688);
   U6 : BUF_X1 port map( A => n630, Z => n632);
   U7 : CLKBUF_X1 port map( A => A(41), Z => n526);
   U8 : CLKBUF_X1 port map( A => n645, Z => n661);
   U9 : BUF_X1 port map( A => A(39), Z => n613);
   U10 : AOI21_X1 port map( B1 => n570, B2 => n676, A => n536, ZN => n527);
   U11 : BUF_X1 port map( A => A(29), Z => n530);
   U12 : NOR2_X1 port map( A1 => n553, A2 => A(44), ZN => net270453);
   U13 : INV_X1 port map( A => n552, ZN => n528);
   U14 : BUF_X1 port map( A => n541, Z => net273387);
   U15 : CLKBUF_X1 port map( A => A(40), Z => n529);
   U16 : INV_X1 port map( A => B(53), ZN => n532);
   U17 : OAI21_X1 port map( B1 => n558, B2 => n559, A => n561, ZN => net278447)
                           ;
   U18 : NAND2_X1 port map( A1 => n560, A2 => net270391, ZN => n559);
   U19 : OR2_X1 port map( A1 => n531, A2 => n602, ZN => n538);
   U20 : NAND2_X1 port map( A1 => n534, A2 => n532, ZN => n531);
   U21 : INV_X1 port map( A => B(44), ZN => n554);
   U22 : INV_X1 port map( A => B(29), ZN => n679);
   U23 : INV_X1 port map( A => B(26), ZN => n683);
   U24 : INV_X1 port map( A => B(33), ZN => n682);
   U25 : INV_X1 port map( A => B(27), ZN => n678);
   U26 : OAI22_X1 port map( A1 => n611, A2 => n688, B1 => n580, B2 => B(51), ZN
                           => n533);
   U27 : OAI21_X1 port map( B1 => n616, B2 => n687, A => B(52), ZN => n534);
   U28 : INV_X1 port map( A => n533, ZN => n535);
   U29 : NAND2_X1 port map( A1 => n537, A2 => n538, ZN => n536);
   U30 : OR2_X1 port map( A1 => A(53), A2 => B(53), ZN => n537);
   U31 : INV_X1 port map( A => B(31), ZN => n668);
   U32 : XNOR2_X1 port map( A => n569, B => n539, ZN => SUM(55));
   U33 : XOR2_X1 port map( A => B(55), B => A(55), Z => n539);
   U34 : AOI21_X1 port map( B1 => net264697, B2 => A(49), A => B(49), ZN => 
                           n587);
   U35 : XNOR2_X1 port map( A => net273589, B => net273387, ZN => SUM(41));
   U36 : INV_X1 port map( A => n540, ZN => n541);
   U37 : INV_X1 port map( A => n541, ZN => net276216);
   U38 : XNOR2_X1 port map( A => A(41), B => B(41), ZN => net273589);
   U39 : INV_X1 port map( A => B(41), ZN => net271782);
   U40 : AND2_X1 port map( A1 => n540, A2 => net271782, ZN => net276201);
   U41 : OAI21_X1 port map( B1 => n529, B2 => B(40), A => n542, ZN => n540);
   U42 : NAND2_X1 port map( A1 => n543, A2 => net276542, ZN => n542);
   U43 : NAND2_X1 port map( A1 => A(40), A2 => B(40), ZN => n543);
   U44 : INV_X1 port map( A => n526, ZN => net276197);
   U45 : NOR2_X1 port map( A1 => B(41), A2 => A(41), ZN => net276208);
   U46 : XNOR2_X1 port map( A => A(40), B => B(40), ZN => net276209);
   U47 : INV_X1 port map( A => net276542, ZN => net276206);
   U48 : BUF_X1 port map( A => n642, Z => n623);
   U49 : BUF_X1 port map( A => n618, Z => n664);
   U50 : XNOR2_X1 port map( A => n591, B => B(48), ZN => SUM(48));
   U51 : NAND2_X1 port map( A1 => n589, A2 => n590, ZN => n591);
   U52 : NAND2_X1 port map( A1 => n592, A2 => A(48), ZN => n590);
   U53 : OR2_X1 port map( A1 => A(48), A2 => n592, ZN => n589);
   U54 : AOI21_X1 port map( B1 => net272775, B2 => B(48), A => net273856, ZN =>
                           net272696);
   U55 : AOI21_X1 port map( B1 => net272775, B2 => B(48), A => net273856, ZN =>
                           n586);
   U56 : OR2_X1 port map( A1 => A(48), A2 => n592, ZN => net272775);
   U57 : AND2_X1 port map( A1 => n592, A2 => A(48), ZN => net273856);
   U58 : AOI21_X1 port map( B1 => n544, B2 => net271092, A => n594, ZN => n592)
                           ;
   U59 : AOI21_X1 port map( B1 => net264695, B2 => A(47), A => B(47), ZN => 
                           n594);
   U60 : INV_X1 port map( A => n593, ZN => net264695);
   U61 : CLKBUF_X1 port map( A => n593, Z => net271092);
   U62 : INV_X1 port map( A => net271092, ZN => net271098);
   U63 : INV_X1 port map( A => A(47), ZN => n544);
   U64 : XNOR2_X1 port map( A => A(47), B => B(47), ZN => n595);
   U65 : OAI21_X1 port map( B1 => n596, B2 => B(46), A => n597, ZN => n593);
   U66 : NOR2_X1 port map( A1 => n599, A2 => net264670, ZN => n596);
   U67 : INV_X1 port map( A => A(46), ZN => net264670);
   U68 : NAND2_X1 port map( A1 => net264670, A2 => net272487, ZN => n597);
   U69 : OR2_X1 port map( A1 => n599, A2 => net264670, ZN => net271700);
   U70 : XNOR2_X1 port map( A => n598, B => B(46), ZN => SUM(46));
   U71 : NAND2_X1 port map( A1 => net271700, A2 => n597, ZN => n598);
   U72 : CLKBUF_X1 port map( A => A(45), Z => n549);
   U73 : XNOR2_X1 port map( A => n535, B => n545, ZN => SUM(52));
   U74 : XNOR2_X1 port map( A => A(52), B => B(52), ZN => n545);
   U75 : OR2_X2 port map( A1 => n602, A2 => n694, ZN => n546);
   U76 : CLKBUF_X1 port map( A => n527, Z => n547);
   U77 : AOI21_X1 port map( B1 => net272159, B2 => n549, A => n548, ZN => n599)
                           ;
   U78 : INV_X1 port map( A => n601, ZN => n548);
   U79 : AOI21_X1 port map( B1 => net272159, B2 => n549, A => n548, ZN => 
                           net272487);
   U80 : OAI21_X1 port map( B1 => A(45), B2 => n600, A => B(45), ZN => n601);
   U81 : NOR2_X1 port map( A1 => net278458, A2 => net270453, ZN => n600);
   U82 : CLKBUF_X1 port map( A => n551, Z => net272159);
   U83 : XNOR2_X1 port map( A => net272159, B => n550, ZN => SUM(45));
   U84 : NOR2_X1 port map( A1 => net278458, A2 => net270453, ZN => n551);
   U85 : XNOR2_X1 port map( A => A(45), B => B(45), ZN => n550);
   U86 : OAI21_X1 port map( B1 => net278437, B2 => n552, A => net278444, ZN => 
                           n553);
   U87 : INV_X1 port map( A => net278447, ZN => n552);
   U88 : OAI21_X1 port map( B1 => net278437, B2 => n552, A => net278444, ZN => 
                           n555);
   U89 : AOI21_X1 port map( B1 => A(44), B2 => n555, A => B(44), ZN => 
                           net278458);
   U90 : XNOR2_X1 port map( A => n528, B => net278453, ZN => SUM(43));
   U91 : XNOR2_X1 port map( A => A(44), B => n554, ZN => net270039);
   U92 : INV_X1 port map( A => n559, ZN => net264690);
   U93 : CLKBUF_X1 port map( A => A(25), Z => n614);
   U94 : CLKBUF_X1 port map( A => A(36), Z => n575);
   U95 : CLKBUF_X1 port map( A => A(38), Z => n556);
   U96 : XNOR2_X1 port map( A => A(37), B => B(37), ZN => n557);
   U97 : XNOR2_X1 port map( A => n557, B => n565, ZN => SUM(37));
   U98 : NAND2_X1 port map( A1 => A(42), A2 => B(42), ZN => n561);
   U99 : XNOR2_X1 port map( A => A(42), B => B(42), ZN => net270279);
   U100 : NOR2_X1 port map( A1 => B(42), A2 => A(42), ZN => n558);
   U101 : XNOR2_X1 port map( A => A(43), B => B(43), ZN => net278453);
   U102 : NAND2_X1 port map( A1 => A(43), A2 => B(43), ZN => net278444);
   U103 : NOR2_X1 port map( A1 => A(43), A2 => B(43), ZN => net278437);
   U104 : AOI21_X1 port map( B1 => n620, B2 => n575, A => B(36), ZN => n562);
   U105 : NOR2_X1 port map( A1 => n622, A2 => n612, ZN => n563);
   U106 : BUF_X1 port map( A => A(34), Z => n564);
   U107 : AND2_X1 port map( A1 => n619, A2 => n566, ZN => net276542);
   U108 : NOR2_X1 port map( A1 => n562, A2 => n680, ZN => n565);
   U109 : OR2_X1 port map( A1 => n630, A2 => A(35), ZN => n631);
   U110 : NAND2_X1 port map( A1 => n524, A2 => n613, ZN => n566);
   U111 : BUF_X1 port map( A => n639, Z => n665);
   U112 : NAND2_X1 port map( A1 => net276197, A2 => net276216, ZN => net270391)
                           ;
   U113 : CLKBUF_X1 port map( A => A(51), Z => n611);
   U114 : CLKBUF_X1 port map( A => n703, Z => n570);
   U115 : CLKBUF_X1 port map( A => A(27), Z => n578);
   U116 : XNOR2_X1 port map( A => net276209, B => net276206, ZN => SUM(40));
   U117 : AND2_X1 port map( A1 => n701, A2 => n671, ZN => n574);
   U118 : NOR2_X1 port map( A1 => n660, A2 => n610, ZN => n588);
   U119 : AND2_X1 port map( A1 => n535, A2 => n616, ZN => n602);
   U120 : XNOR2_X1 port map( A => n632, B => n603, ZN => SUM(35));
   U121 : XNOR2_X1 port map( A => A(35), B => B(35), ZN => n603);
   U122 : CLKBUF_X1 port map( A => A(26), Z => n604);
   U123 : INV_X1 port map( A => n608, ZN => n605);
   U124 : AND2_X1 port map( A1 => n705, A2 => n618, ZN => n680);
   U125 : OAI21_X1 port map( B1 => n702, B2 => n578, A => B(27), ZN => n606);
   U126 : CLKBUF_X1 port map( A => A(35), Z => n607);
   U127 : OAI21_X1 port map( B1 => n665, B2 => n615, A => n698, ZN => n608);
   U128 : XOR2_X1 port map( A => A(49), B => B(49), Z => n675);
   U129 : NAND2_X1 port map( A1 => n681, A2 => n655, ZN => n609);
   U130 : OR2_X1 port map( A1 => n610, A2 => n660, ZN => n658);
   U131 : NOR2_X1 port map( A1 => B(25), A2 => A(25), ZN => n610);
   U132 : AND2_X1 port map( A1 => n621, A2 => n711, ZN => n612);
   U133 : INV_X1 port map( A => n555, ZN => net273386);
   U134 : CLKBUF_X1 port map( A => A(32), Z => n615);
   U135 : CLKBUF_X1 port map( A => A(52), Z => n616);
   U136 : CLKBUF_X1 port map( A => A(30), Z => n617);
   U137 : AOI22_X1 port map( A1 => n632, A2 => n607, B1 => n631, B2 => B(35), 
                           ZN => n618);
   U138 : INV_X1 port map( A => n627, ZN => n620);
   U139 : OAI21_X1 port map( B1 => n617, B2 => n661, A => n700, ZN => n642);
   U140 : OAI22_X1 port map( A1 => n604, A2 => n667, B1 => n657, B2 => B(26), 
                           ZN => n626);
   U141 : OAI21_X1 port map( B1 => n697, B2 => n666, A => B(33), ZN => n641);
   U142 : AND2_X1 port map( A1 => n704, A2 => net272696, ZN => n647);
   U143 : NOR2_X1 port map( A1 => n587, A2 => n647, ZN => n583);
   U144 : CLKBUF_X1 port map( A => n568, Z => n653);
   U145 : INV_X1 port map( A => n707, ZN => n666);
   U146 : CLKBUF_X1 port map( A => n588, Z => n667);
   U147 : NOR2_X1 port map( A1 => n686, A2 => n696, ZN => n621);
   U148 : XNOR2_X1 port map( A => A(31), B => n668, ZN => n644);
   U149 : INV_X1 port map( A => n523, ZN => n669);
   U151 : XOR2_X1 port map( A => A(34), B => B(34), Z => n635);
   U152 : OR2_X1 port map( A1 => n696, A2 => n686, ZN => n670);
   U153 : OR2_X1 port map( A1 => n609, A2 => A(28), ZN => n671);
   U154 : NAND2_X1 port map( A1 => n701, A2 => n671, ZN => n648);
   U155 : AND2_X1 port map( A1 => n673, A2 => n637, ZN => n672);
   U156 : OR2_X1 port map( A1 => n707, A2 => n636, ZN => n673);
   U157 : NAND2_X1 port map( A1 => n641, A2 => n673, ZN => n634);
   U158 : OR2_X1 port map( A1 => n648, A2 => n708, ZN => n674);
   U159 : NAND2_X1 port map( A1 => n649, A2 => n674, ZN => n645);
   U160 : XNOR2_X1 port map( A => n675, B => net272696, ZN => SUM(49));
   U161 : INV_X1 port map( A => n546, ZN => n676);
   U162 : BUF_X1 port map( A => n583, Z => n677);
   U163 : XNOR2_X1 port map( A => A(27), B => n678, ZN => n656);
   U164 : XNOR2_X1 port map( A => A(29), B => n679, ZN => n650);
   U165 : NOR2_X1 port map( A1 => n628, A2 => n680, ZN => n624);
   U166 : OR2_X1 port map( A1 => n626, A2 => n709, ZN => n681);
   U167 : NAND2_X1 port map( A1 => n606, A2 => n681, ZN => n651);
   U168 : XNOR2_X1 port map( A => A(33), B => n682, ZN => n638);
   U169 : XNOR2_X1 port map( A => A(26), B => n683, ZN => n659);
   U170 : XNOR2_X1 port map( A => n684, B => n621, ZN => SUM(38));
   U171 : XNOR2_X1 port map( A => A(38), B => n711, ZN => n684);
   U172 : XNOR2_X1 port map( A => net270039, B => net273386, ZN => SUM(44));
   U177 : XNOR2_X1 port map( A => n665, B => n685, ZN => SUM(32));
   U178 : XNOR2_X1 port map( A => A(32), B => B(32), ZN => n685);
   U179 : AND2_X1 port map( A1 => A(37), A2 => n565, ZN => n686);
   U180 : INV_X1 port map( A => n579, ZN => n687);
   U181 : CLKBUF_X1 port map( A => A(50), Z => n689);
   U182 : XNOR2_X1 port map( A => net270279, B => net264690, ZN => SUM(42));
   U183 : INV_X1 port map( A => A(29), ZN => n708);
   U184 : INV_X1 port map( A => A(36), ZN => n705);
   U185 : INV_X1 port map( A => A(49), ZN => n704);
   U186 : INV_X1 port map( A => n525, ZN => n710);
   U187 : XNOR2_X1 port map( A => n705, B => B(36), ZN => n629);
   U188 : XNOR2_X1 port map( A => n690, B => n661, ZN => SUM(30));
   U189 : XNOR2_X1 port map( A => A(30), B => B(30), ZN => n690);
   U190 : XNOR2_X1 port map( A => n691, B => n609, ZN => SUM(28));
   U191 : XNOR2_X1 port map( A => A(28), B => B(28), ZN => n691);
   U192 : XNOR2_X1 port map( A => n692, B => n524, ZN => SUM(39));
   U193 : XNOR2_X1 port map( A => A(39), B => B(39), ZN => n692);
   U194 : XNOR2_X1 port map( A => A(51), B => B(51), ZN => n581);
   U195 : XNOR2_X1 port map( A => n693, B => n614, ZN => SUM(25));
   U196 : XNOR2_X1 port map( A => carry_25_port, B => B(25), ZN => n693);
   U197 : XNOR2_X1 port map( A => n608, B => n638, ZN => SUM(33));
   U198 : INV_X1 port map( A => n577, ZN => n694);
   U199 : OAI21_X1 port map( B1 => n687, B2 => n616, A => B(52), ZN => n577);
   U200 : XNOR2_X1 port map( A => n623, B => n644, ZN => SUM(31));
   U201 : XNOR2_X1 port map( A => A(23), B => B(23), ZN => n568);
   U202 : OAI22_X1 port map( A1 => n604, A2 => n667, B1 => n657, B2 => B(26), 
                           ZN => n654);
   U203 : AND2_X1 port map( A1 => A(26), A2 => n588, ZN => n657);
   U204 : INV_X1 port map( A => B(23), ZN => n712);
   U205 : INV_X1 port map( A => B(38), ZN => n711);
   U206 : AOI22_X1 port map( A1 => B(22), A2 => A(22), B1 => n662, B2 => 
                           carry_22_port, ZN => n567);
   U207 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U208 : XNOR2_X1 port map( A => A(54), B => B(54), ZN => n573);
   U209 : XNOR2_X1 port map( A => A(50), B => B(50), ZN => n585);
   U210 : XNOR2_X1 port map( A => n635, B => n672, ZN => SUM(34));
   U211 : INV_X1 port map( A => A(33), ZN => n707);
   U212 : OAI21_X1 port map( B1 => n669, B2 => n623, A => n643, ZN => n639);
   U213 : OAI21_X1 port map( B1 => n699, B2 => n523, A => B(31), ZN => n643);
   U214 : OAI22_X1 port map( A1 => n712, A2 => n710, B1 => n567, B2 => n568, ZN
                           => n663);
   U215 : AOI22_X1 port map( A1 => n632, A2 => n607, B1 => n631, B2 => B(35), 
                           ZN => n627);
   U216 : AOI21_X1 port map( B1 => n706, B2 => n672, A => n633, ZN => n630);
   U217 : INV_X1 port map( A => n642, ZN => n699);
   U218 : OAI21_X1 port map( B1 => n574, B2 => n530, A => B(29), ZN => n649);
   U219 : INV_X1 port map( A => n564, ZN => n706);
   U220 : OAI21_X1 port map( B1 => n563, B2 => n613, A => B(39), ZN => n619);
   U221 : AOI21_X1 port map( B1 => n670, B2 => B(38), A => n556, ZN => n622);
   U222 : INV_X1 port map( A => n636, ZN => n697);
   U223 : INV_X1 port map( A => n652, ZN => n701);
   U224 : AOI21_X1 port map( B1 => A(28), B2 => n651, A => B(28), ZN => n652);
   U225 : OAI21_X1 port map( B1 => n666, B2 => n605, A => B(33), ZN => n637);
   U226 : XNOR2_X1 port map( A => n546, B => n576, ZN => SUM(53));
   U227 : INV_X1 port map( A => n654, ZN => n702);
   U228 : OAI21_X1 port map( B1 => n665, B2 => n615, A => n698, ZN => n636);
   U229 : XNOR2_X1 port map( A => net271098, B => n595, ZN => SUM(47));
   U230 : AOI21_X1 port map( B1 => n570, B2 => n676, A => n536, ZN => n571);
   U231 : XNOR2_X1 port map( A => n688, B => n581, ZN => SUM(51));
   U232 : OAI22_X1 port map( A1 => n611, A2 => n688, B1 => n580, B2 => B(51), 
                           ZN => n579);
   U233 : AND2_X1 port map( A1 => n695, A2 => A(51), ZN => n580);
   U234 : INV_X1 port map( A => n586, ZN => net264697);
   U235 : INV_X1 port map( A => n625, ZN => n696);
   U236 : AOI21_X1 port map( B1 => n634, B2 => n564, A => B(34), ZN => n633);
   U237 : INV_X1 port map( A => n640, ZN => n698);
   U238 : INV_X1 port map( A => n646, ZN => n700);
   U239 : INV_X1 port map( A => A(27), ZN => n709);
   U240 : OAI21_X1 port map( B1 => n702, B2 => n578, A => B(27), ZN => n655);
   U241 : INV_X1 port map( A => A(53), ZN => n703);
   U242 : XNOR2_X1 port map( A => n656, B => n626, ZN => SUM(27));
   U243 : OAI21_X1 port map( B1 => n624, B2 => A(37), A => B(37), ZN => n625);
   U244 : AOI21_X1 port map( B1 => n639, B2 => A(32), A => B(32), ZN => n640);
   U245 : AOI21_X1 port map( B1 => A(30), B2 => n645, A => B(30), ZN => n646);
   U246 : XNOR2_X1 port map( A => n650, B => n648, ZN => SUM(29));
   U247 : XNOR2_X1 port map( A => n659, B => n658, ZN => SUM(26));
   U248 : AOI21_X1 port map( B1 => A(25), B2 => B(25), A => carry_25_port, ZN 
                           => n660);
   U249 : XNOR2_X1 port map( A => n571, B => n573, ZN => SUM(54));
   U250 : OAI22_X1 port map( A1 => A(54), A2 => n547, B1 => B(54), B2 => n572, 
                           ZN => n569);
   U251 : AND2_X1 port map( A1 => n527, A2 => A(54), ZN => n572);
   U252 : XNOR2_X1 port map( A => n677, B => n585, ZN => SUM(50));
   U253 : INV_X1 port map( A => n582, ZN => n695);
   U254 : OAI22_X1 port map( A1 => n677, A2 => n689, B1 => n584, B2 => B(50), 
                           ZN => n582);
   U255 : AND2_X1 port map( A1 => n583, A2 => A(50), ZN => n584);
   U256 : AOI21_X1 port map( B1 => n620, B2 => n575, A => B(36), ZN => n628);
   U257 : XNOR2_X1 port map( A => n629, B => n664, ZN => SUM(36));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT54_DW01_add_0 is

   port( A, B : in std_logic_vector (53 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (53 downto 0);  CO : out std_logic);

end RCA_NBIT54_DW01_add_0;

architecture SYN_rpl of RCA_NBIT54_DW01_add_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_51_port, carry_16_port, carry_15_port, carry_14_port, 
      carry_13_port, carry_12_port, carry_11_port, carry_10_port, carry_9_port,
      carry_8_port, carry_7_port, carry_6_port, carry_5_port, carry_4_port, 
      carry_3_port, carry_2_port, n1, carry_49_port, carry_48_port, n597, n598,
      n599, n600, n601, n602, n605, n607, n610, n611, n613, n616, n617, n633, 
      n634, n638, n654, n655, n657, n658, n661, n665, n666, n669, n670, n671, 
      n673, n681, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, 
      n694, n695, n696, n697, net264620, net264633, net264637, net264651, 
      net270741, net272018, net272316, net272575, net273024, net273669, 
      net274032, net275383, net275382, net275840, net276458, net276618, n667, 
      n664, n663, n660, net279581, net287700, n612, net276671, net275808, 
      net271122, net264619, n644, n640, n639, n636, net274118, net271892, 
      net264618, n647, n643, n642, n653, n652, n649, n648, n646, n645, n630, 
      n627, net276376, net271129, net264621, n629, n628, n624, net275392, 
      net272776, n625, n621, n552, n553, n554, n555, n556, n557, n558, n559, 
      n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, 
      n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, 
      n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, 
      n596, n603, n604, n606, n608, n609, n614, n615, n618, n619, n620, n622, 
      n623, n626, n631, n632, n635, n637, n641, n650, n651, n656, n659, n662, 
      n668, n672, n674, n675, n676, n677, n678, n679, n680, n682, n683, n698, 
      n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, 
      n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, 
      n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, 
      n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, 
      n747, n748, n749 : std_logic;

begin
   
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U1_48 : FA_X1 port map( A => A(48), B => B(48), CI => carry_48_port, CO => 
                           carry_49_port, S => SUM(48));
   U148 : XOR2_X1 port map( A => n598, B => carry_49_port, Z => SUM(49));
   U176 : XOR2_X1 port map( A => n684, B => n686, Z => SUM(20));
   U177 : XOR2_X1 port map( A => B(20), B => A(20), Z => n686);
   U178 : XOR2_X1 port map( A => B(19), B => A(19), Z => n689);
   U179 : XOR2_X1 port map( A => B(18), B => A(18), Z => n692);
   U180 : XOR2_X1 port map( A => B(17), B => A(17), Z => n695);
   U181 : XOR2_X1 port map( A => A(16), B => n697, Z => SUM(16));
   U182 : XOR2_X1 port map( A => carry_16_port, B => B(16), Z => n697);
   U183 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : BUF_X1 port map( A => n674, Z => n552);
   U2 : BUF_X1 port map( A => A(46), Z => n712);
   U3 : INV_X1 port map( A => B(22), ZN => n580);
   U4 : BUF_X1 port map( A => A(36), Z => n622);
   U5 : OR2_X1 port map( A1 => net272575, A2 => net264651, ZN => n707);
   U6 : INV_X1 port map( A => B(23), ZN => n579);
   U7 : XNOR2_X1 port map( A => n582, B => B(21), ZN => n577);
   U8 : XNOR2_X1 port map( A => B(22), B => n564, ZN => n576);
   U9 : XNOR2_X1 port map( A => n577, B => n571, ZN => SUM(21));
   U10 : INV_X1 port map( A => B(51), ZN => n729);
   U11 : AND2_X1 port map( A1 => n651, A2 => n672, ZN => n553);
   U12 : BUF_X1 port map( A => n600, Z => n710);
   U13 : AND2_X1 port map( A1 => n569, A2 => n568, ZN => n554);
   U14 : OR2_X2 port map( A1 => n655, A2 => net273669, ZN => n608);
   U15 : BUF_X1 port map( A => n648, Z => n604);
   U16 : CLKBUF_X1 port map( A => n572, Z => n555);
   U17 : CLKBUF_X1 port map( A => n666, Z => net276458);
   U18 : BUF_X1 port map( A => A(39), Z => net276376);
   U19 : AND2_X1 port map( A1 => n746, A2 => n637, ZN => net272316);
   U20 : OAI21_X1 port map( B1 => A(42), B2 => n680, A => B(42), ZN => n556);
   U21 : NAND2_X1 port map( A1 => n572, A2 => n584, ZN => n568);
   U22 : NAND2_X1 port map( A1 => n581, A2 => n580, ZN => n569);
   U23 : INV_X1 port map( A => net264618, ZN => n557);
   U24 : AOI22_X1 port map( A1 => net272776, A2 => n560, B1 => n625, B2 => 
                           B(40), ZN => n558);
   U25 : INV_X1 port map( A => B(43), ZN => n702);
   U26 : INV_X1 port map( A => B(45), ZN => n727);
   U27 : INV_X1 port map( A => B(33), ZN => n609);
   U28 : INV_X1 port map( A => B(49), ZN => n728);
   U29 : INV_X1 port map( A => B(39), ZN => n587);
   U30 : INV_X1 port map( A => B(34), ZN => n614);
   U31 : INV_X1 port map( A => B(36), ZN => n619);
   U32 : NAND2_X1 port map( A1 => n670, A2 => n717, ZN => n666);
   U33 : NOR2_X1 port map( A1 => net272316, A2 => n616, ZN => n612);
   U34 : XNOR2_X1 port map( A => n733, B => n705, ZN => SUM(30));
   U35 : XNOR2_X1 port map( A => n561, B => net275392, ZN => SUM(41));
   U36 : INV_X1 port map( A => n558, ZN => net275392);
   U37 : XNOR2_X1 port map( A => A(41), B => B(41), ZN => n561);
   U38 : AOI22_X1 port map( A1 => net272776, A2 => n560, B1 => n625, B2 => 
                           B(40), ZN => n621);
   U39 : OR2_X1 port map( A1 => A(40), A2 => n624, ZN => n625);
   U40 : CLKBUF_X1 port map( A => A(40), Z => n560);
   U41 : BUF_X1 port map( A => n624, Z => net272776);
   U42 : XNOR2_X1 port map( A => net272776, B => n559, ZN => SUM(40));
   U43 : NAND2_X1 port map( A1 => A(41), A2 => B(41), ZN => net275383);
   U44 : NOR2_X1 port map( A1 => A(41), A2 => B(41), ZN => net275382);
   U45 : XNOR2_X1 port map( A => A(40), B => B(40), ZN => n559);
   U46 : CLKBUF_X1 port map( A => A(24), Z => n562);
   U47 : AOI21_X1 port map( B1 => n615, B2 => n622, A => B(36), ZN => n563);
   U48 : INV_X1 port map( A => n681, ZN => n570);
   U49 : INV_X1 port map( A => n570, ZN => n582);
   U50 : NAND2_X1 port map( A1 => A(22), A2 => n564, ZN => n581);
   U51 : XNOR2_X1 port map( A => n583, B => n576, ZN => SUM(22));
   U52 : INV_X1 port map( A => A(22), ZN => n572);
   U53 : XNOR2_X1 port map( A => A(23), B => B(23), ZN => n578);
   U54 : INV_X1 port map( A => A(23), ZN => n573);
   U55 : NAND2_X1 port map( A1 => B(21), A2 => n570, ZN => n565);
   U56 : OAI21_X1 port map( B1 => B(21), B2 => n570, A => A(21), ZN => n566);
   U57 : INV_X1 port map( A => n555, ZN => n583);
   U58 : NAND2_X1 port map( A1 => n565, A2 => n566, ZN => n564);
   U59 : AND2_X1 port map( A1 => n565, A2 => n566, ZN => n584);
   U60 : AOI21_X1 port map( B1 => A(24), B2 => n585, A => B(24), ZN => n673);
   U61 : XNOR2_X1 port map( A => n578, B => n554, ZN => SUM(23));
   U62 : OAI21_X1 port map( B1 => n573, B2 => n567, A => n579, ZN => n575);
   U63 : AND2_X1 port map( A1 => n575, A2 => n574, ZN => net273024);
   U64 : AND2_X1 port map( A1 => n575, A2 => n574, ZN => n585);
   U65 : INV_X1 port map( A => A(21), ZN => n571);
   U66 : NAND2_X1 port map( A1 => n569, A2 => n568, ZN => n567);
   U67 : NAND2_X1 port map( A1 => n573, A2 => n567, ZN => n574);
   U68 : OAI21_X1 port map( B1 => net264621, B2 => net271129, A => n628, ZN => 
                           n624);
   U69 : OAI21_X1 port map( B1 => n586, B2 => A(39), A => B(39), ZN => n628);
   U70 : INV_X1 port map( A => n627, ZN => n586);
   U71 : BUF_X1 port map( A => n627, Z => net271129);
   U72 : XNOR2_X1 port map( A => n629, B => net271129, ZN => SUM(39));
   U73 : INV_X1 port map( A => net276376, ZN => net264621);
   U74 : XNOR2_X1 port map( A => A(39), B => n587, ZN => n629);
   U75 : OAI21_X1 port map( B1 => n591, B2 => n590, A => n588, ZN => n627);
   U76 : INV_X1 port map( A => n630, ZN => n588);
   U77 : AOI21_X1 port map( B1 => net272018, B2 => A(38), A => B(38), ZN => 
                           n630);
   U78 : BUF_X1 port map( A => net272018, Z => n590);
   U79 : XNOR2_X1 port map( A => n589, B => n590, ZN => SUM(38));
   U80 : CLKBUF_X1 port map( A => A(38), Z => n591);
   U81 : XNOR2_X1 port map( A => A(38), B => B(38), ZN => n589);
   U82 : OAI21_X1 port map( B1 => n594, B2 => n557, A => B(33), ZN => n646);
   U83 : NAND2_X1 port map( A1 => n646, A2 => net271892, ZN => n643);
   U84 : AND2_X1 port map( A1 => n646, A2 => net271892, ZN => net275808);
   U85 : INV_X1 port map( A => n645, ZN => n594);
   U86 : OAI21_X1 port map( B1 => n604, B2 => n596, A => n593, ZN => n645);
   U87 : INV_X1 port map( A => n649, ZN => n593);
   U88 : OAI21_X1 port map( B1 => n604, B2 => n596, A => n593, ZN => net274118)
                           ;
   U89 : AOI21_X1 port map( B1 => n648, B2 => A(32), A => B(32), ZN => n649);
   U90 : CLKBUF_X1 port map( A => A(32), Z => n596);
   U91 : XNOR2_X1 port map( A => n604, B => n595, ZN => SUM(32));
   U92 : INV_X1 port map( A => A(33), ZN => net264618);
   U93 : XNOR2_X1 port map( A => A(33), B => n609, ZN => n647);
   U94 : OAI21_X1 port map( B1 => n608, B2 => n592, A => n652, ZN => n648);
   U95 : OAI21_X1 port map( B1 => n603, B2 => n606, A => B(31), ZN => n652);
   U96 : NOR2_X1 port map( A1 => net273669, A2 => n655, ZN => n603);
   U97 : INV_X1 port map( A => n606, ZN => n592);
   U98 : BUF_X1 port map( A => A(31), Z => n606);
   U99 : XNOR2_X1 port map( A => A(32), B => B(32), ZN => n595);
   U100 : XNOR2_X1 port map( A => n608, B => n653, ZN => SUM(31));
   U101 : XOR2_X1 port map( A => A(31), B => B(31), Z => n653);
   U102 : AOI21_X1 port map( B1 => n643, B2 => A(34), A => B(34), ZN => n642);
   U103 : AOI21_X1 port map( B1 => net264619, B2 => net275808, A => n642, ZN =>
                           n639);
   U104 : XNOR2_X1 port map( A => A(34), B => n614, ZN => n644);
   U105 : CLKBUF_X1 port map( A => A(34), Z => net276671);
   U106 : OR2_X1 port map( A1 => net274118, A2 => net264618, ZN => net271892);
   U107 : XNOR2_X1 port map( A => net274118, B => n647, ZN => SUM(33));
   U108 : AOI21_X1 port map( B1 => n615, B2 => n622, A => B(36), ZN => n623);
   U109 : NOR2_X1 port map( A1 => n563, A2 => net279581, ZN => n633);
   U110 : INV_X1 port map( A => n622, ZN => net264620);
   U111 : INV_X1 port map( A => n636, ZN => n615);
   U112 : AOI22_X1 port map( A1 => net271122, A2 => n620, B1 => n640, B2 => 
                           B(35), ZN => n636);
   U113 : CLKBUF_X1 port map( A => A(35), Z => n620);
   U114 : AOI22_X1 port map( A1 => net271122, A2 => n620, B1 => n640, B2 => 
                           B(35), ZN => net276618);
   U115 : BUF_X1 port map( A => n639, Z => net271122);
   U116 : XNOR2_X1 port map( A => net271122, B => n618, ZN => SUM(35));
   U117 : XNOR2_X1 port map( A => A(36), B => n619, ZN => n638);
   U118 : OR2_X1 port map( A1 => n639, A2 => A(35), ZN => n640);
   U119 : XNOR2_X1 port map( A => A(35), B => B(35), ZN => n618);
   U120 : INV_X1 port map( A => net276671, ZN => net264619);
   U121 : XNOR2_X1 port map( A => n644, B => net275808, ZN => SUM(34));
   U122 : CLKBUF_X1 port map( A => n632, Z => n626);
   U123 : XNOR2_X1 port map( A => n602, B => n730, ZN => SUM(53));
   U124 : XNOR2_X1 port map( A => n631, B => n626, ZN => SUM(44));
   U125 : XNOR2_X1 port map( A => A(44), B => B(44), ZN => n631);
   U126 : NOR2_X1 port map( A1 => n616, A2 => net272316, ZN => n632);
   U127 : AND2_X1 port map( A1 => A(44), A2 => n632, ZN => net272575);
   U128 : OAI21_X1 port map( B1 => n612, B2 => A(44), A => B(44), ZN => n613);
   U129 : CLKBUF_X1 port map( A => net276618, Z => net287700);
   U130 : CLKBUF_X1 port map( A => A(51), Z => n635);
   U131 : BUF_X1 port map( A => A(29), Z => n714);
   U132 : AND2_X1 port map( A1 => net276618, A2 => net264620, ZN => net279581);
   U133 : AND2_X1 port map( A1 => n698, A2 => n699, ZN => n637);
   U134 : AOI22_X1 port map( A1 => n607, A2 => carry_51_port, B1 => n635, B2 =>
                           B(51), ZN => n641);
   U135 : XNOR2_X1 port map( A => n668, B => n656, ZN => SUM(28));
   U136 : XNOR2_X1 port map( A => A(28), B => B(28), ZN => n656);
   U137 : BUF_X1 port map( A => n660, Z => n668);
   U138 : CLKBUF_X1 port map( A => A(28), Z => net274032);
   U139 : AOI21_X1 port map( B1 => n660, B2 => A(28), A => B(28), ZN => n661);
   U140 : NAND2_X1 port map( A1 => n664, A2 => n659, ZN => n660);
   U141 : OR2_X1 port map( A1 => n663, A2 => n650, ZN => n659);
   U142 : INV_X1 port map( A => A(27), ZN => n650);
   U143 : INV_X1 port map( A => n650, ZN => n662);
   U144 : NAND2_X1 port map( A1 => n651, A2 => n672, ZN => n663);
   U145 : INV_X1 port map( A => n667, ZN => n651);
   U146 : AND2_X1 port map( A1 => n651, A2 => n672, ZN => net275840);
   U147 : AOI21_X1 port map( B1 => n666, B2 => A(26), A => B(26), ZN => n667);
   U149 : OAI21_X1 port map( B1 => net275840, B2 => n662, A => B(27), ZN => 
                           n664);
   U150 : XNOR2_X1 port map( A => A(27), B => B(27), ZN => n665);
   U151 : OR2_X1 port map( A1 => A(26), A2 => n666, ZN => n672);
   U152 : XNOR2_X1 port map( A => A(26), B => B(26), ZN => net270741);
   U153 : BUF_X1 port map( A => n739, Z => n708);
   U154 : AOI21_X1 port map( B1 => net287700, B2 => net264620, A => n623, ZN =>
                           n674);
   U155 : OR2_X1 port map( A1 => n747, A2 => n676, ZN => n675);
   U156 : XNOR2_X1 port map( A => n597, B => n718, ZN => SUM(50));
   U157 : CLKBUF_X1 port map( A => n657, Z => n676);
   U158 : BUF_X1 port map( A => A(30), Z => n679);
   U159 : OAI21_X1 port map( B1 => net275382, B2 => n621, A => net275383, ZN =>
                           n677);
   U160 : CLKBUF_X1 port map( A => A(47), Z => n678);
   U161 : XNOR2_X1 port map( A => n617, B => n637, ZN => SUM(43));
   U162 : OAI21_X1 port map( B1 => A(42), B2 => n680, A => B(42), ZN => n698);
   U163 : NAND2_X1 port map( A1 => n677, A2 => A(42), ZN => n699);
   U164 : XNOR2_X1 port map( A => n682, B => n700, ZN => SUM(42));
   U165 : OAI21_X1 port map( B1 => n621, B2 => net275382, A => net275383, ZN =>
                           n680);
   U166 : XNOR2_X1 port map( A => n677, B => B(42), ZN => n682);
   U167 : CLKBUF_X1 port map( A => A(42), Z => n700);
   U168 : NAND2_X1 port map( A1 => n556, A2 => n699, ZN => n683);
   U169 : NAND2_X1 port map( A1 => n634, A2 => n701, ZN => net272018);
   U170 : NAND2_X1 port map( A1 => n674, A2 => A(37), ZN => n701);
   U171 : XNOR2_X1 port map( A => A(51), B => B(51), ZN => n713);
   U172 : NOR2_X1 port map( A1 => n705, A2 => n679, ZN => net273669);
   U173 : OR2_X1 port map( A1 => n676, A2 => n747, ZN => n711);
   U174 : XNOR2_X1 port map( A => A(43), B => n702, ZN => n617);
   U175 : INV_X1 port map( A => n735, ZN => n703);
   U184 : XNOR2_X1 port map( A => n704, B => n738, ZN => SUM(29));
   U185 : XNOR2_X1 port map( A => A(29), B => B(29), ZN => n704);
   U186 : NAND2_X1 port map( A1 => n711, A2 => n658, ZN => n705);
   U187 : OR2_X1 port map( A1 => net264651, A2 => net272575, ZN => n706);
   U188 : XNOR2_X1 port map( A => n709, B => net273024, ZN => SUM(24));
   U189 : XNOR2_X1 port map( A => A(24), B => B(24), ZN => n709);
   U190 : NAND2_X1 port map( A1 => n658, A2 => n675, ZN => n654);
   U191 : XNOR2_X1 port map( A => n713, B => carry_51_port, ZN => SUM(51));
   U192 : INV_X1 port map( A => n707, ZN => n715);
   U193 : NOR2_X1 port map( A1 => n707, A2 => A(45), ZN => n716);
   U194 : NOR2_X1 port map( A1 => n716, A2 => n610, ZN => n600);
   U195 : OR2_X1 port map( A1 => n748, A2 => n669, ZN => n717);
   U196 : XOR2_X1 port map( A => A(50), B => B(50), Z => n718);
   U197 : NAND2_X1 port map( A1 => n736, A2 => A(50), ZN => n719);
   U198 : NAND2_X1 port map( A1 => n736, A2 => B(50), ZN => n720);
   U199 : NAND2_X1 port map( A1 => A(50), A2 => B(50), ZN => n721);
   U200 : NAND3_X1 port map( A1 => n719, A2 => n720, A3 => n721, ZN => 
                           carry_51_port);
   U201 : XNOR2_X1 port map( A => n737, B => n722, ZN => SUM(47));
   U202 : XNOR2_X1 port map( A => A(47), B => B(47), ZN => n722);
   U203 : XNOR2_X1 port map( A => n723, B => n552, ZN => SUM(37));
   U204 : XNOR2_X1 port map( A => A(37), B => B(37), ZN => n723);
   U205 : NAND2_X1 port map( A1 => n737, A2 => n678, ZN => n724);
   U206 : NAND2_X1 port map( A1 => n737, A2 => B(47), ZN => n725);
   U207 : NAND2_X1 port map( A1 => A(47), A2 => B(47), ZN => n726);
   U208 : NAND3_X1 port map( A1 => n725, A2 => n724, A3 => n726, ZN => 
                           carry_48_port);
   U209 : XNOR2_X1 port map( A => A(45), B => n727, ZN => n611);
   U210 : XNOR2_X1 port map( A => net276458, B => net270741, ZN => SUM(26));
   U211 : XNOR2_X1 port map( A => A(49), B => n728, ZN => n598);
   U212 : XNOR2_X1 port map( A => A(51), B => n729, ZN => n607);
   U213 : XNOR2_X1 port map( A => B(53), B => A(53), ZN => n730);
   U214 : CLKBUF_X1 port map( A => A(49), Z => n731);
   U215 : XOR2_X1 port map( A => n641, B => n732, Z => SUM(52));
   U216 : XOR2_X1 port map( A => B(52), B => n745, Z => n732);
   U217 : XNOR2_X1 port map( A => A(30), B => B(30), ZN => n733);
   U218 : INV_X1 port map( A => A(25), ZN => n748);
   U219 : XNOR2_X1 port map( A => n553, B => n665, ZN => SUM(27));
   U220 : XNOR2_X1 port map( A => n611, B => n715, ZN => SUM(45));
   U221 : XNOR2_X1 port map( A => n734, B => n710, ZN => SUM(46));
   U222 : XNOR2_X1 port map( A => A(46), B => B(46), ZN => n734);
   U223 : INV_X1 port map( A => n714, ZN => n747);
   U224 : OAI21_X1 port map( B1 => A(52), B2 => n735, A => B(52), ZN => n605);
   U225 : INV_X1 port map( A => A(52), ZN => n745);
   U226 : OAI21_X1 port map( B1 => A(20), B2 => n684, A => n740, ZN => n681);
   U227 : INV_X1 port map( A => n685, ZN => n740);
   U228 : AOI21_X1 port map( B1 => n684, B2 => A(20), A => B(20), ZN => n685);
   U229 : OAI22_X1 port map( A1 => A(18), A2 => n742, B1 => B(18), B2 => n690, 
                           ZN => n687);
   U230 : AND2_X1 port map( A1 => n742, A2 => A(18), ZN => n690);
   U231 : INV_X1 port map( A => n691, ZN => n742);
   U232 : OAI22_X1 port map( A1 => A(17), A2 => n743, B1 => B(17), B2 => n693, 
                           ZN => n691);
   U233 : AND2_X1 port map( A1 => n743, A2 => A(17), ZN => n693);
   U234 : INV_X1 port map( A => n694, ZN => n743);
   U235 : OAI21_X1 port map( B1 => n687, B2 => n749, A => n688, ZN => n684);
   U236 : INV_X1 port map( A => A(19), ZN => n749);
   U237 : OAI21_X1 port map( B1 => n741, B2 => A(19), A => B(19), ZN => n688);
   U238 : INV_X1 port map( A => n687, ZN => n741);
   U239 : OAI21_X1 port map( B1 => B(16), B2 => A(16), A => n744, ZN => n694);
   U240 : INV_X1 port map( A => n696, ZN => n744);
   U241 : AOI21_X1 port map( B1 => A(16), B2 => B(16), A => carry_16_port, ZN 
                           => n696);
   U242 : XNOR2_X1 port map( A => n694, B => n695, ZN => SUM(17));
   U243 : XNOR2_X1 port map( A => n691, B => n692, ZN => SUM(18));
   U244 : XNOR2_X1 port map( A => n687, B => n689, ZN => SUM(19));
   U245 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U246 : OAI21_X1 port map( B1 => net274032, B2 => n668, A => net264637, ZN =>
                           n657);
   U247 : XNOR2_X1 port map( A => A(25), B => B(25), ZN => n671);
   U248 : INV_X1 port map( A => n661, ZN => net264637);
   U249 : INV_X1 port map( A => A(43), ZN => n746);
   U250 : OAI21_X1 port map( B1 => n714, B2 => n738, A => B(29), ZN => n658);
   U251 : OAI21_X1 port map( B1 => n739, B2 => A(25), A => B(25), ZN => n670);
   U252 : INV_X1 port map( A => n669, ZN => n739);
   U253 : OAI21_X1 port map( B1 => n703, B2 => n745, A => n605, ZN => n602);
   U254 : INV_X1 port map( A => n641, ZN => n735);
   U255 : INV_X1 port map( A => n597, ZN => n736);
   U256 : XNOR2_X1 port map( A => n671, B => n708, ZN => SUM(25));
   U257 : AOI21_X1 port map( B1 => A(45), B2 => n706, A => B(45), ZN => n610);
   U258 : INV_X1 port map( A => n673, ZN => net264633);
   U259 : AOI22_X1 port map( A1 => B(49), A2 => n731, B1 => n598, B2 => 
                           carry_49_port, ZN => n597);
   U260 : INV_X1 port map( A => n599, ZN => n737);
   U261 : AOI21_X1 port map( B1 => A(43), B2 => n683, A => B(43), ZN => n616);
   U262 : XNOR2_X1 port map( A => net276618, B => n638, ZN => SUM(36));
   U263 : INV_X1 port map( A => n657, ZN => n738);
   U264 : OAI21_X1 port map( B1 => n562, B2 => net273024, A => net264633, ZN =>
                           n669);
   U265 : INV_X1 port map( A => n613, ZN => net264651);
   U266 : AOI22_X1 port map( A1 => n710, A2 => n712, B1 => n601, B2 => B(46), 
                           ZN => n599);
   U267 : OR2_X1 port map( A1 => n600, A2 => A(46), ZN => n601);
   U268 : OAI21_X1 port map( B1 => n633, B2 => A(37), A => B(37), ZN => n634);
   U269 : AOI21_X1 port map( B1 => n679, B2 => n654, A => B(30), ZN => n655);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT52_DW01_add_0 is

   port( A, B : in std_logic_vector (51 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (51 downto 0);  CO : out std_logic);

end RCA_NBIT52_DW01_add_0;

architecture SYN_rpl of RCA_NBIT52_DW01_add_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_18_port, carry_17_port, carry_16_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_10_port
      , carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, n1, n586, n588, n589, n590, 
      n591, n593, n594, n595, n596, n597, n603, n606, n620, n624, n627, n645, 
      n677, n680, n681, n682, n683, n684, net264596, net270022, net271069, 
      net271621, net271690, net271720, net272082, net272213, net272365, 
      net272472, net272919, net273792, net274030, net275693, net275676, 
      net275668, net275667, net275652, net275647, net275643, net275641, 
      net276573, net276693, n658, net274721, n679, net264601, n612, n608, 
      net272480, net272479, net272285, net264574, net275685, net275665, 
      net275664, net275663, net271193, net264594, n633, n631, n630, n626, 
      net264600, n615, n611, net287683, net271948, net270519, net270509, 
      net264572, n642, n641, n639, n638, n637, n636, n632, net273613, net271609
      , net270507, net264589, net264570, n654, n653, n651, n650, n649, n648, 
      n644, n621, n618, n614, n542, n543, n544, n545, n546, n547, n548, n549, 
      n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, 
      n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, 
      n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, 
      n587, n592, n598, n599, n600, n601, n602, n604, n605, n607, n609, n610, 
      n613, n616, n617, n619, n622, n623, n625, n628, n629, n634, n635, n640, 
      n643, n646, n647, n652, n655, n656, n657, n659, n660, n661, n662, n663, 
      n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, 
      n676, n678, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, 
      n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, 
      n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, 
      n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, 
      n731, n732 : std_logic;

begin
   
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U144 : XOR2_X1 port map( A => B(50), B => A(50), Z => n590);
   U145 : XOR2_X1 port map( A => n591, B => n552, Z => SUM(49));
   U176 : XOR2_X1 port map( A => B(19), B => n718, Z => n682);
   U177 : XOR2_X1 port map( A => A(18), B => n684, Z => SUM(18));
   U178 : XOR2_X1 port map( A => carry_18_port, B => B(18), Z => n684);
   U179 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : CLKBUF_X1 port map( A => n569, Z => n542);
   U2 : AND2_X2 port map( A1 => net272285, A2 => net264574, ZN => net272082);
   U3 : INV_X1 port map( A => B(22), ZN => n668);
   U4 : INV_X1 port map( A => B(49), ZN => n717);
   U5 : INV_X1 port map( A => B(23), ZN => n664);
   U6 : INV_X1 port map( A => B(24), ZN => n698);
   U7 : OR2_X1 port map( A1 => n634, A2 => net275647, ZN => net275664);
   U8 : AND2_X1 port map( A1 => n713, A2 => n712, ZN => n589);
   U9 : AND2_X1 port map( A1 => n674, A2 => n673, ZN => net275643);
   U10 : INV_X1 port map( A => B(44), ZN => net272479);
   U11 : XOR2_X1 port map( A => A(21), B => B(21), Z => n543);
   U12 : CLKBUF_X1 port map( A => n573, Z => n544);
   U13 : CLKBUF_X1 port map( A => net270519, Z => net287683);
   U14 : CLKBUF_X1 port map( A => A(34), Z => n617);
   U15 : CLKBUF_X1 port map( A => n568, Z => n545);
   U16 : XNOR2_X1 port map( A => A(25), B => n699, ZN => n700);
   U17 : INV_X1 port map( A => B(25), ZN => n699);
   U18 : XNOR2_X1 port map( A => A(32), B => B(32), ZN => n598);
   U19 : CLKBUF_X1 port map( A => n638, Z => net270519);
   U20 : CLKBUF_X1 port map( A => A(48), Z => n546);
   U21 : BUF_X1 port map( A => n628, Z => n547);
   U22 : BUF_X1 port map( A => A(44), Z => n553);
   U23 : BUF_X1 port map( A => n680, Z => n705);
   U24 : OR2_X1 port map( A1 => n555, A2 => net264594, ZN => n548);
   U25 : BUF_X2 port map( A => A(33), Z => n622);
   U26 : AOI22_X1 port map( A1 => net287683, A2 => n622, B1 => n592, B2 => 
                           B(33), ZN => n549);
   U27 : AOI22_X1 port map( A1 => net287683, A2 => n622, B1 => n592, B2 => 
                           B(33), ZN => n562);
   U28 : BUF_X1 port map( A => n599, Z => net270507);
   U29 : BUF_X1 port map( A => net264589, Z => n600);
   U30 : NAND2_X1 port map( A1 => n665, A2 => n664, ZN => n672);
   U31 : AOI21_X1 port map( B1 => n574, B2 => n579, A => net264600, ZN => n550)
                           ;
   U32 : NOR2_X1 port map( A1 => n606, A2 => net272082, ZN => n551);
   U33 : AOI21_X1 port map( B1 => n730, B2 => n710, A => n594, ZN => n552);
   U34 : BUF_X1 port map( A => A(39), Z => n573);
   U35 : AND2_X1 port map( A1 => n659, A2 => n657, ZN => n554);
   U36 : AND2_X1 port map( A1 => n657, A2 => n659, ZN => n676);
   U37 : AND2_X1 port map( A1 => n563, A2 => net271193, ZN => n555);
   U38 : AOI21_X1 port map( B1 => n727, B2 => n706, A => B(46), ZN => n556);
   U39 : CLKBUF_X1 port map( A => A(29), Z => n607);
   U40 : INV_X1 port map( A => B(34), ZN => n557);
   U41 : XNOR2_X1 port map( A => A(34), B => n557, ZN => n637);
   U42 : AND2_X1 port map( A1 => net264596, A2 => net271690, ZN => n558);
   U43 : NAND2_X1 port map( A1 => n558, A2 => A(38), ZN => n716);
   U44 : NAND2_X1 port map( A1 => n600, A2 => n607, ZN => n559);
   U45 : NAND2_X1 port map( A1 => n650, A2 => B(29), ZN => n560);
   U46 : NAND2_X1 port map( A1 => n560, A2 => n559, ZN => n561);
   U47 : INV_X1 port map( A => B(46), ZN => n688);
   U48 : INV_X1 port map( A => B(27), ZN => net275693);
   U49 : AOI22_X1 port map( A1 => net287683, A2 => n622, B1 => n592, B2 => 
                           B(33), ZN => n623);
   U50 : AOI21_X1 port map( B1 => n562, B2 => n616, A => n636, ZN => n563);
   U51 : BUF_X1 port map( A => n639, Z => n592);
   U52 : NAND2_X1 port map( A1 => net270519, A2 => n622, ZN => n564);
   U53 : NAND2_X1 port map( A1 => n639, A2 => B(33), ZN => n565);
   U54 : NAND2_X1 port map( A1 => n565, A2 => n564, ZN => n566);
   U55 : AOI21_X1 port map( B1 => n553, B2 => n583, A => B(44), ZN => n606);
   U56 : AOI21_X1 port map( B1 => n566, B2 => A(34), A => B(34), ZN => n636);
   U57 : OAI21_X1 port map( B1 => n606, B2 => net272082, A => n708, ZN => n603)
                           ;
   U58 : INV_X1 port map( A => B(45), ZN => n708);
   U59 : XNOR2_X1 port map( A => n690, B => n687, ZN => SUM(46));
   U60 : XNOR2_X1 port map( A => n572, B => n574, ZN => SUM(41));
   U61 : CLKBUF_X1 port map( A => n614, Z => n574);
   U62 : AOI21_X1 port map( B1 => n574, B2 => n579, A => net264600, ZN => n611)
                           ;
   U63 : XNOR2_X1 port map( A => A(41), B => B(41), ZN => n572);
   U64 : NOR2_X1 port map( A1 => n618, A2 => n578, ZN => n614);
   U65 : OAI21_X1 port map( B1 => n614, B2 => A(41), A => B(41), ZN => n615);
   U66 : AND2_X1 port map( A1 => n571, A2 => n567, ZN => n578);
   U67 : INV_X1 port map( A => B(40), ZN => n567);
   U68 : XNOR2_X1 port map( A => A(40), B => n567, ZN => net271621);
   U69 : AOI21_X1 port map( B1 => n577, B2 => n573, A => n568, ZN => n571);
   U70 : INV_X1 port map( A => n621, ZN => n568);
   U71 : AOI21_X1 port map( B1 => n577, B2 => n544, A => n545, ZN => net273792)
                           ;
   U72 : OR2_X1 port map( A1 => n575, A2 => n568, ZN => n576);
   U73 : OAI21_X1 port map( B1 => n620, B2 => A(39), A => B(39), ZN => n621);
   U74 : AND2_X1 port map( A1 => n569, A2 => n573, ZN => n575);
   U75 : BUF_X1 port map( A => n569, Z => n577);
   U76 : BUF_X1 port map( A => n620, Z => n569);
   U77 : XNOR2_X1 port map( A => n542, B => n570, ZN => SUM(39));
   U78 : AOI21_X1 port map( B1 => n576, B2 => B(40), A => A(40), ZN => n618);
   U79 : CLKBUF_X1 port map( A => A(41), Z => n579);
   U80 : XNOR2_X1 port map( A => A(39), B => B(39), ZN => n570);
   U81 : NAND2_X1 port map( A1 => net275667, A2 => n698, ZN => n580);
   U82 : CLKBUF_X1 port map( A => A(47), Z => n581);
   U83 : NAND2_X1 port map( A1 => n608, A2 => n587, ZN => n584);
   U84 : OAI21_X1 port map( B1 => n608, B2 => n587, A => B(43), ZN => n585);
   U85 : XNOR2_X1 port map( A => n608, B => n582, ZN => SUM(43));
   U86 : NAND2_X1 port map( A1 => n584, A2 => n585, ZN => n583);
   U87 : AND2_X1 port map( A1 => n585, A2 => n584, ZN => net272285);
   U88 : XNOR2_X1 port map( A => A(44), B => net272479, ZN => net272480);
   U89 : INV_X1 port map( A => n553, ZN => net264574);
   U90 : NOR2_X1 port map( A1 => net272082, A2 => n606, ZN => net272919);
   U91 : XNOR2_X1 port map( A => A(43), B => B(43), ZN => n582);
   U92 : CLKBUF_X1 port map( A => A(43), Z => n587);
   U93 : BUF_X1 port map( A => n593, Z => n710);
   U94 : XNOR2_X1 port map( A => n613, B => n598, ZN => SUM(32));
   U95 : XNOR2_X1 port map( A => A(20), B => n667, ZN => n679);
   U96 : INV_X1 port map( A => B(20), ZN => n667);
   U97 : XNOR2_X1 port map( A => n586, B => n720, ZN => SUM(51));
   U98 : AOI22_X1 port map( A1 => n600, A2 => n607, B1 => n650, B2 => B(29), ZN
                           => n599);
   U99 : AOI21_X1 port map( B1 => net270507, B2 => n601, A => n648, ZN => n644)
                           ;
   U100 : NAND2_X1 port map( A1 => n644, A2 => net271069, ZN => net272365);
   U101 : XNOR2_X1 port map( A => n644, B => net271720, ZN => SUM(31));
   U102 : OAI21_X1 port map( B1 => n644, B2 => net271069, A => B(31), ZN => 
                           n645);
   U103 : AOI21_X1 port map( B1 => n561, B2 => A(30), A => B(30), ZN => n648);
   U104 : INV_X1 port map( A => A(30), ZN => n601);
   U105 : XNOR2_X1 port map( A => n649, B => net270507, ZN => SUM(30));
   U106 : XOR2_X1 port map( A => A(30), B => B(30), Z => n649);
   U107 : OR2_X1 port map( A1 => net264589, A2 => A(29), ZN => n650);
   U108 : INV_X1 port map( A => n651, ZN => net264589);
   U109 : AOI22_X1 port map( A1 => n605, A2 => n604, B1 => n654, B2 => B(28), 
                           ZN => n651);
   U110 : OR2_X1 port map( A1 => n653, A2 => A(28), ZN => n654);
   U111 : NOR2_X1 port map( A1 => net275685, A2 => net271609, ZN => n653);
   U112 : AND2_X1 port map( A1 => net264570, A2 => net273613, ZN => net271609);
   U113 : AND2_X1 port map( A1 => net275665, A2 => net275664, ZN => net273613);
   U114 : INV_X1 port map( A => A(27), ZN => net264570);
   U115 : AND2_X1 port map( A1 => net264570, A2 => net276693, ZN => n609);
   U116 : CLKBUF_X1 port map( A => A(28), Z => n604);
   U117 : XNOR2_X1 port map( A => n600, B => n610, ZN => SUM(29));
   U118 : XNOR2_X1 port map( A => A(29), B => B(29), ZN => n610);
   U119 : XNOR2_X1 port map( A => n602, B => n605, ZN => SUM(28));
   U120 : XNOR2_X1 port map( A => A(28), B => B(28), ZN => n602);
   U121 : NOR2_X1 port map( A1 => n609, A2 => net275685, ZN => n605);
   U122 : AND2_X1 port map( A1 => net275665, A2 => net275664, ZN => net276693);
   U123 : CLKBUF_X1 port map( A => n619, Z => n613);
   U124 : XNOR2_X1 port map( A => A(45), B => B(45), ZN => n689);
   U125 : AOI21_X1 port map( B1 => n623, B2 => n616, A => n636, ZN => n632);
   U126 : OAI21_X1 port map( B1 => n632, B2 => A(35), A => B(35), ZN => n633);
   U127 : INV_X1 port map( A => n617, ZN => n616);
   U128 : XNOR2_X1 port map( A => net270519, B => net271948, ZN => SUM(33));
   U129 : XNOR2_X1 port map( A => n549, B => n637, ZN => SUM(34));
   U130 : OR2_X1 port map( A1 => n638, A2 => A(33), ZN => n639);
   U131 : XNOR2_X1 port map( A => A(33), B => B(33), ZN => net271948);
   U132 : NOR2_X1 port map( A1 => n642, A2 => net270509, ZN => n638);
   U133 : AND2_X1 port map( A1 => net264572, A2 => n641, ZN => net270509);
   U134 : INV_X1 port map( A => A(32), ZN => net264572);
   U135 : AND2_X1 port map( A1 => n645, A2 => net272365, ZN => n641);
   U136 : AOI21_X1 port map( B1 => n619, B2 => A(32), A => B(32), ZN => n642);
   U137 : NAND2_X1 port map( A1 => n645, A2 => net272365, ZN => n619);
   U138 : INV_X1 port map( A => n611, ZN => net264601);
   U139 : INV_X1 port map( A => n615, ZN => net264600);
   U140 : NOR2_X1 port map( A1 => n630, A2 => n629, ZN => n626);
   U141 : OR2_X1 port map( A1 => n626, A2 => A(37), ZN => net271690);
   U142 : CLKBUF_X1 port map( A => n626, Z => net276573);
   U143 : AOI21_X1 port map( B1 => n626, B2 => A(37), A => B(37), ZN => n627);
   U146 : AND2_X1 port map( A1 => n628, A2 => n625, ZN => n629);
   U147 : INV_X1 port map( A => A(36), ZN => n625);
   U148 : AOI21_X1 port map( B1 => n548, B2 => A(36), A => B(36), ZN => n630);
   U149 : INV_X1 port map( A => n633, ZN => net264594);
   U150 : AOI21_X1 port map( B1 => n563, B2 => net271193, A => net264594, ZN =>
                           n628);
   U151 : CLKBUF_X1 port map( A => A(35), Z => net271193);
   U152 : XNOR2_X1 port map( A => n563, B => net272213, ZN => SUM(35));
   U153 : XNOR2_X1 port map( A => n547, B => n631, ZN => SUM(36));
   U154 : XOR2_X1 port map( A => A(36), B => B(36), Z => n631);
   U155 : AOI21_X1 port map( B1 => A(27), B2 => net275663, A => B(27), ZN => 
                           net275685);
   U156 : NAND2_X1 port map( A1 => n635, A2 => net275664, ZN => net275663);
   U157 : NAND2_X1 port map( A1 => net275668, A2 => B(26), ZN => n635);
   U158 : NAND2_X1 port map( A1 => net275668, A2 => B(26), ZN => net275665);
   U159 : INV_X1 port map( A => A(26), ZN => n634);
   U160 : XNOR2_X1 port map( A => net275652, B => n634, ZN => SUM(26));
   U161 : XNOR2_X1 port map( A => A(27), B => net275693, ZN => n658);
   U162 : XNOR2_X1 port map( A => net272480, B => net272285, ZN => SUM(44));
   U163 : AOI21_X1 port map( B1 => n550, B2 => n640, A => n612, ZN => n608);
   U164 : AOI21_X1 port map( B1 => net264601, B2 => A(42), A => B(42), ZN => 
                           n612);
   U165 : INV_X1 port map( A => A(42), ZN => n640);
   U166 : XNOR2_X1 port map( A => n643, B => n550, ZN => SUM(42));
   U167 : XOR2_X1 port map( A => A(42), B => B(42), Z => n643);
   U168 : NAND2_X1 port map( A1 => n677, A2 => A(20), ZN => n669);
   U169 : INV_X1 port map( A => n677, ZN => n661);
   U170 : INV_X1 port map( A => net274721, ZN => n670);
   U171 : OAI21_X1 port map( B1 => n685, B2 => n670, A => B(21), ZN => n656);
   U172 : NAND2_X1 port map( A1 => n656, A2 => n655, ZN => n652);
   U173 : NAND2_X1 port map( A1 => A(22), A2 => n652, ZN => n671);
   U174 : NAND2_X1 port map( A1 => n685, A2 => n670, ZN => n655);
   U175 : INV_X1 port map( A => A(20), ZN => n662);
   U180 : AND2_X1 port map( A1 => n656, A2 => n655, ZN => n675);
   U181 : NAND2_X1 port map( A1 => n671, A2 => n668, ZN => n659);
   U182 : NAND2_X1 port map( A1 => n663, A2 => n675, ZN => n657);
   U183 : INV_X1 port map( A => n675, ZN => net272472);
   U184 : XNOR2_X1 port map( A => A(23), B => B(23), ZN => n666);
   U185 : NAND2_X1 port map( A1 => n678, A2 => B(23), ZN => n674);
   U186 : INV_X1 port map( A => A(23), ZN => n665);
   U187 : NAND2_X1 port map( A1 => n669, A2 => n667, ZN => n647);
   U188 : NAND2_X1 port map( A1 => n661, A2 => n662, ZN => n646);
   U189 : NAND2_X1 port map( A1 => n647, A2 => n646, ZN => net274721);
   U190 : INV_X1 port map( A => A(22), ZN => n663);
   U191 : XNOR2_X1 port map( A => n661, B => n679, ZN => SUM(20));
   U192 : CLKBUF_X1 port map( A => A(23), Z => n678);
   U193 : CLKBUF_X1 port map( A => A(21), Z => n685);
   U194 : NAND2_X1 port map( A1 => n674, A2 => n673, ZN => n660);
   U195 : NAND2_X1 port map( A1 => A(24), A2 => n660, ZN => net275667);
   U196 : XNOR2_X1 port map( A => n666, B => n554, ZN => SUM(23));
   U197 : NAND2_X1 port map( A1 => n672, A2 => n676, ZN => n673);
   U198 : XNOR2_X1 port map( A => A(22), B => B(22), ZN => net270022);
   U199 : CLKBUF_X1 port map( A => net274721, Z => net274030);
   U200 : INV_X1 port map( A => A(48), ZN => n686);
   U201 : XNOR2_X1 port map( A => n658, B => net276693, ZN => SUM(27));
   U202 : AOI22_X1 port map( A1 => n551, A2 => B(45), B1 => n603, B2 => n691, 
                           ZN => n687);
   U203 : XNOR2_X1 port map( A => A(46), B => n688, ZN => n690);
   U204 : XNOR2_X1 port map( A => n689, B => net272919, ZN => SUM(45));
   U205 : CLKBUF_X1 port map( A => A(45), Z => n691);
   U206 : XNOR2_X1 port map( A => n697, B => net275676, ZN => SUM(24));
   U207 : INV_X1 port map( A => net275643, ZN => net275676);
   U208 : INV_X1 port map( A => A(25), ZN => n694);
   U209 : XNOR2_X1 port map( A => A(24), B => B(24), ZN => n697);
   U210 : INV_X1 port map( A => A(24), ZN => net275641);
   U211 : NAND2_X1 port map( A1 => n580, A2 => n693, ZN => n692);
   U212 : NAND2_X1 port map( A1 => n701, A2 => n694, ZN => n695);
   U213 : OAI21_X1 port map( B1 => n694, B2 => n692, A => n699, ZN => n696);
   U214 : NAND2_X1 port map( A1 => net275647, A2 => n634, ZN => net275668);
   U215 : NAND2_X1 port map( A1 => n695, A2 => n696, ZN => net275647);
   U216 : XNOR2_X1 port map( A => n702, B => B(26), ZN => net275652);
   U217 : XNOR2_X1 port map( A => n700, B => n701, ZN => SUM(25));
   U218 : NAND2_X1 port map( A1 => net275643, A2 => net275641, ZN => n693);
   U219 : NAND2_X1 port map( A1 => n693, A2 => n580, ZN => n701);
   U220 : NAND2_X1 port map( A1 => n695, A2 => n703, ZN => n702);
   U221 : OAI21_X1 port map( B1 => n694, B2 => n692, A => n699, ZN => n703);
   U222 : AOI22_X1 port map( A1 => n551, A2 => B(45), B1 => n603, B2 => n691, 
                           ZN => n704);
   U223 : INV_X1 port map( A => n731, ZN => n706);
   U224 : NOR2_X1 port map( A1 => n556, A2 => n709, ZN => n707);
   U225 : AND2_X1 port map( A1 => n704, A2 => n731, ZN => n709);
   U226 : NOR2_X1 port map( A1 => n556, A2 => n709, ZN => n596);
   U227 : XNOR2_X1 port map( A => n707, B => n711, ZN => SUM(47));
   U228 : XNOR2_X1 port map( A => B(47), B => A(47), ZN => n711);
   U229 : XNOR2_X1 port map( A => A(35), B => B(35), ZN => net272213);
   U230 : NAND2_X1 port map( A1 => B(49), A2 => n719, ZN => n712);
   U231 : NAND2_X1 port map( A1 => n591, A2 => n552, ZN => n713);
   U232 : AND2_X1 port map( A1 => net264596, A2 => net271690, ZN => n714);
   U233 : CLKBUF_X1 port map( A => A(31), Z => net271069);
   U234 : XNOR2_X1 port map( A => n715, B => n558, ZN => SUM(38));
   U235 : XNOR2_X1 port map( A => A(38), B => B(38), ZN => n715);
   U236 : XNOR2_X1 port map( A => A(31), B => B(31), ZN => net271720);
   U237 : NAND2_X1 port map( A1 => n624, A2 => n716, ZN => n620);
   U238 : XNOR2_X1 port map( A => net271621, B => net273792, ZN => SUM(40));
   U239 : XNOR2_X1 port map( A => A(49), B => n717, ZN => n591);
   U240 : INV_X1 port map( A => n732, ZN => n718);
   U241 : CLKBUF_X1 port map( A => A(49), Z => n719);
   U242 : NOR2_X1 port map( A1 => n723, A2 => n726, ZN => n593);
   U243 : XOR2_X1 port map( A => B(51), B => A(51), Z => n720);
   U244 : XNOR2_X1 port map( A => net276573, B => n721, ZN => SUM(37));
   U245 : XNOR2_X1 port map( A => A(37), B => B(37), ZN => n721);
   U246 : OR2_X1 port map( A1 => n726, A2 => n723, ZN => n722);
   U247 : AND2_X1 port map( A1 => n707, A2 => n581, ZN => n723);
   U248 : INV_X1 port map( A => n546, ZN => n730);
   U249 : XNOR2_X1 port map( A => net270022, B => net272472, ZN => SUM(22));
   U250 : XNOR2_X1 port map( A => n686, B => B(48), ZN => n595);
   U251 : INV_X1 port map( A => n683, ZN => n729);
   U252 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U253 : XNOR2_X1 port map( A => n543, B => net274030, ZN => SUM(21));
   U254 : OAI21_X1 port map( B1 => n596, B2 => n581, A => B(47), ZN => n597);
   U255 : INV_X1 port map( A => A(19), ZN => n732);
   U256 : OAI21_X1 port map( B1 => n728, B2 => A(19), A => B(19), ZN => n681);
   U257 : XNOR2_X1 port map( A => n705, B => n682, ZN => SUM(19));
   U258 : OAI21_X1 port map( B1 => n705, B2 => n732, A => n681, ZN => n677);
   U259 : INV_X1 port map( A => n680, ZN => n728);
   U260 : OAI21_X1 port map( B1 => B(18), B2 => A(18), A => n729, ZN => n680);
   U261 : AOI21_X1 port map( B1 => A(18), B2 => B(18), A => carry_18_port, ZN 
                           => n683);
   U262 : AOI21_X1 port map( B1 => n725, B2 => A(50), A => B(50), ZN => n588);
   U263 : INV_X1 port map( A => n597, ZN => n726);
   U264 : OAI21_X1 port map( B1 => n714, B2 => A(38), A => B(38), ZN => n624);
   U265 : INV_X1 port map( A => n588, ZN => n724);
   U266 : INV_X1 port map( A => n627, ZN => net264596);
   U267 : OAI21_X1 port map( B1 => A(50), B2 => n725, A => n724, ZN => n586);
   U268 : AOI21_X1 port map( B1 => n722, B2 => n546, A => B(48), ZN => n594);
   U269 : INV_X1 port map( A => A(46), ZN => n731);
   U270 : XNOR2_X1 port map( A => n589, B => n590, ZN => SUM(50));
   U271 : INV_X1 port map( A => n589, ZN => n725);
   U272 : XNOR2_X1 port map( A => n593, B => n595, ZN => SUM(48));
   U273 : INV_X1 port map( A => n704, ZN => n727);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT50_DW01_add_0 is

   port( A, B : in std_logic_vector (49 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (49 downto 0);  CO : out std_logic);

end RCA_NBIT50_DW01_add_0;

architecture SYN_rpl of RCA_NBIT50_DW01_add_0 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_15_port, carry_14_port, carry_13_port, carry_12_port, 
      carry_11_port, carry_10_port, carry_9_port, carry_8_port, carry_7_port, 
      carry_6_port, carry_5_port, carry_4_port, carry_3_port, carry_2_port, n1,
      carry_44_port, carry_16_port, carry_43_port, carry_42_port, net76696, 
      n506, n507, n508, n509, n510, n511, n513, n517, n518, n519, n522, n523, 
      n526, n528, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, 
      n541, n543, n544, n546, n547, n549, n550, n551, n552, n553, n556, n564, 
      n569, n573, n576, n578, n585, n588, n589, n590, n591, n592, net264533, 
      net264542, net264544, net264547, net264556, net269882, net272303, 
      net272512, net272842, net273614, net275721, net275802, net276032, 
      net279674, net280979, net280944, net280938, n529, n525, net282889, 
      net279641, net269896, net279610, net276012, net270558, net270556, 
      net270424, net264534, n565, n563, n561, n559, n558, n557, net272302, 
      net264540, n587, n586, n584, n583, n582, n580, n577, n466, n467, n468, 
      n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, 
      n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, 
      n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, 
      n505, n512, n514, n515, n516, n520, n521, n524, n527, n530, n542, n545, 
      n548, n554, n555, n560, n562, n566, n567, n568, n570, n571, n572, n574, 
      n575, n579, n581, n593, n594, n595, n596, n597, n598, n599, n600, n601, 
      n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, 
      n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, 
      n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, 
      n638, n639, n640, n641 : std_logic;

begin
   
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_44 : FA_X1 port map( A => A(44), B => B(44), CI => carry_44_port, CO => 
                           net76696, S => SUM(44));
   U1_41 : FA_X1 port map( A => A(41), B => B(41), CI => n477, CO => 
                           carry_42_port, S => SUM(41));
   U1_43 : FA_X1 port map( A => A(43), B => B(43), CI => carry_43_port, CO => 
                           carry_44_port, S => SUM(43));
   U1_42 : FA_X1 port map( A => A(42), B => B(42), CI => carry_42_port, CO => 
                           carry_43_port, S => SUM(42));
   U131 : XOR2_X1 port map( A => B(49), B => A(49), Z => n509);
   U157 : XOR2_X1 port map( A => B(17), B => n612, Z => n590);
   U158 : XOR2_X1 port map( A => n620, B => n592, Z => SUM(16));
   U159 : XOR2_X1 port map( A => carry_16_port, B => B(16), Z => n592);
   U160 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U155 : XOR2_X1 port map( A => n587, B => n488, Z => SUM(18));
   U1 : BUF_X1 port map( A => A(36), Z => n600);
   U2 : CLKBUF_X1 port map( A => n525, Z => n520);
   U3 : BUF_X1 port map( A => n472, Z => n466);
   U4 : BUF_X1 port map( A => n582, Z => n487);
   U5 : AOI22_X1 port map( A1 => net282889, A2 => n501, B1 => n565, B2 => B(25)
                           , ZN => n561);
   U6 : OR2_X1 port map( A1 => n564, A2 => A(25), ZN => n565);
   U7 : OAI221_X1 port map( B1 => net264544, B2 => n512, C1 => net264544, C2 =>
                           n514, A => net280938, ZN => net282889);
   U8 : CLKBUF_X1 port map( A => A(26), Z => n467);
   U9 : BUF_X2 port map( A => A(45), Z => n605);
   U10 : AND2_X1 port map( A1 => n566, A2 => n567, ZN => net264544);
   U11 : BUF_X1 port map( A => n549, Z => n527);
   U12 : CLKBUF_X1 port map( A => A(46), Z => n595);
   U13 : BUF_X1 port map( A => n470, Z => n468);
   U14 : OAI21_X1 port map( B1 => n521, B2 => n520, A => net264556, ZN => n469)
                           ;
   U15 : AOI22_X1 port map( A1 => n575, A2 => n466, B1 => n579, B2 => n574, ZN 
                           => n470);
   U16 : AOI21_X1 port map( B1 => n497, B2 => n467, A => B(26), ZN => n471);
   U17 : INV_X1 port map( A => B(37), ZN => n473);
   U18 : CLKBUF_X1 port map( A => n588, Z => n615);
   U19 : OAI21_X1 port map( B1 => B(45), B2 => n605, A => n629, ZN => n472);
   U20 : XNOR2_X1 port map( A => A(37), B => n473, ZN => n515);
   U21 : NAND2_X1 port map( A1 => n475, A2 => n603, ZN => n474);
   U22 : OAI21_X1 port map( B1 => n597, B2 => net273614, A => B(39), ZN => n475
                           );
   U23 : BUF_X1 port map( A => n585, Z => n488);
   U24 : AND2_X1 port map( A1 => n631, A2 => n480, ZN => n476);
   U25 : INV_X1 port map( A => B(19), ZN => n486);
   U26 : INV_X1 port map( A => B(46), ZN => n574);
   U27 : BUF_X1 port map( A => n537, Z => n604);
   U28 : AND2_X1 port map( A1 => n631, A2 => n480, ZN => n479);
   U29 : NAND2_X1 port map( A1 => n506, A2 => n478, ZN => n477);
   U30 : NAND2_X1 port map( A1 => n474, A2 => A(40), ZN => n478);
   U31 : INV_X1 port map( A => n476, ZN => n528);
   U32 : INV_X1 port map( A => B(21), ZN => n485);
   U33 : INV_X1 port map( A => B(18), ZN => n490);
   U34 : OR2_X1 port map( A1 => n600, A2 => n531, ZN => n480);
   U35 : INV_X1 port map( A => B(26), ZN => net270556);
   U36 : BUF_X1 port map( A => A(22), Z => net275721);
   U37 : OAI21_X1 port map( B1 => n491, B2 => n492, A => B(21), ZN => n577);
   U38 : OAI21_X1 port map( B1 => n576, B2 => n482, A => n577, ZN => n573);
   U39 : BUF_X1 port map( A => A(21), Z => n492);
   U40 : INV_X1 port map( A => n492, ZN => n482);
   U41 : AND2_X1 port map( A1 => net264540, A2 => net272302, ZN => n491);
   U42 : INV_X1 port map( A => n580, ZN => net264540);
   U43 : NAND2_X1 port map( A1 => net264540, A2 => net272302, ZN => n576);
   U44 : AOI21_X1 port map( B1 => n493, B2 => A(20), A => B(20), ZN => n580);
   U45 : OAI21_X1 port map( B1 => n487, B2 => n481, A => n583, ZN => n493);
   U46 : INV_X1 port map( A => A(19), ZN => n481);
   U47 : XNOR2_X1 port map( A => n487, B => n584, ZN => SUM(19));
   U48 : XNOR2_X1 port map( A => A(21), B => n485, ZN => n578);
   U49 : OR2_X1 port map( A1 => A(20), A2 => n493, ZN => net272302);
   U50 : XNOR2_X1 port map( A => A(20), B => B(20), ZN => net269896);
   U51 : OAI21_X1 port map( B1 => n484, B2 => A(19), A => B(19), ZN => n583);
   U52 : INV_X1 port map( A => n582, ZN => n484);
   U53 : XNOR2_X1 port map( A => A(19), B => n486, ZN => n584);
   U54 : OAI21_X1 port map( B1 => n489, B2 => n488, A => n483, ZN => n582);
   U55 : INV_X1 port map( A => n586, ZN => n483);
   U56 : AOI21_X1 port map( B1 => n585, B2 => A(18), A => B(18), ZN => n586);
   U57 : CLKBUF_X1 port map( A => A(18), Z => n489);
   U58 : CLKBUF_X1 port map( A => n493, Z => net279641);
   U59 : XNOR2_X1 port map( A => A(18), B => n490, ZN => n587);
   U60 : AOI21_X1 port map( B1 => n500, B2 => n499, A => n498, ZN => n494);
   U61 : CLKBUF_X1 port map( A => n547, Z => n495);
   U62 : AOI21_X1 port map( B1 => n500, B2 => n499, A => n498, ZN => n496);
   U63 : XNOR2_X1 port map( A => n494, B => n557, ZN => SUM(28));
   U64 : XOR2_X1 port map( A => A(28), B => B(28), Z => n557);
   U65 : INV_X1 port map( A => n559, ZN => n498);
   U66 : OAI21_X1 port map( B1 => n502, B2 => n558, A => B(27), ZN => n559);
   U67 : NOR2_X1 port map( A1 => n504, A2 => n471, ZN => n558);
   U68 : AND2_X1 port map( A1 => net264534, A2 => n561, ZN => n504);
   U69 : INV_X1 port map( A => A(26), ZN => net264534);
   U70 : AOI21_X1 port map( B1 => n561, B2 => net264534, A => net279610, ZN => 
                           net276012);
   U71 : BUF_X1 port map( A => A(27), Z => n502);
   U72 : CLKBUF_X1 port map( A => n502, Z => n499);
   U73 : BUF_X1 port map( A => net276012, Z => n500);
   U74 : INV_X1 port map( A => A(28), ZN => net264533);
   U75 : AOI21_X1 port map( B1 => net264547, B2 => net279674, A => B(28), ZN =>
                           n556);
   U76 : AOI21_X1 port map( B1 => net264547, B2 => net279674, A => B(28), ZN =>
                           net276032);
   U77 : XNOR2_X1 port map( A => A(27), B => B(27), ZN => net270558);
   U78 : AOI21_X1 port map( B1 => n497, B2 => n467, A => B(26), ZN => net279610
                           );
   U79 : INV_X1 port map( A => n503, ZN => n497);
   U80 : AOI22_X1 port map( A1 => net282889, A2 => n501, B1 => n565, B2 => 
                           B(25), ZN => n503);
   U81 : CLKBUF_X1 port map( A => A(25), Z => n501);
   U82 : XNOR2_X1 port map( A => n563, B => n561, ZN => SUM(26));
   U83 : XNOR2_X1 port map( A => A(26), B => net270556, ZN => n563);
   U84 : XNOR2_X1 port map( A => net270558, B => net276012, ZN => SUM(27));
   U85 : XNOR2_X1 port map( A => net270424, B => net282889, ZN => SUM(25));
   U86 : XNOR2_X1 port map( A => A(25), B => B(25), ZN => net270424);
   U87 : CLKBUF_X1 port map( A => n641, Z => n505);
   U88 : XNOR2_X1 port map( A => net269896, B => net279641, ZN => SUM(20));
   U89 : BUF_X1 port map( A => n573, Z => net272303);
   U90 : INV_X1 port map( A => B(24), ZN => n514);
   U91 : XNOR2_X1 port map( A => A(24), B => n514, ZN => n569);
   U92 : OAI221_X1 port map( B1 => net280979, B2 => n512, C1 => net280979, C2 
                           => n514, A => net280938, ZN => n564);
   U93 : INV_X1 port map( A => A(24), ZN => n512);
   U94 : XNOR2_X1 port map( A => n516, B => n520, ZN => SUM(38));
   U95 : OAI21_X1 port map( B1 => n520, B2 => n521, A => net264556, ZN => n522)
                           ;
   U96 : XNOR2_X1 port map( A => A(38), B => B(38), ZN => n516);
   U97 : OAI21_X1 port map( B1 => n524, B2 => n528, A => n529, ZN => n525);
   U98 : AOI21_X1 port map( B1 => n525, B2 => A(38), A => B(38), ZN => n526);
   U99 : OAI21_X1 port map( B1 => n479, B2 => A(37), A => B(37), ZN => n529);
   U100 : XNOR2_X1 port map( A => n515, B => n528, ZN => SUM(37));
   U101 : INV_X1 port map( A => A(37), ZN => n524);
   U102 : CLKBUF_X1 port map( A => A(38), Z => n521);
   U103 : BUF_X1 port map( A => A(39), Z => n597);
   U104 : NOR2_X1 port map( A1 => n573, A2 => B(22), ZN => n542);
   U105 : NOR2_X1 port map( A1 => n542, A2 => n530, ZN => net264542);
   U106 : NAND2_X1 port map( A1 => A(24), A2 => B(24), ZN => net280938);
   U107 : INV_X1 port map( A => net272512, ZN => n555);
   U108 : INV_X1 port map( A => A(23), ZN => n548);
   U109 : NOR2_X1 port map( A1 => A(22), A2 => B(22), ZN => n530);
   U110 : INV_X1 port map( A => net272303, ZN => net280944);
   U111 : NAND2_X1 port map( A1 => B(22), A2 => net275721, ZN => n560);
   U112 : NOR2_X1 port map( A1 => net275721, A2 => B(22), ZN => n545);
   U113 : XNOR2_X1 port map( A => A(22), B => B(22), ZN => net269882);
   U114 : OAI211_X1 port map( C1 => n545, C2 => net280944, A => n548, B => n560
                           , ZN => n562);
   U115 : NAND2_X1 port map( A1 => n562, A2 => B(23), ZN => n566);
   U116 : AND2_X1 port map( A1 => n566, A2 => n567, ZN => net280979);
   U117 : XNOR2_X1 port map( A => n555, B => n554, ZN => SUM(23));
   U118 : XNOR2_X1 port map( A => A(23), B => B(23), ZN => n554);
   U119 : OR2_X1 port map( A1 => n548, A2 => net272512, ZN => n567);
   U120 : CLKBUF_X1 port map( A => n544, Z => n617);
   U121 : INV_X1 port map( A => net264533, ZN => net279674);
   U122 : NOR2_X1 port map( A1 => n556, A2 => net272842, ZN => n568);
   U123 : BUF_X1 port map( A => A(47), Z => n570);
   U124 : BUF_X1 port map( A => A(29), Z => n613);
   U125 : INV_X1 port map( A => n595, ZN => n575);
   U126 : AND2_X1 port map( A1 => n494, A2 => net264533, ZN => net272842);
   U127 : OAI22_X1 port map( A1 => n622, A2 => n604, B1 => B(34), B2 => n538, 
                           ZN => n571);
   U128 : XNOR2_X1 port map( A => A(46), B => n574, ZN => n518);
   U129 : AOI22_X1 port map( A1 => n575, A2 => n466, B1 => n579, B2 => n574, ZN
                           => n572);
   U130 : NAND2_X1 port map( A1 => n593, A2 => n595, ZN => n579);
   U132 : CLKBUF_X1 port map( A => A(32), Z => n609);
   U133 : XNOR2_X1 port map( A => n581, B => n605, ZN => SUM(45));
   U134 : XNOR2_X1 port map( A => net76696, B => B(45), ZN => n581);
   U135 : INV_X1 port map( A => n517, ZN => n593);
   U136 : OAI21_X1 port map( B1 => n552, B2 => n613, A => B(29), ZN => n594);
   U137 : CLKBUF_X1 port map( A => A(31), Z => n596);
   U138 : INV_X1 port map( A => n534, ZN => n598);
   U139 : INV_X1 port map( A => n469, ZN => net275802);
   U140 : OAI22_X1 port map( A1 => n570, A2 => n468, B1 => B(47), B2 => n513, 
                           ZN => n599);
   U141 : XNOR2_X1 port map( A => n611, B => n601, ZN => SUM(32));
   U142 : XNOR2_X1 port map( A => A(32), B => B(32), ZN => n601);
   U143 : NAND2_X1 port map( A1 => n610, A2 => n594, ZN => n602);
   U144 : AND2_X1 port map( A1 => n553, A2 => n610, ZN => n549);
   U145 : NAND2_X1 port map( A1 => n597, A2 => net275802, ZN => n603);
   U146 : NAND2_X1 port map( A1 => n523, A2 => n603, ZN => n507);
   U147 : INV_X1 port map( A => n522, ZN => net273614);
   U148 : XNOR2_X1 port map( A => A(39), B => B(39), ZN => n623);
   U149 : OAI21_X1 port map( B1 => n615, B2 => n641, A => n589, ZN => n585);
   U150 : XNOR2_X1 port map( A => n470, B => n624, ZN => SUM(47));
   U151 : AND2_X1 port map( A1 => n549, A2 => n638, ZN => n606);
   U152 : NOR2_X1 port map( A1 => n606, A2 => n550, ZN => n547);
   U153 : OAI21_X1 port map( B1 => n609, B2 => n611, A => n634, ZN => n607);
   U154 : NOR2_X1 port map( A1 => net276032, A2 => net272842, ZN => n552);
   U156 : XNOR2_X1 port map( A => n633, B => n608, ZN => SUM(33));
   U161 : XNOR2_X1 port map( A => A(33), B => B(33), ZN => n608);
   U162 : XOR2_X1 port map( A => A(40), B => B(40), Z => n627);
   U163 : NAND2_X1 port map( A1 => n568, A2 => n613, ZN => n610);
   U164 : OAI21_X1 port map( B1 => net272303, B2 => net275721, A => net264542, 
                           ZN => net272512);
   U165 : INV_X1 port map( A => n617, ZN => n611);
   U166 : INV_X1 port map( A => n505, ZN => n612);
   U167 : XOR2_X1 port map( A => A(30), B => B(30), Z => n551);
   U168 : XNOR2_X1 port map( A => A(35), B => B(35), ZN => n536);
   U169 : CLKBUF_X1 port map( A => A(16), Z => n614);
   U170 : XNOR2_X1 port map( A => n616, B => n568, ZN => SUM(29));
   U171 : XNOR2_X1 port map( A => A(29), B => B(29), ZN => n616);
   U172 : INV_X1 port map( A => n632, ZN => n618);
   U173 : AND2_X1 port map( A1 => n640, A2 => n607, ZN => n619);
   U174 : NOR2_X1 port map( A1 => n541, A2 => n619, ZN => n537);
   U175 : CLKBUF_X1 port map( A => n614, Z => n620);
   U176 : XNOR2_X1 port map( A => n508, B => n509, ZN => SUM(49));
   U177 : INV_X1 port map( A => n540, ZN => n621);
   U178 : CLKBUF_X1 port map( A => A(34), Z => n622);
   U179 : XNOR2_X1 port map( A => n623, B => net275802, ZN => SUM(39));
   U180 : OAI22_X1 port map( A1 => n570, A2 => n468, B1 => n513, B2 => B(47), 
                           ZN => n511);
   U181 : AND2_X1 port map( A1 => n572, A2 => n570, ZN => n513);
   U182 : INV_X1 port map( A => n607, ZN => n633);
   U183 : AND2_X1 port map( A1 => n628, A2 => A(48), ZN => n510);
   U184 : XNOR2_X1 port map( A => B(47), B => A(47), ZN => n624);
   U185 : XOR2_X1 port map( A => n599, B => n625, Z => SUM(48));
   U186 : XNOR2_X1 port map( A => B(48), B => A(48), ZN => n625);
   U187 : XNOR2_X1 port map( A => n495, B => n626, ZN => SUM(31));
   U188 : XNOR2_X1 port map( A => A(31), B => B(31), ZN => n626);
   U189 : INV_X1 port map( A => n496, ZN => net264547);
   U190 : INV_X1 port map( A => n588, ZN => n636);
   U191 : INV_X1 port map( A => A(33), ZN => n640);
   U192 : XNOR2_X1 port map( A => n472, B => n518, ZN => SUM(46));
   U193 : XNOR2_X1 port map( A => n627, B => n630, ZN => SUM(40));
   U194 : INV_X1 port map( A => n526, ZN => net264556);
   U195 : OAI21_X1 port map( B1 => B(45), B2 => n605, A => n629, ZN => n517);
   U196 : INV_X1 port map( A => n519, ZN => n629);
   U197 : AOI21_X1 port map( B1 => A(45), B2 => B(45), A => net76696, ZN => 
                           n519);
   U198 : XNOR2_X1 port map( A => net269882, B => net272303, ZN => SUM(22));
   U199 : OAI22_X1 port map( A1 => n510, A2 => B(48), B1 => n628, B2 => A(48), 
                           ZN => n508);
   U200 : AOI21_X1 port map( B1 => A(16), B2 => B(16), A => carry_16_port, ZN 
                           => n591);
   U201 : XNOR2_X1 port map( A => n615, B => n590, ZN => SUM(17));
   U202 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U203 : XNOR2_X1 port map( A => n531, B => n533, ZN => SUM(36));
   U204 : XNOR2_X1 port map( A => A(34), B => B(34), ZN => n539);
   U205 : AOI21_X1 port map( B1 => n635, B2 => A(32), A => B(32), ZN => n543);
   U206 : XNOR2_X1 port map( A => A(36), B => B(36), ZN => n533);
   U207 : AOI21_X1 port map( B1 => n531, B2 => n600, A => B(36), ZN => n532);
   U208 : INV_X1 port map( A => n474, ZN => n630);
   U209 : OAI21_X1 port map( B1 => n507, B2 => A(40), A => B(40), ZN => n506);
   U210 : INV_X1 port map( A => n571, ZN => n632);
   U211 : INV_X1 port map( A => n544, ZN => n635);
   U212 : OR2_X1 port map( A1 => A(31), A2 => B(31), ZN => n546);
   U213 : OAI21_X1 port map( B1 => net273614, B2 => n597, A => B(39), ZN => 
                           n523);
   U214 : INV_X1 port map( A => A(30), ZN => n638);
   U215 : AOI22_X1 port map( A1 => n596, A2 => B(31), B1 => n546, B2 => n547, 
                           ZN => n544);
   U216 : OAI21_X1 port map( B1 => n552, B2 => n613, A => B(29), ZN => n553);
   U217 : XNOR2_X1 port map( A => n569, B => net264544, ZN => SUM(24));
   U218 : XNOR2_X1 port map( A => n576, B => n578, ZN => SUM(21));
   U219 : INV_X1 port map( A => A(35), ZN => n639);
   U220 : AOI21_X1 port map( B1 => A(30), B2 => n602, A => B(30), ZN => n550);
   U221 : AOI21_X1 port map( B1 => n621, B2 => A(33), A => B(33), ZN => n541);
   U222 : INV_X1 port map( A => A(17), ZN => n641);
   U223 : INV_X1 port map( A => n511, ZN => n628);
   U224 : OAI21_X1 port map( B1 => n609, B2 => n611, A => n634, ZN => n540);
   U225 : INV_X1 port map( A => n543, ZN => n634);
   U226 : OAI21_X1 port map( B1 => n636, B2 => A(17), A => B(17), ZN => n589);
   U227 : XNOR2_X1 port map( A => n536, B => n632, ZN => SUM(35));
   U228 : INV_X1 port map( A => n532, ZN => n631);
   U229 : OAI21_X1 port map( B1 => B(16), B2 => n614, A => n637, ZN => n588);
   U230 : INV_X1 port map( A => n591, ZN => n637);
   U231 : OAI22_X1 port map( A1 => n622, A2 => n604, B1 => n538, B2 => B(34), 
                           ZN => n534);
   U232 : AND2_X1 port map( A1 => n537, A2 => A(34), ZN => n538);
   U233 : OAI21_X1 port map( B1 => n618, B2 => n639, A => n535, ZN => n531);
   U234 : OAI21_X1 port map( B1 => n598, B2 => A(35), A => B(35), ZN => n535);
   U235 : XNOR2_X1 port map( A => n604, B => n539, ZN => SUM(34));
   U236 : XNOR2_X1 port map( A => n527, B => n551, ZN => SUM(30));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT48_DW01_add_0 is

   port( A, B : in std_logic_vector (47 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (47 downto 0);  CO : out std_logic);

end RCA_NBIT48_DW01_add_0;

architecture SYN_rpl of RCA_NBIT48_DW01_add_0 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_14_port, carry_13_port, carry_12_port, carry_11_port, 
      carry_10_port, carry_9_port, carry_8_port, carry_7_port, carry_6_port, 
      carry_5_port, carry_4_port, carry_3_port, carry_2_port, n1, n554, n555, 
      n556, n559, n560, n562, n563, n565, n566, n568, n569, n571, n572, n574, 
      n575, n577, n578, n580, n581, n583, n584, n586, n587, n589, n590, n592, 
      n593, n596, n604, n607, n608, n611, n637, n641, n643, n644, n646, n647, 
      n649, n650, n652, n653, net264480, net264508, net270458, net270516, 
      net270769, net271055, net271478, net276011, net271728, net264500, 
      net279549, net279539, net279508, net279507, net279503, net279500, 
      net279490, net279489, net279488, net288445, net270456, net264503, n614, 
      n610, net271625, n626, net274277, net274244, net274177, net273969, 
      net273960, net271811, net271340, net270610, net264490, n623, n619, 
      net276125, net273126, net272305, net271455, n620, n617, n613, net279521, 
      net279520, net279512, net279504, net271806, net271341, net270885, n629, 
      n605, n602, n601, n600, n599, n595, n510, n511, n512, n513, n514, n515, 
      n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, 
      n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, 
      n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, 
      n552, n553, n557, n558, n561, n564, n567, n570, n573, n576, n579, n582, 
      n585, n588, n591, n594, n597, n598, n603, n606, n609, n612, n615, n616, 
      n618, n621, n622, n624, n625, n627, n628, n630, n631, n632, n633, n634, 
      n635, n636, n638, n639, n640, n642, n645, n648, n651, n654, n655, n656, 
      n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, 
      n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, 
      n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, 
      n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, 
      n705, n706, n707, n708, n709, n710 : std_logic;

begin
   
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U121 : XOR2_X1 port map( A => B(47), B => A(47), Z => n555);
   U176 : XOR2_X1 port map( A => n683, B => n650, Z => SUM(15));
   U177 : XOR2_X1 port map( A => B(15), B => n658, Z => n650);
   U178 : XOR2_X1 port map( A => n682, B => n653, Z => SUM(14));
   U179 : XOR2_X1 port map( A => carry_14_port, B => B(14), Z => n653);
   U180 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U144 : XOR2_X1 port map( A => A(32), B => B(32), Z => n600);
   U1 : BUF_X1 port map( A => A(24), Z => net273969);
   U2 : OAI21_X1 port map( B1 => n594, B2 => n655, A => B(18), ZN => n510);
   U3 : OR2_X2 port map( A1 => n637, A2 => n511, ZN => net279490);
   U4 : AND2_X1 port map( A1 => A(19), A2 => B(19), ZN => n511);
   U5 : INV_X1 port map( A => B(22), ZN => n547);
   U6 : BUF_X1 port map( A => n583, Z => n630);
   U7 : INV_X1 port map( A => B(40), ZN => n631);
   U8 : INV_X1 port map( A => B(42), ZN => n524);
   U9 : INV_X1 port map( A => B(44), ZN => n523);
   U10 : INV_X1 port map( A => B(20), ZN => net279512);
   U11 : BUF_X1 port map( A => A(15), Z => n658);
   U12 : AOI21_X1 port map( B1 => n527, B2 => n539, A => B(32), ZN => n512);
   U13 : CLKBUF_X1 port map( A => n601, Z => n541);
   U14 : OR2_X1 port map( A1 => n601, A2 => n542, ZN => n602);
   U15 : CLKBUF_X1 port map( A => A(45), Z => n667);
   U16 : CLKBUF_X1 port map( A => n607, Z => n690);
   U17 : BUF_X1 port map( A => n574, Z => n672);
   U18 : AOI22_X1 port map( A1 => n541, A2 => n544, B1 => n602, B2 => B(31), ZN
                           => n513);
   U19 : OAI21_X1 port map( B1 => n706, B2 => n615, A => n575, ZN => n514);
   U20 : CLKBUF_X1 port map( A => A(41), Z => n515);
   U21 : NOR2_X1 port map( A1 => n599, A2 => n535, ZN => n516);
   U22 : INV_X1 port map( A => n519, ZN => n517);
   U23 : BUF_X1 port map( A => n613, Z => net272305);
   U24 : OAI21_X1 port map( B1 => n665, B2 => n688, A => B(42), ZN => n518);
   U25 : AOI21_X1 port map( B1 => n690, B2 => n638, A => n701, ZN => n519);
   U26 : INV_X1 port map( A => n635, ZN => n520);
   U27 : CLKBUF_X1 port map( A => n580, Z => n558);
   U28 : AOI22_X1 port map( A1 => net271811, A2 => net270610, B1 => n626, B2 =>
                           B(23), ZN => n521);
   U29 : NAND2_X1 port map( A1 => n518, A2 => n679, ZN => n522);
   U30 : INV_X1 port map( A => net279488, ZN => n609);
   U31 : BUF_X1 port map( A => A(38), Z => n654);
   U32 : BUF_X1 port map( A => A(33), Z => net271478);
   U33 : XNOR2_X1 port map( A => A(44), B => n523, ZN => n531);
   U34 : XNOR2_X1 port map( A => A(42), B => n524, ZN => n612);
   U35 : NAND2_X1 port map( A1 => n541, A2 => n542, ZN => n525);
   U36 : NAND2_X1 port map( A1 => n602, A2 => B(31), ZN => n526);
   U37 : NAND2_X1 port map( A1 => n525, A2 => n526, ZN => n527);
   U38 : INV_X1 port map( A => B(19), ZN => n621);
   U39 : NOR2_X1 port map( A1 => n584, A2 => B(37), ZN => n528);
   U40 : NOR2_X1 port map( A1 => n630, A2 => n639, ZN => n529);
   U41 : NOR2_X1 port map( A1 => n528, A2 => n529, ZN => n530);
   U42 : XNOR2_X1 port map( A => n562, B => n531, ZN => SUM(44));
   U43 : INV_X1 port map( A => B(34), ZN => n668);
   U44 : INV_X1 port map( A => B(28), ZN => n603);
   U45 : INV_X1 port map( A => B(29), ZN => n633);
   U46 : XNOR2_X1 port map( A => A(16), B => B(16), ZN => n591);
   U47 : NOR2_X1 port map( A1 => n512, A2 => n535, ZN => n595);
   U48 : OR2_X1 port map( A1 => n595, A2 => net271478, ZN => net270458);
   U49 : XNOR2_X1 port map( A => n595, B => net270516, ZN => SUM(33));
   U50 : AOI21_X1 port map( B1 => n516, B2 => net271478, A => B(33), ZN => n596
                           );
   U51 : AND2_X1 port map( A1 => n533, A2 => n543, ZN => n535);
   U52 : INV_X1 port map( A => A(32), ZN => n533);
   U53 : INV_X1 port map( A => n533, ZN => n539);
   U54 : AOI21_X1 port map( B1 => n527, B2 => n539, A => B(32), ZN => n599);
   U55 : CLKBUF_X1 port map( A => A(31), Z => n542);
   U56 : CLKBUF_X1 port map( A => n542, Z => n544);
   U57 : AOI22_X1 port map( A1 => n541, A2 => n544, B1 => n602, B2 => B(31), ZN
                           => n543);
   U58 : XNOR2_X1 port map( A => n513, B => n600, ZN => SUM(32));
   U59 : XNOR2_X1 port map( A => A(31), B => B(31), ZN => n536);
   U60 : NOR2_X1 port map( A1 => n605, A2 => n537, ZN => n601);
   U61 : XNOR2_X1 port map( A => n601, B => n536, ZN => SUM(31));
   U62 : AND2_X1 port map( A1 => n519, A2 => n532, ZN => n537);
   U63 : INV_X1 port map( A => A(30), ZN => n532);
   U64 : INV_X1 port map( A => n532, ZN => n540);
   U65 : AOI21_X1 port map( B1 => n534, B2 => n540, A => B(30), ZN => n605);
   U66 : INV_X1 port map( A => n604, ZN => n534);
   U67 : XNOR2_X1 port map( A => n517, B => n538, ZN => SUM(30));
   U68 : XNOR2_X1 port map( A => A(30), B => B(30), ZN => n538);
   U69 : AOI21_X1 port map( B1 => net270885, B2 => net271806, A => n629, ZN => 
                           net271341);
   U70 : BUF_X1 port map( A => net271341, Z => net271811);
   U71 : XNOR2_X1 port map( A => net271625, B => net271341, ZN => SUM(23));
   U72 : OR2_X1 port map( A1 => net271341, A2 => A(23), ZN => n626);
   U73 : AOI21_X1 port map( B1 => A(22), B2 => n552, A => B(22), ZN => n629);
   U74 : NAND2_X1 port map( A1 => net279521, A2 => net279520, ZN => n552);
   U75 : INV_X1 port map( A => A(22), ZN => net271806);
   U76 : INV_X1 port map( A => net271806, ZN => net279549);
   U77 : AND2_X1 port map( A1 => net279521, A2 => net279520, ZN => net270885);
   U78 : XNOR2_X1 port map( A => net270885, B => n547, ZN => net279507);
   U79 : NAND2_X1 port map( A1 => n550, A2 => n549, ZN => net279520);
   U80 : AND2_X1 port map( A1 => net279503, A2 => net279504, ZN => n549);
   U81 : OAI21_X1 port map( B1 => net279488, B2 => n553, A => net279512, ZN => 
                           net279504);
   U82 : OAI21_X1 port map( B1 => n553, B2 => n606, A => net279512, ZN => n551)
                           ;
   U83 : INV_X1 port map( A => A(20), ZN => n553);
   U84 : XNOR2_X1 port map( A => net279500, B => net279512, ZN => net288445);
   U85 : BUF_X1 port map( A => A(21), Z => n550);
   U86 : INV_X1 port map( A => n550, ZN => net279539);
   U87 : NAND2_X1 port map( A1 => n548, A2 => B(21), ZN => net279521);
   U88 : NAND2_X1 port map( A1 => n545, A2 => n546, ZN => n548);
   U89 : INV_X1 port map( A => A(21), ZN => n546);
   U90 : NAND2_X1 port map( A1 => n551, A2 => net279503, ZN => n545);
   U91 : INV_X1 port map( A => A(20), ZN => net279500);
   U92 : XNOR2_X1 port map( A => n545, B => B(21), ZN => net279508);
   U93 : CLKBUF_X1 port map( A => A(25), Z => n564);
   U94 : NAND2_X1 port map( A1 => n560, A2 => n557, ZN => n632);
   U95 : NAND2_X1 port map( A1 => n667, A2 => n666, ZN => n557);
   U96 : CLKBUF_X1 port map( A => n580, Z => n671);
   U97 : INV_X1 port map( A => n562, ZN => n561);
   U98 : CLKBUF_X1 port map( A => A(25), Z => net273126);
   U99 : CLKBUF_X1 port map( A => A(28), Z => n567);
   U100 : BUF_X1 port map( A => A(26), Z => n585);
   U101 : OAI21_X1 port map( B1 => n662, B2 => n674, A => n510, ZN => n570);
   U102 : XNOR2_X1 port map( A => net271455, B => net272305, ZN => SUM(27));
   U103 : XNOR2_X1 port map( A => A(27), B => B(27), ZN => net271455);
   U104 : NOR2_X1 port map( A1 => n617, A2 => n576, ZN => n613);
   U105 : OAI21_X1 port map( B1 => n613, B2 => A(27), A => B(27), ZN => n614);
   U106 : AND2_X1 port map( A1 => n613, A2 => A(27), ZN => net270456);
   U107 : NOR2_X1 port map( A1 => n588, A2 => n585, ZN => n576);
   U108 : NAND2_X1 port map( A1 => n579, A2 => n620, ZN => n588);
   U109 : OAI21_X1 port map( B1 => n564, B2 => n619, A => B(25), ZN => n620);
   U110 : NAND2_X1 port map( A1 => net274244, A2 => n564, ZN => n579);
   U111 : OAI21_X1 port map( B1 => n619, B2 => net273126, A => B(25), ZN => 
                           net276125);
   U112 : AOI21_X1 port map( B1 => n582, B2 => n585, A => B(26), ZN => n617);
   U113 : NAND2_X1 port map( A1 => net276125, A2 => n579, ZN => n582);
   U114 : XNOR2_X1 port map( A => A(25), B => B(25), ZN => net271055);
   U115 : XNOR2_X1 port map( A => A(26), B => B(26), ZN => n573);
   U116 : XNOR2_X1 port map( A => n582, B => n573, ZN => SUM(26));
   U117 : AOI21_X1 port map( B1 => net264490, B2 => net271340, A => n623, ZN =>
                           net274244);
   U118 : BUF_X1 port map( A => n521, Z => net271340);
   U119 : AOI21_X1 port map( B1 => net264490, B2 => net271340, A => n623, ZN =>
                           net276011);
   U120 : AOI21_X1 port map( B1 => net264490, B2 => net271340, A => net274277, 
                           ZN => n619);
   U122 : INV_X1 port map( A => net273969, ZN => net264490);
   U123 : AOI21_X1 port map( B1 => net273969, B2 => net274177, A => B(24), ZN 
                           => net274277);
   U124 : AOI21_X1 port map( B1 => net273969, B2 => net274177, A => B(24), ZN 
                           => n623);
   U125 : INV_X1 port map( A => net273960, ZN => net274177);
   U126 : AOI22_X1 port map( A1 => net271811, A2 => net270610, B1 => n626, B2 
                           => B(23), ZN => net273960);
   U127 : CLKBUF_X1 port map( A => A(23), Z => net270610);
   U128 : XNOR2_X1 port map( A => A(24), B => B(24), ZN => net271728);
   U129 : XNOR2_X1 port map( A => A(23), B => B(23), ZN => net271625);
   U130 : INV_X1 port map( A => n521, ZN => net264500);
   U131 : XNOR2_X1 port map( A => n591, B => n520, ZN => SUM(16));
   U132 : XNOR2_X1 port map( A => n570, B => B(19), ZN => n618);
   U133 : BUF_X1 port map( A => A(18), Z => n594);
   U134 : XNOR2_X1 port map( A => n598, B => n610, ZN => SUM(28));
   U135 : XNOR2_X1 port map( A => A(28), B => n603, ZN => n598);
   U136 : NOR2_X1 port map( A1 => net264503, A2 => net270456, ZN => n610);
   U137 : AND2_X1 port map( A1 => n610, A2 => net264480, ZN => net270769);
   U138 : INV_X1 port map( A => n614, ZN => net264503);
   U139 : OR2_X1 port map( A1 => net264503, A2 => net270456, ZN => n597);
   U140 : INV_X1 port map( A => A(28), ZN => net264480);
   U141 : AOI21_X1 port map( B1 => n597, B2 => n567, A => B(28), ZN => n611);
   U142 : XNOR2_X1 port map( A => net288445, B => n609, ZN => SUM(20));
   U143 : NAND2_X1 port map( A1 => net279490, A2 => net279489, ZN => n606);
   U145 : NAND2_X1 port map( A1 => n606, A2 => net279500, ZN => net279503);
   U146 : NAND2_X1 port map( A1 => net279490, A2 => net279489, ZN => net279488)
                           ;
   U147 : NAND2_X1 port map( A1 => n616, A2 => n621, ZN => net279489);
   U148 : XNOR2_X1 port map( A => n612, B => n568, ZN => SUM(42));
   U149 : INV_X1 port map( A => n697, ZN => n615);
   U150 : INV_X1 port map( A => A(19), ZN => n616);
   U151 : INV_X1 port map( A => n616, ZN => n622);
   U152 : XNOR2_X1 port map( A => net279508, B => net279539, ZN => SUM(21));
   U153 : XNOR2_X1 port map( A => net279507, B => net279549, ZN => SUM(22));
   U154 : XNOR2_X1 port map( A => n618, B => n622, ZN => SUM(19));
   U155 : XNOR2_X1 port map( A => net271728, B => net264500, ZN => SUM(24));
   U156 : OR2_X2 port map( A1 => n566, A2 => n624, ZN => n562);
   U157 : NOR2_X1 port map( A1 => n565, A2 => A(43), ZN => n624);
   U158 : INV_X1 port map( A => n706, ZN => n625);
   U159 : OAI21_X1 port map( B1 => n634, B2 => n561, A => B(44), ZN => n627);
   U160 : XNOR2_X1 port map( A => n690, B => n628, ZN => SUM(29));
   U161 : XOR2_X1 port map( A => A(29), B => n633, Z => n628);
   U162 : BUF_X1 port map( A => n577, Z => n660);
   U163 : XNOR2_X1 port map( A => A(40), B => n631, ZN => n695);
   U164 : XNOR2_X1 port map( A => A(18), B => B(18), ZN => n648);
   U165 : XNOR2_X1 port map( A => n554, B => n555, ZN => SUM(47));
   U166 : INV_X1 port map( A => n704, ZN => n634);
   U167 : OAI22_X1 port map( A1 => n658, A2 => n683, B1 => n649, B2 => B(15), 
                           ZN => n635);
   U168 : OAI21_X1 port map( B1 => n675, B2 => n676, A => n700, ZN => n636);
   U169 : CLKBUF_X1 port map( A => A(29), Z => n638);
   U170 : CLKBUF_X1 port map( A => A(37), Z => n639);
   U171 : NOR2_X1 port map( A1 => n652, A2 => n640, ZN => n673);
   U172 : NOR2_X1 port map( A1 => A(14), A2 => B(14), ZN => n640);
   U173 : AND2_X1 port map( A1 => n702, A2 => n656, ZN => n642);
   U174 : AND2_X1 port map( A1 => n702, A2 => n656, ZN => n645);
   U175 : AND2_X1 port map( A1 => n702, A2 => n656, ZN => n655);
   U181 : XNOR2_X1 port map( A => n648, B => n645, ZN => SUM(18));
   U182 : CLKBUF_X1 port map( A => n643, Z => n651);
   U183 : INV_X1 port map( A => n642, ZN => n662);
   U184 : OR2_X1 port map( A1 => n643, A2 => A(17), ZN => n656);
   U185 : INV_X1 port map( A => n709, ZN => n657);
   U186 : CLKBUF_X1 port map( A => n589, Z => n676);
   U187 : AND2_X1 port map( A1 => n636, A2 => n708, ZN => n659);
   U188 : NOR2_X1 port map( A1 => n587, A2 => n659, ZN => n583);
   U189 : OAI21_X1 port map( B1 => n675, B2 => n676, A => n700, ZN => n586);
   U190 : OR2_X1 port map( A1 => n635, A2 => n710, ZN => n661);
   U191 : NAND2_X1 port map( A1 => n647, A2 => n661, ZN => n643);
   U192 : XNOR2_X1 port map( A => n558, B => n663, ZN => SUM(38));
   U193 : XOR2_X1 port map( A => A(38), B => B(38), Z => n663);
   U194 : INV_X1 port map( A => n708, ZN => n664);
   U195 : AND2_X1 port map( A1 => n696, A2 => n680, ZN => n665);
   U196 : NAND2_X1 port map( A1 => n627, A2 => n678, ZN => n666);
   U197 : XNOR2_X1 port map( A => A(34), B => n668, ZN => n689);
   U198 : XNOR2_X1 port map( A => n669, B => n666, ZN => SUM(45));
   U199 : XNOR2_X1 port map( A => A(45), B => B(45), ZN => n669);
   U200 : XNOR2_X1 port map( A => n522, B => n670, ZN => SUM(43));
   U201 : XNOR2_X1 port map( A => B(43), B => A(43), ZN => n670);
   U202 : OAI22_X1 port map( A1 => n639, A2 => n630, B1 => n584, B2 => B(37), 
                           ZN => n580);
   U203 : INV_X1 port map( A => n594, ZN => n674);
   U204 : CLKBUF_X1 port map( A => n686, Z => n675);
   U205 : BUF_X1 port map( A => A(35), Z => n686);
   U206 : XNOR2_X1 port map( A => n677, B => n651, ZN => SUM(17));
   U207 : XNOR2_X1 port map( A => A(17), B => B(17), ZN => n677);
   U208 : OR2_X1 port map( A1 => n562, A2 => n704, ZN => n678);
   U209 : NAND2_X1 port map( A1 => n563, A2 => n678, ZN => n559);
   U210 : OR2_X1 port map( A1 => n568, A2 => n705, ZN => n679);
   U211 : NAND2_X1 port map( A1 => n569, A2 => n679, ZN => n565);
   U212 : OR2_X1 port map( A1 => n571, A2 => n515, ZN => n680);
   U213 : NAND2_X1 port map( A1 => n696, A2 => n680, ZN => n568);
   U214 : XNOR2_X1 port map( A => n681, B => n632, ZN => SUM(46));
   U215 : XNOR2_X1 port map( A => B(46), B => A(46), ZN => n681);
   U216 : XNOR2_X1 port map( A => B(35), B => A(35), ZN => n687);
   U217 : CLKBUF_X1 port map( A => A(14), Z => n682);
   U218 : BUF_X1 port map( A => n673, Z => n683);
   U219 : AND2_X1 port map( A1 => net264508, A2 => net270458, ZN => n684);
   U220 : XNOR2_X1 port map( A => n636, B => n685, ZN => SUM(36));
   U221 : XOR2_X1 port map( A => A(36), B => B(36), Z => n685);
   U222 : XNOR2_X1 port map( A => net271055, B => net276011, ZN => SUM(25));
   U223 : XNOR2_X1 port map( A => n589, B => n687, ZN => SUM(35));
   U224 : INV_X1 port map( A => n705, ZN => n688);
   U225 : XNOR2_X1 port map( A => n592, B => n689, ZN => SUM(34));
   U226 : NOR2_X1 port map( A1 => n611, A2 => net270769, ZN => n607);
   U227 : XNOR2_X1 port map( A => n514, B => n691, ZN => SUM(41));
   U228 : XNOR2_X1 port map( A => A(41), B => B(41), ZN => n691);
   U229 : XNOR2_X1 port map( A => A(33), B => B(33), ZN => net270516);
   U230 : OR2_X1 port map( A1 => n592, A2 => n709, ZN => n692);
   U231 : NAND2_X1 port map( A1 => n593, A2 => n692, ZN => n589);
   U232 : NAND2_X1 port map( A1 => net264508, A2 => net270458, ZN => n592);
   U233 : XNOR2_X1 port map( A => n630, B => n693, ZN => SUM(37));
   U234 : XNOR2_X1 port map( A => A(37), B => B(37), ZN => n693);
   U235 : XNOR2_X1 port map( A => n660, B => n694, ZN => SUM(39));
   U236 : XNOR2_X1 port map( A => A(39), B => B(39), ZN => n694);
   U237 : INV_X1 port map( A => n644, ZN => n702);
   U238 : INV_X1 port map( A => A(34), ZN => n709);
   U239 : OAI22_X1 port map( A1 => n556, A2 => B(46), B1 => n632, B2 => A(46), 
                           ZN => n554);
   U240 : AND2_X1 port map( A1 => A(46), A2 => n632, ZN => n556);
   U241 : INV_X1 port map( A => n654, ZN => n707);
   U242 : INV_X1 port map( A => n590, ZN => n700);
   U243 : INV_X1 port map( A => n572, ZN => n696);
   U244 : INV_X1 port map( A => A(36), ZN => n708);
   U245 : XNOR2_X1 port map( A => n672, B => n695, ZN => SUM(40));
   U246 : AOI21_X1 port map( B1 => A(14), B2 => B(14), A => carry_14_port, ZN 
                           => n652);
   U247 : INV_X1 port map( A => A(44), ZN => n704);
   U248 : OAI21_X1 port map( B1 => n561, B2 => n634, A => B(44), ZN => n563);
   U249 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U250 : INV_X1 port map( A => A(40), ZN => n706);
   U251 : AOI21_X1 port map( B1 => n699, B2 => n664, A => B(36), ZN => n587);
   U252 : INV_X1 port map( A => n586, ZN => n699);
   U253 : INV_X1 port map( A => n596, ZN => net264508);
   U254 : OAI22_X1 port map( A1 => n658, A2 => n683, B1 => n649, B2 => B(15), 
                           ZN => n646);
   U255 : AND2_X1 port map( A1 => n673, A2 => A(15), ZN => n649);
   U256 : AOI21_X1 port map( B1 => n577, B2 => A(39), A => B(39), ZN => n578);
   U257 : INV_X1 port map( A => n574, ZN => n697);
   U258 : OAI21_X1 port map( B1 => n707, B2 => n671, A => n581, ZN => n577);
   U259 : AOI21_X1 port map( B1 => n690, B2 => n638, A => n701, ZN => n604);
   U260 : OAI21_X1 port map( B1 => n703, B2 => A(16), A => B(16), ZN => n647);
   U261 : INV_X1 port map( A => n646, ZN => n703);
   U262 : OAI21_X1 port map( B1 => n530, B2 => n654, A => B(38), ZN => n581);
   U263 : OAI21_X1 port map( B1 => n697, B2 => n625, A => B(40), ZN => n575);
   U264 : OAI21_X1 port map( B1 => n706, B2 => n615, A => n575, ZN => n571);
   U265 : OAI21_X1 port map( B1 => A(39), B2 => n660, A => n698, ZN => n574);
   U266 : INV_X1 port map( A => n578, ZN => n698);
   U267 : INV_X1 port map( A => A(42), ZN => n705);
   U268 : AOI21_X1 port map( B1 => n565, B2 => A(43), A => B(43), ZN => n566);
   U269 : OAI21_X1 port map( B1 => n665, B2 => n688, A => B(42), ZN => n569);
   U270 : OAI21_X1 port map( B1 => n674, B2 => n662, A => n641, ZN => n637);
   U271 : OAI21_X1 port map( B1 => n594, B2 => n655, A => B(18), ZN => n641);
   U272 : AOI21_X1 port map( B1 => A(17), B2 => n643, A => B(17), ZN => n644);
   U273 : OAI21_X1 port map( B1 => n684, B2 => n657, A => B(34), ZN => n593);
   U274 : INV_X1 port map( A => A(16), ZN => n710);
   U275 : OAI21_X1 port map( B1 => n559, B2 => n667, A => B(45), ZN => n560);
   U276 : AOI21_X1 port map( B1 => n571, B2 => n515, A => B(41), ZN => n572);
   U277 : AND2_X1 port map( A1 => n583, A2 => A(37), ZN => n584);
   U278 : AOI21_X1 port map( B1 => n589, B2 => n686, A => B(35), ZN => n590);
   U279 : INV_X1 port map( A => n608, ZN => n701);
   U280 : OAI21_X1 port map( B1 => n607, B2 => A(29), A => B(29), ZN => n608);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT46_DW01_add_0 is

   port( A, B : in std_logic_vector (45 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (45 downto 0);  CO : out std_logic);

end RCA_NBIT46_DW01_add_0;

architecture SYN_rpl of RCA_NBIT46_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_12_port, carry_11_port, carry_10_port, carry_9_port, 
      carry_8_port, carry_7_port, carry_6_port, carry_5_port, carry_4_port, 
      carry_3_port, carry_2_port, n1, n572, n574, n575, n577, n578, n580, n581,
      n583, n584, n586, n587, n589, n590, n592, n593, n595, n596, n598, n599, 
      n601, n602, n604, n605, n607, n608, n609, n610, n611, n613, n614, n615, 
      n616, n617, n619, n620, n623, n630, n631, n633, n635, n656, n658, n661, 
      n662, n663, n664, n667, n669, n670, n671, net264428, net264441, net264455
      , net271501, net272296, net273275, net273495, net274023, n659, n657, n655
      , n645, n643, n640, net279625, net279645, net287642, net273517, net273029
      , n653, n651, net282809, net276162, net271509, net271502, net271241, 
      net264429, n632, n629, n628, n626, n625, n622, net271346, net264451, n650
      , n647, n646, n644, net274026, net271508, net264454, net264453, n641, 
      n638, n637, n634, n525, n526, n527, n528, n529, n530, n531, n532, n533, 
      n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, 
      n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, 
      n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, 
      n570, n571, n573, n576, n579, n582, n585, n588, n591, n594, n597, n600, 
      n603, n606, n612, n618, n621, n624, n627, n636, n639, n642, n648, n649, 
      n652, n654, n660, n665, n666, n668, n672, n673, n674, n675, n676, n677, 
      n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, 
      n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, 
      n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, 
      n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, 
      n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, 
      n738, n739 : std_logic;

begin
   
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U180 : XOR2_X1 port map( A => B(13), B => n570, Z => n669);
   U181 : XOR2_X1 port map( A => n693, B => n671, Z => SUM(12));
   U182 : XOR2_X1 port map( A => carry_12_port, B => B(12), Z => n671);
   U183 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : BUF_X1 port map( A => n661, Z => n525);
   U2 : CLKBUF_X1 port map( A => A(24), Z => n526);
   U3 : AND2_X2 port map( A1 => n631, A2 => net264428, ZN => n541);
   U4 : AND2_X1 port map( A1 => n705, A2 => n584, ZN => n642);
   U5 : AND2_X1 port map( A1 => n624, A2 => n728, ZN => n535);
   U6 : INV_X1 port map( A => B(41), ZN => n711);
   U7 : OR2_X1 port map( A1 => n625, A2 => net264429, ZN => net271502);
   U8 : INV_X1 port map( A => B(35), ZN => n530);
   U9 : CLKBUF_X1 port map( A => A(35), Z => n527);
   U10 : BUF_X1 port map( A => n592, Z => n678);
   U11 : CLKBUF_X1 port map( A => A(17), Z => n528);
   U12 : OAI21_X1 port map( B1 => n721, B2 => n688, A => B(41), ZN => n529);
   U13 : XNOR2_X1 port map( A => A(35), B => n530, ZN => n690);
   U14 : CLKBUF_X1 port map( A => n704, Z => n531);
   U15 : AND2_X1 port map( A1 => n729, A2 => n680, ZN => n532);
   U16 : AND2_X1 port map( A1 => n729, A2 => n680, ZN => n648);
   U17 : CLKBUF_X1 port map( A => A(41), Z => n688);
   U18 : BUF_X1 port map( A => A(36), Z => n683);
   U19 : BUF_X1 port map( A => A(22), Z => n549);
   U20 : NAND2_X1 port map( A1 => n534, A2 => n540, ZN => n555);
   U21 : OR2_X1 port map( A1 => net273029, A2 => n653, ZN => n533);
   U22 : BUF_X1 port map( A => n618, Z => n687);
   U23 : NOR2_X1 port map( A1 => n653, A2 => net273029, ZN => n534);
   U24 : OR2_X1 port map( A1 => n561, A2 => net271509, ZN => n564);
   U25 : NOR2_X1 port map( A1 => n667, A2 => B(13), ZN => n536);
   U26 : NOR2_X1 port map( A1 => n704, A2 => n570, ZN => n537);
   U27 : NOR2_X1 port map( A1 => n537, A2 => n536, ZN => n538);
   U28 : BUF_X1 port map( A => A(13), Z => n570);
   U29 : INV_X1 port map( A => B(15), ZN => n700);
   U30 : INV_X1 port map( A => B(17), ZN => n582);
   U31 : XNOR2_X1 port map( A => B(43), B => A(43), ZN => n689);
   U32 : CLKBUF_X1 port map( A => n592, Z => n597);
   U33 : INV_X1 port map( A => B(19), ZN => n556);
   U34 : INV_X1 port map( A => B(42), ZN => n709);
   U35 : INV_X1 port map( A => B(21), ZN => n553);
   U36 : INV_X1 port map( A => B(23), ZN => n550);
   U37 : INV_X1 port map( A => B(27), ZN => n565);
   U38 : XNOR2_X1 port map( A => n572, B => n539, ZN => SUM(45));
   U39 : XOR2_X1 port map( A => B(45), B => A(45), Z => n539);
   U40 : NAND2_X1 port map( A1 => n650, A2 => n555, ZN => n646);
   U41 : NAND2_X1 port map( A1 => net273495, A2 => n656, ZN => net274023);
   U42 : BUF_X1 port map( A => A(19), Z => n540);
   U43 : BUF_X1 port map( A => n538, Z => n649);
   U44 : BUF_X1 port map( A => A(16), Z => n588);
   U45 : BUF_X1 port map( A => A(18), Z => n569);
   U46 : AND2_X1 port map( A1 => net264455, A2 => net271501, ZN => n542);
   U47 : XNOR2_X1 port map( A => n551, B => n544, ZN => SUM(24));
   U48 : XNOR2_X1 port map( A => A(24), B => B(24), ZN => n544);
   U49 : BUF_X1 port map( A => n634, Z => n551);
   U50 : OR2_X1 port map( A1 => n526, A2 => n634, ZN => net271501);
   U51 : AOI21_X1 port map( B1 => n634, B2 => n526, A => B(24), ZN => n635);
   U52 : NAND2_X1 port map( A1 => n638, A2 => n547, ZN => n634);
   U53 : OAI21_X1 port map( B1 => net264454, B2 => n546, A => B(23), ZN => n638
                           );
   U54 : INV_X1 port map( A => n543, ZN => n546);
   U55 : INV_X1 port map( A => A(23), ZN => n543);
   U56 : OR2_X1 port map( A1 => net274026, A2 => n543, ZN => n547);
   U57 : INV_X1 port map( A => n637, ZN => net264454);
   U58 : OAI21_X1 port map( B1 => net271508, B2 => n549, A => net264453, ZN => 
                           n637);
   U59 : INV_X1 port map( A => n641, ZN => net264453);
   U60 : OAI21_X1 port map( B1 => n549, B2 => net271508, A => net264453, ZN => 
                           net274026);
   U61 : AOI21_X1 port map( B1 => n640, B2 => A(22), A => B(22), ZN => n641);
   U62 : BUF_X1 port map( A => n640, Z => net271508);
   U63 : XNOR2_X1 port map( A => n545, B => net271508, ZN => SUM(22));
   U64 : XNOR2_X1 port map( A => A(23), B => n550, ZN => n548);
   U65 : XNOR2_X1 port map( A => A(22), B => B(22), ZN => n545);
   U66 : XNOR2_X1 port map( A => net274026, B => n548, ZN => SUM(23));
   U67 : AOI21_X1 port map( B1 => n559, B2 => n558, A => B(21), ZN => n644);
   U68 : NOR2_X1 port map( A1 => n644, A2 => n554, ZN => n640);
   U69 : INV_X1 port map( A => n552, ZN => n558);
   U70 : INV_X1 port map( A => A(21), ZN => n552);
   U71 : AND2_X1 port map( A1 => n643, A2 => n552, ZN => n554);
   U72 : AND2_X1 port map( A1 => net264451, A2 => n557, ZN => n559);
   U73 : INV_X1 port map( A => n647, ZN => net264451);
   U74 : NAND2_X1 port map( A1 => net264451, A2 => n557, ZN => n643);
   U75 : AOI21_X1 port map( B1 => n646, B2 => net271346, A => B(20), ZN => n647
                           );
   U76 : BUF_X1 port map( A => A(20), Z => net271346);
   U77 : OR2_X1 port map( A1 => net271346, A2 => n646, ZN => n557);
   U78 : XNOR2_X1 port map( A => A(21), B => n553, ZN => n645);
   U79 : OAI21_X1 port map( B1 => n534, B2 => n540, A => B(19), ZN => n650);
   U80 : OAI21_X1 port map( B1 => n540, B2 => n534, A => B(19), ZN => n560);
   U81 : XNOR2_X1 port map( A => A(20), B => B(20), ZN => net273517);
   U82 : NAND2_X1 port map( A1 => n555, A2 => n560, ZN => net287642);
   U83 : XNOR2_X1 port map( A => A(19), B => n556, ZN => n651);
   U84 : XNOR2_X1 port map( A => n562, B => n622, ZN => SUM(28));
   U85 : NAND2_X1 port map( A1 => net282809, A2 => net271502, ZN => n622);
   U86 : OAI21_X1 port map( B1 => n564, B2 => net271241, A => B(27), ZN => 
                           net282809);
   U87 : INV_X1 port map( A => net264429, ZN => net271241);
   U88 : OAI21_X1 port map( B1 => n564, B2 => net271241, A => B(27), ZN => n626
                           );
   U89 : INV_X1 port map( A => A(27), ZN => net264429);
   U90 : XNOR2_X1 port map( A => A(28), B => B(28), ZN => n562);
   U91 : NAND2_X1 port map( A1 => net271502, A2 => n626, ZN => net279645);
   U92 : INV_X1 port map( A => n629, ZN => n561);
   U93 : NOR2_X1 port map( A1 => net271509, A2 => n561, ZN => n625);
   U94 : OAI21_X1 port map( B1 => n628, B2 => net276162, A => B(26), ZN => n629
                           );
   U95 : BUF_X1 port map( A => A(26), Z => net276162);
   U96 : AND2_X1 port map( A1 => net279625, A2 => net276162, ZN => net271509);
   U97 : NOR2_X1 port map( A1 => n567, A2 => n541, ZN => n628);
   U98 : AOI21_X1 port map( B1 => net272296, B2 => n566, A => B(25), ZN => n567
                           );
   U99 : CLKBUF_X1 port map( A => A(25), Z => n566);
   U100 : AOI21_X1 port map( B1 => net272296, B2 => n566, A => B(25), ZN => 
                           n632);
   U101 : XNOR2_X1 port map( A => A(27), B => n565, ZN => n563);
   U102 : CLKBUF_X1 port map( A => A(28), Z => net273275);
   U103 : AOI21_X1 port map( B1 => net279645, B2 => net273275, A => B(28), ZN 
                           => n623);
   U104 : XNOR2_X1 port map( A => n625, B => n563, ZN => SUM(27));
   U105 : XNOR2_X1 port map( A => A(26), B => B(26), ZN => n630);
   U106 : NOR2_X1 port map( A1 => n632, A2 => n541, ZN => net279625);
   U107 : XNOR2_X1 port map( A => A(25), B => B(25), ZN => n633);
   U108 : INV_X1 port map( A => A(25), ZN => net264428);
   U109 : XNOR2_X1 port map( A => net273517, B => net287642, ZN => SUM(20));
   U110 : AOI21_X1 port map( B1 => net274023, B2 => n569, A => B(18), ZN => 
                           n653);
   U111 : NOR2_X1 port map( A1 => net274023, A2 => n569, ZN => net273029);
   U112 : XNOR2_X1 port map( A => n651, B => n533, ZN => SUM(19));
   U113 : XNOR2_X1 port map( A => net274023, B => n568, ZN => SUM(18));
   U114 : XNOR2_X1 port map( A => A(18), B => B(18), ZN => n568);
   U115 : BUF_X1 port map( A => A(34), Z => n639);
   U116 : CLKBUF_X1 port map( A => A(15), Z => n691);
   U117 : BUF_X1 port map( A => A(40), Z => n666);
   U118 : BUF_X1 port map( A => A(32), Z => n576);
   U119 : CLKBUF_X1 port map( A => A(42), Z => n571);
   U120 : OAI21_X1 port map( B1 => n701, B2 => n535, A => B(33), ZN => n573);
   U121 : XNOR2_X1 port map( A => n643, B => n645, ZN => SUM(21));
   U122 : XNOR2_X1 port map( A => n657, B => n655, ZN => SUM(17));
   U123 : XNOR2_X1 port map( A => A(17), B => n582, ZN => n657);
   U124 : NAND2_X1 port map( A1 => n579, A2 => n591, ZN => n655);
   U125 : OR2_X1 port map( A1 => n655, A2 => net264441, ZN => net273495);
   U126 : INV_X1 port map( A => n659, ZN => n579);
   U127 : AND2_X1 port map( A1 => n579, A2 => n591, ZN => n594);
   U128 : AOI21_X1 port map( B1 => n658, B2 => n588, A => B(16), ZN => n659);
   U129 : OR2_X1 port map( A1 => n588, A2 => n658, ZN => n591);
   U130 : INV_X1 port map( A => A(17), ZN => net264441);
   U131 : OAI21_X1 port map( B1 => n594, B2 => n528, A => B(17), ZN => n656);
   U132 : XNOR2_X1 port map( A => n658, B => n585, ZN => SUM(16));
   U133 : XNOR2_X1 port map( A => A(16), B => B(16), ZN => n585);
   U134 : CLKBUF_X1 port map( A => A(39), Z => n600);
   U135 : NAND2_X1 port map( A1 => n573, A2 => n697, ZN => n603);
   U136 : OAI21_X1 port map( B1 => n600, B2 => n723, A => B(39), ZN => n606);
   U137 : AOI22_X1 port map( A1 => n673, A2 => A(43), B1 => n578, B2 => B(43), 
                           ZN => n612);
   U138 : NAND2_X1 port map( A1 => n706, A2 => n606, ZN => n618);
   U139 : OAI21_X1 port map( B1 => n660, B2 => n597, A => n724, ZN => n621);
   U140 : OR2_X1 port map( A1 => n576, A2 => n684, ZN => n624);
   U141 : NAND2_X1 port map( A1 => n624, A2 => n728, ZN => n607);
   U142 : OR2_X1 port map( A1 => n619, A2 => n739, ZN => n627);
   U143 : NAND2_X1 port map( A1 => n620, A2 => n627, ZN => n616);
   U144 : NOR2_X1 port map( A1 => n682, A2 => n623, ZN => n636);
   U145 : OAI21_X1 port map( B1 => n679, B2 => n527, A => B(35), ZN => n602);
   U146 : OR2_X1 port map( A1 => n601, A2 => n736, ZN => n652);
   U147 : NAND2_X1 port map( A1 => n602, A2 => n652, ZN => n598);
   U148 : OR2_X1 port map( A1 => n661, A2 => n731, ZN => n654);
   U149 : NAND2_X1 port map( A1 => n662, A2 => n654, ZN => n658);
   U150 : XNOR2_X1 port map( A => n725, B => n719, ZN => SUM(37));
   U151 : CLKBUF_X1 port map( A => A(38), Z => n660);
   U152 : INV_X1 port map( A => n738, ZN => n665);
   U153 : BUF_X1 port map( A => n616, Z => n668);
   U154 : XNOR2_X1 port map( A => n672, B => n649, ZN => SUM(14));
   U155 : XNOR2_X1 port map( A => A(14), B => B(14), ZN => n672);
   U156 : CLKBUF_X1 port map( A => n577, Z => n673);
   U157 : OAI22_X1 port map( A1 => n698, A2 => n649, B1 => n664, B2 => B(14), 
                           ZN => n674);
   U158 : OAI21_X1 port map( B1 => n665, B2 => n532, A => B(31), ZN => n675);
   U159 : OAI21_X1 port map( B1 => n710, B2 => n687, A => n722, ZN => n676);
   U160 : INV_X1 port map( A => n739, ZN => n677);
   U161 : AND2_X1 port map( A1 => n696, A2 => n727, ZN => n679);
   U162 : OR2_X1 port map( A1 => A(30), A2 => n616, ZN => n680);
   U163 : NAND2_X1 port map( A1 => n729, A2 => n680, ZN => n613);
   U164 : NOR2_X1 port map( A1 => n670, A2 => n681, ZN => n686);
   U165 : NOR2_X1 port map( A1 => A(12), A2 => B(12), ZN => n681);
   U166 : OR2_X1 port map( A1 => n623, A2 => n682, ZN => n619);
   U167 : NOR2_X1 port map( A1 => net273275, A2 => net279645, ZN => n682);
   U168 : NAND2_X1 port map( A1 => n675, A2 => n695, ZN => n684);
   U169 : INV_X1 port map( A => n732, ZN => n685);
   U170 : XNOR2_X1 port map( A => n577, B => n689, ZN => SUM(43));
   U171 : AND2_X1 port map( A1 => net264455, A2 => net271501, ZN => net272296);
   U172 : XNOR2_X1 port map( A => n690, B => n601, ZN => SUM(35));
   U173 : XNOR2_X1 port map( A => A(36), B => B(36), ZN => n692);
   U174 : XNOR2_X1 port map( A => n692, B => n598, ZN => SUM(36));
   U175 : CLKBUF_X1 port map( A => A(12), Z => n693);
   U176 : AOI22_X1 port map( A1 => n673, A2 => A(43), B1 => n578, B2 => B(43), 
                           ZN => n575);
   U177 : OR2_X1 port map( A1 => n577, A2 => A(43), ZN => n578);
   U178 : NAND2_X1 port map( A1 => net264455, A2 => net271501, ZN => n631);
   U179 : OR2_X1 port map( A1 => n595, A2 => n732, ZN => n694);
   U184 : NAND2_X1 port map( A1 => n596, A2 => n694, ZN => n592);
   U185 : OR2_X1 port map( A1 => n613, A2 => n738, ZN => n695);
   U186 : NAND2_X1 port map( A1 => n695, A2 => n614, ZN => n610);
   U187 : OR2_X1 port map( A1 => n603, A2 => n639, ZN => n696);
   U188 : NAND2_X1 port map( A1 => n696, A2 => n727, ZN => n601);
   U189 : OR2_X1 port map( A1 => n607, A2 => n737, ZN => n697);
   U190 : NAND2_X1 port map( A1 => n608, A2 => n697, ZN => n604);
   U191 : OAI22_X1 port map( A1 => n698, A2 => n649, B1 => B(14), B2 => n664, 
                           ZN => n661);
   U192 : CLKBUF_X1 port map( A => A(14), Z => n698);
   U193 : INV_X1 port map( A => n531, ZN => n699);
   U194 : BUF_X1 port map( A => n686, Z => n704);
   U195 : XNOR2_X1 port map( A => A(15), B => n700, ZN => n663);
   U196 : INV_X1 port map( A => n737, ZN => n701);
   U197 : XNOR2_X1 port map( A => n702, B => n684, ZN => SUM(32));
   U198 : XNOR2_X1 port map( A => A(32), B => B(32), ZN => n702);
   U199 : XNOR2_X1 port map( A => n678, B => n703, ZN => SUM(38));
   U200 : XNOR2_X1 port map( A => A(38), B => B(38), ZN => n703);
   U201 : OR2_X1 port map( A1 => n734, A2 => n583, ZN => n705);
   U202 : NAND2_X1 port map( A1 => n529, A2 => n705, ZN => n581);
   U203 : OR2_X1 port map( A1 => n733, A2 => n621, ZN => n706);
   U204 : NAND2_X1 port map( A1 => n590, A2 => n706, ZN => n586);
   U205 : OR2_X1 port map( A1 => n683, A2 => n598, ZN => n707);
   U206 : NAND2_X1 port map( A1 => n707, A2 => n726, ZN => n595);
   U207 : XNOR2_X1 port map( A => n621, B => n708, ZN => SUM(39));
   U208 : XNOR2_X1 port map( A => B(39), B => n733, ZN => n708);
   U209 : XNOR2_X1 port map( A => n709, B => A(42), ZN => n717);
   U210 : CLKBUF_X1 port map( A => n666, Z => n710);
   U211 : XNOR2_X1 port map( A => A(41), B => n711, ZN => n715);
   U212 : XNOR2_X1 port map( A => n712, B => n668, ZN => SUM(30));
   U213 : XNOR2_X1 port map( A => A(30), B => B(30), ZN => n712);
   U214 : XNOR2_X1 port map( A => n603, B => n713, ZN => SUM(34));
   U215 : XNOR2_X1 port map( A => A(34), B => B(34), ZN => n713);
   U216 : XNOR2_X1 port map( A => n612, B => n714, ZN => SUM(44));
   U217 : XOR2_X1 port map( A => B(44), B => A(44), Z => n714);
   U218 : XNOR2_X1 port map( A => n715, B => n583, ZN => SUM(41));
   U219 : XNOR2_X1 port map( A => n636, B => n716, ZN => SUM(29));
   U220 : XNOR2_X1 port map( A => A(29), B => B(29), ZN => n716);
   U221 : XNOR2_X1 port map( A => n642, B => n717, ZN => SUM(42));
   U222 : INV_X1 port map( A => n571, ZN => n735);
   U223 : AND2_X1 port map( A1 => n720, A2 => A(44), ZN => n574);
   U224 : OAI22_X1 port map( A1 => n574, A2 => B(44), B1 => A(44), B2 => n720, 
                           ZN => n572);
   U225 : INV_X1 port map( A => A(39), ZN => n733);
   U226 : INV_X1 port map( A => n575, ZN => n720);
   U227 : INV_X1 port map( A => A(29), ZN => n739);
   U228 : OAI21_X1 port map( B1 => n636, B2 => n677, A => B(29), ZN => n620);
   U229 : AND2_X1 port map( A1 => n686, A2 => A(13), ZN => n667);
   U230 : AOI21_X1 port map( B1 => n642, B2 => n735, A => n580, ZN => n577);
   U231 : XNOR2_X1 port map( A => n618, B => n718, ZN => SUM(40));
   U232 : XNOR2_X1 port map( A => A(40), B => B(40), ZN => n718);
   U233 : OAI21_X1 port map( B1 => n660, B2 => n597, A => n724, ZN => n589);
   U234 : INV_X1 port map( A => n605, ZN => n727);
   U235 : XNOR2_X1 port map( A => B(37), B => A(37), ZN => n719);
   U236 : INV_X1 port map( A => A(33), ZN => n737);
   U237 : INV_X1 port map( A => A(37), ZN => n732);
   U238 : OAI21_X1 port map( B1 => n725, B2 => n685, A => B(37), ZN => n596);
   U239 : INV_X1 port map( A => n617, ZN => n729);
   U240 : XNOR2_X1 port map( A => n699, B => n669, ZN => SUM(13));
   U241 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U242 : AOI21_X1 port map( B1 => n604, B2 => n639, A => B(34), ZN => n605);
   U243 : INV_X1 port map( A => n599, ZN => n726);
   U244 : INV_X1 port map( A => A(15), ZN => n731);
   U245 : XNOR2_X1 port map( A => A(31), B => B(31), ZN => n615);
   U246 : INV_X1 port map( A => A(31), ZN => n738);
   U247 : INV_X1 port map( A => A(35), ZN => n736);
   U248 : AOI21_X1 port map( B1 => n592, B2 => A(38), A => B(38), ZN => n593);
   U249 : XNOR2_X1 port map( A => A(33), B => B(33), ZN => n609);
   U250 : INV_X1 port map( A => A(41), ZN => n734);
   U251 : XNOR2_X1 port map( A => net279625, B => n630, ZN => SUM(26));
   U252 : XNOR2_X1 port map( A => n615, B => n648, ZN => SUM(31));
   U253 : OAI21_X1 port map( B1 => n665, B2 => n532, A => B(31), ZN => n614);
   U254 : OAI21_X1 port map( B1 => n710, B2 => n687, A => n722, ZN => n583);
   U255 : AOI21_X1 port map( B1 => n581, B2 => n571, A => B(42), ZN => n580);
   U256 : INV_X1 port map( A => n587, ZN => n722);
   U257 : AOI21_X1 port map( B1 => n598, B2 => n683, A => B(36), ZN => n599);
   U258 : XNOR2_X1 port map( A => n542, B => n633, ZN => SUM(25));
   U259 : XNOR2_X1 port map( A => n535, B => n609, ZN => SUM(33));
   U260 : OAI21_X1 port map( B1 => n730, B2 => n691, A => B(15), ZN => n662);
   U261 : INV_X1 port map( A => n674, ZN => n730);
   U262 : XNOR2_X1 port map( A => n525, B => n663, ZN => SUM(15));
   U263 : AOI21_X1 port map( B1 => n586, B2 => n666, A => B(40), ZN => n587);
   U264 : OAI21_X1 port map( B1 => n721, B2 => n688, A => B(41), ZN => n584);
   U265 : OAI21_X1 port map( B1 => n723, B2 => n600, A => B(39), ZN => n590);
   U266 : INV_X1 port map( A => n593, ZN => n724);
   U267 : AOI21_X1 port map( B1 => n616, B2 => A(30), A => B(30), ZN => n617);
   U268 : INV_X1 port map( A => n676, ZN => n721);
   U269 : INV_X1 port map( A => n589, ZN => n723);
   U270 : INV_X1 port map( A => n595, ZN => n725);
   U271 : INV_X1 port map( A => n611, ZN => n728);
   U272 : INV_X1 port map( A => n635, ZN => net264455);
   U273 : OAI21_X1 port map( B1 => n701, B2 => n535, A => B(33), ZN => n608);
   U274 : AOI21_X1 port map( B1 => A(12), B2 => B(12), A => carry_12_port, ZN 
                           => n670);
   U275 : AOI21_X1 port map( B1 => n610, B2 => n576, A => B(32), ZN => n611);
   U276 : AND2_X1 port map( A1 => n538, A2 => A(14), ZN => n664);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT44_DW01_add_0 is

   port( A, B : in std_logic_vector (43 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (43 downto 0);  CO : out std_logic);

end RCA_NBIT44_DW01_add_0;

architecture SYN_rpl of RCA_NBIT44_DW01_add_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal n1, carry_9_port, carry_8_port, carry_7_port, carry_6_port, 
      carry_5_port, carry_4_port, carry_3_port, carry_2_port, carry_10_port, 
      carry_14_port, carry_13_port, n567, n568, n569, n570, n571, n572, n574, 
      n576, n577, n578, n584, n586, n587, n589, n590, n591, n592, n593, n595, 
      n596, n598, n599, n601, n602, n604, n605, n607, n608, n610, n611, n614, 
      n617, n627, n654, n657, n658, net264387, net264411, net269626, net270354,
      net270783, net271576, net272996, net273304, net273973, net274038, 
      net274148, net275938, net280436, net280411, net280410, net280405, 
      net270423, net274008, net274045, net272977, net272080, net271392, 
      net271381, net271018, n623, n620, n619, n616, net280491, n631, net273863,
      net269661, net273953, net273769, n644, n523, n524, n525, n526, n527, n528
      , n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
      n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, 
      n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, 
      n565, n566, n573, n575, n579, n580, n581, n582, n583, n585, n588, n594, 
      n597, n600, n603, n606, n609, n612, n613, n615, n618, n621, n622, n624, 
      n625, n626, n628, n629, n630, n632, n633, n634, n635, n636, n637, n638, 
      n639, n640, n641, n642, n643, n645, n646, n647, n648, n649, n650, n651, 
      n652, n653, n655, n656, n659, n660, n661, n662, n663, n664, n665, n666, 
      n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, 
      n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, 
      n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, 
      n703, n704, n705, n706, n707 : std_logic;

begin
   
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => n658, CO => 
                           carry_13_port, S => SUM(12));
   U116 : XOR2_X1 port map( A => B(43), B => A(43), Z => n570);
   U166 : XOR2_X1 port map( A => n568, B => n567, Z => SUM(11));
   U168 : XOR2_X1 port map( A => carry_10_port, B => n657, Z => SUM(10));
   U169 : XOR2_X1 port map( A => A(10), B => B(10), Z => n657);
   U170 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : INV_X1 port map( A => n703, ZN => n523);
   U2 : BUF_X1 port map( A => n610, Z => n524);
   U3 : OR2_X1 port map( A1 => B(20), A2 => n552, ZN => n544);
   U4 : INV_X1 port map( A => B(22), ZN => n579);
   U5 : INV_X1 port map( A => B(16), ZN => n633);
   U6 : INV_X1 port map( A => B(39), ZN => n538);
   U7 : INV_X1 port map( A => B(14), ZN => n630);
   U8 : INV_X1 port map( A => B(21), ZN => n550);
   U9 : AND2_X1 port map( A1 => n566, A2 => n573, ZN => net274008);
   U10 : INV_X1 port map( A => B(13), ZN => n530);
   U11 : INV_X1 port map( A => B(23), ZN => net280491);
   U12 : INV_X1 port map( A => B(36), ZN => n672);
   U13 : OR2_X1 port map( A1 => n677, A2 => n537, ZN => n652);
   U14 : OAI21_X1 port map( B1 => n588, B2 => n558, A => B(23), ZN => n525);
   U15 : OAI21_X1 port map( B1 => n557, B2 => net280410, A => net280411, ZN => 
                           n526);
   U16 : OAI21_X1 port map( B1 => n549, B2 => net272996, A => B(21), ZN => n527
                           );
   U17 : BUF_X1 port map( A => A(21), Z => net272996);
   U18 : AOI21_X1 port map( B1 => n600, B2 => n606, A => B(26), ZN => n528);
   U19 : BUF_X1 port map( A => n604, Z => n683);
   U20 : CLKBUF_X1 port map( A => n607, Z => n666);
   U21 : NOR2_X1 port map( A1 => n644, A2 => net273769, ZN => n529);
   U22 : XNOR2_X1 port map( A => A(13), B => n530, ZN => n531);
   U23 : XOR2_X1 port map( A => carry_13_port, B => n531, Z => SUM(13));
   U24 : NAND2_X1 port map( A1 => carry_13_port, A2 => A(13), ZN => n532);
   U25 : NAND2_X1 port map( A1 => carry_13_port, A2 => B(13), ZN => n533);
   U26 : NAND2_X1 port map( A1 => A(13), A2 => B(13), ZN => n534);
   U27 : NAND3_X1 port map( A1 => n532, A2 => n533, A3 => n534, ZN => 
                           carry_14_port);
   U28 : CLKBUF_X1 port map( A => A(19), Z => n535);
   U29 : BUF_X1 port map( A => n626, Z => n641);
   U30 : CLKBUF_X1 port map( A => n625, Z => n536);
   U31 : INV_X1 port map( A => B(15), ZN => net273304);
   U32 : BUF_X1 port map( A => A(25), Z => net272080);
   U33 : INV_X1 port map( A => B(41), ZN => n659);
   U34 : AND2_X1 port map( A1 => n621, A2 => n622, ZN => n612);
   U35 : AOI21_X1 port map( B1 => n539, B2 => n676, A => n538, ZN => n537);
   U36 : OR2_X1 port map( A1 => n584, A2 => n682, ZN => n539);
   U37 : INV_X1 port map( A => B(30), ZN => n648);
   U38 : OAI21_X1 port map( B1 => n549, B2 => net272996, A => B(21), ZN => n553
                           );
   U39 : NAND2_X1 port map( A1 => n544, A2 => n545, ZN => n543);
   U40 : XNOR2_X1 port map( A => n551, B => n543, ZN => SUM(21));
   U41 : NAND2_X1 port map( A1 => n548, A2 => n547, ZN => n545);
   U42 : AND2_X1 port map( A1 => n544, A2 => n545, ZN => n549);
   U43 : NAND2_X1 port map( A1 => n542, A2 => n541, ZN => n540);
   U44 : NAND2_X1 port map( A1 => n540, A2 => B(20), ZN => n548);
   U45 : XNOR2_X1 port map( A => n546, B => n552, ZN => SUM(20));
   U46 : XNOR2_X1 port map( A => A(21), B => n550, ZN => n551);
   U47 : NAND2_X1 port map( A1 => n535, A2 => n529, ZN => n541);
   U48 : OAI21_X1 port map( B1 => net273863, B2 => A(19), A => B(19), ZN => 
                           n542);
   U49 : XNOR2_X1 port map( A => A(19), B => B(19), ZN => net269661);
   U50 : XNOR2_X1 port map( A => A(20), B => B(20), ZN => n546);
   U51 : INV_X1 port map( A => A(20), ZN => n547);
   U52 : NAND2_X1 port map( A1 => n542, A2 => n541, ZN => n552);
   U53 : BUF_X1 port map( A => A(28), Z => n618);
   U54 : AOI21_X1 port map( B1 => n619, B2 => n597, A => n620, ZN => n554);
   U55 : AOI21_X1 port map( B1 => n619, B2 => n597, A => n528, ZN => n616);
   U56 : OAI21_X1 port map( B1 => n543, B2 => net264387, A => n527, ZN => n555)
                           ;
   U57 : AOI21_X1 port map( B1 => net273953, B2 => n556, A => B(18), ZN => n644
                           );
   U58 : NOR2_X1 port map( A1 => n644, A2 => net273769, ZN => net273863);
   U59 : BUF_X1 port map( A => A(18), Z => net273953);
   U60 : NOR2_X1 port map( A1 => net273953, A2 => n556, ZN => net273769);
   U61 : OAI21_X1 port map( B1 => n557, B2 => net280410, A => net280411, ZN => 
                           n556);
   U62 : CLKBUF_X1 port map( A => net280405, Z => n557);
   U63 : XNOR2_X1 port map( A => A(18), B => B(18), ZN => net270783);
   U64 : XNOR2_X1 port map( A => net280405, B => B(17), ZN => net280436);
   U65 : XNOR2_X1 port map( A => net269661, B => n529, ZN => SUM(19));
   U66 : AND2_X1 port map( A1 => n561, A2 => n560, ZN => n558);
   U67 : NAND2_X1 port map( A1 => n581, A2 => n588, ZN => n564);
   U68 : CLKBUF_X1 port map( A => A(40), Z => n559);
   U69 : INV_X1 port map( A => A(22), ZN => n563);
   U70 : NAND2_X1 port map( A1 => n580, A2 => n579, ZN => n561);
   U71 : NAND2_X1 port map( A1 => n562, A2 => n563, ZN => n560);
   U72 : NAND2_X1 port map( A1 => n631, A2 => A(22), ZN => n580);
   U73 : XNOR2_X1 port map( A => net269626, B => n555, ZN => SUM(22));
   U74 : INV_X1 port map( A => n631, ZN => n562);
   U75 : OAI21_X1 port map( B1 => n588, B2 => n558, A => B(23), ZN => n565);
   U76 : INV_X1 port map( A => net273973, ZN => n581);
   U77 : NAND2_X1 port map( A1 => n583, A2 => n594, ZN => n573);
   U78 : OAI21_X1 port map( B1 => net275938, B2 => n594, A => n575, ZN => n566)
                           ;
   U79 : OAI21_X1 port map( B1 => n594, B2 => n583, A => n575, ZN => n582);
   U80 : INV_X1 port map( A => B(24), ZN => n575);
   U81 : XNOR2_X1 port map( A => A(24), B => n575, ZN => n627);
   U82 : AND2_X1 port map( A1 => n525, A2 => n564, ZN => net275938);
   U83 : AND2_X1 port map( A1 => n565, A2 => n564, ZN => n583);
   U84 : AND2_X1 port map( A1 => n582, A2 => n573, ZN => n585);
   U85 : XNOR2_X1 port map( A => net270423, B => n585, ZN => SUM(25));
   U86 : CLKBUF_X1 port map( A => A(23), Z => n588);
   U87 : NAND2_X1 port map( A1 => net274008, A2 => net272080, ZN => net271018);
   U88 : INV_X1 port map( A => A(24), ZN => n594);
   U89 : NAND2_X1 port map( A1 => n561, A2 => n560, ZN => net273973);
   U90 : XNOR2_X1 port map( A => A(23), B => net280491, ZN => net274148);
   U91 : OAI21_X1 port map( B1 => n543, B2 => net264387, A => n553, ZN => n631)
                           ;
   U92 : XNOR2_X1 port map( A => net272977, B => n603, ZN => SUM(27));
   U93 : XNOR2_X1 port map( A => A(27), B => B(27), ZN => n603);
   U94 : BUF_X1 port map( A => n554, Z => net272977);
   U95 : OAI21_X1 port map( B1 => n616, B2 => A(27), A => B(27), ZN => n617);
   U96 : AND2_X1 port map( A1 => n554, A2 => A(27), ZN => net270354);
   U97 : AOI21_X1 port map( B1 => n600, B2 => n606, A => B(26), ZN => n620);
   U98 : BUF_X1 port map( A => A(26), Z => n606);
   U99 : NAND2_X1 port map( A1 => net271018, A2 => n623, ZN => n600);
   U100 : OAI21_X1 port map( B1 => net272080, B2 => net274008, A => B(25), ZN 
                           => n623);
   U101 : OAI21_X1 port map( B1 => net272080, B2 => net274008, A => B(25), ZN 
                           => net274045);
   U102 : INV_X1 port map( A => A(26), ZN => n597);
   U103 : INV_X1 port map( A => net271392, ZN => n619);
   U104 : XNOR2_X1 port map( A => A(26), B => B(26), ZN => net271381);
   U105 : NAND2_X1 port map( A1 => net271018, A2 => net274045, ZN => net271392)
                           ;
   U106 : XNOR2_X1 port map( A => A(25), B => B(25), ZN => net270423);
   U107 : XNOR2_X1 port map( A => net271392, B => net271381, ZN => SUM(26));
   U108 : BUF_X1 port map( A => A(15), Z => n609);
   U109 : INV_X1 port map( A => carry_14_port, ZN => n636);
   U110 : BUF_X1 port map( A => A(33), Z => n655);
   U111 : XNOR2_X1 port map( A => n613, B => n685, ZN => SUM(38));
   U112 : NOR2_X1 port map( A1 => n674, A2 => n693, ZN => n613);
   U113 : OR2_X1 port map( A1 => n674, A2 => n693, ZN => n615);
   U114 : OR2_X1 port map( A1 => n674, A2 => n693, ZN => n667);
   U115 : XNOR2_X1 port map( A => net271576, B => n639, ZN => SUM(14));
   U117 : INV_X1 port map( A => A(14), ZN => n632);
   U118 : INV_X1 port map( A => n632, ZN => n639);
   U119 : NAND2_X1 port map( A1 => A(14), A2 => B(14), ZN => n638);
   U120 : OAI21_X1 port map( B1 => n612, B2 => n609, A => B(15), ZN => n626);
   U121 : NAND2_X1 port map( A1 => n641, A2 => n536, ZN => n624);
   U122 : NAND2_X1 port map( A1 => n612, A2 => n609, ZN => n625);
   U123 : NAND2_X1 port map( A1 => A(17), A2 => B(17), ZN => net280411);
   U124 : NOR2_X1 port map( A1 => A(17), A2 => B(17), ZN => net280410);
   U125 : INV_X1 port map( A => A(17), ZN => n634);
   U126 : XNOR2_X1 port map( A => net280436, B => n634, ZN => SUM(17));
   U127 : NAND2_X1 port map( A1 => n629, A2 => n628, ZN => net280405);
   U128 : XNOR2_X1 port map( A => net270783, B => n526, ZN => SUM(18));
   U129 : OAI21_X1 port map( B1 => n640, B2 => n633, A => n637, ZN => n629);
   U130 : XNOR2_X1 port map( A => n635, B => n624, ZN => SUM(16));
   U131 : AND2_X1 port map( A1 => n626, A2 => n625, ZN => n640);
   U132 : NAND2_X1 port map( A1 => n640, A2 => n633, ZN => n628);
   U133 : NAND2_X1 port map( A1 => n630, A2 => n632, ZN => n621);
   U134 : NAND2_X1 port map( A1 => n638, A2 => n636, ZN => n622);
   U135 : NAND2_X1 port map( A1 => n621, A2 => n622, ZN => net274038);
   U136 : XNOR2_X1 port map( A => A(16), B => B(16), ZN => n635);
   U137 : INV_X1 port map( A => A(16), ZN => n637);
   U138 : XNOR2_X1 port map( A => A(29), B => B(29), ZN => n642);
   U139 : XNOR2_X1 port map( A => n666, B => n680, ZN => SUM(30));
   U140 : XNOR2_X1 port map( A => n656, B => n576, ZN => SUM(41));
   U141 : OR2_X1 port map( A1 => n593, A2 => n649, ZN => n589);
   U142 : XNOR2_X1 port map( A => n524, B => n642, ZN => SUM(29));
   U143 : NOR2_X1 port map( A1 => n649, A2 => n593, ZN => n643);
   U144 : XNOR2_X1 port map( A => n651, B => n645, ZN => SUM(34));
   U145 : XOR2_X1 port map( A => A(34), B => B(34), Z => n645);
   U146 : NOR2_X1 port map( A1 => n646, A2 => net270354, ZN => n660);
   U147 : OR2_X1 port map( A1 => A(28), A2 => net264411, ZN => n646);
   U148 : BUF_X1 port map( A => A(32), Z => n678);
   U149 : NOR2_X1 port map( A1 => n673, A2 => n590, ZN => n647);
   U150 : BUF_X1 port map( A => n598, Z => n664);
   U151 : BUF_X1 port map( A => n601, Z => n665);
   U152 : XNOR2_X1 port map( A => A(30), B => n648, ZN => n680);
   U153 : NOR2_X1 port map( A1 => n592, A2 => n687, ZN => n649);
   U154 : XNOR2_X1 port map( A => n665, B => n650, ZN => SUM(32));
   U155 : XOR2_X1 port map( A => A(32), B => B(32), Z => n650);
   U156 : AOI21_X1 port map( B1 => n664, B2 => n655, A => n695, ZN => n651);
   U157 : XNOR2_X1 port map( A => n569, B => n570, ZN => SUM(43));
   U158 : XNOR2_X1 port map( A => net273973, B => net274148, ZN => SUM(23));
   U159 : NOR2_X1 port map( A1 => n584, A2 => n682, ZN => n653);
   U160 : AOI21_X1 port map( B1 => n700, B2 => n577, A => n578, ZN => n656);
   U161 : XNOR2_X1 port map( A => n699, B => n659, ZN => n576);
   U162 : NOR2_X1 port map( A1 => n614, A2 => n660, ZN => n610);
   U163 : XNOR2_X1 port map( A => A(33), B => B(33), ZN => n668);
   U164 : XNOR2_X1 port map( A => n661, B => n683, ZN => SUM(31));
   U165 : XNOR2_X1 port map( A => A(31), B => B(31), ZN => n661);
   U167 : CLKBUF_X1 port map( A => A(11), Z => n679);
   U171 : OR2_X1 port map( A1 => net264411, A2 => net270354, ZN => n662);
   U172 : OR2_X1 port map( A1 => net264411, A2 => net270354, ZN => n684);
   U173 : XNOR2_X1 port map( A => A(15), B => net273304, ZN => n654);
   U174 : AND2_X1 port map( A1 => n651, A2 => n703, ZN => n663);
   U175 : NOR2_X1 port map( A1 => n596, A2 => n663, ZN => n592);
   U176 : XNOR2_X1 port map( A => n664, B => n668, ZN => SUM(33));
   U177 : XNOR2_X1 port map( A => A(28), B => B(28), ZN => n675);
   U178 : BUF_X1 port map( A => A(35), Z => n687);
   U179 : AND2_X1 port map( A1 => n698, A2 => n670, ZN => n669);
   U180 : OR2_X1 port map( A1 => A(29), A2 => n610, ZN => n670);
   U181 : NAND2_X1 port map( A1 => n698, A2 => n670, ZN => n607);
   U182 : XNOR2_X1 port map( A => n592, B => n671, ZN => SUM(35));
   U183 : XNOR2_X1 port map( A => B(35), B => A(35), ZN => n671);
   U184 : XNOR2_X1 port map( A => A(36), B => n672, ZN => n591);
   U185 : AND2_X1 port map( A1 => n702, A2 => n589, ZN => n673);
   U186 : NOR2_X1 port map( A1 => n590, A2 => n673, ZN => n586);
   U187 : AND2_X1 port map( A1 => n647, A2 => A(37), ZN => n674);
   U188 : XNOR2_X1 port map( A => n675, B => n662, ZN => SUM(28));
   U189 : NOR2_X1 port map( A1 => n539, A2 => n676, ZN => n677);
   U190 : NOR2_X1 port map( A1 => n677, A2 => n537, ZN => n577);
   U191 : INV_X1 port map( A => A(39), ZN => n676);
   U192 : NOR2_X1 port map( A1 => n615, A2 => A(38), ZN => n682);
   U193 : INV_X1 port map( A => n701, ZN => n681);
   U194 : XNOR2_X1 port map( A => carry_14_port, B => B(14), ZN => net271576);
   U195 : XNOR2_X1 port map( A => n654, B => net274038, ZN => SUM(15));
   U196 : XNOR2_X1 port map( A => net275938, B => n627, ZN => SUM(24));
   U197 : XNOR2_X1 port map( A => n591, B => n589, ZN => SUM(36));
   U198 : XNOR2_X1 port map( A => n701, B => B(38), ZN => n685);
   U199 : XNOR2_X1 port map( A => n647, B => n686, ZN => SUM(37));
   U200 : XNOR2_X1 port map( A => A(37), B => B(37), ZN => n686);
   U201 : XNOR2_X1 port map( A => A(11), B => B(11), ZN => n568);
   U202 : OAI21_X1 port map( B1 => n692, B2 => n699, A => n574, ZN => n572);
   U203 : XNOR2_X1 port map( A => n577, B => n688, ZN => SUM(40));
   U204 : XNOR2_X1 port map( A => B(40), B => n700, ZN => n688);
   U205 : OR2_X1 port map( A1 => n607, A2 => n705, ZN => n689);
   U206 : NAND2_X1 port map( A1 => n608, A2 => n689, ZN => n604);
   U207 : XNOR2_X1 port map( A => n653, B => n690, ZN => SUM(39));
   U208 : XNOR2_X1 port map( A => A(39), B => B(39), ZN => n690);
   U209 : INV_X1 port map( A => A(41), ZN => n699);
   U210 : INV_X1 port map( A => A(40), ZN => n700);
   U211 : XNOR2_X1 port map( A => n572, B => n691, ZN => SUM(42));
   U212 : XNOR2_X1 port map( A => B(42), B => A(42), ZN => n691);
   U213 : OAI22_X1 port map( A1 => n571, A2 => B(42), B1 => n572, B2 => A(42), 
                           ZN => n569);
   U214 : AND2_X1 port map( A1 => A(42), A2 => n572, ZN => n571);
   U215 : INV_X1 port map( A => A(36), ZN => n702);
   U216 : INV_X1 port map( A => A(34), ZN => n703);
   U217 : OAI21_X1 port map( B1 => n656, B2 => A(41), A => B(41), ZN => n574);
   U218 : XNOR2_X1 port map( A => A(22), B => B(22), ZN => net269626);
   U219 : AOI22_X1 port map( A1 => B(10), A2 => A(10), B1 => n657, B2 => 
                           carry_10_port, ZN => n567);
   U220 : INV_X1 port map( A => A(38), ZN => n701);
   U221 : INV_X1 port map( A => A(30), ZN => n705);
   U222 : INV_X1 port map( A => B(11), ZN => n707);
   U223 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U224 : INV_X1 port map( A => n656, ZN => n692);
   U225 : AOI21_X1 port map( B1 => n652, B2 => n559, A => B(40), ZN => n578);
   U226 : OAI21_X1 port map( B1 => n669, B2 => A(30), A => B(30), ZN => n608);
   U227 : AOI21_X1 port map( B1 => n684, B2 => n618, A => B(28), ZN => n614);
   U228 : OAI21_X1 port map( B1 => n586, B2 => A(37), A => B(37), ZN => n587);
   U229 : INV_X1 port map( A => n678, ZN => n704);
   U230 : INV_X1 port map( A => n605, ZN => n697);
   U231 : AOI21_X1 port map( B1 => n664, B2 => n655, A => n695, ZN => n595);
   U232 : INV_X1 port map( A => n599, ZN => n695);
   U233 : AOI21_X1 port map( B1 => n592, B2 => n687, A => B(35), ZN => n593);
   U234 : INV_X1 port map( A => n679, ZN => n706);
   U235 : INV_X1 port map( A => n595, ZN => n694);
   U236 : OAI21_X1 port map( B1 => n683, B2 => A(31), A => n697, ZN => n601);
   U237 : AOI21_X1 port map( B1 => n604, B2 => A(31), A => B(31), ZN => n605);
   U238 : INV_X1 port map( A => n611, ZN => n698);
   U239 : OAI21_X1 port map( B1 => n696, B2 => n678, A => B(32), ZN => n602);
   U240 : INV_X1 port map( A => net272996, ZN => net264387);
   U241 : AOI21_X1 port map( B1 => n694, B2 => n523, A => B(34), ZN => n596);
   U242 : AOI21_X1 port map( B1 => n643, B2 => A(36), A => B(36), ZN => n590);
   U243 : AOI21_X1 port map( B1 => n667, B2 => n681, A => B(38), ZN => n584);
   U244 : INV_X1 port map( A => n587, ZN => n693);
   U245 : OAI22_X1 port map( A1 => n707, A2 => n706, B1 => n568, B2 => n567, ZN
                           => n658);
   U246 : OAI21_X1 port map( B1 => n598, B2 => A(33), A => B(33), ZN => n599);
   U247 : OAI21_X1 port map( B1 => n665, B2 => n704, A => n602, ZN => n598);
   U248 : INV_X1 port map( A => n601, ZN => n696);
   U249 : AOI21_X1 port map( B1 => n610, B2 => A(29), A => B(29), ZN => n611);
   U250 : INV_X1 port map( A => n617, ZN => net264411);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT42_DW01_add_0 is

   port( A, B : in std_logic_vector (41 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (41 downto 0);  CO : out std_logic);

end RCA_NBIT42_DW01_add_0;

architecture SYN_rpl of RCA_NBIT42_DW01_add_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_39_port, carry_38_port, carry_37_port, carry_36_port, 
      carry_35_port, carry_32_port, carry_31_port, carry_30_port, carry_29_port
      , carry_28_port, carry_23_port, n430, n432, n436, n437, n438, n439, n440,
      n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, 
      n453, n454, n455, n456, n458, n460, n461, n462, n464, n465, n470, n471, 
      n485, n486, n487, n500, n501, n502, n503, n504, n505, n506, n507, n508, 
      n509, net264371, net264374, net270977, net271166, net271263, net271313, 
      net271387, net271611, net272691, net272728, net273128, net273759, 
      net274170, net275426, net276108, net276120, net273947, net272692, 
      net287657, net273047, net271701, net264369, net264348, n473, net293635, 
      net271383, n483, n482, n480, n477, n476, net274012, net271395, n469, n389
      , n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
      n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, 
      n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, 
      n426, n427, n428, n429, n431, n433, n434, n435, n457, n459, n463, n466, 
      n467, n468, n472, n474, n475, n478, n479, n481, n484, n488, n489, n490, 
      n491, n492, n493, n494, n495, n496, n497, n498, n499, n510, n511, n512, 
      n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, 
      n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, 
      n537, n538, n539, n540, n541 : std_logic;

begin
   
   U1_38 : FA_X1 port map( A => A(38), B => B(38), CI => carry_38_port, CO => 
                           carry_39_port, S => SUM(38));
   U1_37 : FA_X1 port map( A => A(37), B => B(37), CI => carry_37_port, CO => 
                           carry_38_port, S => SUM(37));
   U1_36 : FA_X1 port map( A => A(36), B => B(36), CI => carry_36_port, CO => 
                           carry_37_port, S => SUM(36));
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => carry_35_port, CO => 
                           carry_36_port, S => SUM(35));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => net264374, CO => 
                           carry_28_port, S => SUM(27));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U117 : XOR2_X1 port map( A => n515, B => n439, Z => SUM(9));
   U118 : XOR2_X1 port map( A => B(9), B => n510, Z => n439);
   U119 : XOR2_X1 port map( A => n442, B => n443, Z => SUM(7));
   U120 : XOR2_X1 port map( A => B(7), B => A(7), Z => n443);
   U121 : XOR2_X1 port map( A => n529, B => n444, Z => SUM(6));
   U122 : XOR2_X1 port map( A => B(6), B => A(6), Z => n444);
   U123 : XOR2_X1 port map( A => B(41), B => A(41), Z => n450);
   U124 : XOR2_X1 port map( A => B(40), B => A(40), Z => n453);
   U125 : XOR2_X1 port map( A => n455, B => n456, Z => SUM(3));
   U126 : XOR2_X1 port map( A => B(3), B => A(3), Z => n456);
   U130 : XOR2_X1 port map( A => A(34), B => B(34), Z => n458);
   U141 : XOR2_X1 port map( A => n470, B => n471, Z => SUM(1));
   U142 : XOR2_X1 port map( A => B(1), B => A(1), Z => n471);
   U152 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : INV_X1 port map( A => B(14), ZN => n414);
   U2 : NAND2_X1 port map( A1 => n431, A2 => n429, ZN => n425);
   U3 : INV_X1 port map( A => B(21), ZN => n413);
   U4 : INV_X1 port map( A => B(11), ZN => n475);
   U5 : INV_X1 port map( A => B(12), ZN => n491);
   U6 : INV_X1 port map( A => B(24), ZN => n433);
   U7 : INV_X1 port map( A => B(26), ZN => n416);
   U8 : INV_X1 port map( A => B(16), ZN => n407);
   U9 : BUF_X1 port map( A => A(21), Z => n412);
   U10 : BUF_X1 port map( A => A(18), Z => net271701);
   U11 : CLKBUF_X1 port map( A => A(16), Z => n389);
   U12 : NAND2_X1 port map( A1 => n421, A2 => n422, ZN => n390);
   U13 : INV_X1 port map( A => n393, ZN => n394);
   U14 : AND2_X1 port map( A1 => n492, A2 => n392, ZN => n391);
   U15 : OR2_X1 port map( A1 => n479, A2 => A(12), ZN => n392);
   U16 : XNOR2_X1 port map( A => n488, B => n484, ZN => SUM(12));
   U17 : OR2_X1 port map( A1 => n430, A2 => n413, ZN => n518);
   U18 : NAND2_X1 port map( A1 => n392, A2 => n492, ZN => n468);
   U19 : INV_X1 port map( A => B(19), ZN => n399);
   U20 : AND2_X1 port map( A1 => n395, A2 => n525, ZN => n393);
   U21 : OR2_X1 port map( A1 => B(32), A2 => A(32), ZN => n395);
   U22 : INV_X1 port map( A => B(33), ZN => n516);
   U23 : BUF_X1 port map( A => n397, Z => n398);
   U24 : XNOR2_X1 port map( A => n420, B => B(25), ZN => n426);
   U25 : XNOR2_X1 port map( A => n397, B => n396, ZN => SUM(20));
   U26 : XNOR2_X1 port map( A => A(20), B => B(20), ZN => n396);
   U27 : NAND2_X1 port map( A1 => net270977, A2 => n469, ZN => n397);
   U28 : OAI21_X1 port map( B1 => net273047, B2 => net271395, A => B(19), ZN =>
                           n469);
   U29 : BUF_X1 port map( A => A(19), Z => net271395);
   U30 : INV_X1 port map( A => net271395, ZN => net264348);
   U31 : OAI21_X1 port map( B1 => net273047, B2 => net271395, A => B(19), ZN =>
                           net274012);
   U32 : INV_X1 port map( A => A(20), ZN => net273759);
   U33 : AOI22_X1 port map( A1 => n398, A2 => net276108, B1 => n432, B2 => 
                           B(20), ZN => net287657);
   U34 : AOI22_X1 port map( A1 => n398, A2 => net276108, B1 => n432, B2 => 
                           B(20), ZN => n430);
   U35 : AND2_X1 port map( A1 => net274012, A2 => net270977, ZN => net274170);
   U36 : XNOR2_X1 port map( A => A(19), B => n399, ZN => net273947);
   U37 : INV_X1 port map( A => n427, ZN => net273128);
   U38 : OR2_X1 port map( A1 => n403, A2 => n404, ZN => n400);
   U39 : XNOR2_X1 port map( A => net271383, B => n410, ZN => SUM(18));
   U40 : OR2_X1 port map( A1 => n403, A2 => n404, ZN => n410);
   U41 : INV_X1 port map( A => n477, ZN => n403);
   U42 : OAI21_X1 port map( B1 => n476, B2 => A(17), A => B(17), ZN => n477);
   U43 : XNOR2_X1 port map( A => A(18), B => B(18), ZN => net271383);
   U44 : AND2_X1 port map( A1 => n476, A2 => A(17), ZN => n404);
   U45 : NOR2_X1 port map( A1 => n480, A2 => n406, ZN => n476);
   U46 : CLKBUF_X1 port map( A => n476, Z => net272691);
   U47 : AND2_X1 port map( A1 => n401, A2 => n408, ZN => n406);
   U48 : INV_X1 port map( A => A(16), ZN => n401);
   U49 : AOI21_X1 port map( B1 => n409, B2 => n389, A => B(16), ZN => n480);
   U50 : OR2_X1 port map( A1 => n402, A2 => net271387, ZN => n409);
   U51 : INV_X1 port map( A => n483, ZN => n402);
   U52 : NOR2_X1 port map( A1 => n402, A2 => net271387, ZN => n408);
   U53 : OAI21_X1 port map( B1 => n482, B2 => A(15), A => B(15), ZN => n483);
   U54 : NOR2_X1 port map( A1 => n486, A2 => net271611, ZN => n482);
   U55 : XNOR2_X1 port map( A => A(17), B => B(17), ZN => net271313);
   U56 : AOI21_X1 port map( B1 => n400, B2 => net271701, A => B(18), ZN => n473
                           );
   U57 : XNOR2_X1 port map( A => n405, B => n408, ZN => SUM(16));
   U58 : XNOR2_X1 port map( A => A(16), B => n407, ZN => n405);
   U59 : XNOR2_X1 port map( A => A(15), B => B(15), ZN => net271166);
   U60 : NOR2_X1 port map( A1 => net271611, A2 => n486, ZN => net293635);
   U61 : INV_X1 port map( A => n473, ZN => net264369);
   U62 : AND2_X1 port map( A1 => net264369, A2 => n411, ZN => net273047);
   U63 : NAND2_X1 port map( A1 => net264369, A2 => n411, ZN => net272692);
   U64 : OR2_X1 port map( A1 => n410, A2 => net271701, ZN => n411);
   U65 : OR2_X1 port map( A1 => net264348, A2 => net272692, ZN => net270977);
   U66 : NAND2_X1 port map( A1 => n421, A2 => n422, ZN => n420);
   U67 : XNOR2_X1 port map( A => net272692, B => net273947, ZN => SUM(19));
   U68 : OAI21_X1 port map( B1 => B(25), B2 => n390, A => A(25), ZN => n429);
   U69 : NAND2_X1 port map( A1 => B(25), A2 => n390, ZN => n431);
   U70 : XNOR2_X1 port map( A => A(21), B => n413, ZN => n415);
   U71 : XNOR2_X1 port map( A => A(14), B => n414, ZN => n487);
   U72 : XNOR2_X1 port map( A => net287657, B => n415, ZN => SUM(21));
   U73 : NAND2_X1 port map( A1 => n417, A2 => n418, ZN => net264374);
   U74 : OAI21_X1 port map( B1 => n419, B2 => n423, A => n428, ZN => n427);
   U75 : NAND2_X1 port map( A1 => n493, A2 => n491, ZN => n492);
   U76 : INV_X1 port map( A => A(11), ZN => n478);
   U77 : NAND2_X1 port map( A1 => n463, A2 => A(11), ZN => n481);
   U78 : CLKBUF_X1 port map( A => A(13), Z => net271263);
   U79 : BUF_X1 port map( A => n434, Z => net276120);
   U80 : XNOR2_X1 port map( A => A(26), B => n416, ZN => n435);
   U81 : NAND2_X1 port map( A1 => A(24), A2 => B(24), ZN => n422);
   U82 : XNOR2_X1 port map( A => A(24), B => n433, ZN => n434);
   U83 : NAND2_X1 port map( A1 => A(26), A2 => B(26), ZN => n418);
   U84 : XNOR2_X1 port map( A => A(26), B => B(26), ZN => n424);
   U85 : NAND2_X1 port map( A1 => A(23), A2 => B(23), ZN => n428);
   U86 : XNOR2_X1 port map( A => A(23), B => B(23), ZN => n423);
   U87 : NAND2_X1 port map( A1 => n427, A2 => n434, ZN => n421);
   U88 : XNOR2_X1 port map( A => carry_23_port, B => n423, ZN => SUM(23));
   U89 : INV_X1 port map( A => carry_23_port, ZN => n419);
   U90 : XNOR2_X1 port map( A => n424, B => n425, ZN => SUM(26));
   U91 : NAND2_X1 port map( A1 => n435, A2 => n425, ZN => n417);
   U92 : XNOR2_X1 port map( A => n426, B => A(25), ZN => SUM(25));
   U93 : XNOR2_X1 port map( A => n479, B => n491, ZN => n488);
   U94 : NAND3_X1 port map( A1 => n517, A2 => n518, A3 => n519, ZN => n457);
   U95 : NAND3_X1 port map( A1 => n517, A2 => n518, A3 => n519, ZN => n459);
   U96 : NAND2_X1 port map( A1 => n472, A2 => n468, ZN => net275426);
   U97 : INV_X1 port map( A => A(13), ZN => n472);
   U98 : NAND2_X1 port map( A1 => A(10), A2 => B(10), ZN => n466);
   U99 : OAI21_X1 port map( B1 => A(10), B2 => B(10), A => net272728, ZN => 
                           n467);
   U100 : XNOR2_X1 port map( A => n494, B => n490, ZN => SUM(10));
   U101 : CLKBUF_X1 port map( A => A(10), Z => n494);
   U102 : NOR2_X1 port map( A1 => A(11), A2 => n463, ZN => n474);
   U103 : OAI21_X1 port map( B1 => n474, B2 => n475, A => n481, ZN => n479);
   U104 : XNOR2_X1 port map( A => net272728, B => B(10), ZN => n490);
   U105 : NAND2_X1 port map( A1 => n467, A2 => n466, ZN => n463);
   U106 : XNOR2_X1 port map( A => n463, B => n475, ZN => n489);
   U107 : NAND2_X1 port map( A1 => n479, A2 => A(12), ZN => n493);
   U108 : INV_X1 port map( A => A(12), ZN => n484);
   U109 : XNOR2_X1 port map( A => n489, B => n478, ZN => SUM(11));
   U110 : XNOR2_X1 port map( A => n459, B => n495, ZN => SUM(22));
   U111 : XNOR2_X1 port map( A => A(22), B => B(22), ZN => n495);
   U112 : CLKBUF_X1 port map( A => A(22), Z => n496);
   U113 : NAND2_X1 port map( A1 => n457, A2 => n496, ZN => n497);
   U114 : NAND2_X1 port map( A1 => n457, A2 => B(22), ZN => n498);
   U115 : NAND2_X1 port map( A1 => n496, A2 => B(22), ZN => n499);
   U116 : NAND3_X1 port map( A1 => n498, A2 => n497, A3 => n499, ZN => 
                           carry_23_port);
   U127 : INV_X1 port map( A => net273759, ZN => net276108);
   U128 : CLKBUF_X1 port map( A => A(9), Z => n510);
   U129 : CLKBUF_X1 port map( A => n438, Z => n515);
   U131 : NAND2_X1 port map( A1 => net274170, A2 => net273759, ZN => n432);
   U132 : AOI22_X1 port map( A1 => n391, A2 => net271263, B1 => net275426, B2 
                           => B(13), ZN => n511);
   U133 : XNOR2_X1 port map( A => n524, B => n458, ZN => SUM(34));
   U134 : XNOR2_X1 port map( A => A(13), B => B(13), ZN => n514);
   U135 : CLKBUF_X1 port map( A => A(32), Z => n512);
   U136 : NAND2_X1 port map( A1 => n513, A2 => n500, ZN => net272728);
   U137 : NAND2_X1 port map( A1 => n438, A2 => A(9), ZN => n513);
   U138 : XNOR2_X1 port map( A => n514, B => n391, ZN => SUM(13));
   U139 : AND2_X1 port map( A1 => n537, A2 => n511, ZN => net271611);
   U140 : AOI22_X1 port map( A1 => n391, A2 => net271263, B1 => net275426, B2 
                           => B(13), ZN => n485);
   U143 : XNOR2_X1 port map( A => A(33), B => n516, ZN => n461);
   U144 : AND2_X1 port map( A1 => net293635, A2 => A(15), ZN => net271387);
   U145 : XNOR2_X1 port map( A => net271313, B => net272691, ZN => SUM(17));
   U146 : NAND2_X1 port map( A1 => net264371, A2 => n412, ZN => n517);
   U147 : NAND2_X1 port map( A1 => n412, A2 => B(21), ZN => n519);
   U148 : XNOR2_X1 port map( A => net271166, B => net293635, ZN => SUM(15));
   U149 : INV_X1 port map( A => A(34), ZN => n535);
   U150 : INV_X1 port map( A => A(8), ZN => n538);
   U151 : INV_X1 port map( A => A(14), ZN => n537);
   U153 : XNOR2_X1 port map( A => n449, B => n450, ZN => SUM(41));
   U154 : OAI22_X1 port map( A1 => n451, A2 => B(40), B1 => n522, B2 => A(40), 
                           ZN => n449);
   U155 : XNOR2_X1 port map( A => n452, B => n453, ZN => SUM(40));
   U156 : INV_X1 port map( A => n452, ZN => n522);
   U157 : AND2_X1 port map( A1 => A(40), A2 => n522, ZN => n451);
   U158 : INV_X1 port map( A => n437, ZN => n524);
   U159 : INV_X1 port map( A => n503, ZN => n529);
   U160 : INV_X1 port map( A => A(33), ZN => n536);
   U161 : XNOR2_X1 port map( A => n512, B => n520, ZN => SUM(32));
   U162 : XNOR2_X1 port map( A => carry_32_port, B => B(32), ZN => n520);
   U163 : AOI21_X1 port map( B1 => n538, B2 => n440, A => n501, ZN => n438);
   U164 : AOI21_X1 port map( B1 => A(8), B2 => n527, A => B(8), ZN => n501);
   U165 : INV_X1 port map( A => n440, ZN => n527);
   U166 : XNOR2_X1 port map( A => A(39), B => n521, ZN => SUM(39));
   U167 : XNOR2_X1 port map( A => carry_39_port, B => B(39), ZN => n521);
   U168 : AOI21_X1 port map( B1 => A(39), B2 => B(39), A => n523, ZN => n452);
   U169 : INV_X1 port map( A => n454, ZN => n523);
   U170 : OAI21_X1 port map( B1 => A(39), B2 => B(39), A => carry_39_port, ZN 
                           => n454);
   U171 : XNOR2_X1 port map( A => B(8), B => n538, ZN => n441);
   U172 : XNOR2_X1 port map( A => A(5), B => B(5), ZN => n446);
   U173 : XNOR2_X1 port map( A => B(2), B => n541, ZN => n465);
   U174 : XNOR2_X1 port map( A => B(4), B => n540, ZN => n448);
   U175 : INV_X1 port map( A => A(2), ZN => n541);
   U176 : INV_X1 port map( A => A(4), ZN => n540);
   U177 : AOI21_X1 port map( B1 => n442, B2 => A(7), A => n528, ZN => n440);
   U178 : INV_X1 port map( A => n502, ZN => n528);
   U179 : OAI21_X1 port map( B1 => n442, B2 => A(7), A => B(7), ZN => n502);
   U180 : AOI21_X1 port map( B1 => n455, B2 => A(3), A => n532, ZN => n447);
   U181 : INV_X1 port map( A => n507, ZN => n532);
   U182 : OAI21_X1 port map( B1 => n455, B2 => A(3), A => B(3), ZN => n507);
   U183 : AOI21_X1 port map( B1 => n540, B2 => n447, A => n506, ZN => n445);
   U184 : AOI21_X1 port map( B1 => n531, B2 => A(4), A => B(4), ZN => n506);
   U185 : INV_X1 port map( A => n447, ZN => n531);
   U186 : AOI21_X1 port map( B1 => n541, B2 => n464, A => n508, ZN => n455);
   U187 : AOI21_X1 port map( B1 => n533, B2 => A(2), A => B(2), ZN => n508);
   U188 : INV_X1 port map( A => n464, ZN => n533);
   U189 : AOI21_X1 port map( B1 => n539, B2 => n503, A => n504, ZN => n442);
   U190 : INV_X1 port map( A => A(6), ZN => n539);
   U191 : AOI21_X1 port map( B1 => n529, B2 => A(6), A => B(6), ZN => n504);
   U192 : AOI21_X1 port map( B1 => n445, B2 => A(5), A => n530, ZN => n503);
   U193 : INV_X1 port map( A => n505, ZN => n530);
   U194 : OAI21_X1 port map( B1 => n445, B2 => A(5), A => B(5), ZN => n505);
   U195 : XNOR2_X1 port map( A => n440, B => n441, ZN => SUM(8));
   U196 : XNOR2_X1 port map( A => n464, B => n465, ZN => SUM(2));
   U197 : XNOR2_X1 port map( A => n447, B => n448, ZN => SUM(4));
   U198 : XNOR2_X1 port map( A => n445, B => n446, ZN => SUM(5));
   U199 : AOI21_X1 port map( B1 => A(1), B2 => B(1), A => n534, ZN => n464);
   U200 : INV_X1 port map( A => n509, ZN => n534);
   U201 : OAI211_X1 port map( C1 => A(1), C2 => B(1), A => A(0), B => B(0), ZN 
                           => n509);
   U202 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n470);
   U203 : XNOR2_X1 port map( A => net273128, B => net276120, ZN => SUM(24));
   U204 : AOI21_X1 port map( B1 => A(32), B2 => B(32), A => carry_32_port, ZN 
                           => n462);
   U205 : OAI21_X1 port map( B1 => n437, B2 => A(34), A => B(34), ZN => n436);
   U206 : XNOR2_X1 port map( A => n461, B => n394, ZN => SUM(33));
   U207 : OAI21_X1 port map( B1 => A(9), B2 => n438, A => B(9), ZN => n500);
   U208 : OAI21_X1 port map( B1 => n524, B2 => n535, A => n436, ZN => 
                           carry_35_port);
   U209 : OAI21_X1 port map( B1 => n394, B2 => n536, A => n460, ZN => n437);
   U210 : OAI21_X1 port map( B1 => n393, B2 => A(33), A => B(33), ZN => n460);
   U211 : INV_X1 port map( A => n462, ZN => n525);
   U212 : XNOR2_X1 port map( A => n487, B => n511, ZN => SUM(14));
   U213 : INV_X1 port map( A => n485, ZN => n526);
   U214 : INV_X1 port map( A => n430, ZN => net264371);
   U215 : AOI21_X1 port map( B1 => n526, B2 => A(14), A => B(14), ZN => n486);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT40_DW01_add_0 is

   port( A, B : in std_logic_vector (39 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (39 downto 0);  CO : out std_logic);

end RCA_NBIT40_DW01_add_0;

architecture SYN_rpl of RCA_NBIT40_DW01_add_0 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_39_port, carry_38_port, carry_37_port, carry_36_port, 
      carry_34_port, carry_33_port, carry_30_port, carry_29_port, carry_28_port
      , carry_6_port, carry_5_port, carry_4_port, carry_3_port, carry_2_port, 
      n1, n392, n393, n396, n397, n398, n399, n400, n401, n402, n403, n404, 
      n405, n407, n411, n412, n416, n417, n419, n432, n440, n444, n446, n447, 
      n448, n451, n456, n457, n458, n459, net264311, net264313, net264331, 
      net271177, net271574, net271642, net271699, net271816, net273116, 
      net273280, net273603, net273719, net274117, net274213, net275813, 
      net271173, n454, n452, n450, net283792, net283791, net285233, net285232, 
      net285370, net287643, net273484, net269658, net285260, net264330, n423, 
      n422, net273117, net270215, net283825, net283793, net283773, net272440, 
      net272323, n437, net285167, net283842, net280555, net279578, net276697, 
      net273656, net273294, net273118, net271335, net264328, net264306, n433, 
      n430, n429, n427, n426, n425, n424, n358, n359, n360, n361, n362, n363, 
      n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, 
      n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, 
      n388, n389, n390, n391, n394, n395, n406, n408, n409, n410, n413, n414, 
      n415, n418, n420, n421, n428, n431, n434, n435, n436, n438, n439, n441, 
      n442, n443, n445, n449, n453, n455, n460, n461, n462, n463, n464, n465, 
      n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, 
      n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, 
      n490, n491, n492, n493, n494, n495, n496, n497 : std_logic;

begin
   
   U1_38 : FA_X1 port map( A => A(38), B => B(38), CI => carry_38_port, CO => 
                           carry_39_port, S => SUM(38));
   U1_37 : FA_X1 port map( A => A(37), B => B(37), CI => carry_37_port, CO => 
                           carry_38_port, S => SUM(37));
   U1_36 : FA_X1 port map( A => A(36), B => B(36), CI => carry_36_port, CO => 
                           carry_37_port, S => SUM(36));
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => n489, CO => 
                           carry_36_port, S => SUM(35));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => n490, CO => 
                           carry_33_port, S => SUM(32));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U101 : XOR2_X1 port map( A => n480, B => n402, Z => SUM(8));
   U103 : XOR2_X1 port map( A => B(7), B => n478, Z => n404);
   U104 : XOR2_X1 port map( A => A(6), B => n405, Z => SUM(6));
   U105 : XOR2_X1 port map( A => carry_6_port, B => B(6), Z => n405);
   U108 : XOR2_X1 port map( A => carry_34_port, B => n393, Z => SUM(34));
   U111 : XOR2_X1 port map( A => carry_30_port, B => n407, Z => SUM(30));
   U130 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : BUF_X1 port map( A => A(10), Z => n358);
   U2 : NAND2_X1 port map( A1 => n413, A2 => n391, ZN => n386);
   U3 : INV_X1 port map( A => B(13), ZN => net271574);
   U4 : XNOR2_X1 port map( A => B(25), B => A(25), ZN => n411);
   U5 : INV_X1 port map( A => B(39), ZN => n470);
   U6 : INV_X1 port map( A => B(26), ZN => n414);
   U7 : AND2_X1 port map( A1 => n492, A2 => n482, ZN => net274117);
   U8 : INV_X1 port map( A => B(14), ZN => n455);
   U9 : INV_X1 port map( A => B(16), ZN => n379);
   U10 : NAND2_X1 port map( A1 => n389, A2 => n390, ZN => n383);
   U11 : INV_X1 port map( A => B(24), ZN => n389);
   U12 : INV_X1 port map( A => B(20), ZN => n373);
   U13 : INV_X1 port map( A => B(34), ZN => n467);
   U14 : INV_X1 port map( A => B(11), ZN => n465);
   U15 : INV_X1 port map( A => B(30), ZN => n485);
   U16 : OAI21_X1 port map( B1 => net285370, B2 => n391, A => n406, ZN => n359)
                           ;
   U17 : OAI21_X1 port map( B1 => n461, B2 => n449, A => n453, ZN => n360);
   U18 : AOI22_X1 port map( A1 => B(20), A2 => A(20), B1 => n424, B2 => n425, 
                           ZN => n361);
   U19 : NAND2_X1 port map( A1 => net264328, A2 => n362, ZN => net279578);
   U20 : AND2_X1 port map( A1 => net273118, A2 => A(19), ZN => n362);
   U21 : NAND2_X1 port map( A1 => B(26), A2 => n408, ZN => n363);
   U22 : INV_X1 port map( A => n361, ZN => n364);
   U23 : NAND2_X1 port map( A1 => n381, A2 => n382, ZN => n365);
   U24 : OR2_X1 port map( A1 => n370, A2 => n412, ZN => n384);
   U25 : OAI21_X1 port map( B1 => net271816, B2 => n464, A => B(11), ZN => n366
                           );
   U26 : OR2_X2 port map( A1 => n394, A2 => net273484, ZN => n410);
   U27 : OR2_X1 port map( A1 => n466, A2 => n454, ZN => n367);
   U28 : BUF_X1 port map( A => n399, Z => n477);
   U29 : NAND2_X1 port map( A1 => n363, A2 => n410, ZN => n368);
   U30 : CLKBUF_X1 port map( A => A(17), Z => net283825);
   U31 : OAI21_X1 port map( B1 => n428, B2 => net274117, A => B(13), ZN => n369
                           );
   U32 : INV_X1 port map( A => B(9), ZN => n487);
   U33 : AND2_X1 port map( A1 => n415, A2 => B(24), ZN => n370);
   U34 : INV_X1 port map( A => B(8), ZN => n471);
   U35 : NAND2_X1 port map( A1 => n422, A2 => n372, ZN => n371);
   U36 : NAND2_X1 port map( A1 => net264330, A2 => n418, ZN => n372);
   U37 : INV_X1 port map( A => B(31), ZN => n484);
   U38 : INV_X1 port map( A => B(19), ZN => n374);
   U39 : NAND2_X1 port map( A1 => n363, A2 => n410, ZN => n375);
   U40 : OAI21_X1 port map( B1 => net285370, B2 => n391, A => n406, ZN => n387)
                           ;
   U41 : INV_X1 port map( A => B(25), ZN => n391);
   U42 : INV_X1 port map( A => A(25), ZN => n406);
   U43 : AND2_X1 port map( A1 => net264331, A2 => net271642, ZN => n439);
   U44 : XNOR2_X1 port map( A => net285167, B => n425, ZN => SUM(20));
   U45 : AND2_X1 port map( A1 => net283842, A2 => net279578, ZN => net285167);
   U46 : OAI21_X1 port map( B1 => net276697, B2 => net273656, A => B(19), ZN =>
                           net283842);
   U47 : INV_X1 port map( A => net264306, ZN => net276697);
   U48 : OAI21_X1 port map( B1 => net273656, B2 => net276697, A => B(19), ZN =>
                           n427);
   U49 : INV_X1 port map( A => A(19), ZN => net264306);
   U50 : XNOR2_X1 port map( A => A(20), B => n373, ZN => n425);
   U51 : AOI22_X1 port map( A1 => B(20), A2 => A(20), B1 => n424, B2 => n425, 
                           ZN => net285260);
   U52 : NAND2_X1 port map( A1 => net279578, A2 => n427, ZN => n424);
   U53 : AND2_X1 port map( A1 => net264328, A2 => net273118, ZN => net273656);
   U54 : INV_X1 port map( A => n430, ZN => net264328);
   U55 : NAND2_X1 port map( A1 => net264328, A2 => net273118, ZN => n426);
   U56 : AOI21_X1 port map( B1 => n429, B2 => A(18), A => B(18), ZN => n430);
   U57 : NOR2_X1 port map( A1 => n433, A2 => net271177, ZN => n429);
   U58 : AOI21_X1 port map( B1 => net273294, B2 => net272323, A => B(17), ZN =>
                           n433);
   U59 : BUF_X1 port map( A => A(17), Z => net273294);
   U60 : AOI21_X1 port map( B1 => net273294, B2 => net272323, A => B(17), ZN =>
                           net280555);
   U61 : XNOR2_X1 port map( A => A(19), B => n374, ZN => net271335);
   U62 : XNOR2_X1 port map( A => n426, B => net271335, ZN => SUM(19));
   U63 : XNOR2_X1 port map( A => A(18), B => B(18), ZN => net270215);
   U64 : OR2_X1 port map( A1 => net273117, A2 => A(18), ZN => net273118);
   U65 : NOR2_X1 port map( A1 => net280555, A2 => net271177, ZN => net273117);
   U66 : XNOR2_X1 port map( A => net283773, B => B(17), ZN => net283793);
   U67 : INV_X1 port map( A => A(17), ZN => net264311);
   U68 : NAND2_X1 port map( A1 => n366, A2 => net271699, ZN => n376);
   U69 : XNOR2_X1 port map( A => net287643, B => n368, ZN => SUM(27));
   U70 : XNOR2_X1 port map( A => net283793, B => net283825, ZN => SUM(17));
   U71 : NAND2_X1 port map( A1 => n378, A2 => n377, ZN => net283773);
   U72 : NAND2_X1 port map( A1 => n381, A2 => n382, ZN => n378);
   U73 : AND2_X1 port map( A1 => n365, A2 => n377, ZN => n432);
   U74 : NAND2_X1 port map( A1 => n365, A2 => n377, ZN => net272323);
   U75 : CLKBUF_X1 port map( A => A(16), Z => n382);
   U76 : NAND2_X1 port map( A1 => n380, A2 => n379, ZN => n381);
   U77 : NAND2_X1 port map( A1 => net283792, A2 => n360, ZN => n380);
   U78 : NAND2_X1 port map( A1 => net272440, A2 => B(16), ZN => n377);
   U79 : XNOR2_X1 port map( A => A(16), B => B(16), ZN => n437);
   U80 : AND2_X1 port map( A1 => net283791, A2 => net283792, ZN => net272440);
   U81 : XNOR2_X1 port map( A => net272440, B => n437, ZN => SUM(16));
   U82 : NAND2_X1 port map( A1 => n359, A2 => n386, ZN => n385);
   U83 : NAND2_X1 port map( A1 => n385, A2 => n394, ZN => n408);
   U84 : INV_X1 port map( A => A(26), ZN => n394);
   U85 : NAND2_X1 port map( A1 => n387, A2 => n386, ZN => net273484);
   U86 : XNOR2_X1 port map( A => A(24), B => B(24), ZN => n395);
   U87 : XNOR2_X1 port map( A => n412, B => n395, ZN => SUM(24));
   U88 : NAND2_X1 port map( A1 => n383, A2 => n384, ZN => net285370);
   U89 : NAND2_X1 port map( A1 => n383, A2 => n384, ZN => n413);
   U90 : NAND2_X1 port map( A1 => n410, A2 => n409, ZN => n388);
   U91 : NAND2_X1 port map( A1 => n375, A2 => B(27), ZN => net285233);
   U92 : NAND2_X1 port map( A1 => A(27), A2 => n388, ZN => net285232);
   U93 : XNOR2_X1 port map( A => A(26), B => n414, ZN => net269658);
   U94 : INV_X1 port map( A => n415, ZN => n390);
   U95 : NAND2_X1 port map( A1 => B(26), A2 => n408, ZN => n409);
   U96 : BUF_X1 port map( A => A(24), Z => n415);
   U97 : XNOR2_X1 port map( A => net273117, B => net270215, ZN => SUM(18));
   U98 : CLKBUF_X1 port map( A => n371, Z => net273116);
   U99 : OR2_X1 port map( A1 => A(22), A2 => n371, ZN => net271642);
   U100 : AOI21_X1 port map( B1 => n371, B2 => A(22), A => B(22), ZN => n419);
   U102 : OAI21_X1 port map( B1 => n364, B2 => n418, A => B(21), ZN => n422);
   U106 : BUF_X1 port map( A => A(21), Z => n418);
   U107 : INV_X1 port map( A => net285260, ZN => net264330);
   U109 : XNOR2_X1 port map( A => net264330, B => n423, ZN => SUM(21));
   U110 : XNOR2_X1 port map( A => A(21), B => B(21), ZN => n423);
   U112 : XNOR2_X1 port map( A => net273484, B => net269658, ZN => SUM(26));
   U113 : XNOR2_X1 port map( A => A(27), B => B(27), ZN => net287643);
   U114 : BUF_X1 port map( A => n420, Z => net273719);
   U115 : NAND2_X1 port map( A1 => n439, A2 => n481, ZN => n473);
   U116 : OAI21_X1 port map( B1 => n477, B2 => n479, A => n456, ZN => n420);
   U117 : XNOR2_X1 port map( A => carry_33_port, B => n421, ZN => SUM(33));
   U118 : XNOR2_X1 port map( A => A(33), B => B(33), ZN => n421);
   U119 : OR2_X1 port map( A1 => n454, A2 => n466, ZN => n450);
   U120 : CLKBUF_X1 port map( A => A(13), Z => n428);
   U121 : NAND2_X1 port map( A1 => n460, A2 => n455, ZN => n431);
   U122 : NAND2_X1 port map( A1 => carry_33_port, A2 => A(33), ZN => n434);
   U123 : NAND2_X1 port map( A1 => carry_33_port, A2 => B(33), ZN => n435);
   U124 : NAND2_X1 port map( A1 => A(33), A2 => B(33), ZN => n436);
   U125 : NAND3_X1 port map( A1 => n434, A2 => n435, A3 => n436, ZN => 
                           carry_34_port);
   U126 : NAND2_X1 port map( A1 => A(27), A2 => B(27), ZN => n438);
   U127 : NAND3_X1 port map( A1 => net285233, A2 => net285232, A3 => n438, ZN 
                           => carry_28_port);
   U128 : NAND2_X1 port map( A1 => n445, A2 => n462, ZN => n443);
   U129 : OAI21_X1 port map( B1 => n461, B2 => n449, A => n453, ZN => net283791
                           );
   U131 : NAND2_X1 port map( A1 => n431, A2 => n443, ZN => net274213);
   U132 : NAND2_X1 port map( A1 => n431, A2 => n443, ZN => n461);
   U133 : NAND2_X1 port map( A1 => n463, A2 => net271173, ZN => n460);
   U134 : INV_X1 port map( A => A(15), ZN => n449);
   U135 : OAI21_X1 port map( B1 => net274117, B2 => n428, A => B(13), ZN => 
                           n442);
   U136 : NAND2_X1 port map( A1 => n442, A2 => n441, ZN => net271173);
   U137 : NAND2_X1 port map( A1 => net274117, A2 => n428, ZN => n441);
   U138 : AND2_X1 port map( A1 => n441, A2 => n369, ZN => n462);
   U139 : INV_X1 port map( A => B(15), ZN => n453);
   U140 : XNOR2_X1 port map( A => A(15), B => n453, ZN => n440);
   U141 : INV_X1 port map( A => n463, ZN => n445);
   U142 : BUF_X1 port map( A => A(14), Z => n463);
   U143 : NAND2_X1 port map( A1 => net274213, A2 => n449, ZN => net283792);
   U144 : NOR2_X1 port map( A1 => n466, A2 => n454, ZN => n464);
   U145 : XNOR2_X1 port map( A => n367, B => n452, ZN => SUM(11));
   U146 : XNOR2_X1 port map( A => A(11), B => n465, ZN => n452);
   U147 : OR2_X1 port map( A1 => n450, A2 => net264313, ZN => net271699);
   U148 : NOR2_X1 port map( A1 => B(10), A2 => n420, ZN => n466);
   U149 : AOI21_X1 port map( B1 => n420, B2 => B(10), A => n358, ZN => n454);
   U150 : INV_X1 port map( A => A(11), ZN => net264313);
   U151 : OAI21_X1 port map( B1 => net271816, B2 => n464, A => B(11), ZN => 
                           n451);
   U152 : XNOR2_X1 port map( A => A(10), B => B(10), ZN => net273280);
   U153 : XNOR2_X1 port map( A => net273603, B => net271173, ZN => SUM(14));
   U154 : XNOR2_X1 port map( A => A(34), B => n467, ZN => n393);
   U155 : CLKBUF_X1 port map( A => A(30), Z => n468);
   U156 : INV_X1 port map( A => net285370, ZN => net275813);
   U157 : XNOR2_X1 port map( A => A(14), B => B(14), ZN => net273603);
   U158 : XNOR2_X1 port map( A => net273116, B => n469, ZN => SUM(22));
   U159 : XNOR2_X1 port map( A => A(22), B => B(22), ZN => n469);
   U160 : XNOR2_X1 port map( A => carry_39_port, B => n470, ZN => n488);
   U161 : XNOR2_X1 port map( A => A(8), B => n471, ZN => n402);
   U162 : CLKBUF_X1 port map( A => A(8), Z => n472);
   U163 : CLKBUF_X1 port map( A => n401, Z => n480);
   U164 : XNOR2_X1 port map( A => net273719, B => net273280, ZN => SUM(10));
   U165 : NAND2_X1 port map( A1 => n416, A2 => n473, ZN => n412);
   U166 : AND2_X1 port map( A1 => net264331, A2 => net271642, ZN => n474);
   U167 : AND2_X1 port map( A1 => n476, A2 => n495, ZN => n475);
   U168 : OR2_X1 port map( A1 => B(6), A2 => A(6), ZN => n476);
   U169 : NAND2_X1 port map( A1 => n476, A2 => n495, ZN => n403);
   U170 : INV_X1 port map( A => n496, ZN => n478);
   U171 : INV_X1 port map( A => net264313, ZN => net271816);
   U172 : NAND2_X1 port map( A1 => net271699, A2 => n451, ZN => n447);
   U173 : INV_X1 port map( A => A(9), ZN => n479);
   U174 : XNOR2_X1 port map( A => A(13), B => net271574, ZN => n446);
   U175 : OAI21_X1 port map( B1 => n403, B2 => n496, A => n458, ZN => n401);
   U176 : INV_X1 port map( A => n497, ZN => n481);
   U177 : OR2_X1 port map( A1 => n376, A2 => A(12), ZN => n482);
   U178 : NAND2_X1 port map( A1 => n492, A2 => n482, ZN => n444);
   U179 : AND2_X1 port map( A1 => net264311, A2 => n432, ZN => net271177);
   U180 : CLKBUF_X1 port map( A => A(31), Z => n483);
   U181 : XNOR2_X1 port map( A => A(31), B => n484, ZN => n397);
   U182 : XNOR2_X1 port map( A => A(30), B => n485, ZN => n407);
   U183 : XNOR2_X1 port map( A => n486, B => n376, ZN => SUM(12));
   U184 : XNOR2_X1 port map( A => B(12), B => A(12), ZN => n486);
   U185 : XNOR2_X1 port map( A => A(9), B => n487, ZN => n400);
   U186 : XOR2_X1 port map( A => n488, B => A(39), Z => SUM(39));
   U187 : AOI21_X1 port map( B1 => A(6), B2 => B(6), A => carry_6_port, ZN => 
                           n459);
   U188 : OAI21_X1 port map( B1 => n475, B2 => A(7), A => B(7), ZN => n458);
   U189 : INV_X1 port map( A => A(7), ZN => n496);
   U190 : INV_X1 port map( A => n398, ZN => n491);
   U191 : AOI22_X1 port map( A1 => B(34), A2 => A(34), B1 => n393, B2 => 
                           carry_34_port, ZN => n392);
   U192 : INV_X1 port map( A => n392, ZN => n489);
   U193 : INV_X1 port map( A => n396, ZN => n490);
   U194 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U195 : OAI21_X1 port map( B1 => n474, B2 => n481, A => B(23), ZN => n416);
   U196 : INV_X1 port map( A => A(23), ZN => n497);
   U197 : AOI22_X1 port map( A1 => B(31), A2 => n483, B1 => n491, B2 => n397, 
                           ZN => n396);
   U198 : XNOR2_X1 port map( A => n397, B => n398, ZN => SUM(31));
   U199 : XNOR2_X1 port map( A => net274213, B => n440, ZN => SUM(15));
   U200 : XNOR2_X1 port map( A => A(23), B => B(23), ZN => n417);
   U201 : XNOR2_X1 port map( A => n439, B => n417, ZN => SUM(23));
   U202 : INV_X1 port map( A => n419, ZN => net264331);
   U203 : XNOR2_X1 port map( A => n446, B => n444, ZN => SUM(13));
   U204 : XNOR2_X1 port map( A => n403, B => n404, ZN => SUM(7));
   U205 : XNOR2_X1 port map( A => n477, B => n400, ZN => SUM(9));
   U206 : INV_X1 port map( A => n399, ZN => n493);
   U207 : AOI21_X1 port map( B1 => n401, B2 => A(8), A => B(8), ZN => n457);
   U208 : AOI21_X1 port map( B1 => n447, B2 => A(12), A => B(12), ZN => n448);
   U209 : OAI21_X1 port map( B1 => n493, B2 => A(9), A => B(9), ZN => n456);
   U210 : INV_X1 port map( A => n459, ZN => n495);
   U211 : INV_X1 port map( A => n448, ZN => n492);
   U212 : OAI21_X1 port map( B1 => n480, B2 => n472, A => n494, ZN => n399);
   U213 : INV_X1 port map( A => n457, ZN => n494);
   U214 : AOI22_X1 port map( A1 => n407, A2 => carry_30_port, B1 => n468, B2 =>
                           B(30), ZN => n398);
   U215 : XNOR2_X1 port map( A => net275813, B => n411, ZN => SUM(25));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT38_DW01_add_0 is

   port( A, B : in std_logic_vector (37 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (37 downto 0);  CO : out std_logic);

end RCA_NBIT38_DW01_add_0;

architecture SYN_rpl of RCA_NBIT38_DW01_add_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_36_port, carry_34_port, carry_33_port, carry_4_port, 
      carry_3_port, carry_2_port, n1, n479, n480, n481, n482, n484, n487, n489,
      n490, n491, n492, n493, n496, n498, n499, n500, n501, n502, n503, n504, 
      n505, n507, n508, n510, n511, n513, n517, n522, n523, n525, n526, n531, 
      n544, n547, n548, n553, n556, n557, n559, n560, n561, n563, n564, n565, 
      n566, n567, n568, net264260, net264281, net269617, net271149, net271141, 
      net271140, net272170, net280507, net274327, n554, n551, n550, net293549, 
      net293534, n545, n542, n541, n540, n539, n538, n537, n536, n535, n534, 
      n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, 
      n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, 
      n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, 
      n471, n472, n473, n474, n475, n476, n477, n478, n483, n485, n486, n488, 
      n494, n495, n497, n506, n509, n512, n514, n515, n516, n518, n519, n520, 
      n521, n524, n527, n528, n529, n530, n532, n533, n543, n546, n549, n552, 
      n555, n558, n562, n569, n570, n571, n572, n573, n574, n575, n576, n577, 
      n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, 
      n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, 
      n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, 
      n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, 
      n626, n627, n628, n629, n630, n631, n632, n633, n634, n635 : std_logic;

begin
   
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => n617, CO => 
                           carry_36_port, S => SUM(35));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => n568, CO => 
                           carry_33_port, S => SUM(32));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U137 : XOR2_X1 port map( A => n573, B => n489, Z => SUM(5));
   U138 : XOR2_X1 port map( A => A(4), B => n490, Z => SUM(4));
   U139 : XOR2_X1 port map( A => carry_4_port, B => B(4), Z => n490);
   U140 : XOR2_X1 port map( A => n491, B => n492, Z => SUM(37));
   U141 : XOR2_X1 port map( A => carry_36_port, B => n493, Z => SUM(36));
   U142 : XOR2_X1 port map( A => A(36), B => B(36), Z => n493);
   U143 : XOR2_X1 port map( A => carry_34_port, B => n480, Z => SUM(34));
   U167 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : AOI21_X1 port map( B1 => n583, B2 => n443, A => B(22), ZN => n435);
   U2 : XNOR2_X1 port map( A => n436, B => n578, ZN => SUM(24));
   U3 : XNOR2_X1 port map( A => A(24), B => B(24), ZN => n436);
   U4 : BUF_X1 port map( A => n471, Z => n437);
   U5 : INV_X1 port map( A => B(19), ZN => n478);
   U6 : INV_X1 port map( A => B(34), ZN => n576);
   U7 : INV_X1 port map( A => B(25), ZN => n612);
   U8 : XNOR2_X1 port map( A => n477, B => net293534, ZN => SUM(18));
   U9 : INV_X1 port map( A => B(29), ZN => n587);
   U10 : CLKBUF_X1 port map( A => A(29), Z => n472);
   U11 : NAND3_X1 port map( A1 => n606, A2 => n607, A3 => n608, ZN => n438);
   U12 : AND2_X1 port map( A1 => n539, A2 => n468, ZN => n439);
   U13 : AOI21_X1 port map( B1 => n530, B2 => n472, A => B(29), ZN => n440);
   U14 : AND2_X1 port map( A1 => n539, A2 => n468, ZN => n537);
   U15 : AND2_X1 port map( A1 => n483, A2 => n485, ZN => n441);
   U16 : CLKBUF_X1 port map( A => A(11), Z => n442);
   U17 : BUF_X1 port map( A => A(22), Z => n443);
   U18 : NAND2_X1 port map( A1 => n542, A2 => net271149, ZN => n444);
   U19 : OR2_X2 port map( A1 => net272170, A2 => net264260, ZN => net271149);
   U20 : NOR2_X1 port map( A1 => n564, A2 => n445, ZN => n454);
   U21 : NOR2_X1 port map( A1 => A(6), A2 => n487, ZN => n445);
   U22 : OAI21_X1 port map( B1 => n621, B2 => n549, A => B(25), ZN => n446);
   U23 : BUF_X1 port map( A => n454, Z => n594);
   U24 : BUF_X1 port map( A => n559, Z => n562);
   U25 : AND2_X1 port map( A1 => n623, A2 => n457, ZN => n447);
   U26 : CLKBUF_X1 port map( A => n552, Z => n448);
   U27 : OR2_X1 port map( A1 => n512, A2 => n631, ZN => n601);
   U28 : BUF_X1 port map( A => n561, Z => n449);
   U29 : BUF_X1 port map( A => n625, Z => n572);
   U30 : BUF_X1 port map( A => n531, Z => net293549);
   U31 : INV_X1 port map( A => n603, ZN => n450);
   U32 : INV_X1 port map( A => n598, ZN => n451);
   U33 : NAND2_X1 port map( A1 => n450, A2 => n451, ZN => n452);
   U34 : NAND2_X1 port map( A1 => n452, A2 => n453, ZN => n584);
   U35 : NOR2_X1 port map( A1 => n627, A2 => n564, ZN => n453);
   U36 : NOR2_X2 port map( A1 => n526, A2 => n528, ZN => n522);
   U37 : NOR2_X1 port map( A1 => n604, A2 => n543, ZN => n455);
   U38 : NOR2_X1 port map( A1 => n455, A2 => n449, ZN => n456);
   U39 : BUF_X1 port map( A => n484, Z => n604);
   U40 : INV_X1 port map( A => B(31), ZN => n611);
   U41 : CLKBUF_X1 port map( A => n556, Z => n602);
   U42 : NAND2_X1 port map( A1 => n623, A2 => n457, ZN => n553);
   U43 : OR2_X1 port map( A1 => A(10), A2 => n556, ZN => n457);
   U44 : INV_X1 port map( A => B(15), ZN => n461);
   U45 : XNOR2_X1 port map( A => n533, B => n509, ZN => SUM(22));
   U46 : XNOR2_X1 port map( A => n536, B => B(17), ZN => SUM(17));
   U47 : NAND2_X1 port map( A1 => n535, A2 => n464, ZN => n536);
   U48 : OR2_X1 port map( A1 => n537, A2 => n458, ZN => n464);
   U49 : INV_X1 port map( A => A(17), ZN => n458);
   U50 : NOR2_X1 port map( A1 => n458, A2 => n439, ZN => n534);
   U51 : NAND2_X1 port map( A1 => n439, A2 => n458, ZN => n535);
   U52 : OAI21_X1 port map( B1 => n534, B2 => B(17), A => n535, ZN => n531);
   U53 : NAND2_X1 port map( A1 => n467, A2 => n463, ZN => n468);
   U54 : CLKBUF_X1 port map( A => A(16), Z => n463);
   U55 : OAI21_X1 port map( B1 => n538, B2 => A(16), A => B(16), ZN => n539);
   U56 : NAND2_X1 port map( A1 => n469, A2 => net271149, ZN => n538);
   U57 : OAI21_X1 port map( B1 => n460, B2 => A(15), A => B(15), ZN => n469);
   U58 : INV_X1 port map( A => n541, ZN => n460);
   U59 : OAI21_X1 port map( B1 => n460, B2 => A(15), A => B(15), ZN => n542);
   U60 : OAI21_X1 port map( B1 => n465, B2 => n466, A => n459, ZN => n541);
   U61 : INV_X1 port map( A => n545, ZN => n459);
   U62 : OAI21_X1 port map( B1 => n465, B2 => n466, A => n459, ZN => net272170)
                           ;
   U63 : AOI21_X1 port map( B1 => n544, B2 => A(14), A => B(14), ZN => n545);
   U64 : BUF_X1 port map( A => n544, Z => n466);
   U65 : XNOR2_X1 port map( A => n466, B => n462, ZN => SUM(14));
   U66 : CLKBUF_X1 port map( A => A(14), Z => n465);
   U67 : XNOR2_X1 port map( A => n444, B => n540, ZN => SUM(16));
   U68 : XNOR2_X1 port map( A => A(16), B => B(16), ZN => n540);
   U69 : NAND2_X1 port map( A1 => n542, A2 => net271149, ZN => n467);
   U70 : INV_X1 port map( A => A(15), ZN => net264260);
   U71 : XNOR2_X1 port map( A => A(15), B => n461, ZN => net269617);
   U72 : XNOR2_X1 port map( A => A(14), B => B(14), ZN => n462);
   U73 : AOI21_X1 port map( B1 => n583, B2 => n443, A => B(22), ZN => n470);
   U74 : AOI21_X1 port map( B1 => n630, B2 => n509, A => n470, ZN => n471);
   U75 : OAI211_X1 port map( C1 => net293549, C2 => n476, A => n474, B => n478,
                           ZN => n485);
   U76 : INV_X1 port map( A => n531, ZN => net293534);
   U77 : OAI211_X1 port map( C1 => net293549, C2 => n473, A => n474, B => n475,
                           ZN => net271141);
   U78 : OAI21_X1 port map( B1 => net293549, B2 => n473, A => n474, ZN => 
                           net280507);
   U79 : XNOR2_X1 port map( A => B(18), B => A(18), ZN => n477);
   U80 : NAND2_X1 port map( A1 => A(18), A2 => B(18), ZN => n474);
   U81 : NOR2_X1 port map( A1 => A(18), A2 => B(18), ZN => n473);
   U82 : NOR2_X1 port map( A1 => B(18), A2 => A(18), ZN => n476);
   U83 : INV_X1 port map( A => A(19), ZN => n475);
   U84 : XNOR2_X1 port map( A => B(19), B => A(19), ZN => net274327);
   U85 : NAND2_X1 port map( A1 => n475, A2 => n478, ZN => n483);
   U86 : XNOR2_X1 port map( A => A(12), B => B(12), ZN => n495);
   U87 : AOI21_X1 port map( B1 => n550, B2 => A(12), A => B(12), ZN => n551);
   U88 : INV_X1 port map( A => n551, ZN => net264281);
   U89 : OR2_X1 port map( A1 => A(12), A2 => n550, ZN => net271140);
   U90 : NAND2_X1 port map( A1 => n554, A2 => n494, ZN => n550);
   U91 : XNOR2_X1 port map( A => n550, B => n495, ZN => SUM(12));
   U92 : OR2_X1 port map( A1 => n553, A2 => n486, ZN => n494);
   U93 : INV_X1 port map( A => A(11), ZN => n486);
   U94 : OAI21_X1 port map( B1 => n447, B2 => n442, A => B(11), ZN => n554);
   U95 : XNOR2_X1 port map( A => n447, B => n488, ZN => SUM(11));
   U96 : XNOR2_X1 port map( A => A(11), B => B(11), ZN => n488);
   U97 : XNOR2_X1 port map( A => net280507, B => net274327, ZN => SUM(19));
   U98 : NAND2_X1 port map( A1 => n446, A2 => n601, ZN => n497);
   U99 : BUF_X1 port map( A => A(30), Z => n521);
   U100 : INV_X1 port map( A => n504, ZN => n506);
   U101 : AND2_X1 port map( A1 => n523, A2 => n519, ZN => n509);
   U102 : OAI21_X1 port map( B1 => n448, B2 => n610, A => n622, ZN => n512);
   U103 : XNOR2_X1 port map( A => n514, B => n512, ZN => SUM(25));
   U104 : XNOR2_X1 port map( A => A(25), B => n612, ZN => n514);
   U105 : AND2_X1 port map( A1 => n504, A2 => n632, ZN => n515);
   U106 : NOR2_X1 port map( A1 => n505, A2 => n515, ZN => n501);
   U107 : BUF_X1 port map( A => n501, Z => n546);
   U108 : NOR2_X1 port map( A1 => n570, A2 => n440, ZN => n516);
   U109 : NOR2_X1 port map( A1 => n499, A2 => n570, ZN => n518);
   U110 : NAND2_X1 port map( A1 => n523, A2 => n519, ZN => n583);
   U111 : NAND2_X1 port map( A1 => n522, A2 => A(21), ZN => n519);
   U112 : CLKBUF_X1 port map( A => A(26), Z => n520);
   U113 : BUF_X1 port map( A => A(24), Z => n552);
   U114 : XNOR2_X1 port map( A => n522, B => n524, ZN => SUM(21));
   U115 : XNOR2_X1 port map( A => A(21), B => B(21), ZN => n524);
   U116 : CLKBUF_X1 port map( A => n581, Z => n527);
   U117 : AND2_X1 port map( A1 => n629, A2 => n525, ZN => n528);
   U118 : BUF_X1 port map( A => A(7), Z => n529);
   U119 : OR2_X1 port map( A1 => n619, A2 => n571, ZN => n530);
   U120 : AOI21_X1 port map( B1 => n630, B2 => n509, A => n435, ZN => n532);
   U121 : XNOR2_X1 port map( A => B(22), B => n630, ZN => n533);
   U122 : CLKBUF_X1 port map( A => A(8), Z => n543);
   U123 : CLKBUF_X1 port map( A => A(25), Z => n549);
   U124 : XNOR2_X1 port map( A => n555, B => n562, ZN => SUM(9));
   U125 : XOR2_X1 port map( A => A(9), B => B(9), Z => n555);
   U126 : XNOR2_X1 port map( A => n558, B => n594, ZN => SUM(7));
   U127 : XNOR2_X1 port map( A => n529, B => B(7), ZN => n558);
   U128 : XNOR2_X1 port map( A => A(8), B => B(8), ZN => n597);
   U129 : XNOR2_X1 port map( A => n603, B => n569, ZN => SUM(6));
   U130 : XNOR2_X1 port map( A => A(6), B => B(6), ZN => n569);
   U131 : AND2_X1 port map( A1 => n634, A2 => n498, ZN => n570);
   U132 : AND2_X1 port map( A1 => A(28), A2 => n501, ZN => n571);
   U133 : NOR2_X1 port map( A1 => n571, A2 => n619, ZN => n498);
   U134 : AND2_X1 port map( A1 => n591, A2 => n620, ZN => n588);
   U135 : INV_X1 port map( A => n565, ZN => n573);
   U136 : XNOR2_X1 port map( A => A(10), B => B(10), ZN => n593);
   U144 : AND2_X1 port map( A1 => n625, A2 => n581, ZN => n574);
   U145 : AND2_X1 port map( A1 => n441, A2 => net271141, ZN => n575);
   U146 : XNOR2_X1 port map( A => A(34), B => n576, ZN => n480);
   U147 : XNOR2_X1 port map( A => n575, B => n577, ZN => SUM(20));
   U148 : XNOR2_X1 port map( A => B(20), B => A(20), ZN => n577);
   U149 : NAND2_X1 port map( A1 => n517, A2 => n579, ZN => n578);
   U150 : NAND2_X1 port map( A1 => n471, A2 => A(23), ZN => n579);
   U151 : XNOR2_X1 port map( A => n547, B => n580, ZN => SUM(13));
   U152 : XOR2_X1 port map( A => A(13), B => B(13), Z => n580);
   U153 : OR2_X1 port map( A1 => B(4), A2 => A(4), ZN => n581);
   U154 : NAND2_X1 port map( A1 => n572, A2 => n527, ZN => n565);
   U155 : AND2_X1 port map( A1 => n600, A2 => n618, ZN => n582);
   U156 : NAND2_X1 port map( A1 => n563, A2 => n584, ZN => n484);
   U157 : OR2_X1 port map( A1 => n559, A2 => n628, ZN => n585);
   U158 : NAND2_X1 port map( A1 => n585, A2 => n560, ZN => n556);
   U159 : INV_X1 port map( A => n633, ZN => n586);
   U160 : XNOR2_X1 port map( A => A(29), B => n587, ZN => n500);
   U161 : AND2_X1 port map( A1 => n441, A2 => net271141, ZN => n589);
   U162 : AND2_X1 port map( A1 => n547, A2 => n635, ZN => n590);
   U163 : NOR2_X1 port map( A1 => n548, A2 => n590, ZN => n544);
   U164 : OR2_X1 port map( A1 => n497, A2 => n520, ZN => n591);
   U165 : NAND2_X1 port map( A1 => n591, A2 => n620, ZN => n504);
   U166 : AND2_X1 port map( A1 => net264281, A2 => net271140, ZN => n592);
   U168 : XNOR2_X1 port map( A => n602, B => n593, ZN => SUM(10));
   U169 : INV_X1 port map( A => n629, ZN => n595);
   U170 : INV_X1 port map( A => n635, ZN => n596);
   U171 : XNOR2_X1 port map( A => n604, B => n597, ZN => SUM(8));
   U172 : CLKBUF_X1 port map( A => A(6), Z => n598);
   U173 : XNOR2_X1 port map( A => n599, B => n506, ZN => SUM(27));
   U174 : XNOR2_X1 port map( A => A(27), B => B(27), ZN => n599);
   U175 : NAND2_X1 port map( A1 => net264281, A2 => net271140, ZN => n547);
   U176 : NAND2_X1 port map( A1 => n441, A2 => net271141, ZN => n525);
   U177 : OR2_X1 port map( A1 => n516, A2 => n521, ZN => n600);
   U178 : NAND2_X1 port map( A1 => n618, A2 => n600, ZN => n481);
   U179 : NAND2_X1 port map( A1 => n511, A2 => n601, ZN => n507);
   U180 : BUF_X1 port map( A => n487, Z => n603);
   U181 : XOR2_X1 port map( A => A(33), B => B(33), Z => n605);
   U182 : XOR2_X1 port map( A => carry_33_port, B => n605, Z => SUM(33));
   U183 : NAND2_X1 port map( A1 => carry_33_port, A2 => A(33), ZN => n606);
   U184 : NAND2_X1 port map( A1 => carry_33_port, A2 => B(33), ZN => n607);
   U185 : NAND2_X1 port map( A1 => A(33), A2 => B(33), ZN => n608);
   U186 : NAND3_X1 port map( A1 => n606, A2 => n607, A3 => n608, ZN => 
                           carry_34_port);
   U187 : OR2_X1 port map( A1 => n481, A2 => n633, ZN => n609);
   U188 : NAND2_X1 port map( A1 => n482, A2 => n609, ZN => n568);
   U189 : CLKBUF_X1 port map( A => n578, Z => n610);
   U190 : XNOR2_X1 port map( A => A(31), B => n611, ZN => n616);
   U191 : XNOR2_X1 port map( A => n516, B => n613, ZN => SUM(30));
   U192 : XNOR2_X1 port map( A => A(30), B => B(30), ZN => n613);
   U193 : XNOR2_X1 port map( A => n437, B => n614, ZN => SUM(23));
   U194 : XNOR2_X1 port map( A => A(23), B => B(23), ZN => n614);
   U195 : INV_X1 port map( A => A(25), ZN => n631);
   U196 : INV_X1 port map( A => A(5), ZN => n626);
   U197 : INV_X1 port map( A => A(29), ZN => n634);
   U198 : INV_X1 port map( A => A(22), ZN => n630);
   U199 : INV_X1 port map( A => A(13), ZN => n635);
   U200 : AOI21_X1 port map( B1 => n592, B2 => n596, A => B(13), ZN => n548);
   U201 : OAI21_X1 port map( B1 => n621, B2 => n549, A => B(25), ZN => n511);
   U202 : OAI21_X1 port map( B1 => n574, B2 => A(5), A => B(5), ZN => n566);
   U203 : XNOR2_X1 port map( A => n497, B => n615, ZN => SUM(26));
   U204 : XNOR2_X1 port map( A => B(26), B => A(26), ZN => n615);
   U205 : OAI21_X1 port map( B1 => n522, B2 => A(21), A => B(21), ZN => n523);
   U206 : XNOR2_X1 port map( A => n481, B => n616, ZN => SUM(31));
   U207 : XNOR2_X1 port map( A => net272170, B => net269617, ZN => SUM(15));
   U208 : INV_X1 port map( A => A(27), ZN => n632);
   U209 : AOI21_X1 port map( B1 => n588, B2 => A(27), A => B(27), ZN => n505);
   U210 : XNOR2_X1 port map( A => B(37), B => A(37), ZN => n491);
   U211 : AOI22_X1 port map( A1 => carry_36_port, A2 => n493, B1 => A(36), B2 
                           => B(36), ZN => n492);
   U212 : AOI22_X1 port map( A1 => B(34), A2 => A(34), B1 => n480, B2 => n438, 
                           ZN => n479);
   U213 : XNOR2_X1 port map( A => A(28), B => B(28), ZN => n503);
   U214 : INV_X1 port map( A => n479, ZN => n617);
   U215 : XNOR2_X1 port map( A => B(5), B => n626, ZN => n489);
   U216 : XNOR2_X1 port map( A => n503, B => n546, ZN => SUM(28));
   U217 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U218 : INV_X1 port map( A => A(20), ZN => n629);
   U219 : OAI21_X1 port map( B1 => n529, B2 => n454, A => B(7), ZN => n563);
   U220 : INV_X1 port map( A => A(7), ZN => n627);
   U221 : INV_X1 port map( A => n510, ZN => n621);
   U222 : OAI21_X1 port map( B1 => n448, B2 => n610, A => n622, ZN => n510);
   U223 : AOI21_X1 port map( B1 => n589, B2 => n595, A => B(20), ZN => n526);
   U224 : INV_X1 port map( A => n502, ZN => n619);
   U225 : OAI21_X1 port map( B1 => n501, B2 => A(28), A => B(28), ZN => n502);
   U226 : AOI21_X1 port map( B1 => n530, B2 => n472, A => B(29), ZN => n499);
   U227 : INV_X1 port map( A => n496, ZN => n618);
   U228 : OAI21_X1 port map( B1 => n582, B2 => n586, A => B(31), ZN => n482);
   U229 : INV_X1 port map( A => A(31), ZN => n633);
   U230 : INV_X1 port map( A => n513, ZN => n622);
   U231 : INV_X1 port map( A => A(9), ZN => n628);
   U232 : OAI21_X1 port map( B1 => n456, B2 => A(9), A => B(9), ZN => n560);
   U233 : AOI21_X1 port map( B1 => n552, B2 => n578, A => B(24), ZN => n513);
   U234 : AOI21_X1 port map( B1 => A(4), B2 => B(4), A => carry_4_port, ZN => 
                           n567);
   U235 : INV_X1 port map( A => n567, ZN => n625);
   U236 : AOI21_X1 port map( B1 => n518, B2 => n521, A => B(30), ZN => n496);
   U237 : XNOR2_X1 port map( A => n500, B => n498, ZN => SUM(29));
   U238 : INV_X1 port map( A => n508, ZN => n620);
   U239 : AOI21_X1 port map( B1 => n507, B2 => n520, A => B(26), ZN => n508);
   U240 : OAI21_X1 port map( B1 => n532, B2 => A(23), A => B(23), ZN => n517);
   U241 : INV_X1 port map( A => n557, ZN => n623);
   U242 : INV_X1 port map( A => n561, ZN => n624);
   U243 : OAI21_X1 port map( B1 => n565, B2 => n626, A => n566, ZN => n487);
   U244 : AOI21_X1 port map( B1 => n556, B2 => A(10), A => B(10), ZN => n557);
   U245 : OAI21_X1 port map( B1 => n543, B2 => n604, A => n624, ZN => n559);
   U246 : AOI21_X1 port map( B1 => n484, B2 => A(8), A => B(8), ZN => n561);
   U247 : AOI21_X1 port map( B1 => n487, B2 => A(6), A => B(6), ZN => n564);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT36_DW01_add_0 is

   port( A, B : in std_logic_vector (35 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (35 downto 0);  CO : out std_logic);

end RCA_NBIT36_DW01_add_0;

architecture SYN_rpl of RCA_NBIT36_DW01_add_0 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X2
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_33_port, n493, n494, n495, n496, n497, n498, n500, n501, n506, 
      n507, n511, n512, n513, n515, n516, n519, n520, n521, n522, n526, n530, 
      n532, n533, n534, n536, n537, n539, n540, n541, n542, n543, n545, n546, 
      n547, n548, n549, n550, n551, n552, n553, n554, n555, n557, n558, n560, 
      n561, n563, n564, n566, n567, n568, n569, n572, n573, n574, n575, n576, 
      n577, n584, n585, net272096, net278119, net274702, net273042, net271163, 
      n580, n504, n1, carry_2_port, net270702, n583, net274157, net273252, 
      net271675, net264210, n581, n446, n447, n448, n449, n450, n451, n452, 
      n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, 
      n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, 
      n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, 
      n489, n490, n491, n492, n499, n502, n503, n505, n508, n509, n510, n514, 
      n517, n518, n523, n524, n525, n527, n528, n529, n531, n535, n538, n544, 
      n556, n559, n562, n565, n570, n571, n578, n579, n582, n586, n587, n588, 
      n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, 
      n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, 
      n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, 
      n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, 
      n637, n638, n_1030 : std_logic;

begin
   
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => n584, CO => n_1030, S 
                           => SUM(35));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => n585, CO => 
                           carry_33_port, S => SUM(32));
   U123 : XOR2_X1 port map( A => B(9), B => A(9), Z => n497);
   U127 : XOR2_X1 port map( A => B(7), B => A(7), Z => n500);
   U134 : XOR2_X1 port map( A => net272096, B => n506, Z => SUM(3));
   U135 : XOR2_X1 port map( A => n494, B => n493, Z => SUM(34));
   U136 : XOR2_X1 port map( A => n627, B => B(34), Z => n494);
   U138 : XOR2_X1 port map( A => A(33), B => B(33), Z => n507);
   U140 : XOR2_X1 port map( A => n626, B => B(31), Z => n496);
   U141 : XOR2_X1 port map( A => net278119, B => n513, Z => SUM(2));
   U148 : XOR2_X1 port map( A => B(27), B => A(27), Z => n520);
   U152 : XOR2_X1 port map( A => B(25), B => A(25), Z => n526);
   U156 : XOR2_X1 port map( A => B(23), B => A(23), Z => n532);
   U157 : XOR2_X1 port map( A => n598, B => n534, Z => SUM(22));
   U158 : XOR2_X1 port map( A => B(22), B => A(22), Z => n534);
   U162 : XOR2_X1 port map( A => B(20), B => A(20), Z => n541);
   U166 : XOR2_X1 port map( A => B(18), B => A(18), Z => n547);
   U167 : XOR2_X1 port map( A => n508, B => n550, Z => SUM(17));
   U168 : XOR2_X1 port map( A => B(17), B => A(17), Z => n550);
   U169 : XOR2_X1 port map( A => n528, B => n553, Z => SUM(16));
   U171 : XOR2_X1 port map( A => B(11), B => A(11), Z => n568);
   U174 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U142 : XOR2_X1 port map( A => carry_2_port, B => n471, Z => n513);
   U1 : AOI21_X1 port map( B1 => n535, B2 => A(10), A => B(10), ZN => n446);
   U2 : INV_X1 port map( A => A(24), ZN => n463);
   U3 : INV_X1 port map( A => B(24), ZN => n464);
   U4 : OR2_X1 port map( A1 => n600, A2 => A(22), ZN => n533);
   U5 : INV_X1 port map( A => B(30), ZN => n492);
   U6 : XNOR2_X1 port map( A => B(26), B => A(26), ZN => n447);
   U7 : OR2_X1 port map( A1 => n590, A2 => n619, ZN => n448);
   U8 : AOI21_X1 port map( B1 => n483, B2 => A(25), A => B(25), ZN => n449);
   U9 : OAI21_X1 port map( B1 => n563, B2 => A(12), A => B(12), ZN => n450);
   U10 : NAND2_X1 port map( A1 => n454, A2 => n452, ZN => n451);
   U11 : AND2_X2 port map( A1 => n566, A2 => n637, ZN => n611);
   U12 : OAI21_X1 port map( B1 => n562, B2 => A(9), A => B(9), ZN => n452);
   U13 : NOR2_X1 port map( A1 => n449, A2 => n529, ZN => n453);
   U14 : CLKBUF_X1 port map( A => n542, Z => n486);
   U15 : OR2_X1 port map( A1 => n572, A2 => n638, ZN => n454);
   U16 : OR2_X1 port map( A1 => n572, A2 => n638, ZN => n518);
   U17 : OR2_X1 port map( A1 => n574, A2 => n589, ZN => n572);
   U18 : INV_X1 port map( A => n577, ZN => n455);
   U19 : OR2_X1 port map( A1 => n501, A2 => A(6), ZN => n595);
   U20 : AND2_X1 port map( A1 => n478, A2 => n558, ZN => n456);
   U21 : AND2_X1 port map( A1 => n478, A2 => n558, ZN => n588);
   U22 : AND2_X1 port map( A1 => n564, A2 => n457, ZN => n616);
   U23 : AND2_X1 port map( A1 => n594, A2 => n636, ZN => n457);
   U24 : INV_X1 port map( A => n507, ZN => n479);
   U25 : OR2_X1 port map( A1 => B(5), A2 => A(5), ZN => n459);
   U26 : NAND2_X1 port map( A1 => n460, A2 => n459, ZN => n458);
   U27 : NOR2_X1 port map( A1 => n580, A2 => net271163, ZN => n460);
   U28 : NOR2_X1 port map( A1 => n519, A2 => n593, ZN => n515);
   U29 : OR2_X2 port map( A1 => n468, A2 => n604, ZN => n566);
   U30 : OR2_X1 port map( A1 => n456, A2 => n477, ZN => n461);
   U31 : AOI21_X1 port map( B1 => n465, B2 => n463, A => n464, ZN => n462);
   U32 : OR2_X1 port map( A1 => n485, A2 => n608, ZN => n465);
   U33 : INV_X1 port map( A => A(30), ZN => n491);
   U34 : INV_X1 port map( A => n496, ZN => n606);
   U35 : XNOR2_X2 port map( A => n554, B => n614, ZN => SUM(15));
   U36 : NOR2_X1 port map( A1 => n616, A2 => n561, ZN => n557);
   U37 : XNOR2_X1 port map( A => net274157, B => net273252, ZN => SUM(4));
   U38 : OAI21_X1 port map( B1 => n581, B2 => net264210, A => n466, ZN => 
                           net273252);
   U39 : INV_X1 port map( A => A(3), ZN => net264210);
   U40 : OAI21_X1 port map( B1 => n581, B2 => net264210, A => n466, ZN => n504)
                           ;
   U41 : XNOR2_X1 port map( A => B(3), B => net264210, ZN => n506);
   U42 : XNOR2_X1 port map( A => A(4), B => B(4), ZN => net274157);
   U43 : OR2_X1 port map( A1 => net270702, A2 => n583, ZN => n581);
   U44 : INV_X1 port map( A => n581, ZN => net272096);
   U45 : OAI21_X1 port map( B1 => net271675, B2 => A(3), A => B(3), ZN => n466)
                           ;
   U46 : NOR2_X1 port map( A1 => net270702, A2 => n583, ZN => net271675);
   U47 : CLKBUF_X1 port map( A => A(4), Z => net274702);
   U48 : CLKBUF_X1 port map( A => B(4), Z => net273042);
   U49 : NOR2_X1 port map( A1 => n480, A2 => A(10), ZN => n467);
   U50 : AOI21_X1 port map( B1 => n535, B2 => A(10), A => B(10), ZN => n468);
   U51 : XNOR2_X1 port map( A => n515, B => n469, ZN => SUM(28));
   U52 : XNOR2_X1 port map( A => B(28), B => A(28), ZN => n469);
   U53 : AOI21_X1 port map( B1 => n499, B2 => n491, A => n492, ZN => n470);
   U54 : NOR2_X1 port map( A1 => B(2), A2 => A(2), ZN => net270702);
   U55 : AOI21_X1 port map( B1 => B(2), B2 => A(2), A => carry_2_port, ZN => 
                           n583);
   U56 : CLKBUF_X1 port map( A => B(2), Z => n471);
   U57 : CLKBUF_X1 port map( A => A(2), Z => net278119);
   U58 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U59 : NAND2_X1 port map( A1 => n458, A2 => n474, ZN => n472);
   U60 : NAND2_X1 port map( A1 => n623, A2 => n473, ZN => n556);
   U61 : AND2_X1 port map( A1 => n559, A2 => A(18), ZN => n473);
   U62 : XNOR2_X1 port map( A => A(5), B => B(5), ZN => n476);
   U63 : NAND2_X1 port map( A1 => A(5), A2 => B(5), ZN => n474);
   U64 : NOR2_X1 port map( A1 => net271163, A2 => n580, ZN => n475);
   U65 : XNOR2_X1 port map( A => n475, B => n476, ZN => SUM(5));
   U66 : NAND2_X1 port map( A1 => n458, A2 => n474, ZN => n501);
   U67 : AOI21_X1 port map( B1 => n504, B2 => net274702, A => net273042, ZN => 
                           n580);
   U68 : NOR2_X1 port map( A1 => net274702, A2 => n504, ZN => net271163);
   U69 : AOI21_X1 port map( B1 => n579, B2 => A(15), A => B(15), ZN => n477);
   U70 : AND2_X1 port map( A1 => n596, A2 => n635, ZN => n478);
   U71 : XNOR2_X1 port map( A => carry_33_port, B => n479, ZN => SUM(33));
   U72 : NAND2_X1 port map( A1 => n454, A2 => n452, ZN => n480);
   U73 : XNOR2_X1 port map( A => n488, B => n481, ZN => SUM(24));
   U74 : XNOR2_X1 port map( A => B(24), B => A(24), ZN => n481);
   U75 : AND2_X1 port map( A1 => n622, A2 => n587, ZN => n482);
   U76 : OR2_X1 port map( A1 => n578, A2 => n462, ZN => n483);
   U77 : AND2_X1 port map( A1 => n450, A2 => n594, ZN => n560);
   U78 : NAND2_X1 port map( A1 => n564, A2 => n594, ZN => n484);
   U79 : AOI21_X1 port map( B1 => n620, B2 => A(23), A => B(23), ZN => n485);
   U80 : CLKBUF_X1 port map( A => n536, Z => n514);
   U81 : XNOR2_X1 port map( A => n525, B => n532, ZN => SUM(23));
   U82 : XNOR2_X1 port map( A => n514, B => n487, ZN => SUM(21));
   U83 : XNOR2_X1 port map( A => B(21), B => A(21), ZN => n487);
   U84 : NOR2_X1 port map( A1 => n485, A2 => n608, ZN => n488);
   U85 : CLKBUF_X1 port map( A => n595, Z => n489);
   U86 : AOI21_X2 port map( B1 => n597, B2 => A(11), A => B(11), ZN => n567);
   U87 : AOI21_X1 port map( B1 => n499, B2 => n491, A => n492, ZN => n490);
   U88 : OR2_X1 port map( A1 => n607, A2 => n512, ZN => n499);
   U89 : NOR2_X1 port map( A1 => n578, A2 => n462, ZN => n502);
   U90 : NOR2_X1 port map( A1 => n512, A2 => n607, ZN => n503);
   U91 : OAI21_X1 port map( B1 => A(9), B2 => n562, A => B(9), ZN => n505);
   U92 : CLKBUF_X1 port map( A => n548, Z => n508);
   U93 : XNOR2_X1 port map( A => n501, B => n509, ZN => SUM(6));
   U94 : XNOR2_X1 port map( A => B(6), B => A(6), ZN => n509);
   U95 : AND2_X1 port map( A1 => n623, A2 => n559, ZN => n510);
   U96 : NOR2_X1 port map( A1 => n619, A2 => n590, ZN => n517);
   U97 : XNOR2_X1 port map( A => n569, B => n523, ZN => SUM(10));
   U98 : XNOR2_X1 port map( A => B(10), B => A(10), ZN => n523);
   U99 : OAI21_X1 port map( B1 => n557, B2 => A(14), A => B(14), ZN => n524);
   U100 : AOI22_X1 port map( A1 => n602, A2 => A(22), B1 => n533, B2 => B(22), 
                           ZN => n525);
   U101 : OR2_X1 port map( A1 => n539, A2 => n633, ZN => n527);
   U102 : NAND2_X1 port map( A1 => n527, A2 => n540, ZN => n536);
   U103 : NOR2_X1 port map( A1 => n456, A2 => n477, ZN => n528);
   U104 : AND2_X1 port map( A1 => n502, A2 => n631, ZN => n529);
   U105 : NOR2_X1 port map( A1 => n449, A2 => n529, ZN => n521);
   U106 : AOI21_X1 port map( B1 => n484, B2 => A(13), A => B(13), ZN => n531);
   U107 : NAND2_X1 port map( A1 => n518, A2 => n573, ZN => n535);
   U108 : NOR2_X1 port map( A1 => n611, A2 => n567, ZN => n538);
   U109 : NOR2_X1 port map( A1 => n567, A2 => n611, ZN => n544);
   U110 : NAND2_X1 port map( A1 => n546, A2 => n556, ZN => n542);
   U111 : OR2_X1 port map( A1 => A(17), A2 => n548, ZN => n559);
   U112 : NAND2_X1 port map( A1 => n623, A2 => n559, ZN => n545);
   U113 : NOR2_X1 port map( A1 => n611, A2 => n567, ZN => n563);
   U114 : NOR2_X1 port map( A1 => n589, A2 => n574, ZN => n562);
   U115 : NAND2_X1 port map( A1 => n489, A2 => n565, ZN => n613);
   U116 : AND2_X1 port map( A1 => n624, A2 => A(7), ZN => n565);
   U117 : AND2_X1 port map( A1 => n612, A2 => n618, ZN => n570);
   U118 : NOR2_X1 port map( A1 => n586, A2 => n470, ZN => n571);
   U119 : NAND2_X1 port map( A1 => n454, A2 => n505, ZN => n569);
   U120 : AND2_X1 port map( A1 => n596, A2 => n558, ZN => n554);
   U121 : AND2_X1 port map( A1 => n488, A2 => A(24), ZN => n578);
   U122 : BUF_X1 port map( A => n598, Z => n602);
   U124 : NAND2_X1 port map( A1 => n596, A2 => n524, ZN => n579);
   U125 : AND2_X1 port map( A1 => n455, A2 => n595, ZN => n582);
   U126 : AOI21_X1 port map( B1 => n484, B2 => A(13), A => B(13), ZN => n561);
   U128 : XNOR2_X1 port map( A => n517, B => n520, ZN => SUM(27));
   U129 : AND2_X1 port map( A1 => n503, A2 => A(30), ZN => n586);
   U130 : NOR2_X1 port map( A1 => n586, A2 => n490, ZN => n495);
   U131 : OR2_X1 port map( A1 => A(19), A2 => n542, ZN => n587);
   U132 : NAND2_X1 port map( A1 => n622, A2 => n587, ZN => n539);
   U133 : NOR2_X1 port map( A1 => n588, A2 => n555, ZN => n552);
   U137 : NOR2_X1 port map( A1 => n498, A2 => A(8), ZN => n589);
   U139 : AND2_X1 port map( A1 => n453, A2 => A(26), ZN => n590);
   U143 : NOR2_X1 port map( A1 => n531, A2 => n616, ZN => n591);
   U144 : NOR2_X1 port map( A1 => n616, A2 => n531, ZN => n592);
   U145 : AND2_X1 port map( A1 => n630, A2 => n517, ZN => n593);
   U146 : NAND2_X1 port map( A1 => n538, A2 => A(12), ZN => n594);
   U147 : NAND2_X1 port map( A1 => n624, A2 => n595, ZN => n575);
   U149 : NAND2_X1 port map( A1 => n591, A2 => A(14), ZN => n596);
   U150 : NOR2_X1 port map( A1 => n446, A2 => n467, ZN => n597);
   U151 : AND2_X1 port map( A1 => n621, A2 => n603, ZN => n598);
   U153 : XNOR2_X1 port map( A => n498, B => n599, ZN => SUM(8));
   U154 : XNOR2_X1 port map( A => B(8), B => A(8), ZN => n599);
   U155 : AND2_X1 port map( A1 => n621, A2 => n603, ZN => n600);
   U159 : XNOR2_X1 port map( A => n486, B => n601, ZN => SUM(19));
   U160 : XNOR2_X1 port map( A => B(19), B => A(19), ZN => n601);
   U161 : OR2_X1 port map( A1 => A(21), A2 => n536, ZN => n603);
   U163 : NOR2_X1 port map( A1 => n451, A2 => A(10), ZN => n604);
   U164 : XNOR2_X1 port map( A => n511, B => n605, ZN => SUM(29));
   U165 : XNOR2_X1 port map( A => n629, B => B(29), ZN => n605);
   U170 : XNOR2_X1 port map( A => n495, B => n606, ZN => SUM(31));
   U172 : XNOR2_X1 port map( A => n545, B => n547, ZN => SUM(18));
   U173 : AND2_X1 port map( A1 => n629, A2 => n511, ZN => n607);
   U175 : AND2_X1 port map( A1 => n525, A2 => n632, ZN => n608);
   U176 : XNOR2_X1 port map( A => n503, B => n609, ZN => SUM(30));
   U177 : XNOR2_X1 port map( A => A(30), B => B(30), ZN => n609);
   U178 : XNOR2_X1 port map( A => n453, B => n447, ZN => SUM(26));
   U179 : XNOR2_X1 port map( A => n544, B => n610, ZN => SUM(12));
   U180 : XNOR2_X1 port map( A => A(12), B => B(12), ZN => n610);
   U181 : XNOR2_X1 port map( A => n539, B => n541, ZN => SUM(20));
   U182 : XNOR2_X1 port map( A => n575, B => n500, ZN => SUM(7));
   U183 : OR2_X1 port map( A1 => A(28), A2 => n515, ZN => n612);
   U184 : NAND2_X1 port map( A1 => n612, A2 => n618, ZN => n511);
   U185 : XNOR2_X1 port map( A => n566, B => n568, ZN => SUM(11));
   U186 : NAND2_X1 port map( A1 => n613, A2 => n576, ZN => n498);
   U187 : XNOR2_X1 port map( A => B(15), B => n635, ZN => n614);
   U188 : XNOR2_X1 port map( A => n560, B => n615, ZN => SUM(13));
   U189 : XNOR2_X1 port map( A => B(13), B => n636, ZN => n615);
   U190 : XNOR2_X1 port map( A => n502, B => n526, ZN => SUM(25));
   U191 : XNOR2_X1 port map( A => n572, B => n497, ZN => SUM(9));
   U192 : INV_X1 port map( A => A(11), ZN => n637);
   U193 : XOR2_X1 port map( A => n592, B => n617, Z => SUM(14));
   U194 : XOR2_X1 port map( A => A(14), B => B(14), Z => n617);
   U195 : XNOR2_X1 port map( A => B(16), B => n634, ZN => n553);
   U196 : INV_X1 port map( A => A(25), ZN => n631);
   U197 : INV_X1 port map( A => A(23), ZN => n632);
   U198 : INV_X1 port map( A => A(27), ZN => n630);
   U199 : INV_X1 port map( A => A(20), ZN => n633);
   U200 : INV_X1 port map( A => A(9), ZN => n638);
   U201 : AOI22_X1 port map( A1 => B(33), A2 => A(33), B1 => n507, B2 => 
                           carry_33_port, ZN => n493);
   U202 : OAI22_X1 port map( A1 => n628, A2 => n626, B1 => n571, B2 => n496, ZN
                           => n585);
   U203 : INV_X1 port map( A => A(13), ZN => n636);
   U204 : INV_X1 port map( A => A(15), ZN => n635);
   U205 : INV_X1 port map( A => A(16), ZN => n634);
   U206 : INV_X1 port map( A => A(34), ZN => n627);
   U207 : INV_X1 port map( A => B(31), ZN => n628);
   U208 : INV_X1 port map( A => A(29), ZN => n629);
   U209 : INV_X1 port map( A => B(34), ZN => n625);
   U210 : OAI22_X1 port map( A1 => n625, A2 => n627, B1 => n493, B2 => n494, ZN
                           => n584);
   U211 : INV_X1 port map( A => A(31), ZN => n626);
   U212 : AOI21_X1 port map( B1 => n448, B2 => A(27), A => B(27), ZN => n519);
   U213 : INV_X1 port map( A => n549, ZN => n623);
   U214 : AOI21_X1 port map( B1 => n548, B2 => A(17), A => B(17), ZN => n549);
   U215 : AOI22_X1 port map( A1 => n602, A2 => A(22), B1 => n533, B2 => B(22), 
                           ZN => n530);
   U216 : OAI21_X1 port map( B1 => n521, B2 => A(26), A => B(26), ZN => n522);
   U217 : INV_X1 port map( A => n516, ZN => n618);
   U218 : OAI21_X1 port map( B1 => n482, B2 => A(20), A => B(20), ZN => n540);
   U219 : AOI21_X1 port map( B1 => n515, B2 => A(28), A => B(28), ZN => n516);
   U220 : OAI21_X1 port map( B1 => n557, B2 => A(14), A => B(14), ZN => n558);
   U221 : OAI21_X1 port map( B1 => n510, B2 => A(18), A => B(18), ZN => n546);
   U222 : INV_X1 port map( A => n522, ZN => n619);
   U223 : AOI21_X1 port map( B1 => n570, B2 => A(29), A => B(29), ZN => n512);
   U224 : AOI21_X1 port map( B1 => n498, B2 => A(8), A => B(8), ZN => n574);
   U225 : INV_X1 port map( A => n530, ZN => n620);
   U226 : INV_X1 port map( A => n543, ZN => n622);
   U227 : OAI21_X1 port map( B1 => n461, B2 => n634, A => n551, ZN => n548);
   U228 : INV_X1 port map( A => n577, ZN => n624);
   U229 : AOI21_X1 port map( B1 => n472, B2 => A(6), A => B(6), ZN => n577);
   U230 : OAI21_X1 port map( B1 => n562, B2 => A(9), A => B(9), ZN => n573);
   U231 : INV_X1 port map( A => n537, ZN => n621);
   U232 : AOI21_X1 port map( B1 => n536, B2 => A(21), A => B(21), ZN => n537);
   U233 : AOI21_X1 port map( B1 => n542, B2 => A(19), A => B(19), ZN => n543);
   U234 : OAI21_X1 port map( B1 => n552, B2 => A(16), A => B(16), ZN => n551);
   U235 : AOI21_X1 port map( B1 => n579, B2 => A(15), A => B(15), ZN => n555);
   U236 : OAI21_X1 port map( B1 => n563, B2 => A(12), A => B(12), ZN => n564);
   U237 : OAI21_X1 port map( B1 => n582, B2 => A(7), A => B(7), ZN => n576);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHMUL_NBIT32_DW01_sub_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end BOOTHMUL_NBIT32_DW01_sub_0;

architecture SYN_rpl of BOOTHMUL_NBIT32_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n96, n97, n98, n99, n100, n102, n103, n104, n106, n107, n108, n110, 
      n111, n112, n114, n115, n116, n118, n119, n120, n122, n123, n124, n95, 
      n101, n105, n109, n113, n117, n121, n125 : std_logic;

begin
   DIFF <= ( DIFF(31), DIFF(30), DIFF(29), DIFF(28), DIFF(27), DIFF(26), 
      DIFF(25), DIFF(24), DIFF(23), DIFF(22), DIFF(21), DIFF(20), DIFF(19), 
      DIFF(18), DIFF(17), DIFF(16), DIFF(15), DIFF(14), DIFF(13), DIFF(12), 
      DIFF(11), DIFF(10), DIFF(9), DIFF(8), DIFF(7), DIFF(6), DIFF(5), DIFF(4),
      DIFF(3), DIFF(2), DIFF(1), DIFF(0) );
   
   U42 : XOR2_X1 port map( A => n96, B => B(30), Z => DIFF(30));
   U43 : XOR2_X1 port map( A => n98, B => B(27), Z => DIFF(27));
   U45 : XOR2_X1 port map( A => n100, B => B(25), Z => DIFF(25));
   U46 : XOR2_X1 port map( A => n102, B => B(23), Z => DIFF(23));
   U48 : XOR2_X1 port map( A => n104, B => B(21), Z => DIFF(21));
   U49 : XOR2_X1 port map( A => n106, B => B(19), Z => DIFF(19));
   U51 : XOR2_X1 port map( A => n108, B => B(17), Z => DIFF(17));
   U52 : XOR2_X1 port map( A => n110, B => B(15), Z => DIFF(15));
   U54 : XOR2_X1 port map( A => n112, B => B(13), Z => DIFF(13));
   U55 : XOR2_X1 port map( A => n114, B => B(11), Z => DIFF(11));
   U57 : XOR2_X1 port map( A => n116, B => B(9), Z => DIFF(9));
   U58 : XOR2_X1 port map( A => n118, B => B(7), Z => DIFF(7));
   U60 : XOR2_X1 port map( A => n120, B => B(5), Z => DIFF(5));
   U61 : XOR2_X1 port map( A => n122, B => B(3), Z => DIFF(3));
   U62 : XOR2_X1 port map( A => B(0), B => B(1), Z => DIFF(1));
   U1 : BUF_X1 port map( A => B(0), Z => DIFF(0));
   U2 : XNOR2_X1 port map( A => n124, B => B(2), ZN => DIFF(2));
   U3 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n124);
   U4 : OR3_X2 port map( A1 => B(0), A2 => B(2), A3 => B(1), ZN => n122);
   U5 : XOR2_X1 port map( A => n95, B => B(31), Z => DIFF(31));
   U6 : OR2_X1 port map( A1 => n96, A2 => B(30), ZN => n95);
   U7 : NAND2_X1 port map( A1 => n97, A2 => n125, ZN => n96);
   U8 : XOR2_X1 port map( A => n97, B => n125, Z => DIFF(29));
   U9 : XNOR2_X1 port map( A => n101, B => B(6), ZN => DIFF(6));
   U10 : NOR2_X1 port map( A1 => n120, A2 => B(5), ZN => n101);
   U11 : XNOR2_X1 port map( A => n105, B => B(14), ZN => DIFF(14));
   U12 : NOR2_X1 port map( A1 => n112, A2 => B(13), ZN => n105);
   U13 : XNOR2_X1 port map( A => n109, B => B(18), ZN => DIFF(18));
   U14 : NOR2_X1 port map( A1 => n108, A2 => B(17), ZN => n109);
   U15 : XNOR2_X1 port map( A => n113, B => B(10), ZN => DIFF(10));
   U16 : NOR2_X1 port map( A1 => n116, A2 => B(9), ZN => n113);
   U17 : XNOR2_X1 port map( A => B(8), B => n119, ZN => DIFF(8));
   U18 : NOR2_X1 port map( A1 => B(7), A2 => n118, ZN => n119);
   U19 : XNOR2_X1 port map( A => B(4), B => n123, ZN => DIFF(4));
   U20 : NOR2_X1 port map( A1 => B(3), A2 => n122, ZN => n123);
   U21 : XNOR2_X1 port map( A => B(12), B => n115, ZN => DIFF(12));
   U22 : NOR2_X1 port map( A1 => B(11), A2 => n114, ZN => n115);
   U23 : XNOR2_X1 port map( A => B(16), B => n111, ZN => DIFF(16));
   U24 : NOR2_X1 port map( A1 => B(15), A2 => n110, ZN => n111);
   U25 : OR3_X1 port map( A1 => B(17), A2 => B(18), A3 => n108, ZN => n106);
   U26 : OR3_X1 port map( A1 => B(13), A2 => B(14), A3 => n112, ZN => n110);
   U27 : OR3_X1 port map( A1 => B(5), A2 => B(6), A3 => n120, ZN => n118);
   U28 : OR3_X1 port map( A1 => B(10), A2 => B(9), A3 => n116, ZN => n114);
   U29 : OR3_X1 port map( A1 => B(15), A2 => B(16), A3 => n110, ZN => n108);
   U30 : OR3_X1 port map( A1 => n122, A2 => B(4), A3 => B(3), ZN => n120);
   U31 : OR3_X1 port map( A1 => B(11), A2 => B(12), A3 => n114, ZN => n112);
   U32 : OR3_X1 port map( A1 => B(7), A2 => B(8), A3 => n118, ZN => n116);
   U33 : NOR3_X1 port map( A1 => B(27), A2 => B(28), A3 => n98, ZN => n97);
   U34 : XNOR2_X1 port map( A => n117, B => B(22), ZN => DIFF(22));
   U35 : NOR2_X1 port map( A1 => n104, A2 => B(21), ZN => n117);
   U36 : XNOR2_X1 port map( A => n121, B => B(26), ZN => DIFF(26));
   U37 : NOR2_X1 port map( A1 => n100, A2 => B(25), ZN => n121);
   U38 : XNOR2_X1 port map( A => B(24), B => n103, ZN => DIFF(24));
   U39 : NOR2_X1 port map( A1 => B(23), A2 => n102, ZN => n103);
   U40 : XNOR2_X1 port map( A => B(20), B => n107, ZN => DIFF(20));
   U41 : NOR2_X1 port map( A1 => B(19), A2 => n106, ZN => n107);
   U44 : XNOR2_X1 port map( A => B(28), B => n99, ZN => DIFF(28));
   U47 : NOR2_X1 port map( A1 => B(27), A2 => n98, ZN => n99);
   U50 : OR3_X1 port map( A1 => B(25), A2 => B(26), A3 => n100, ZN => n98);
   U53 : OR3_X1 port map( A1 => B(21), A2 => B(22), A3 => n104, ZN => n102);
   U56 : OR3_X1 port map( A1 => B(23), A2 => B(24), A3 => n102, ZN => n100);
   U59 : OR3_X1 port map( A1 => B(19), A2 => B(20), A3 => n106, ZN => n104);
   U63 : INV_X1 port map( A => B(29), ZN => n125);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT64 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64;

architecture SYN_DIRECT of RCA_NBIT64 is

   component RCA_NBIT64_DW01_add_0
      port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (63 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1065 : std_logic;

begin
   
   Co <= '0';
   n1 <= '0';
   add_95 : RCA_NBIT64_DW01_add_0 port map( A(63) => A(63), A(62) => A(62), 
                           A(61) => A(61), A(60) => A(60), A(59) => A(59), 
                           A(58) => A(58), A(57) => A(57), A(56) => A(56), 
                           A(55) => A(55), A(54) => A(54), A(53) => A(53), 
                           A(52) => A(52), A(51) => A(51), A(50) => A(50), 
                           A(49) => A(49), A(48) => A(48), A(47) => A(47), 
                           A(46) => A(46), A(45) => A(45), A(44) => A(44), 
                           A(43) => A(43), A(42) => A(42), A(41) => A(41), 
                           A(40) => A(40), A(39) => A(39), A(38) => A(38), 
                           A(37) => A(37), A(36) => A(36), A(35) => A(35), 
                           A(34) => A(34), A(33) => A(33), A(32) => A(32), 
                           A(31) => A(31), A(30) => A(30), A(29) => A(29), 
                           A(28) => A(28), A(27) => A(27), A(26) => A(26), 
                           A(25) => A(25), A(24) => A(24), A(23) => A(23), 
                           A(22) => A(22), A(21) => A(21), A(20) => A(20), 
                           A(19) => A(19), A(18) => A(18), A(17) => A(17), 
                           A(16) => A(16), A(15) => A(15), A(14) => A(14), 
                           A(13) => A(13), A(12) => A(12), A(11) => A(11), 
                           A(10) => A(10), A(9) => A(9), A(8) => A(8), A(7) => 
                           A(7), A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3)
                           => A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(63) => B(63), B(62) => B(62), B(61) => B(61), 
                           B(60) => B(60), B(59) => B(59), B(58) => B(58), 
                           B(57) => B(57), B(56) => B(56), B(55) => B(55), 
                           B(54) => B(54), B(53) => B(53), B(52) => B(52), 
                           B(51) => B(51), B(50) => B(50), B(49) => B(49), 
                           B(48) => B(48), B(47) => B(47), B(46) => B(46), 
                           B(45) => B(45), B(44) => B(44), B(43) => B(43), 
                           B(42) => B(42), B(41) => B(41), B(40) => B(40), 
                           B(39) => B(39), B(38) => B(38), B(37) => B(37), 
                           B(36) => B(36), B(35) => B(35), B(34) => B(34), 
                           B(33) => B(33), B(32) => B(32), B(31) => B(31), 
                           B(30) => B(30), B(29) => B(29), B(28) => B(28), 
                           B(27) => B(27), B(26) => B(26), B(25) => B(25), 
                           B(24) => B(24), B(23) => B(23), B(22) => B(22), 
                           B(21) => B(21), B(20) => B(20), B(19) => B(19), 
                           B(18) => B(18), B(17) => B(17), B(16) => B(16), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => B(0), CI => n1, SUM(63) 
                           => S(63), SUM(62) => S(62), SUM(61) => S(61), 
                           SUM(60) => S(60), SUM(59) => S(59), SUM(58) => S(58)
                           , SUM(57) => S(57), SUM(56) => S(56), SUM(55) => 
                           S(55), SUM(54) => S(54), SUM(53) => S(53), SUM(52) 
                           => S(52), SUM(51) => S(51), SUM(50) => S(50), 
                           SUM(49) => S(49), SUM(48) => S(48), SUM(47) => S(47)
                           , SUM(46) => S(46), SUM(45) => S(45), SUM(44) => 
                           S(44), SUM(43) => S(43), SUM(42) => S(42), SUM(41) 
                           => S(41), SUM(40) => S(40), SUM(39) => S(39), 
                           SUM(38) => S(38), SUM(37) => S(37), SUM(36) => S(36)
                           , SUM(35) => S(35), SUM(34) => S(34), SUM(33) => 
                           S(33), SUM(32) => S(32), SUM(31) => S(31), SUM(30) 
                           => S(30), SUM(29) => S(29), SUM(28) => S(28), 
                           SUM(27) => S(27), SUM(26) => S(26), SUM(25) => S(25)
                           , SUM(24) => S(24), SUM(23) => S(23), SUM(22) => 
                           S(22), SUM(21) => S(21), SUM(20) => S(20), SUM(19) 
                           => S(19), SUM(18) => S(18), SUM(17) => S(17), 
                           SUM(16) => S(16), SUM(15) => S(15), SUM(14) => S(14)
                           , SUM(13) => S(13), SUM(12) => S(12), SUM(11) => 
                           S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) => 
                           S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5)
                           , SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1065);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT62 is

   port( A, B : in std_logic_vector (61 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (61 downto 0);  Co : out std_logic);

end RCA_NBIT62;

architecture SYN_DIRECT of RCA_NBIT62 is

   component RCA_NBIT62_DW01_add_0
      port( A, B : in std_logic_vector (61 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (61 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1066 : std_logic;

begin
   
   Co <= '0';
   n1 <= '0';
   add_95 : RCA_NBIT62_DW01_add_0 port map( A(61) => A(61), A(60) => A(60), 
                           A(59) => A(59), A(58) => A(58), A(57) => A(57), 
                           A(56) => A(56), A(55) => A(55), A(54) => A(54), 
                           A(53) => A(53), A(52) => A(52), A(51) => A(51), 
                           A(50) => A(50), A(49) => A(49), A(48) => A(48), 
                           A(47) => A(47), A(46) => A(46), A(45) => A(45), 
                           A(44) => A(44), A(43) => A(43), A(42) => A(42), 
                           A(41) => A(41), A(40) => A(40), A(39) => A(39), 
                           A(38) => A(38), A(37) => A(37), A(36) => A(36), 
                           A(35) => A(35), A(34) => A(34), A(33) => A(33), 
                           A(32) => A(32), A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(61) => B(61), B(60) => B(60), 
                           B(59) => B(59), B(58) => B(58), B(57) => B(57), 
                           B(56) => B(56), B(55) => B(55), B(54) => B(54), 
                           B(53) => B(53), B(52) => B(52), B(51) => B(51), 
                           B(50) => B(50), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => n1, SUM(61) => S(61), 
                           SUM(60) => S(60), SUM(59) => S(59), SUM(58) => S(58)
                           , SUM(57) => S(57), SUM(56) => S(56), SUM(55) => 
                           S(55), SUM(54) => S(54), SUM(53) => S(53), SUM(52) 
                           => S(52), SUM(51) => S(51), SUM(50) => S(50), 
                           SUM(49) => S(49), SUM(48) => S(48), SUM(47) => S(47)
                           , SUM(46) => S(46), SUM(45) => S(45), SUM(44) => 
                           S(44), SUM(43) => S(43), SUM(42) => S(42), SUM(41) 
                           => S(41), SUM(40) => S(40), SUM(39) => S(39), 
                           SUM(38) => S(38), SUM(37) => S(37), SUM(36) => S(36)
                           , SUM(35) => S(35), SUM(34) => S(34), SUM(33) => 
                           S(33), SUM(32) => S(32), SUM(31) => S(31), SUM(30) 
                           => S(30), SUM(29) => S(29), SUM(28) => S(28), 
                           SUM(27) => S(27), SUM(26) => S(26), SUM(25) => S(25)
                           , SUM(24) => S(24), SUM(23) => S(23), SUM(22) => 
                           S(22), SUM(21) => S(21), SUM(20) => S(20), SUM(19) 
                           => S(19), SUM(18) => S(18), SUM(17) => S(17), 
                           SUM(16) => S(16), SUM(15) => S(15), SUM(14) => S(14)
                           , SUM(13) => S(13), SUM(12) => S(12), SUM(11) => 
                           S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) => 
                           S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5)
                           , SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1066);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT60 is

   port( A, B : in std_logic_vector (59 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (59 downto 0);  Co : out std_logic);

end RCA_NBIT60;

architecture SYN_DIRECT of RCA_NBIT60 is

   component RCA_NBIT60_DW01_add_0
      port( A, B : in std_logic_vector (59 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (59 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1067 : std_logic;

begin
   
   Co <= '0';
   n1 <= '0';
   add_95 : RCA_NBIT60_DW01_add_0 port map( A(59) => A(59), A(58) => A(58), 
                           A(57) => A(57), A(56) => A(56), A(55) => A(55), 
                           A(54) => A(54), A(53) => A(53), A(52) => A(52), 
                           A(51) => A(51), A(50) => A(50), A(49) => A(49), 
                           A(48) => A(48), A(47) => A(47), A(46) => A(46), 
                           A(45) => A(45), A(44) => A(44), A(43) => A(43), 
                           A(42) => A(42), A(41) => A(41), A(40) => A(40), 
                           A(39) => A(39), A(38) => A(38), A(37) => A(37), 
                           A(36) => A(36), A(35) => A(35), A(34) => A(34), 
                           A(33) => A(33), A(32) => A(32), A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(59) => B(59), 
                           B(58) => B(58), B(57) => B(57), B(56) => B(56), 
                           B(55) => B(55), B(54) => B(54), B(53) => B(53), 
                           B(52) => B(52), B(51) => B(51), B(50) => B(50), 
                           B(49) => B(49), B(48) => B(48), B(47) => B(47), 
                           B(46) => B(46), B(45) => B(45), B(44) => B(44), 
                           B(43) => B(43), B(42) => B(42), B(41) => B(41), 
                           B(40) => B(40), B(39) => B(39), B(38) => B(38), 
                           B(37) => B(37), B(36) => B(36), B(35) => B(35), 
                           B(34) => B(34), B(33) => B(33), B(32) => B(32), 
                           B(31) => B(31), B(30) => B(30), B(29) => B(29), 
                           B(28) => B(28), B(27) => B(27), B(26) => B(26), 
                           B(25) => B(25), B(24) => B(24), B(23) => B(23), 
                           B(22) => B(22), B(21) => B(21), B(20) => B(20), 
                           B(19) => B(19), B(18) => B(18), B(17) => B(17), 
                           B(16) => B(16), B(15) => B(15), B(14) => B(14), 
                           B(13) => B(13), B(12) => B(12), B(11) => B(11), 
                           B(10) => B(10), B(9) => B(9), B(8) => B(8), B(7) => 
                           B(7), B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3)
                           => B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), 
                           CI => n1, SUM(59) => S(59), SUM(58) => S(58), 
                           SUM(57) => S(57), SUM(56) => S(56), SUM(55) => S(55)
                           , SUM(54) => S(54), SUM(53) => S(53), SUM(52) => 
                           S(52), SUM(51) => S(51), SUM(50) => S(50), SUM(49) 
                           => S(49), SUM(48) => S(48), SUM(47) => S(47), 
                           SUM(46) => S(46), SUM(45) => S(45), SUM(44) => S(44)
                           , SUM(43) => S(43), SUM(42) => S(42), SUM(41) => 
                           S(41), SUM(40) => S(40), SUM(39) => S(39), SUM(38) 
                           => S(38), SUM(37) => S(37), SUM(36) => S(36), 
                           SUM(35) => S(35), SUM(34) => S(34), SUM(33) => S(33)
                           , SUM(32) => S(32), SUM(31) => S(31), SUM(30) => 
                           S(30), SUM(29) => S(29), SUM(28) => S(28), SUM(27) 
                           => S(27), SUM(26) => S(26), SUM(25) => S(25), 
                           SUM(24) => S(24), SUM(23) => S(23), SUM(22) => S(22)
                           , SUM(21) => S(21), SUM(20) => S(20), SUM(19) => 
                           S(19), SUM(18) => S(18), SUM(17) => S(17), SUM(16) 
                           => S(16), SUM(15) => S(15), SUM(14) => S(14), 
                           SUM(13) => S(13), SUM(12) => S(12), SUM(11) => S(11)
                           , SUM(10) => S(10), SUM(9) => S(9), SUM(8) => S(8), 
                           SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5), 
                           SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1067);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT58 is

   port( A, B : in std_logic_vector (57 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (57 downto 0);  Co : out std_logic);

end RCA_NBIT58;

architecture SYN_DIRECT of RCA_NBIT58 is

   component RCA_NBIT58_DW01_add_0
      port( A, B : in std_logic_vector (57 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (57 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1068 : std_logic;

begin
   
   Co <= '0';
   n1 <= '0';
   add_95 : RCA_NBIT58_DW01_add_0 port map( A(57) => A(57), A(56) => A(56), 
                           A(55) => A(55), A(54) => A(54), A(53) => A(53), 
                           A(52) => A(52), A(51) => A(51), A(50) => A(50), 
                           A(49) => A(49), A(48) => A(48), A(47) => A(47), 
                           A(46) => A(46), A(45) => A(45), A(44) => A(44), 
                           A(43) => A(43), A(42) => A(42), A(41) => A(41), 
                           A(40) => A(40), A(39) => A(39), A(38) => A(38), 
                           A(37) => A(37), A(36) => A(36), A(35) => A(35), 
                           A(34) => A(34), A(33) => A(33), A(32) => A(32), 
                           A(31) => A(31), A(30) => A(30), A(29) => A(29), 
                           A(28) => A(28), A(27) => A(27), A(26) => A(26), 
                           A(25) => A(25), A(24) => A(24), A(23) => A(23), 
                           A(22) => A(22), A(21) => A(21), A(20) => A(20), 
                           A(19) => A(19), A(18) => A(18), A(17) => A(17), 
                           A(16) => A(16), A(15) => A(15), A(14) => A(14), 
                           A(13) => A(13), A(12) => A(12), A(11) => A(11), 
                           A(10) => A(10), A(9) => A(9), A(8) => A(8), A(7) => 
                           A(7), A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3)
                           => A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(57) => B(57), B(56) => B(56), B(55) => B(55), 
                           B(54) => B(54), B(53) => B(53), B(52) => B(52), 
                           B(51) => B(51), B(50) => B(50), B(49) => B(49), 
                           B(48) => B(48), B(47) => B(47), B(46) => B(46), 
                           B(45) => B(45), B(44) => B(44), B(43) => B(43), 
                           B(42) => B(42), B(41) => B(41), B(40) => B(40), 
                           B(39) => B(39), B(38) => B(38), B(37) => B(37), 
                           B(36) => B(36), B(35) => B(35), B(34) => B(34), 
                           B(33) => B(33), B(32) => B(32), B(31) => B(31), 
                           B(30) => B(30), B(29) => B(29), B(28) => B(28), 
                           B(27) => B(27), B(26) => B(26), B(25) => B(25), 
                           B(24) => B(24), B(23) => B(23), B(22) => B(22), 
                           B(21) => B(21), B(20) => B(20), B(19) => B(19), 
                           B(18) => B(18), B(17) => B(17), B(16) => B(16), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => B(0), CI => n1, SUM(57) 
                           => S(57), SUM(56) => S(56), SUM(55) => S(55), 
                           SUM(54) => S(54), SUM(53) => S(53), SUM(52) => S(52)
                           , SUM(51) => S(51), SUM(50) => S(50), SUM(49) => 
                           S(49), SUM(48) => S(48), SUM(47) => S(47), SUM(46) 
                           => S(46), SUM(45) => S(45), SUM(44) => S(44), 
                           SUM(43) => S(43), SUM(42) => S(42), SUM(41) => S(41)
                           , SUM(40) => S(40), SUM(39) => S(39), SUM(38) => 
                           S(38), SUM(37) => S(37), SUM(36) => S(36), SUM(35) 
                           => S(35), SUM(34) => S(34), SUM(33) => S(33), 
                           SUM(32) => S(32), SUM(31) => S(31), SUM(30) => S(30)
                           , SUM(29) => S(29), SUM(28) => S(28), SUM(27) => 
                           S(27), SUM(26) => S(26), SUM(25) => S(25), SUM(24) 
                           => S(24), SUM(23) => S(23), SUM(22) => S(22), 
                           SUM(21) => S(21), SUM(20) => S(20), SUM(19) => S(19)
                           , SUM(18) => S(18), SUM(17) => S(17), SUM(16) => 
                           S(16), SUM(15) => S(15), SUM(14) => S(14), SUM(13) 
                           => S(13), SUM(12) => S(12), SUM(11) => S(11), 
                           SUM(10) => S(10), SUM(9) => S(9), SUM(8) => S(8), 
                           SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5), 
                           SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1068);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT56 is

   port( A, B : in std_logic_vector (55 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (55 downto 0);  Co : out std_logic);

end RCA_NBIT56;

architecture SYN_DIRECT of RCA_NBIT56 is

   component RCA_NBIT56_DW01_add_0
      port( A, B : in std_logic_vector (55 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (55 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1069 : std_logic;

begin
   
   Co <= '0';
   n1 <= '0';
   add_95 : RCA_NBIT56_DW01_add_0 port map( A(55) => A(55), A(54) => A(54), 
                           A(53) => A(53), A(52) => A(52), A(51) => A(51), 
                           A(50) => A(50), A(49) => A(49), A(48) => A(48), 
                           A(47) => A(47), A(46) => A(46), A(45) => A(45), 
                           A(44) => A(44), A(43) => A(43), A(42) => A(42), 
                           A(41) => A(41), A(40) => A(40), A(39) => A(39), 
                           A(38) => A(38), A(37) => A(37), A(36) => A(36), 
                           A(35) => A(35), A(34) => A(34), A(33) => A(33), 
                           A(32) => A(32), A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(55) => B(55), B(54) => B(54), 
                           B(53) => B(53), B(52) => B(52), B(51) => B(51), 
                           B(50) => B(50), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => n1, SUM(55) => S(55), 
                           SUM(54) => S(54), SUM(53) => S(53), SUM(52) => S(52)
                           , SUM(51) => S(51), SUM(50) => S(50), SUM(49) => 
                           S(49), SUM(48) => S(48), SUM(47) => S(47), SUM(46) 
                           => S(46), SUM(45) => S(45), SUM(44) => S(44), 
                           SUM(43) => S(43), SUM(42) => S(42), SUM(41) => S(41)
                           , SUM(40) => S(40), SUM(39) => S(39), SUM(38) => 
                           S(38), SUM(37) => S(37), SUM(36) => S(36), SUM(35) 
                           => S(35), SUM(34) => S(34), SUM(33) => S(33), 
                           SUM(32) => S(32), SUM(31) => S(31), SUM(30) => S(30)
                           , SUM(29) => S(29), SUM(28) => S(28), SUM(27) => 
                           S(27), SUM(26) => S(26), SUM(25) => S(25), SUM(24) 
                           => S(24), SUM(23) => S(23), SUM(22) => S(22), 
                           SUM(21) => S(21), SUM(20) => S(20), SUM(19) => S(19)
                           , SUM(18) => S(18), SUM(17) => S(17), SUM(16) => 
                           S(16), SUM(15) => S(15), SUM(14) => S(14), SUM(13) 
                           => S(13), SUM(12) => S(12), SUM(11) => S(11), 
                           SUM(10) => S(10), SUM(9) => S(9), SUM(8) => S(8), 
                           SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5), 
                           SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1069);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT54 is

   port( A, B : in std_logic_vector (53 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (53 downto 0);  Co : out std_logic);

end RCA_NBIT54;

architecture SYN_DIRECT of RCA_NBIT54 is

   component RCA_NBIT54_DW01_add_0
      port( A, B : in std_logic_vector (53 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (53 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1070 : std_logic;

begin
   
   Co <= '0';
   n1 <= '0';
   add_95 : RCA_NBIT54_DW01_add_0 port map( A(53) => A(53), A(52) => A(52), 
                           A(51) => A(51), A(50) => A(50), A(49) => A(49), 
                           A(48) => A(48), A(47) => A(47), A(46) => A(46), 
                           A(45) => A(45), A(44) => A(44), A(43) => A(43), 
                           A(42) => A(42), A(41) => A(41), A(40) => A(40), 
                           A(39) => A(39), A(38) => A(38), A(37) => A(37), 
                           A(36) => A(36), A(35) => A(35), A(34) => A(34), 
                           A(33) => A(33), A(32) => A(32), A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(53) => B(53), 
                           B(52) => B(52), B(51) => B(51), B(50) => B(50), 
                           B(49) => B(49), B(48) => B(48), B(47) => B(47), 
                           B(46) => B(46), B(45) => B(45), B(44) => B(44), 
                           B(43) => B(43), B(42) => B(42), B(41) => B(41), 
                           B(40) => B(40), B(39) => B(39), B(38) => B(38), 
                           B(37) => B(37), B(36) => B(36), B(35) => B(35), 
                           B(34) => B(34), B(33) => B(33), B(32) => B(32), 
                           B(31) => B(31), B(30) => B(30), B(29) => B(29), 
                           B(28) => B(28), B(27) => B(27), B(26) => B(26), 
                           B(25) => B(25), B(24) => B(24), B(23) => B(23), 
                           B(22) => B(22), B(21) => B(21), B(20) => B(20), 
                           B(19) => B(19), B(18) => B(18), B(17) => B(17), 
                           B(16) => B(16), B(15) => B(15), B(14) => B(14), 
                           B(13) => B(13), B(12) => B(12), B(11) => B(11), 
                           B(10) => B(10), B(9) => B(9), B(8) => B(8), B(7) => 
                           B(7), B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3)
                           => B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), 
                           CI => n1, SUM(53) => S(53), SUM(52) => S(52), 
                           SUM(51) => S(51), SUM(50) => S(50), SUM(49) => S(49)
                           , SUM(48) => S(48), SUM(47) => S(47), SUM(46) => 
                           S(46), SUM(45) => S(45), SUM(44) => S(44), SUM(43) 
                           => S(43), SUM(42) => S(42), SUM(41) => S(41), 
                           SUM(40) => S(40), SUM(39) => S(39), SUM(38) => S(38)
                           , SUM(37) => S(37), SUM(36) => S(36), SUM(35) => 
                           S(35), SUM(34) => S(34), SUM(33) => S(33), SUM(32) 
                           => S(32), SUM(31) => S(31), SUM(30) => S(30), 
                           SUM(29) => S(29), SUM(28) => S(28), SUM(27) => S(27)
                           , SUM(26) => S(26), SUM(25) => S(25), SUM(24) => 
                           S(24), SUM(23) => S(23), SUM(22) => S(22), SUM(21) 
                           => S(21), SUM(20) => S(20), SUM(19) => S(19), 
                           SUM(18) => S(18), SUM(17) => S(17), SUM(16) => S(16)
                           , SUM(15) => S(15), SUM(14) => S(14), SUM(13) => 
                           S(13), SUM(12) => S(12), SUM(11) => S(11), SUM(10) 
                           => S(10), SUM(9) => S(9), SUM(8) => S(8), SUM(7) => 
                           S(7), SUM(6) => S(6), SUM(5) => S(5), SUM(4) => S(4)
                           , SUM(3) => S(3), SUM(2) => S(2), SUM(1) => S(1), 
                           SUM(0) => S(0), CO => n_1070);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT52 is

   port( A, B : in std_logic_vector (51 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (51 downto 0);  Co : out std_logic);

end RCA_NBIT52;

architecture SYN_DIRECT of RCA_NBIT52 is

   component RCA_NBIT52_DW01_add_0
      port( A, B : in std_logic_vector (51 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (51 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1071 : std_logic;

begin
   
   Co <= '0';
   n1 <= '0';
   add_95 : RCA_NBIT52_DW01_add_0 port map( A(51) => A(51), A(50) => A(50), 
                           A(49) => A(49), A(48) => A(48), A(47) => A(47), 
                           A(46) => A(46), A(45) => A(45), A(44) => A(44), 
                           A(43) => A(43), A(42) => A(42), A(41) => A(41), 
                           A(40) => A(40), A(39) => A(39), A(38) => A(38), 
                           A(37) => A(37), A(36) => A(36), A(35) => A(35), 
                           A(34) => A(34), A(33) => A(33), A(32) => A(32), 
                           A(31) => A(31), A(30) => A(30), A(29) => A(29), 
                           A(28) => A(28), A(27) => A(27), A(26) => A(26), 
                           A(25) => A(25), A(24) => A(24), A(23) => A(23), 
                           A(22) => A(22), A(21) => A(21), A(20) => A(20), 
                           A(19) => A(19), A(18) => A(18), A(17) => A(17), 
                           A(16) => A(16), A(15) => A(15), A(14) => A(14), 
                           A(13) => A(13), A(12) => A(12), A(11) => A(11), 
                           A(10) => A(10), A(9) => A(9), A(8) => A(8), A(7) => 
                           A(7), A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3)
                           => A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(51) => B(51), B(50) => B(50), B(49) => B(49), 
                           B(48) => B(48), B(47) => B(47), B(46) => B(46), 
                           B(45) => B(45), B(44) => B(44), B(43) => B(43), 
                           B(42) => B(42), B(41) => B(41), B(40) => B(40), 
                           B(39) => B(39), B(38) => B(38), B(37) => B(37), 
                           B(36) => B(36), B(35) => B(35), B(34) => B(34), 
                           B(33) => B(33), B(32) => B(32), B(31) => B(31), 
                           B(30) => B(30), B(29) => B(29), B(28) => B(28), 
                           B(27) => B(27), B(26) => B(26), B(25) => B(25), 
                           B(24) => B(24), B(23) => B(23), B(22) => B(22), 
                           B(21) => B(21), B(20) => B(20), B(19) => B(19), 
                           B(18) => B(18), B(17) => B(17), B(16) => B(16), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => B(0), CI => n1, SUM(51) 
                           => S(51), SUM(50) => S(50), SUM(49) => S(49), 
                           SUM(48) => S(48), SUM(47) => S(47), SUM(46) => S(46)
                           , SUM(45) => S(45), SUM(44) => S(44), SUM(43) => 
                           S(43), SUM(42) => S(42), SUM(41) => S(41), SUM(40) 
                           => S(40), SUM(39) => S(39), SUM(38) => S(38), 
                           SUM(37) => S(37), SUM(36) => S(36), SUM(35) => S(35)
                           , SUM(34) => S(34), SUM(33) => S(33), SUM(32) => 
                           S(32), SUM(31) => S(31), SUM(30) => S(30), SUM(29) 
                           => S(29), SUM(28) => S(28), SUM(27) => S(27), 
                           SUM(26) => S(26), SUM(25) => S(25), SUM(24) => S(24)
                           , SUM(23) => S(23), SUM(22) => S(22), SUM(21) => 
                           S(21), SUM(20) => S(20), SUM(19) => S(19), SUM(18) 
                           => S(18), SUM(17) => S(17), SUM(16) => S(16), 
                           SUM(15) => S(15), SUM(14) => S(14), SUM(13) => S(13)
                           , SUM(12) => S(12), SUM(11) => S(11), SUM(10) => 
                           S(10), SUM(9) => S(9), SUM(8) => S(8), SUM(7) => 
                           S(7), SUM(6) => S(6), SUM(5) => S(5), SUM(4) => S(4)
                           , SUM(3) => S(3), SUM(2) => S(2), SUM(1) => S(1), 
                           SUM(0) => S(0), CO => n_1071);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT50 is

   port( A, B : in std_logic_vector (49 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (49 downto 0);  Co : out std_logic);

end RCA_NBIT50;

architecture SYN_DIRECT of RCA_NBIT50 is

   component RCA_NBIT50_DW01_add_0
      port( A, B : in std_logic_vector (49 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (49 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1072 : std_logic;

begin
   
   Co <= '0';
   n1 <= '0';
   add_95 : RCA_NBIT50_DW01_add_0 port map( A(49) => A(49), A(48) => A(48), 
                           A(47) => A(47), A(46) => A(46), A(45) => A(45), 
                           A(44) => A(44), A(43) => A(43), A(42) => A(42), 
                           A(41) => A(41), A(40) => A(40), A(39) => A(39), 
                           A(38) => A(38), A(37) => A(37), A(36) => A(36), 
                           A(35) => A(35), A(34) => A(34), A(33) => A(33), 
                           A(32) => A(32), A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => n1, SUM(49) => S(49), 
                           SUM(48) => S(48), SUM(47) => S(47), SUM(46) => S(46)
                           , SUM(45) => S(45), SUM(44) => S(44), SUM(43) => 
                           S(43), SUM(42) => S(42), SUM(41) => S(41), SUM(40) 
                           => S(40), SUM(39) => S(39), SUM(38) => S(38), 
                           SUM(37) => S(37), SUM(36) => S(36), SUM(35) => S(35)
                           , SUM(34) => S(34), SUM(33) => S(33), SUM(32) => 
                           S(32), SUM(31) => S(31), SUM(30) => S(30), SUM(29) 
                           => S(29), SUM(28) => S(28), SUM(27) => S(27), 
                           SUM(26) => S(26), SUM(25) => S(25), SUM(24) => S(24)
                           , SUM(23) => S(23), SUM(22) => S(22), SUM(21) => 
                           S(21), SUM(20) => S(20), SUM(19) => S(19), SUM(18) 
                           => S(18), SUM(17) => S(17), SUM(16) => S(16), 
                           SUM(15) => S(15), SUM(14) => S(14), SUM(13) => S(13)
                           , SUM(12) => S(12), SUM(11) => S(11), SUM(10) => 
                           S(10), SUM(9) => S(9), SUM(8) => S(8), SUM(7) => 
                           S(7), SUM(6) => S(6), SUM(5) => S(5), SUM(4) => S(4)
                           , SUM(3) => S(3), SUM(2) => S(2), SUM(1) => S(1), 
                           SUM(0) => S(0), CO => n_1072);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT48 is

   port( A, B : in std_logic_vector (47 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (47 downto 0);  Co : out std_logic);

end RCA_NBIT48;

architecture SYN_DIRECT of RCA_NBIT48 is

   component RCA_NBIT48_DW01_add_0
      port( A, B : in std_logic_vector (47 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (47 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1073 : std_logic;

begin
   
   Co <= '0';
   n1 <= '0';
   add_95 : RCA_NBIT48_DW01_add_0 port map( A(47) => A(47), A(46) => A(46), 
                           A(45) => A(45), A(44) => A(44), A(43) => A(43), 
                           A(42) => A(42), A(41) => A(41), A(40) => A(40), 
                           A(39) => A(39), A(38) => A(38), A(37) => A(37), 
                           A(36) => A(36), A(35) => A(35), A(34) => A(34), 
                           A(33) => A(33), A(32) => A(32), A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(47) => B(47), 
                           B(46) => B(46), B(45) => B(45), B(44) => B(44), 
                           B(43) => B(43), B(42) => B(42), B(41) => B(41), 
                           B(40) => B(40), B(39) => B(39), B(38) => B(38), 
                           B(37) => B(37), B(36) => B(36), B(35) => B(35), 
                           B(34) => B(34), B(33) => B(33), B(32) => B(32), 
                           B(31) => B(31), B(30) => B(30), B(29) => B(29), 
                           B(28) => B(28), B(27) => B(27), B(26) => B(26), 
                           B(25) => B(25), B(24) => B(24), B(23) => B(23), 
                           B(22) => B(22), B(21) => B(21), B(20) => B(20), 
                           B(19) => B(19), B(18) => B(18), B(17) => B(17), 
                           B(16) => B(16), B(15) => B(15), B(14) => B(14), 
                           B(13) => B(13), B(12) => B(12), B(11) => B(11), 
                           B(10) => B(10), B(9) => B(9), B(8) => B(8), B(7) => 
                           B(7), B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3)
                           => B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), 
                           CI => n1, SUM(47) => S(47), SUM(46) => S(46), 
                           SUM(45) => S(45), SUM(44) => S(44), SUM(43) => S(43)
                           , SUM(42) => S(42), SUM(41) => S(41), SUM(40) => 
                           S(40), SUM(39) => S(39), SUM(38) => S(38), SUM(37) 
                           => S(37), SUM(36) => S(36), SUM(35) => S(35), 
                           SUM(34) => S(34), SUM(33) => S(33), SUM(32) => S(32)
                           , SUM(31) => S(31), SUM(30) => S(30), SUM(29) => 
                           S(29), SUM(28) => S(28), SUM(27) => S(27), SUM(26) 
                           => S(26), SUM(25) => S(25), SUM(24) => S(24), 
                           SUM(23) => S(23), SUM(22) => S(22), SUM(21) => S(21)
                           , SUM(20) => S(20), SUM(19) => S(19), SUM(18) => 
                           S(18), SUM(17) => S(17), SUM(16) => S(16), SUM(15) 
                           => S(15), SUM(14) => S(14), SUM(13) => S(13), 
                           SUM(12) => S(12), SUM(11) => S(11), SUM(10) => S(10)
                           , SUM(9) => S(9), SUM(8) => S(8), SUM(7) => S(7), 
                           SUM(6) => S(6), SUM(5) => S(5), SUM(4) => S(4), 
                           SUM(3) => S(3), SUM(2) => S(2), SUM(1) => S(1), 
                           SUM(0) => S(0), CO => n_1073);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT46 is

   port( A, B : in std_logic_vector (45 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (45 downto 0);  Co : out std_logic);

end RCA_NBIT46;

architecture SYN_DIRECT of RCA_NBIT46 is

   component RCA_NBIT46_DW01_add_0
      port( A, B : in std_logic_vector (45 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (45 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1074 : std_logic;

begin
   
   Co <= '0';
   n1 <= '0';
   add_95 : RCA_NBIT46_DW01_add_0 port map( A(45) => A(45), A(44) => A(44), 
                           A(43) => A(43), A(42) => A(42), A(41) => A(41), 
                           A(40) => A(40), A(39) => A(39), A(38) => A(38), 
                           A(37) => A(37), A(36) => A(36), A(35) => A(35), 
                           A(34) => A(34), A(33) => A(33), A(32) => A(32), 
                           A(31) => A(31), A(30) => A(30), A(29) => A(29), 
                           A(28) => A(28), A(27) => A(27), A(26) => A(26), 
                           A(25) => A(25), A(24) => A(24), A(23) => A(23), 
                           A(22) => A(22), A(21) => A(21), A(20) => A(20), 
                           A(19) => A(19), A(18) => A(18), A(17) => A(17), 
                           A(16) => A(16), A(15) => A(15), A(14) => A(14), 
                           A(13) => A(13), A(12) => A(12), A(11) => A(11), 
                           A(10) => A(10), A(9) => A(9), A(8) => A(8), A(7) => 
                           A(7), A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3)
                           => A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(45) => B(45), B(44) => B(44), B(43) => B(43), 
                           B(42) => B(42), B(41) => B(41), B(40) => B(40), 
                           B(39) => B(39), B(38) => B(38), B(37) => B(37), 
                           B(36) => B(36), B(35) => B(35), B(34) => B(34), 
                           B(33) => B(33), B(32) => B(32), B(31) => B(31), 
                           B(30) => B(30), B(29) => B(29), B(28) => B(28), 
                           B(27) => B(27), B(26) => B(26), B(25) => B(25), 
                           B(24) => B(24), B(23) => B(23), B(22) => B(22), 
                           B(21) => B(21), B(20) => B(20), B(19) => B(19), 
                           B(18) => B(18), B(17) => B(17), B(16) => B(16), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => B(0), CI => n1, SUM(45) 
                           => S(45), SUM(44) => S(44), SUM(43) => S(43), 
                           SUM(42) => S(42), SUM(41) => S(41), SUM(40) => S(40)
                           , SUM(39) => S(39), SUM(38) => S(38), SUM(37) => 
                           S(37), SUM(36) => S(36), SUM(35) => S(35), SUM(34) 
                           => S(34), SUM(33) => S(33), SUM(32) => S(32), 
                           SUM(31) => S(31), SUM(30) => S(30), SUM(29) => S(29)
                           , SUM(28) => S(28), SUM(27) => S(27), SUM(26) => 
                           S(26), SUM(25) => S(25), SUM(24) => S(24), SUM(23) 
                           => S(23), SUM(22) => S(22), SUM(21) => S(21), 
                           SUM(20) => S(20), SUM(19) => S(19), SUM(18) => S(18)
                           , SUM(17) => S(17), SUM(16) => S(16), SUM(15) => 
                           S(15), SUM(14) => S(14), SUM(13) => S(13), SUM(12) 
                           => S(12), SUM(11) => S(11), SUM(10) => S(10), SUM(9)
                           => S(9), SUM(8) => S(8), SUM(7) => S(7), SUM(6) => 
                           S(6), SUM(5) => S(5), SUM(4) => S(4), SUM(3) => S(3)
                           , SUM(2) => S(2), SUM(1) => S(1), SUM(0) => S(0), CO
                           => n_1074);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT44 is

   port( A, B : in std_logic_vector (43 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (43 downto 0);  Co : out std_logic);

end RCA_NBIT44;

architecture SYN_DIRECT of RCA_NBIT44 is

   component RCA_NBIT44_DW01_add_0
      port( A, B : in std_logic_vector (43 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (43 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1075 : std_logic;

begin
   
   Co <= '0';
   n1 <= '0';
   add_95 : RCA_NBIT44_DW01_add_0 port map( A(43) => A(43), A(42) => A(42), 
                           A(41) => A(41), A(40) => A(40), A(39) => A(39), 
                           A(38) => A(38), A(37) => A(37), A(36) => A(36), 
                           A(35) => A(35), A(34) => A(34), A(33) => A(33), 
                           A(32) => A(32), A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => n1, SUM(43) => S(43), 
                           SUM(42) => S(42), SUM(41) => S(41), SUM(40) => S(40)
                           , SUM(39) => S(39), SUM(38) => S(38), SUM(37) => 
                           S(37), SUM(36) => S(36), SUM(35) => S(35), SUM(34) 
                           => S(34), SUM(33) => S(33), SUM(32) => S(32), 
                           SUM(31) => S(31), SUM(30) => S(30), SUM(29) => S(29)
                           , SUM(28) => S(28), SUM(27) => S(27), SUM(26) => 
                           S(26), SUM(25) => S(25), SUM(24) => S(24), SUM(23) 
                           => S(23), SUM(22) => S(22), SUM(21) => S(21), 
                           SUM(20) => S(20), SUM(19) => S(19), SUM(18) => S(18)
                           , SUM(17) => S(17), SUM(16) => S(16), SUM(15) => 
                           S(15), SUM(14) => S(14), SUM(13) => S(13), SUM(12) 
                           => S(12), SUM(11) => S(11), SUM(10) => S(10), SUM(9)
                           => S(9), SUM(8) => S(8), SUM(7) => S(7), SUM(6) => 
                           S(6), SUM(5) => S(5), SUM(4) => S(4), SUM(3) => S(3)
                           , SUM(2) => S(2), SUM(1) => S(1), SUM(0) => S(0), CO
                           => n_1075);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT42 is

   port( A, B : in std_logic_vector (41 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (41 downto 0);  Co : out std_logic);

end RCA_NBIT42;

architecture SYN_DIRECT of RCA_NBIT42 is

   component RCA_NBIT42_DW01_add_0
      port( A, B : in std_logic_vector (41 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (41 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1076 : std_logic;

begin
   
   Co <= '0';
   n1 <= '0';
   add_95 : RCA_NBIT42_DW01_add_0 port map( A(41) => A(41), A(40) => A(40), 
                           A(39) => A(39), A(38) => A(38), A(37) => A(37), 
                           A(36) => A(36), A(35) => A(35), A(34) => A(34), 
                           A(33) => A(33), A(32) => A(32), A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(41) => B(41), 
                           B(40) => B(40), B(39) => B(39), B(38) => B(38), 
                           B(37) => B(37), B(36) => B(36), B(35) => B(35), 
                           B(34) => B(34), B(33) => B(33), B(32) => B(32), 
                           B(31) => B(31), B(30) => B(30), B(29) => B(29), 
                           B(28) => B(28), B(27) => B(27), B(26) => B(26), 
                           B(25) => B(25), B(24) => B(24), B(23) => B(23), 
                           B(22) => B(22), B(21) => B(21), B(20) => B(20), 
                           B(19) => B(19), B(18) => B(18), B(17) => B(17), 
                           B(16) => B(16), B(15) => B(15), B(14) => B(14), 
                           B(13) => B(13), B(12) => B(12), B(11) => B(11), 
                           B(10) => B(10), B(9) => B(9), B(8) => B(8), B(7) => 
                           B(7), B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3)
                           => B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), 
                           CI => n1, SUM(41) => S(41), SUM(40) => S(40), 
                           SUM(39) => S(39), SUM(38) => S(38), SUM(37) => S(37)
                           , SUM(36) => S(36), SUM(35) => S(35), SUM(34) => 
                           S(34), SUM(33) => S(33), SUM(32) => S(32), SUM(31) 
                           => S(31), SUM(30) => S(30), SUM(29) => S(29), 
                           SUM(28) => S(28), SUM(27) => S(27), SUM(26) => S(26)
                           , SUM(25) => S(25), SUM(24) => S(24), SUM(23) => 
                           S(23), SUM(22) => S(22), SUM(21) => S(21), SUM(20) 
                           => S(20), SUM(19) => S(19), SUM(18) => S(18), 
                           SUM(17) => S(17), SUM(16) => S(16), SUM(15) => S(15)
                           , SUM(14) => S(14), SUM(13) => S(13), SUM(12) => 
                           S(12), SUM(11) => S(11), SUM(10) => S(10), SUM(9) =>
                           S(9), SUM(8) => S(8), SUM(7) => S(7), SUM(6) => S(6)
                           , SUM(5) => S(5), SUM(4) => S(4), SUM(3) => S(3), 
                           SUM(2) => S(2), SUM(1) => S(1), SUM(0) => S(0), CO 
                           => n_1076);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT40 is

   port( A, B : in std_logic_vector (39 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (39 downto 0);  Co : out std_logic);

end RCA_NBIT40;

architecture SYN_DIRECT of RCA_NBIT40 is

   component RCA_NBIT40_DW01_add_0
      port( A, B : in std_logic_vector (39 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (39 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1077 : std_logic;

begin
   
   Co <= '0';
   n1 <= '0';
   add_95 : RCA_NBIT40_DW01_add_0 port map( A(39) => A(39), A(38) => A(38), 
                           A(37) => A(37), A(36) => A(36), A(35) => A(35), 
                           A(34) => A(34), A(33) => A(33), A(32) => A(32), 
                           A(31) => A(31), A(30) => A(30), A(29) => A(29), 
                           A(28) => A(28), A(27) => A(27), A(26) => A(26), 
                           A(25) => A(25), A(24) => A(24), A(23) => A(23), 
                           A(22) => A(22), A(21) => A(21), A(20) => A(20), 
                           A(19) => A(19), A(18) => A(18), A(17) => A(17), 
                           A(16) => A(16), A(15) => A(15), A(14) => A(14), 
                           A(13) => A(13), A(12) => A(12), A(11) => A(11), 
                           A(10) => A(10), A(9) => A(9), A(8) => A(8), A(7) => 
                           A(7), A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3)
                           => A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(39) => B(39), B(38) => B(38), B(37) => B(37), 
                           B(36) => B(36), B(35) => B(35), B(34) => B(34), 
                           B(33) => B(33), B(32) => B(32), B(31) => B(31), 
                           B(30) => B(30), B(29) => B(29), B(28) => B(28), 
                           B(27) => B(27), B(26) => B(26), B(25) => B(25), 
                           B(24) => B(24), B(23) => B(23), B(22) => B(22), 
                           B(21) => B(21), B(20) => B(20), B(19) => B(19), 
                           B(18) => B(18), B(17) => B(17), B(16) => B(16), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => B(0), CI => n1, SUM(39) 
                           => S(39), SUM(38) => S(38), SUM(37) => S(37), 
                           SUM(36) => S(36), SUM(35) => S(35), SUM(34) => S(34)
                           , SUM(33) => S(33), SUM(32) => S(32), SUM(31) => 
                           S(31), SUM(30) => S(30), SUM(29) => S(29), SUM(28) 
                           => S(28), SUM(27) => S(27), SUM(26) => S(26), 
                           SUM(25) => S(25), SUM(24) => S(24), SUM(23) => S(23)
                           , SUM(22) => S(22), SUM(21) => S(21), SUM(20) => 
                           S(20), SUM(19) => S(19), SUM(18) => S(18), SUM(17) 
                           => S(17), SUM(16) => S(16), SUM(15) => S(15), 
                           SUM(14) => S(14), SUM(13) => S(13), SUM(12) => S(12)
                           , SUM(11) => S(11), SUM(10) => S(10), SUM(9) => S(9)
                           , SUM(8) => S(8), SUM(7) => S(7), SUM(6) => S(6), 
                           SUM(5) => S(5), SUM(4) => S(4), SUM(3) => S(3), 
                           SUM(2) => S(2), SUM(1) => S(1), SUM(0) => S(0), CO 
                           => n_1077);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT38 is

   port( A, B : in std_logic_vector (37 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (37 downto 0);  Co : out std_logic);

end RCA_NBIT38;

architecture SYN_DIRECT of RCA_NBIT38 is

   component RCA_NBIT38_DW01_add_0
      port( A, B : in std_logic_vector (37 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (37 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1078 : std_logic;

begin
   
   Co <= '0';
   n1 <= '0';
   add_95 : RCA_NBIT38_DW01_add_0 port map( A(37) => A(37), A(36) => A(36), 
                           A(35) => A(35), A(34) => A(34), A(33) => A(33), 
                           A(32) => A(32), A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => n1, SUM(37) => S(37), 
                           SUM(36) => S(36), SUM(35) => S(35), SUM(34) => S(34)
                           , SUM(33) => S(33), SUM(32) => S(32), SUM(31) => 
                           S(31), SUM(30) => S(30), SUM(29) => S(29), SUM(28) 
                           => S(28), SUM(27) => S(27), SUM(26) => S(26), 
                           SUM(25) => S(25), SUM(24) => S(24), SUM(23) => S(23)
                           , SUM(22) => S(22), SUM(21) => S(21), SUM(20) => 
                           S(20), SUM(19) => S(19), SUM(18) => S(18), SUM(17) 
                           => S(17), SUM(16) => S(16), SUM(15) => S(15), 
                           SUM(14) => S(14), SUM(13) => S(13), SUM(12) => S(12)
                           , SUM(11) => S(11), SUM(10) => S(10), SUM(9) => S(9)
                           , SUM(8) => S(8), SUM(7) => S(7), SUM(6) => S(6), 
                           SUM(5) => S(5), SUM(4) => S(4), SUM(3) => S(3), 
                           SUM(2) => S(2), SUM(1) => S(1), SUM(0) => S(0), CO 
                           => n_1078);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT36 is

   port( A, B : in std_logic_vector (35 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (35 downto 0);  Co : out std_logic);

end RCA_NBIT36;

architecture SYN_DIRECT of RCA_NBIT36 is

   component RCA_NBIT36_DW01_add_0
      port( A, B : in std_logic_vector (35 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (35 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1079 : std_logic;

begin
   
   Co <= '0';
   n1 <= '0';
   add_95 : RCA_NBIT36_DW01_add_0 port map( A(35) => A(35), A(34) => A(34), 
                           A(33) => A(33), A(32) => A(32), A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(35) => B(35), 
                           B(34) => B(34), B(33) => B(33), B(32) => B(32), 
                           B(31) => B(31), B(30) => B(30), B(29) => B(29), 
                           B(28) => B(28), B(27) => B(27), B(26) => B(26), 
                           B(25) => B(25), B(24) => B(24), B(23) => B(23), 
                           B(22) => B(22), B(21) => B(21), B(20) => B(20), 
                           B(19) => B(19), B(18) => B(18), B(17) => B(17), 
                           B(16) => B(16), B(15) => B(15), B(14) => B(14), 
                           B(13) => B(13), B(12) => B(12), B(11) => B(11), 
                           B(10) => B(10), B(9) => B(9), B(8) => B(8), B(7) => 
                           B(7), B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3)
                           => B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), 
                           CI => n1, SUM(35) => S(35), SUM(34) => S(34), 
                           SUM(33) => S(33), SUM(32) => S(32), SUM(31) => S(31)
                           , SUM(30) => S(30), SUM(29) => S(29), SUM(28) => 
                           S(28), SUM(27) => S(27), SUM(26) => S(26), SUM(25) 
                           => S(25), SUM(24) => S(24), SUM(23) => S(23), 
                           SUM(22) => S(22), SUM(21) => S(21), SUM(20) => S(20)
                           , SUM(19) => S(19), SUM(18) => S(18), SUM(17) => 
                           S(17), SUM(16) => S(16), SUM(15) => S(15), SUM(14) 
                           => S(14), SUM(13) => S(13), SUM(12) => S(12), 
                           SUM(11) => S(11), SUM(10) => S(10), SUM(9) => S(9), 
                           SUM(8) => S(8), SUM(7) => S(7), SUM(6) => S(6), 
                           SUM(5) => S(5), SUM(4) => S(4), SUM(3) => S(3), 
                           SUM(2) => S(2), SUM(1) => S(1), SUM(0) => S(0), CO 
                           => n_1079);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT64_i30 is

   port( A_s, A_ns, B : in std_logic_vector (63 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (63 downto 0));

end BOOTHENC_NBIT64_i30;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT64_i30 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, O_63_port, O_62_port, O_61_port, O_60_port, O_59_port,
      O_58_port, O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, 
      O_52_port, O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, 
      O_46_port, O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, 
      O_40_port, O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, 
      O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, 
      O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, 
      O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, 
      O_16_port, O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, 
      O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, 
      O_3_port, O_2_port, O_1_port, n128, n129, n130, n131, n132, n133, n134, 
      n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, 
      n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, 
      n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, 
      n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, 
      n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, 
      n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, 
      n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, 
      n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, 
      n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, 
      n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, 
      n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, 
      n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, 
      n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, 
      n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, 
      n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, 
      n1235, n1236 : std_logic;

begin
   O <= ( O_63_port, O_62_port, O_61_port, O_60_port, O_59_port, O_58_port, 
      O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, O_52_port, 
      O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, O_46_port, 
      O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, O_40_port, 
      O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, 
      O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, 
      O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, 
      O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, O_16_port, 
      O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, O_10_port, 
      O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, O_3_port, 
      O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(61), A_s(60), A_s(59), A_s(58), A_s(57), A_s(56), A_s(55), 
      A_s(54), A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), 
      A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), 
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   A_nso <= ( A_ns(61), A_ns(60), A_ns(59), A_ns(58), A_ns(57), A_ns(56), 
      A_ns(55), A_ns(54), A_ns(53), A_ns(52), A_ns(51), A_ns(50), A_ns(49), 
      A_ns(48), A_ns(47), A_ns(46), A_ns(45), A_ns(44), A_ns(43), A_ns(42), 
      A_ns(41), A_ns(40), A_ns(39), A_ns(38), A_ns(37), A_ns(36), A_ns(35), 
      A_ns(34), A_ns(33), A_ns(32), A_ns(31), A_ns(30), A_ns(29), A_ns(28), 
      A_ns(27), A_ns(26), A_ns(25), A_ns(24), A_ns(23), A_ns(22), A_ns(21), 
      A_ns(20), A_ns(19), A_ns(18), A_ns(17), A_ns(16), A_ns(15), A_ns(14), 
      A_ns(13), A_ns(12), A_ns(11), A_ns(10), A_ns(9), A_ns(8), A_ns(7), 
      A_ns(6), A_ns(5), A_ns(4), A_ns(3), A_ns(2), A_ns(1), A_ns(0), 
      X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U257 : XOR2_X1 port map( A => B(29), B => B(30), Z => n194);
   U258 : NAND3_X1 port map( A1 => B(30), A2 => n1236, A3 => B(29), ZN => n128)
                           ;
   U2 : OAI221_X1 port map( B1 => n1104, B2 => n1173, C1 => n1101, C2 => n1139,
                           A => n136, ZN => O_61_port);
   U3 : AOI22_X1 port map( A1 => A_ns(62), A2 => n1095, B1 => A_s(62), B2 => 
                           n1089, ZN => n134);
   U4 : BUF_X1 port map( A => n1235, Z => n1092);
   U5 : BUF_X1 port map( A => n1235, Z => n1093);
   U6 : BUF_X1 port map( A => n1234, Z => n1086);
   U7 : BUF_X1 port map( A => n1234, Z => n1087);
   U8 : BUF_X1 port map( A => n1235, Z => n1094);
   U9 : BUF_X1 port map( A => n1234, Z => n1088);
   U10 : BUF_X1 port map( A => n1234, Z => n1089);
   U11 : BUF_X1 port map( A => n1235, Z => n1095);
   U12 : BUF_X1 port map( A => n1235, Z => n1091);
   U13 : BUF_X1 port map( A => n1234, Z => n1085);
   U14 : OAI221_X1 port map( B1 => n1104, B2 => n1175, C1 => n1101, C2 => n1141
                           , A => n134, ZN => O_63_port);
   U15 : OAI221_X1 port map( B1 => n1107, B2 => n1144, C1 => n1098, C2 => n1110
                           , A => n168, ZN => O_32_port);
   U16 : AOI22_X1 port map( A1 => A_ns(31), A2 => n1092, B1 => A_s(31), B2 => 
                           n1086, ZN => n168);
   U17 : OAI221_X1 port map( B1 => n1106, B2 => n1148, C1 => n1099, C2 => n1114
                           , A => n164, ZN => O_36_port);
   U18 : AOI22_X1 port map( A1 => A_ns(35), A2 => n1093, B1 => A_s(35), B2 => 
                           n1087, ZN => n164);
   U19 : OAI221_X1 port map( B1 => n1106, B2 => n1150, C1 => n1099, C2 => n1116
                           , A => n162, ZN => O_38_port);
   U20 : AOI22_X1 port map( A1 => A_ns(37), A2 => n1093, B1 => A_s(37), B2 => 
                           n1087, ZN => n162);
   U21 : OAI221_X1 port map( B1 => n1106, B2 => n1147, C1 => n1099, C2 => n1113
                           , A => n165, ZN => O_35_port);
   U22 : AOI22_X1 port map( A1 => A_ns(34), A2 => n1093, B1 => A_s(34), B2 => 
                           n1087, ZN => n165);
   U23 : OAI221_X1 port map( B1 => n1106, B2 => n1149, C1 => n1099, C2 => n1115
                           , A => n163, ZN => O_37_port);
   U24 : AOI22_X1 port map( A1 => A_ns(36), A2 => n1093, B1 => A_s(36), B2 => 
                           n1087, ZN => n163);
   U25 : OAI221_X1 port map( B1 => n1106, B2 => n1151, C1 => n1099, C2 => n1117
                           , A => n161, ZN => O_39_port);
   U26 : AOI22_X1 port map( A1 => A_ns(38), A2 => n1093, B1 => A_s(38), B2 => 
                           n1087, ZN => n161);
   U27 : OAI221_X1 port map( B1 => n1106, B2 => n1153, C1 => n1099, C2 => n1119
                           , A => n158, ZN => O_41_port);
   U28 : AOI22_X1 port map( A1 => A_ns(40), A2 => n1093, B1 => A_s(40), B2 => 
                           n1087, ZN => n158);
   U29 : OAI221_X1 port map( B1 => n1106, B2 => n1155, C1 => n1099, C2 => n1121
                           , A => n156, ZN => O_43_port);
   U30 : AOI22_X1 port map( A1 => A_ns(42), A2 => n1093, B1 => A_s(42), B2 => 
                           n1087, ZN => n156);
   U31 : OAI221_X1 port map( B1 => n1106, B2 => n1152, C1 => n1099, C2 => n1118
                           , A => n159, ZN => O_40_port);
   U32 : AOI22_X1 port map( A1 => A_ns(39), A2 => n1093, B1 => A_s(39), B2 => 
                           n1087, ZN => n159);
   U33 : OAI221_X1 port map( B1 => n1107, B2 => n1146, C1 => n1098, C2 => n1112
                           , A => n166, ZN => O_34_port);
   U34 : AOI22_X1 port map( A1 => A_ns(33), A2 => n1093, B1 => A_s(33), B2 => 
                           n1087, ZN => n166);
   U35 : OAI221_X1 port map( B1 => n1107, B2 => n1143, C1 => n1098, C2 => n1142
                           , A => n169, ZN => O_31_port);
   U36 : AOI22_X1 port map( A1 => A_ns(30), A2 => n1092, B1 => A_s(30), B2 => 
                           n1086, ZN => n169);
   U37 : OAI221_X1 port map( B1 => n1107, B2 => n1145, C1 => n1098, C2 => n1111
                           , A => n167, ZN => O_33_port);
   U38 : AOI22_X1 port map( A1 => A_ns(32), A2 => n1093, B1 => A_s(32), B2 => 
                           n1087, ZN => n167);
   U39 : BUF_X1 port map( A => n1103, Z => n1098);
   U40 : OAI221_X1 port map( B1 => n1106, B2 => n1156, C1 => n1099, C2 => n1122
                           , A => n155, ZN => O_44_port);
   U41 : AOI22_X1 port map( A1 => A_ns(43), A2 => n1094, B1 => A_s(43), B2 => 
                           n1088, ZN => n155);
   U42 : INV_X1 port map( A => n183, ZN => n1235);
   U43 : OAI221_X1 port map( B1 => n1106, B2 => n1154, C1 => n1099, C2 => n1120
                           , A => n157, ZN => O_42_port);
   U44 : AOI22_X1 port map( A1 => A_ns(41), A2 => n1093, B1 => A_s(41), B2 => 
                           n1087, ZN => n157);
   U45 : INV_X1 port map( A => n182, ZN => n1234);
   U46 : OAI221_X1 port map( B1 => n1105, B2 => n1160, C1 => n1100, C2 => n1126
                           , A => n151, ZN => O_48_port);
   U47 : AOI22_X1 port map( A1 => A_ns(47), A2 => n1094, B1 => A_s(47), B2 => 
                           n1088, ZN => n151);
   U48 : OAI221_X1 port map( B1 => n1105, B2 => n1166, C1 => n1100, C2 => n1132
                           , A => n144, ZN => O_54_port);
   U49 : AOI22_X1 port map( A1 => A_ns(53), A2 => n1094, B1 => A_s(53), B2 => 
                           n1088, ZN => n144);
   U50 : OAI221_X1 port map( B1 => n1105, B2 => n1158, C1 => n1099, C2 => n1124
                           , A => n153, ZN => O_46_port);
   U51 : AOI22_X1 port map( A1 => A_ns(45), A2 => n1094, B1 => A_s(45), B2 => 
                           n1088, ZN => n153);
   U52 : OAI221_X1 port map( B1 => n1105, B2 => n1165, C1 => n1100, C2 => n1131
                           , A => n145, ZN => O_53_port);
   U53 : AOI22_X1 port map( A1 => A_ns(52), A2 => n1094, B1 => A_s(52), B2 => 
                           n1088, ZN => n145);
   U54 : OAI221_X1 port map( B1 => n1105, B2 => n1168, C1 => n1100, C2 => n1134
                           , A => n142, ZN => O_56_port);
   U55 : AOI22_X1 port map( A1 => A_ns(55), A2 => n1095, B1 => A_s(55), B2 => 
                           n1089, ZN => n142);
   U56 : BUF_X1 port map( A => n1102, Z => n1099);
   U57 : OAI221_X1 port map( B1 => n1106, B2 => n1157, C1 => n1099, C2 => n1123
                           , A => n154, ZN => O_45_port);
   U58 : AOI22_X1 port map( A1 => A_ns(44), A2 => n1094, B1 => A_s(44), B2 => 
                           n1088, ZN => n154);
   U59 : OAI221_X1 port map( B1 => n1105, B2 => n1159, C1 => n1100, C2 => n1125
                           , A => n152, ZN => O_47_port);
   U60 : AOI22_X1 port map( A1 => A_ns(46), A2 => n1094, B1 => A_s(46), B2 => 
                           n1088, ZN => n152);
   U61 : OAI221_X1 port map( B1 => n1105, B2 => n1161, C1 => n1100, C2 => n1127
                           , A => n150, ZN => O_49_port);
   U62 : AOI22_X1 port map( A1 => A_ns(48), A2 => n1094, B1 => A_s(48), B2 => 
                           n1088, ZN => n150);
   U63 : OAI221_X1 port map( B1 => n1105, B2 => n1162, C1 => n1100, C2 => n1128
                           , A => n148, ZN => O_50_port);
   U64 : AOI22_X1 port map( A1 => A_ns(49), A2 => n1094, B1 => A_s(49), B2 => 
                           n1088, ZN => n148);
   U65 : OAI221_X1 port map( B1 => n1105, B2 => n1163, C1 => n1100, C2 => n1129
                           , A => n147, ZN => O_51_port);
   U66 : AOI22_X1 port map( A1 => A_ns(50), A2 => n1094, B1 => A_s(50), B2 => 
                           n1088, ZN => n147);
   U67 : OAI221_X1 port map( B1 => n1105, B2 => n1164, C1 => n1100, C2 => n1130
                           , A => n146, ZN => O_52_port);
   U68 : AOI22_X1 port map( A1 => A_ns(51), A2 => n1094, B1 => A_s(51), B2 => 
                           n1088, ZN => n146);
   U69 : OAI221_X1 port map( B1 => n1105, B2 => n1167, C1 => n1100, C2 => n1133
                           , A => n143, ZN => O_55_port);
   U70 : AOI22_X1 port map( A1 => A_ns(54), A2 => n1095, B1 => A_s(54), B2 => 
                           n1089, ZN => n143);
   U71 : OAI221_X1 port map( B1 => n1104, B2 => n1169, C1 => n1100, C2 => n1135
                           , A => n141, ZN => O_57_port);
   U72 : AOI22_X1 port map( A1 => A_ns(56), A2 => n1095, B1 => A_s(56), B2 => 
                           n1089, ZN => n141);
   U73 : OAI221_X1 port map( B1 => n1104, B2 => n1170, C1 => n1100, C2 => n1136
                           , A => n140, ZN => O_58_port);
   U74 : AOI22_X1 port map( A1 => A_ns(57), A2 => n1095, B1 => A_s(57), B2 => 
                           n1089, ZN => n140);
   U75 : OAI221_X1 port map( B1 => n1104, B2 => n1171, C1 => n1101, C2 => n1137
                           , A => n139, ZN => O_59_port);
   U76 : AOI22_X1 port map( A1 => A_ns(58), A2 => n1095, B1 => A_s(58), B2 => 
                           n1089, ZN => n139);
   U77 : BUF_X1 port map( A => n1102, Z => n1100);
   U78 : OAI221_X1 port map( B1 => n1104, B2 => n1172, C1 => n1101, C2 => n1138
                           , A => n137, ZN => O_60_port);
   U79 : AOI22_X1 port map( A1 => A_ns(59), A2 => n1095, B1 => A_s(59), B2 => 
                           n1089, ZN => n137);
   U80 : AOI22_X1 port map( A1 => A_ns(60), A2 => n1095, B1 => A_s(60), B2 => 
                           n1089, ZN => n136);
   U81 : OAI221_X1 port map( B1 => n1104, B2 => n1174, C1 => n1101, C2 => n1140
                           , A => n135, ZN => O_62_port);
   U82 : AOI22_X1 port map( A1 => A_ns(61), A2 => n1095, B1 => A_s(61), B2 => 
                           n1089, ZN => n135);
   U83 : BUF_X1 port map( A => n1102, Z => n1101);
   U84 : BUF_X1 port map( A => n1103, Z => n1097);
   U85 : BUF_X1 port map( A => n128, Z => n1107);
   U86 : NAND2_X1 port map( A1 => n194, A2 => n1236, ZN => n182);
   U87 : NAND2_X1 port map( A1 => n194, A2 => n182, ZN => n183);
   U88 : BUF_X1 port map( A => n129, Z => n1103);
   U89 : BUF_X1 port map( A => n128, Z => n1106);
   U90 : BUF_X1 port map( A => n129, Z => n1102);
   U91 : BUF_X1 port map( A => n128, Z => n1105);
   U92 : BUF_X1 port map( A => n128, Z => n1104);
   U93 : BUF_X1 port map( A => n128, Z => n1108);
   U94 : OAI221_X1 port map( B1 => n1108, B2 => n1215, C1 => n1097, C2 => n1213
                           , A => n180, ZN => O_21_port);
   U95 : INV_X1 port map( A => A_s(19), ZN => n1215);
   U96 : INV_X1 port map( A => A_ns(19), ZN => n1213);
   U97 : OAI221_X1 port map( B1 => n1108, B2 => n1218, C1 => n1097, C2 => n1216
                           , A => n179, ZN => O_22_port);
   U98 : INV_X1 port map( A => A_s(20), ZN => n1218);
   U99 : INV_X1 port map( A => A_ns(20), ZN => n1216);
   U100 : OAI221_X1 port map( B1 => n1108, B2 => n1219, C1 => n1098, C2 => 
                           n1217, A => n178, ZN => O_23_port);
   U101 : INV_X1 port map( A => A_s(21), ZN => n1219);
   U102 : INV_X1 port map( A => A_ns(21), ZN => n1217);
   U103 : OAI221_X1 port map( B1 => n1107, B2 => n1222, C1 => n1098, C2 => 
                           n1220, A => n177, ZN => O_24_port);
   U104 : INV_X1 port map( A => A_s(22), ZN => n1222);
   U105 : INV_X1 port map( A => A_ns(22), ZN => n1220);
   U106 : OAI221_X1 port map( B1 => n1107, B2 => n1223, C1 => n1098, C2 => 
                           n1221, A => n176, ZN => O_25_port);
   U107 : INV_X1 port map( A => A_s(23), ZN => n1223);
   U108 : INV_X1 port map( A => A_ns(23), ZN => n1221);
   U109 : OAI221_X1 port map( B1 => n1107, B2 => n1226, C1 => n1098, C2 => 
                           n1224, A => n175, ZN => O_26_port);
   U110 : INV_X1 port map( A => A_s(24), ZN => n1226);
   U111 : INV_X1 port map( A => A_ns(24), ZN => n1224);
   U112 : OAI221_X1 port map( B1 => n1107, B2 => n1227, C1 => n1098, C2 => 
                           n1225, A => n174, ZN => O_27_port);
   U113 : INV_X1 port map( A => A_s(25), ZN => n1227);
   U114 : INV_X1 port map( A => A_ns(25), ZN => n1225);
   U115 : OAI221_X1 port map( B1 => n1107, B2 => n1230, C1 => n1098, C2 => 
                           n1228, A => n173, ZN => O_28_port);
   U116 : INV_X1 port map( A => A_s(26), ZN => n1230);
   U117 : OAI221_X1 port map( B1 => n1107, B2 => n1233, C1 => n1098, C2 => 
                           n1232, A => n170, ZN => O_30_port);
   U118 : INV_X1 port map( A => A_s(28), ZN => n1233);
   U119 : INV_X1 port map( A => A_ns(28), ZN => n1232);
   U120 : AOI22_X1 port map( A1 => A_ns(29), A2 => n1092, B1 => A_s(29), B2 => 
                           n1086, ZN => n170);
   U121 : INV_X1 port map( A => B(31), ZN => n1236);
   U122 : OAI221_X1 port map( B1 => n1108, B2 => n1203, C1 => n1097, C2 => 
                           n1201, A => n188, ZN => O_15_port);
   U123 : INV_X1 port map( A => A_s(13), ZN => n1203);
   U124 : INV_X1 port map( A => A_ns(13), ZN => n1201);
   U125 : OAI221_X1 port map( B1 => n1108, B2 => n1206, C1 => n1097, C2 => 
                           n1204, A => n187, ZN => O_16_port);
   U126 : INV_X1 port map( A => A_s(14), ZN => n1206);
   U127 : INV_X1 port map( A => A_ns(14), ZN => n1204);
   U128 : OAI221_X1 port map( B1 => n1108, B2 => n1207, C1 => n1097, C2 => 
                           n1205, A => n186, ZN => O_17_port);
   U129 : INV_X1 port map( A => A_s(15), ZN => n1207);
   U130 : INV_X1 port map( A => A_ns(15), ZN => n1205);
   U131 : OAI221_X1 port map( B1 => n1108, B2 => n1210, C1 => n1097, C2 => 
                           n1208, A => n185, ZN => O_18_port);
   U132 : INV_X1 port map( A => A_s(16), ZN => n1210);
   U133 : INV_X1 port map( A => A_ns(16), ZN => n1208);
   U134 : OAI221_X1 port map( B1 => n1108, B2 => n1211, C1 => n1097, C2 => 
                           n1209, A => n184, ZN => O_19_port);
   U135 : INV_X1 port map( A => A_s(17), ZN => n1211);
   U136 : INV_X1 port map( A => A_ns(17), ZN => n1209);
   U137 : OAI221_X1 port map( B1 => n1108, B2 => n1214, C1 => n1097, C2 => 
                           n1212, A => n181, ZN => O_20_port);
   U138 : INV_X1 port map( A => A_s(18), ZN => n1214);
   U139 : INV_X1 port map( A => A_ns(18), ZN => n1212);
   U140 : OR3_X1 port map( A1 => B(29), A2 => B(30), A3 => n1236, ZN => n129);
   U141 : OAI221_X1 port map( B1 => n1104, B2 => n1187, C1 => n1101, C2 => 
                           n1185, A => n132, ZN => O_7_port);
   U142 : INV_X1 port map( A => A_s(5), ZN => n1187);
   U143 : INV_X1 port map( A => A_ns(5), ZN => n1185);
   U144 : OAI221_X1 port map( B1 => n1104, B2 => n1190, C1 => n1101, C2 => 
                           n1188, A => n131, ZN => O_8_port);
   U145 : INV_X1 port map( A => A_s(6), ZN => n1190);
   U146 : INV_X1 port map( A => A_ns(6), ZN => n1188);
   U147 : OAI221_X1 port map( B1 => n1104, B2 => n1191, C1 => n1101, C2 => 
                           n1189, A => n130, ZN => O_9_port);
   U148 : INV_X1 port map( A => A_s(7), ZN => n1191);
   U149 : INV_X1 port map( A => A_ns(7), ZN => n1189);
   U150 : OAI221_X1 port map( B1 => n1194, B2 => n1109, C1 => n1192, C2 => 
                           n1097, A => n193, ZN => O_10_port);
   U151 : INV_X1 port map( A => A_ns(8), ZN => n1192);
   U152 : INV_X1 port map( A => A_s(8), ZN => n1194);
   U153 : OAI221_X1 port map( B1 => n1109, B2 => n1195, C1 => n1097, C2 => 
                           n1193, A => n192, ZN => O_11_port);
   U154 : INV_X1 port map( A => A_s(9), ZN => n1195);
   U155 : INV_X1 port map( A => A_ns(9), ZN => n1193);
   U156 : OAI221_X1 port map( B1 => n1108, B2 => n1198, C1 => n1097, C2 => 
                           n1196, A => n191, ZN => O_12_port);
   U157 : INV_X1 port map( A => A_s(10), ZN => n1198);
   U158 : INV_X1 port map( A => A_ns(10), ZN => n1196);
   U159 : OAI221_X1 port map( B1 => n1108, B2 => n1199, C1 => n1097, C2 => 
                           n1197, A => n190, ZN => O_13_port);
   U160 : INV_X1 port map( A => A_s(11), ZN => n1199);
   U161 : INV_X1 port map( A => A_ns(11), ZN => n1197);
   U162 : OAI221_X1 port map( B1 => n1108, B2 => n1202, C1 => n1097, C2 => 
                           n1200, A => n189, ZN => O_14_port);
   U163 : INV_X1 port map( A => A_s(12), ZN => n1202);
   U164 : INV_X1 port map( A => A_ns(12), ZN => n1200);
   U165 : OAI22_X1 port map( A1 => n182, A2 => n1178, B1 => n183, B2 => n1176, 
                           ZN => O_1_port);
   U166 : OAI221_X1 port map( B1 => n1107, B2 => n1178, C1 => n1098, C2 => 
                           n1176, A => n171, ZN => O_2_port);
   U167 : AOI22_X1 port map( A1 => A_ns(1), A2 => n1092, B1 => A_s(1), B2 => 
                           n1086, ZN => n171);
   U168 : OAI221_X1 port map( B1 => n1106, B2 => n1179, C1 => n1099, C2 => 
                           n1177, A => n160, ZN => O_3_port);
   U169 : INV_X1 port map( A => A_s(1), ZN => n1179);
   U170 : INV_X1 port map( A => A_ns(1), ZN => n1177);
   U171 : OAI221_X1 port map( B1 => n1105, B2 => n1182, C1 => n1100, C2 => 
                           n1180, A => n149, ZN => O_4_port);
   U172 : INV_X1 port map( A => A_s(2), ZN => n1182);
   U173 : INV_X1 port map( A => A_ns(2), ZN => n1180);
   U174 : OAI221_X1 port map( B1 => n1104, B2 => n1183, C1 => n1101, C2 => 
                           n1181, A => n138, ZN => O_5_port);
   U175 : INV_X1 port map( A => A_s(3), ZN => n1183);
   U176 : INV_X1 port map( A => A_ns(3), ZN => n1181);
   U177 : OAI221_X1 port map( B1 => n1104, B2 => n1186, C1 => n1101, C2 => 
                           n1184, A => n133, ZN => O_6_port);
   U178 : INV_X1 port map( A => A_s(4), ZN => n1186);
   U179 : INV_X1 port map( A => A_ns(4), ZN => n1184);
   U180 : OAI221_X1 port map( B1 => n1107, B2 => n1231, C1 => n1098, C2 => 
                           n1229, A => n172, ZN => O_29_port);
   U181 : INV_X1 port map( A => A_s(27), ZN => n1231);
   U182 : INV_X1 port map( A => A_ns(27), ZN => n1229);
   U183 : AOI22_X1 port map( A1 => A_ns(28), A2 => n1092, B1 => A_s(28), B2 => 
                           n1086, ZN => n172);
   U184 : INV_X1 port map( A => A_ns(0), ZN => n1176);
   U185 : INV_X1 port map( A => A_s(0), ZN => n1178);
   U186 : AOI22_X1 port map( A1 => A_ns(2), A2 => n1093, B1 => A_s(2), B2 => 
                           n1087, ZN => n160);
   U187 : AOI22_X1 port map( A1 => A_ns(3), A2 => n1094, B1 => A_s(3), B2 => 
                           n1088, ZN => n149);
   U188 : AOI22_X1 port map( A1 => A_ns(4), A2 => n1095, B1 => A_s(4), B2 => 
                           n1089, ZN => n138);
   U189 : AOI22_X1 port map( A1 => A_ns(5), A2 => n1095, B1 => A_s(5), B2 => 
                           n1089, ZN => n133);
   U190 : AOI22_X1 port map( A1 => A_ns(6), A2 => n1095, B1 => A_s(6), B2 => 
                           n1089, ZN => n132);
   U191 : AOI22_X1 port map( A1 => A_ns(7), A2 => n1096, B1 => A_s(7), B2 => 
                           n1090, ZN => n131);
   U192 : AOI22_X1 port map( A1 => A_ns(8), A2 => n1096, B1 => A_s(8), B2 => 
                           n1090, ZN => n130);
   U193 : AOI22_X1 port map( A1 => A_ns(9), A2 => n1091, B1 => A_s(9), B2 => 
                           n1085, ZN => n193);
   U194 : AOI22_X1 port map( A1 => A_ns(10), A2 => n1091, B1 => A_s(10), B2 => 
                           n1085, ZN => n192);
   U195 : AOI22_X1 port map( A1 => A_ns(11), A2 => n1091, B1 => A_s(11), B2 => 
                           n1085, ZN => n191);
   U196 : AOI22_X1 port map( A1 => A_ns(12), A2 => n1091, B1 => A_s(12), B2 => 
                           n1085, ZN => n190);
   U197 : AOI22_X1 port map( A1 => A_ns(13), A2 => n1091, B1 => A_s(13), B2 => 
                           n1085, ZN => n189);
   U198 : AOI22_X1 port map( A1 => A_ns(14), A2 => n1091, B1 => A_s(14), B2 => 
                           n1085, ZN => n188);
   U199 : AOI22_X1 port map( A1 => A_ns(15), A2 => n1091, B1 => A_s(15), B2 => 
                           n1085, ZN => n187);
   U200 : AOI22_X1 port map( A1 => A_ns(16), A2 => n1091, B1 => A_s(16), B2 => 
                           n1085, ZN => n186);
   U201 : AOI22_X1 port map( A1 => A_ns(17), A2 => n1091, B1 => A_s(17), B2 => 
                           n1085, ZN => n185);
   U202 : AOI22_X1 port map( A1 => A_ns(18), A2 => n1091, B1 => A_s(18), B2 => 
                           n1085, ZN => n184);
   U203 : AOI22_X1 port map( A1 => A_ns(19), A2 => n1091, B1 => A_s(19), B2 => 
                           n1085, ZN => n181);
   U204 : AOI22_X1 port map( A1 => A_ns(20), A2 => n1091, B1 => A_s(20), B2 => 
                           n1085, ZN => n180);
   U205 : AOI22_X1 port map( A1 => A_ns(21), A2 => n1092, B1 => A_s(21), B2 => 
                           n1086, ZN => n179);
   U206 : AOI22_X1 port map( A1 => A_ns(22), A2 => n1092, B1 => A_s(22), B2 => 
                           n1086, ZN => n178);
   U207 : AOI22_X1 port map( A1 => A_ns(23), A2 => n1092, B1 => A_s(23), B2 => 
                           n1086, ZN => n177);
   U208 : AOI22_X1 port map( A1 => A_ns(24), A2 => n1092, B1 => A_s(24), B2 => 
                           n1086, ZN => n176);
   U209 : AOI22_X1 port map( A1 => A_ns(25), A2 => n1092, B1 => A_s(25), B2 => 
                           n1086, ZN => n175);
   U210 : AOI22_X1 port map( A1 => A_ns(26), A2 => n1092, B1 => A_s(26), B2 => 
                           n1086, ZN => n174);
   U211 : AOI22_X1 port map( A1 => A_ns(27), A2 => n1092, B1 => A_s(27), B2 => 
                           n1086, ZN => n173);
   U212 : INV_X1 port map( A => A_ns(26), ZN => n1228);
   U213 : CLKBUF_X1 port map( A => n1234, Z => n1090);
   U214 : CLKBUF_X1 port map( A => n1235, Z => n1096);
   U215 : CLKBUF_X1 port map( A => n128, Z => n1109);
   U216 : INV_X1 port map( A => A_ns(30), ZN => n1110);
   U217 : INV_X1 port map( A => A_ns(31), ZN => n1111);
   U218 : INV_X1 port map( A => A_ns(32), ZN => n1112);
   U219 : INV_X1 port map( A => A_ns(33), ZN => n1113);
   U220 : INV_X1 port map( A => A_ns(34), ZN => n1114);
   U221 : INV_X1 port map( A => A_ns(35), ZN => n1115);
   U222 : INV_X1 port map( A => A_ns(36), ZN => n1116);
   U223 : INV_X1 port map( A => A_ns(37), ZN => n1117);
   U224 : INV_X1 port map( A => A_ns(38), ZN => n1118);
   U225 : INV_X1 port map( A => A_ns(39), ZN => n1119);
   U226 : INV_X1 port map( A => A_ns(40), ZN => n1120);
   U227 : INV_X1 port map( A => A_ns(41), ZN => n1121);
   U228 : INV_X1 port map( A => A_ns(42), ZN => n1122);
   U229 : INV_X1 port map( A => A_ns(43), ZN => n1123);
   U230 : INV_X1 port map( A => A_ns(44), ZN => n1124);
   U231 : INV_X1 port map( A => A_ns(45), ZN => n1125);
   U232 : INV_X1 port map( A => A_ns(46), ZN => n1126);
   U233 : INV_X1 port map( A => A_ns(47), ZN => n1127);
   U234 : INV_X1 port map( A => A_ns(48), ZN => n1128);
   U235 : INV_X1 port map( A => A_ns(49), ZN => n1129);
   U236 : INV_X1 port map( A => A_ns(50), ZN => n1130);
   U237 : INV_X1 port map( A => A_ns(51), ZN => n1131);
   U238 : INV_X1 port map( A => A_ns(52), ZN => n1132);
   U239 : INV_X1 port map( A => A_ns(53), ZN => n1133);
   U240 : INV_X1 port map( A => A_ns(54), ZN => n1134);
   U241 : INV_X1 port map( A => A_ns(55), ZN => n1135);
   U242 : INV_X1 port map( A => A_ns(56), ZN => n1136);
   U243 : INV_X1 port map( A => A_ns(57), ZN => n1137);
   U244 : INV_X1 port map( A => A_ns(58), ZN => n1138);
   U245 : INV_X1 port map( A => A_ns(59), ZN => n1139);
   U246 : INV_X1 port map( A => A_ns(60), ZN => n1140);
   U247 : INV_X1 port map( A => A_ns(61), ZN => n1141);
   U248 : INV_X1 port map( A => A_ns(29), ZN => n1142);
   U249 : INV_X1 port map( A => A_s(29), ZN => n1143);
   U250 : INV_X1 port map( A => A_s(30), ZN => n1144);
   U251 : INV_X1 port map( A => A_s(31), ZN => n1145);
   U252 : INV_X1 port map( A => A_s(32), ZN => n1146);
   U253 : INV_X1 port map( A => A_s(33), ZN => n1147);
   U254 : INV_X1 port map( A => A_s(34), ZN => n1148);
   U255 : INV_X1 port map( A => A_s(35), ZN => n1149);
   U256 : INV_X1 port map( A => A_s(36), ZN => n1150);
   U259 : INV_X1 port map( A => A_s(37), ZN => n1151);
   U260 : INV_X1 port map( A => A_s(38), ZN => n1152);
   U261 : INV_X1 port map( A => A_s(39), ZN => n1153);
   U262 : INV_X1 port map( A => A_s(40), ZN => n1154);
   U263 : INV_X1 port map( A => A_s(41), ZN => n1155);
   U264 : INV_X1 port map( A => A_s(42), ZN => n1156);
   U265 : INV_X1 port map( A => A_s(43), ZN => n1157);
   U266 : INV_X1 port map( A => A_s(44), ZN => n1158);
   U267 : INV_X1 port map( A => A_s(45), ZN => n1159);
   U268 : INV_X1 port map( A => A_s(46), ZN => n1160);
   U269 : INV_X1 port map( A => A_s(47), ZN => n1161);
   U270 : INV_X1 port map( A => A_s(48), ZN => n1162);
   U271 : INV_X1 port map( A => A_s(49), ZN => n1163);
   U272 : INV_X1 port map( A => A_s(50), ZN => n1164);
   U273 : INV_X1 port map( A => A_s(51), ZN => n1165);
   U274 : INV_X1 port map( A => A_s(52), ZN => n1166);
   U275 : INV_X1 port map( A => A_s(53), ZN => n1167);
   U276 : INV_X1 port map( A => A_s(54), ZN => n1168);
   U277 : INV_X1 port map( A => A_s(55), ZN => n1169);
   U278 : INV_X1 port map( A => A_s(56), ZN => n1170);
   U279 : INV_X1 port map( A => A_s(57), ZN => n1171);
   U280 : INV_X1 port map( A => A_s(58), ZN => n1172);
   U281 : INV_X1 port map( A => A_s(59), ZN => n1173);
   U282 : INV_X1 port map( A => A_s(60), ZN => n1174);
   U283 : INV_X1 port map( A => A_s(61), ZN => n1175);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT62_i28 is

   port( A_s, A_ns, B : in std_logic_vector (61 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (61 downto 0));

end BOOTHENC_NBIT62_i28;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT62_i28 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, O_61_port, O_60_port, O_59_port, O_58_port, O_57_port,
      O_56_port, O_55_port, O_54_port, O_53_port, O_52_port, O_51_port, 
      O_50_port, O_49_port, O_48_port, O_47_port, O_46_port, O_45_port, 
      O_44_port, O_43_port, O_42_port, O_41_port, O_40_port, O_39_port, 
      O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, O_33_port, 
      O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, O_27_port, 
      O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, O_21_port, 
      O_20_port, O_19_port, O_18_port, O_17_port, O_16_port, O_15_port, 
      O_14_port, O_13_port, O_12_port, O_11_port, O_10_port, O_9_port, O_8_port
      , O_7_port, O_6_port, O_5_port, O_4_port, O_3_port, O_2_port, O_1_port, 
      n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, 
      n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, 
      n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, 
      n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, 
      n184, n185, n186, n187, n188, n1059, n1060, n1061, n1062, n1063, n1064, 
      n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, 
      n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, 
      n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, 
      n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, 
      n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, 
      n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, 
      n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, 
      n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, 
      n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, 
      n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, 
      n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, 
      n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, 
      n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, 
      n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, 
      n1205, n1206, n1207, n1208, n1209 : std_logic;

begin
   O <= ( O_61_port, O_60_port, O_59_port, O_58_port, O_57_port, O_56_port, 
      O_55_port, O_54_port, O_53_port, O_52_port, O_51_port, O_50_port, 
      O_49_port, O_48_port, O_47_port, O_46_port, O_45_port, O_44_port, 
      O_43_port, O_42_port, O_41_port, O_40_port, O_39_port, O_38_port, 
      O_37_port, O_36_port, O_35_port, O_34_port, O_33_port, O_32_port, 
      O_31_port, O_30_port, O_29_port, O_28_port, O_27_port, O_26_port, 
      O_25_port, O_24_port, O_23_port, O_22_port, O_21_port, O_20_port, 
      O_19_port, O_18_port, O_17_port, O_16_port, O_15_port, O_14_port, 
      O_13_port, O_12_port, O_11_port, O_10_port, O_9_port, O_8_port, O_7_port,
      O_6_port, O_5_port, O_4_port, O_3_port, O_2_port, O_1_port, X_Logic0_port
      );
   A_so <= ( A_s(59), A_s(58), A_s(57), A_s(56), A_s(55), A_s(54), A_s(53), 
      A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), A_s(46), A_s(45), 
      A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), A_s(38), A_s(37), 
      A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), A_s(30), A_s(29), 
      A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), A_s(22), A_s(21), 
      A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), A_s(14), A_s(13), 
      A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), A_s(6), A_s(5), A_s(4)
      , A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, X_Logic0_port );
   A_nso <= ( A_ns(59), A_ns(58), A_ns(57), A_ns(56), A_ns(55), A_ns(54), 
      A_ns(53), A_ns(52), A_ns(51), A_ns(50), A_ns(49), A_ns(48), A_ns(47), 
      A_ns(46), A_ns(45), A_ns(44), A_ns(43), A_ns(42), A_ns(41), A_ns(40), 
      A_ns(39), A_ns(38), A_ns(37), A_ns(36), A_ns(35), A_ns(34), A_ns(33), 
      A_ns(32), A_ns(31), A_ns(30), A_ns(29), A_ns(28), A_ns(27), A_ns(26), 
      A_ns(25), A_ns(24), A_ns(23), A_ns(22), A_ns(21), A_ns(20), A_ns(19), 
      A_ns(18), A_ns(17), A_ns(16), A_ns(15), A_ns(14), A_ns(13), A_ns(12), 
      A_ns(11), A_ns(10), A_ns(9), A_ns(8), A_ns(7), A_ns(6), A_ns(5), A_ns(4),
      A_ns(3), A_ns(2), A_ns(1), A_ns(0), X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U249 : XOR2_X1 port map( A => B(27), B => B(28), Z => n188);
   U250 : NAND3_X1 port map( A1 => B(28), A2 => n1209, A3 => B(27), ZN => n124)
                           ;
   U2 : OAI221_X1 port map( B1 => n1082, B2 => n1148, C1 => n1076, C2 => n1114,
                           A => n135, ZN => O_57_port);
   U3 : OAI221_X1 port map( B1 => n1082, B2 => n1150, C1 => n1077, C2 => n1116,
                           A => n133, ZN => O_59_port);
   U4 : AOI22_X1 port map( A1 => A_ns(56), A2 => n1072, B1 => A_s(56), B2 => 
                           n1065, ZN => n135);
   U5 : AOI22_X1 port map( A1 => A_ns(60), A2 => n1072, B1 => A_s(60), B2 => 
                           n1065, ZN => n130);
   U6 : BUF_X1 port map( A => n1066, Z => n1069);
   U7 : BUF_X1 port map( A => n1059, Z => n1062);
   U8 : BUF_X1 port map( A => n1066, Z => n1070);
   U9 : BUF_X1 port map( A => n1059, Z => n1063);
   U10 : BUF_X1 port map( A => n1067, Z => n1071);
   U11 : BUF_X1 port map( A => n1060, Z => n1064);
   U12 : BUF_X1 port map( A => n1067, Z => n1072);
   U13 : BUF_X1 port map( A => n1060, Z => n1065);
   U14 : BUF_X1 port map( A => n1066, Z => n1068);
   U15 : BUF_X1 port map( A => n1059, Z => n1061);
   U16 : OAI221_X1 port map( B1 => n1082, B2 => n1152, C1 => n1077, C2 => n1118
                           , A => n130, ZN => O_61_port);
   U17 : OAI221_X1 port map( B1 => n1082, B2 => n1149, C1 => n1076, C2 => n1115
                           , A => n134, ZN => O_58_port);
   U18 : AOI22_X1 port map( A1 => A_ns(57), A2 => n1072, B1 => A_s(57), B2 => 
                           n1065, ZN => n134);
   U19 : OAI221_X1 port map( B1 => n1085, B2 => n1122, C1 => n1074, C2 => n1088
                           , A => n163, ZN => O_31_port);
   U20 : AOI22_X1 port map( A1 => A_ns(30), A2 => n1069, B1 => A_s(30), B2 => 
                           n1062, ZN => n163);
   U21 : OAI221_X1 port map( B1 => n1085, B2 => n1120, C1 => n1074, C2 => n1119
                           , A => n166, ZN => O_29_port);
   U22 : AOI22_X1 port map( A1 => A_ns(28), A2 => n1069, B1 => A_s(28), B2 => 
                           n1062, ZN => n166);
   U23 : OAI221_X1 port map( B1 => n1085, B2 => n1121, C1 => n1074, C2 => n1087
                           , A => n164, ZN => O_30_port);
   U24 : AOI22_X1 port map( A1 => A_ns(29), A2 => n1069, B1 => A_s(29), B2 => 
                           n1062, ZN => n164);
   U25 : OAI221_X1 port map( B1 => n1085, B2 => n1123, C1 => n1074, C2 => n1089
                           , A => n162, ZN => O_32_port);
   U26 : AOI22_X1 port map( A1 => A_ns(31), A2 => n1069, B1 => A_s(31), B2 => 
                           n1062, ZN => n162);
   U27 : OAI221_X1 port map( B1 => n1084, B2 => n1124, C1 => n1074, C2 => n1090
                           , A => n161, ZN => O_33_port);
   U28 : AOI22_X1 port map( A1 => A_ns(32), A2 => n1070, B1 => A_s(32), B2 => 
                           n1063, ZN => n161);
   U29 : BUF_X1 port map( A => n1207, Z => n1059);
   U30 : BUF_X1 port map( A => n1208, Z => n1066);
   U31 : OAI221_X1 port map( B1 => n1084, B2 => n1125, C1 => n1074, C2 => n1091
                           , A => n160, ZN => O_34_port);
   U32 : AOI22_X1 port map( A1 => A_ns(33), A2 => n1070, B1 => A_s(33), B2 => 
                           n1063, ZN => n160);
   U33 : OAI221_X1 port map( B1 => n1084, B2 => n1127, C1 => n1075, C2 => n1093
                           , A => n158, ZN => O_36_port);
   U34 : AOI22_X1 port map( A1 => A_ns(35), A2 => n1070, B1 => A_s(35), B2 => 
                           n1063, ZN => n158);
   U35 : OAI221_X1 port map( B1 => n1084, B2 => n1130, C1 => n1075, C2 => n1096
                           , A => n155, ZN => O_39_port);
   U36 : AOI22_X1 port map( A1 => A_ns(38), A2 => n1070, B1 => A_s(38), B2 => 
                           n1063, ZN => n155);
   U37 : OAI221_X1 port map( B1 => n1084, B2 => n1129, C1 => n1075, C2 => n1095
                           , A => n156, ZN => O_38_port);
   U38 : AOI22_X1 port map( A1 => A_ns(37), A2 => n1070, B1 => A_s(37), B2 => 
                           n1063, ZN => n156);
   U39 : OAI221_X1 port map( B1 => n1084, B2 => n1132, C1 => n1075, C2 => n1098
                           , A => n152, ZN => O_41_port);
   U40 : AOI22_X1 port map( A1 => A_ns(40), A2 => n1070, B1 => A_s(40), B2 => 
                           n1063, ZN => n152);
   U41 : OAI221_X1 port map( B1 => n1084, B2 => n1131, C1 => n1075, C2 => n1097
                           , A => n153, ZN => O_40_port);
   U42 : AOI22_X1 port map( A1 => A_ns(39), A2 => n1070, B1 => A_s(39), B2 => 
                           n1063, ZN => n153);
   U43 : OAI221_X1 port map( B1 => n1084, B2 => n1126, C1 => n1075, C2 => n1092
                           , A => n159, ZN => O_35_port);
   U44 : AOI22_X1 port map( A1 => A_ns(34), A2 => n1070, B1 => A_s(34), B2 => 
                           n1063, ZN => n159);
   U45 : OAI221_X1 port map( B1 => n1084, B2 => n1133, C1 => n1075, C2 => n1099
                           , A => n151, ZN => O_42_port);
   U46 : AOI22_X1 port map( A1 => A_ns(41), A2 => n1070, B1 => A_s(41), B2 => 
                           n1063, ZN => n151);
   U47 : OAI221_X1 port map( B1 => n1083, B2 => n1135, C1 => n1075, C2 => n1101
                           , A => n149, ZN => O_44_port);
   U48 : AOI22_X1 port map( A1 => A_ns(43), A2 => n1071, B1 => A_s(43), B2 => 
                           n1064, ZN => n149);
   U49 : OAI221_X1 port map( B1 => n1083, B2 => n1137, C1 => n1075, C2 => n1103
                           , A => n147, ZN => O_46_port);
   U50 : AOI22_X1 port map( A1 => A_ns(45), A2 => n1071, B1 => A_s(45), B2 => 
                           n1064, ZN => n147);
   U51 : OAI221_X1 port map( B1 => n1083, B2 => n1139, C1 => n1076, C2 => n1105
                           , A => n145, ZN => O_48_port);
   U52 : AOI22_X1 port map( A1 => A_ns(47), A2 => n1071, B1 => A_s(47), B2 => 
                           n1064, ZN => n145);
   U53 : OAI221_X1 port map( B1 => n1084, B2 => n1128, C1 => n1075, C2 => n1094
                           , A => n157, ZN => O_37_port);
   U54 : AOI22_X1 port map( A1 => A_ns(36), A2 => n1070, B1 => A_s(36), B2 => 
                           n1063, ZN => n157);
   U55 : OAI221_X1 port map( B1 => n1084, B2 => n1134, C1 => n1075, C2 => n1100
                           , A => n150, ZN => O_43_port);
   U56 : AOI22_X1 port map( A1 => A_ns(42), A2 => n1070, B1 => A_s(42), B2 => 
                           n1063, ZN => n150);
   U57 : OAI221_X1 port map( B1 => n1083, B2 => n1136, C1 => n1075, C2 => n1102
                           , A => n148, ZN => O_45_port);
   U58 : AOI22_X1 port map( A1 => A_ns(44), A2 => n1071, B1 => A_s(44), B2 => 
                           n1064, ZN => n148);
   U59 : OAI221_X1 port map( B1 => n1083, B2 => n1138, C1 => n1076, C2 => n1104
                           , A => n146, ZN => O_47_port);
   U60 : AOI22_X1 port map( A1 => A_ns(46), A2 => n1071, B1 => A_s(46), B2 => 
                           n1064, ZN => n146);
   U61 : OAI221_X1 port map( B1 => n1083, B2 => n1140, C1 => n1076, C2 => n1106
                           , A => n144, ZN => O_49_port);
   U62 : AOI22_X1 port map( A1 => A_ns(48), A2 => n1071, B1 => A_s(48), B2 => 
                           n1064, ZN => n144);
   U63 : OAI221_X1 port map( B1 => n1083, B2 => n1142, C1 => n1076, C2 => n1108
                           , A => n141, ZN => O_51_port);
   U64 : AOI22_X1 port map( A1 => A_ns(50), A2 => n1071, B1 => A_s(50), B2 => 
                           n1064, ZN => n141);
   U65 : OAI221_X1 port map( B1 => n1082, B2 => n1147, C1 => n1076, C2 => n1113
                           , A => n136, ZN => O_56_port);
   U66 : AOI22_X1 port map( A1 => A_ns(55), A2 => n1072, B1 => A_s(55), B2 => 
                           n1065, ZN => n136);
   U67 : OAI221_X1 port map( B1 => n1082, B2 => n1146, C1 => n1076, C2 => n1112
                           , A => n137, ZN => O_55_port);
   U68 : AOI22_X1 port map( A1 => A_ns(54), A2 => n1072, B1 => A_s(54), B2 => 
                           n1065, ZN => n137);
   U69 : OAI221_X1 port map( B1 => n1083, B2 => n1144, C1 => n1076, C2 => n1110
                           , A => n139, ZN => O_53_port);
   U70 : AOI22_X1 port map( A1 => A_ns(52), A2 => n1071, B1 => A_s(52), B2 => 
                           n1064, ZN => n139);
   U71 : OAI221_X1 port map( B1 => n1083, B2 => n1141, C1 => n1076, C2 => n1107
                           , A => n142, ZN => O_50_port);
   U72 : AOI22_X1 port map( A1 => A_ns(49), A2 => n1071, B1 => A_s(49), B2 => 
                           n1064, ZN => n142);
   U73 : OAI221_X1 port map( B1 => n1083, B2 => n1143, C1 => n1076, C2 => n1109
                           , A => n140, ZN => O_52_port);
   U74 : AOI22_X1 port map( A1 => A_ns(51), A2 => n1071, B1 => A_s(51), B2 => 
                           n1064, ZN => n140);
   U75 : OAI221_X1 port map( B1 => n1083, B2 => n1145, C1 => n1076, C2 => n1111
                           , A => n138, ZN => O_54_port);
   U76 : AOI22_X1 port map( A1 => A_ns(53), A2 => n1071, B1 => A_s(53), B2 => 
                           n1064, ZN => n138);
   U77 : AOI22_X1 port map( A1 => A_ns(58), A2 => n1072, B1 => A_s(58), B2 => 
                           n1065, ZN => n133);
   U78 : OAI221_X1 port map( B1 => n1082, B2 => n1151, C1 => n1077, C2 => n1117
                           , A => n131, ZN => O_60_port);
   U79 : AOI22_X1 port map( A1 => A_ns(59), A2 => n1072, B1 => A_s(59), B2 => 
                           n1065, ZN => n131);
   U80 : BUF_X1 port map( A => n1207, Z => n1060);
   U81 : BUF_X1 port map( A => n1208, Z => n1067);
   U82 : INV_X1 port map( A => n176, ZN => n1207);
   U83 : INV_X1 port map( A => n177, ZN => n1208);
   U84 : BUF_X1 port map( A => n1081, Z => n1085);
   U85 : BUF_X1 port map( A => n1080, Z => n1084);
   U86 : BUF_X1 port map( A => n1079, Z => n1074);
   U87 : BUF_X1 port map( A => n1078, Z => n1075);
   U88 : BUF_X1 port map( A => n1080, Z => n1083);
   U89 : BUF_X1 port map( A => n1078, Z => n1076);
   U90 : BUF_X1 port map( A => n1080, Z => n1082);
   U91 : BUF_X1 port map( A => n1078, Z => n1077);
   U92 : BUF_X1 port map( A => n1081, Z => n1086);
   U93 : BUF_X1 port map( A => n1079, Z => n1073);
   U94 : NAND2_X1 port map( A1 => n188, A2 => n1209, ZN => n176);
   U95 : NAND2_X1 port map( A1 => n188, A2 => n176, ZN => n177);
   U96 : BUF_X1 port map( A => n124, Z => n1080);
   U97 : BUF_X1 port map( A => n125, Z => n1078);
   U98 : BUF_X1 port map( A => n124, Z => n1081);
   U99 : BUF_X1 port map( A => n125, Z => n1079);
   U100 : OAI221_X1 port map( B1 => n1085, B2 => n1206, C1 => n1074, C2 => 
                           n1205, A => n167, ZN => O_28_port);
   U101 : INV_X1 port map( A => A_s(26), ZN => n1206);
   U102 : INV_X1 port map( A => A_ns(26), ZN => n1205);
   U103 : AOI22_X1 port map( A1 => A_ns(27), A2 => n1069, B1 => A_s(27), B2 => 
                           n1062, ZN => n167);
   U104 : OAI221_X1 port map( B1 => n1086, B2 => n1192, C1 => n1073, C2 => 
                           n1190, A => n174, ZN => O_21_port);
   U105 : INV_X1 port map( A => A_s(19), ZN => n1192);
   U106 : INV_X1 port map( A => A_ns(19), ZN => n1190);
   U107 : OAI221_X1 port map( B1 => n1085, B2 => n1195, C1 => n1073, C2 => 
                           n1193, A => n173, ZN => O_22_port);
   U108 : INV_X1 port map( A => A_s(20), ZN => n1195);
   U109 : INV_X1 port map( A => A_ns(20), ZN => n1193);
   U110 : OAI221_X1 port map( B1 => n1085, B2 => n1196, C1 => n1074, C2 => 
                           n1194, A => n172, ZN => O_23_port);
   U111 : INV_X1 port map( A => A_s(21), ZN => n1196);
   U112 : INV_X1 port map( A => A_ns(21), ZN => n1194);
   U113 : OAI221_X1 port map( B1 => n1085, B2 => n1199, C1 => n1074, C2 => 
                           n1197, A => n171, ZN => O_24_port);
   U114 : INV_X1 port map( A => A_s(22), ZN => n1199);
   U115 : INV_X1 port map( A => A_ns(22), ZN => n1197);
   U116 : OAI221_X1 port map( B1 => n1085, B2 => n1200, C1 => n1074, C2 => 
                           n1198, A => n170, ZN => O_25_port);
   U117 : INV_X1 port map( A => A_s(23), ZN => n1200);
   U118 : INV_X1 port map( A => A_ns(23), ZN => n1198);
   U119 : OAI221_X1 port map( B1 => n1085, B2 => n1203, C1 => n1074, C2 => 
                           n1201, A => n169, ZN => O_26_port);
   U120 : INV_X1 port map( A => A_s(24), ZN => n1203);
   U121 : OAI221_X1 port map( B1 => n1085, B2 => n1204, C1 => n1074, C2 => 
                           n1202, A => n168, ZN => O_27_port);
   U122 : INV_X1 port map( A => A_s(25), ZN => n1204);
   U123 : INV_X1 port map( A => B(29), ZN => n1209);
   U124 : OAI221_X1 port map( B1 => n1086, B2 => n1180, C1 => n1073, C2 => 
                           n1178, A => n182, ZN => O_15_port);
   U125 : INV_X1 port map( A => A_s(13), ZN => n1180);
   U126 : INV_X1 port map( A => A_ns(13), ZN => n1178);
   U127 : OAI221_X1 port map( B1 => n1086, B2 => n1183, C1 => n1073, C2 => 
                           n1181, A => n181, ZN => O_16_port);
   U128 : INV_X1 port map( A => A_s(14), ZN => n1183);
   U129 : INV_X1 port map( A => A_ns(14), ZN => n1181);
   U130 : OAI221_X1 port map( B1 => n1086, B2 => n1184, C1 => n1073, C2 => 
                           n1182, A => n180, ZN => O_17_port);
   U131 : INV_X1 port map( A => A_s(15), ZN => n1184);
   U132 : INV_X1 port map( A => A_ns(15), ZN => n1182);
   U133 : OAI221_X1 port map( B1 => n1086, B2 => n1187, C1 => n1073, C2 => 
                           n1185, A => n179, ZN => O_18_port);
   U134 : INV_X1 port map( A => A_s(16), ZN => n1187);
   U135 : INV_X1 port map( A => A_ns(16), ZN => n1185);
   U136 : OAI221_X1 port map( B1 => n1086, B2 => n1188, C1 => n1073, C2 => 
                           n1186, A => n178, ZN => O_19_port);
   U137 : INV_X1 port map( A => A_s(17), ZN => n1188);
   U138 : INV_X1 port map( A => A_ns(17), ZN => n1186);
   U139 : OAI221_X1 port map( B1 => n1086, B2 => n1191, C1 => n1073, C2 => 
                           n1189, A => n175, ZN => O_20_port);
   U140 : INV_X1 port map( A => A_s(18), ZN => n1191);
   U141 : INV_X1 port map( A => A_ns(18), ZN => n1189);
   U142 : OR3_X1 port map( A1 => B(27), A2 => B(28), A3 => n1209, ZN => n125);
   U143 : OAI221_X1 port map( B1 => n1082, B2 => n1164, C1 => n1077, C2 => 
                           n1162, A => n128, ZN => O_7_port);
   U144 : INV_X1 port map( A => A_s(5), ZN => n1164);
   U145 : INV_X1 port map( A => A_ns(5), ZN => n1162);
   U146 : OAI221_X1 port map( B1 => n1082, B2 => n1167, C1 => n1077, C2 => 
                           n1165, A => n127, ZN => O_8_port);
   U147 : INV_X1 port map( A => A_s(6), ZN => n1167);
   U148 : INV_X1 port map( A => A_ns(6), ZN => n1165);
   U149 : OAI221_X1 port map( B1 => n1082, B2 => n1168, C1 => n1077, C2 => 
                           n1166, A => n126, ZN => O_9_port);
   U150 : INV_X1 port map( A => A_s(7), ZN => n1168);
   U151 : INV_X1 port map( A => A_ns(7), ZN => n1166);
   U152 : OAI221_X1 port map( B1 => n1171, B2 => n1086, C1 => n1169, C2 => 
                           n1073, A => n187, ZN => O_10_port);
   U153 : INV_X1 port map( A => A_ns(8), ZN => n1169);
   U154 : INV_X1 port map( A => A_s(8), ZN => n1171);
   U155 : OAI221_X1 port map( B1 => n1086, B2 => n1172, C1 => n1073, C2 => 
                           n1170, A => n186, ZN => O_11_port);
   U156 : INV_X1 port map( A => A_s(9), ZN => n1172);
   U157 : INV_X1 port map( A => A_ns(9), ZN => n1170);
   U158 : OAI221_X1 port map( B1 => n1086, B2 => n1175, C1 => n1073, C2 => 
                           n1173, A => n185, ZN => O_12_port);
   U159 : INV_X1 port map( A => A_s(10), ZN => n1175);
   U160 : INV_X1 port map( A => A_ns(10), ZN => n1173);
   U161 : OAI221_X1 port map( B1 => n1086, B2 => n1176, C1 => n1073, C2 => 
                           n1174, A => n184, ZN => O_13_port);
   U162 : INV_X1 port map( A => A_s(11), ZN => n1176);
   U163 : INV_X1 port map( A => A_ns(11), ZN => n1174);
   U164 : OAI221_X1 port map( B1 => n1086, B2 => n1179, C1 => n1073, C2 => 
                           n1177, A => n183, ZN => O_14_port);
   U165 : INV_X1 port map( A => A_s(12), ZN => n1179);
   U166 : INV_X1 port map( A => A_ns(12), ZN => n1177);
   U167 : OAI22_X1 port map( A1 => n176, A2 => n1155, B1 => n177, B2 => n1153, 
                           ZN => O_1_port);
   U168 : OAI221_X1 port map( B1 => n1085, B2 => n1155, C1 => n1074, C2 => 
                           n1153, A => n165, ZN => O_2_port);
   U169 : AOI22_X1 port map( A1 => A_ns(1), A2 => n1069, B1 => A_s(1), B2 => 
                           n1062, ZN => n165);
   U170 : OAI221_X1 port map( B1 => n1084, B2 => n1156, C1 => n1075, C2 => 
                           n1154, A => n154, ZN => O_3_port);
   U171 : INV_X1 port map( A => A_s(1), ZN => n1156);
   U172 : INV_X1 port map( A => A_ns(1), ZN => n1154);
   U173 : OAI221_X1 port map( B1 => n1083, B2 => n1159, C1 => n1076, C2 => 
                           n1157, A => n143, ZN => O_4_port);
   U174 : INV_X1 port map( A => A_s(2), ZN => n1159);
   U175 : INV_X1 port map( A => A_ns(2), ZN => n1157);
   U176 : OAI221_X1 port map( B1 => n1082, B2 => n1160, C1 => n1077, C2 => 
                           n1158, A => n132, ZN => O_5_port);
   U177 : INV_X1 port map( A => A_s(3), ZN => n1160);
   U178 : INV_X1 port map( A => A_ns(3), ZN => n1158);
   U179 : OAI221_X1 port map( B1 => n1082, B2 => n1163, C1 => n1077, C2 => 
                           n1161, A => n129, ZN => O_6_port);
   U180 : INV_X1 port map( A => A_s(4), ZN => n1163);
   U181 : INV_X1 port map( A => A_ns(4), ZN => n1161);
   U182 : INV_X1 port map( A => A_ns(0), ZN => n1153);
   U183 : INV_X1 port map( A => A_s(0), ZN => n1155);
   U184 : AOI22_X1 port map( A1 => A_ns(2), A2 => n1070, B1 => A_s(2), B2 => 
                           n1063, ZN => n154);
   U185 : AOI22_X1 port map( A1 => A_ns(3), A2 => n1071, B1 => A_s(3), B2 => 
                           n1064, ZN => n143);
   U186 : AOI22_X1 port map( A1 => A_ns(4), A2 => n1072, B1 => A_s(4), B2 => 
                           n1065, ZN => n132);
   U187 : AOI22_X1 port map( A1 => A_ns(5), A2 => n1072, B1 => A_s(5), B2 => 
                           n1065, ZN => n129);
   U188 : AOI22_X1 port map( A1 => A_ns(6), A2 => n1072, B1 => A_s(6), B2 => 
                           n1065, ZN => n128);
   U189 : AOI22_X1 port map( A1 => A_ns(7), A2 => n1072, B1 => A_s(7), B2 => 
                           n1065, ZN => n127);
   U190 : AOI22_X1 port map( A1 => A_ns(8), A2 => n1072, B1 => A_s(8), B2 => 
                           n1065, ZN => n126);
   U191 : AOI22_X1 port map( A1 => A_ns(9), A2 => n1068, B1 => A_s(9), B2 => 
                           n1061, ZN => n187);
   U192 : AOI22_X1 port map( A1 => A_ns(10), A2 => n1068, B1 => A_s(10), B2 => 
                           n1061, ZN => n186);
   U193 : AOI22_X1 port map( A1 => A_ns(11), A2 => n1068, B1 => A_s(11), B2 => 
                           n1061, ZN => n185);
   U194 : AOI22_X1 port map( A1 => A_ns(12), A2 => n1068, B1 => A_s(12), B2 => 
                           n1061, ZN => n184);
   U195 : AOI22_X1 port map( A1 => A_ns(13), A2 => n1068, B1 => A_s(13), B2 => 
                           n1061, ZN => n183);
   U196 : AOI22_X1 port map( A1 => A_ns(14), A2 => n1068, B1 => A_s(14), B2 => 
                           n1061, ZN => n182);
   U197 : AOI22_X1 port map( A1 => A_ns(15), A2 => n1068, B1 => A_s(15), B2 => 
                           n1061, ZN => n181);
   U198 : AOI22_X1 port map( A1 => A_ns(16), A2 => n1068, B1 => A_s(16), B2 => 
                           n1061, ZN => n180);
   U199 : AOI22_X1 port map( A1 => A_ns(17), A2 => n1068, B1 => A_s(17), B2 => 
                           n1061, ZN => n179);
   U200 : AOI22_X1 port map( A1 => A_ns(18), A2 => n1068, B1 => A_s(18), B2 => 
                           n1061, ZN => n178);
   U201 : AOI22_X1 port map( A1 => A_ns(19), A2 => n1068, B1 => A_s(19), B2 => 
                           n1061, ZN => n175);
   U202 : AOI22_X1 port map( A1 => A_ns(20), A2 => n1068, B1 => A_s(20), B2 => 
                           n1061, ZN => n174);
   U203 : AOI22_X1 port map( A1 => A_ns(21), A2 => n1069, B1 => A_s(21), B2 => 
                           n1062, ZN => n173);
   U204 : AOI22_X1 port map( A1 => A_ns(22), A2 => n1069, B1 => A_s(22), B2 => 
                           n1062, ZN => n172);
   U205 : AOI22_X1 port map( A1 => A_ns(23), A2 => n1069, B1 => A_s(23), B2 => 
                           n1062, ZN => n171);
   U206 : AOI22_X1 port map( A1 => A_ns(24), A2 => n1069, B1 => A_s(24), B2 => 
                           n1062, ZN => n170);
   U207 : AOI22_X1 port map( A1 => A_ns(25), A2 => n1069, B1 => A_s(25), B2 => 
                           n1062, ZN => n169);
   U208 : AOI22_X1 port map( A1 => A_ns(26), A2 => n1069, B1 => A_s(26), B2 => 
                           n1062, ZN => n168);
   U209 : INV_X1 port map( A => A_ns(24), ZN => n1201);
   U210 : INV_X1 port map( A => A_ns(25), ZN => n1202);
   U211 : INV_X1 port map( A => A_ns(28), ZN => n1087);
   U212 : INV_X1 port map( A => A_ns(29), ZN => n1088);
   U213 : INV_X1 port map( A => A_ns(30), ZN => n1089);
   U214 : INV_X1 port map( A => A_ns(31), ZN => n1090);
   U215 : INV_X1 port map( A => A_ns(32), ZN => n1091);
   U216 : INV_X1 port map( A => A_ns(33), ZN => n1092);
   U217 : INV_X1 port map( A => A_ns(34), ZN => n1093);
   U218 : INV_X1 port map( A => A_ns(35), ZN => n1094);
   U219 : INV_X1 port map( A => A_ns(36), ZN => n1095);
   U220 : INV_X1 port map( A => A_ns(37), ZN => n1096);
   U221 : INV_X1 port map( A => A_ns(38), ZN => n1097);
   U222 : INV_X1 port map( A => A_ns(39), ZN => n1098);
   U223 : INV_X1 port map( A => A_ns(40), ZN => n1099);
   U224 : INV_X1 port map( A => A_ns(41), ZN => n1100);
   U225 : INV_X1 port map( A => A_ns(42), ZN => n1101);
   U226 : INV_X1 port map( A => A_ns(43), ZN => n1102);
   U227 : INV_X1 port map( A => A_ns(44), ZN => n1103);
   U228 : INV_X1 port map( A => A_ns(45), ZN => n1104);
   U229 : INV_X1 port map( A => A_ns(46), ZN => n1105);
   U230 : INV_X1 port map( A => A_ns(47), ZN => n1106);
   U231 : INV_X1 port map( A => A_ns(48), ZN => n1107);
   U232 : INV_X1 port map( A => A_ns(49), ZN => n1108);
   U233 : INV_X1 port map( A => A_ns(50), ZN => n1109);
   U234 : INV_X1 port map( A => A_ns(51), ZN => n1110);
   U235 : INV_X1 port map( A => A_ns(52), ZN => n1111);
   U236 : INV_X1 port map( A => A_ns(53), ZN => n1112);
   U237 : INV_X1 port map( A => A_ns(54), ZN => n1113);
   U238 : INV_X1 port map( A => A_ns(55), ZN => n1114);
   U239 : INV_X1 port map( A => A_ns(56), ZN => n1115);
   U240 : INV_X1 port map( A => A_ns(57), ZN => n1116);
   U241 : INV_X1 port map( A => A_ns(58), ZN => n1117);
   U242 : INV_X1 port map( A => A_ns(59), ZN => n1118);
   U243 : INV_X1 port map( A => A_ns(27), ZN => n1119);
   U244 : INV_X1 port map( A => A_s(27), ZN => n1120);
   U245 : INV_X1 port map( A => A_s(28), ZN => n1121);
   U246 : INV_X1 port map( A => A_s(29), ZN => n1122);
   U247 : INV_X1 port map( A => A_s(30), ZN => n1123);
   U248 : INV_X1 port map( A => A_s(31), ZN => n1124);
   U251 : INV_X1 port map( A => A_s(32), ZN => n1125);
   U252 : INV_X1 port map( A => A_s(33), ZN => n1126);
   U253 : INV_X1 port map( A => A_s(34), ZN => n1127);
   U254 : INV_X1 port map( A => A_s(35), ZN => n1128);
   U255 : INV_X1 port map( A => A_s(36), ZN => n1129);
   U256 : INV_X1 port map( A => A_s(37), ZN => n1130);
   U257 : INV_X1 port map( A => A_s(38), ZN => n1131);
   U258 : INV_X1 port map( A => A_s(39), ZN => n1132);
   U259 : INV_X1 port map( A => A_s(40), ZN => n1133);
   U260 : INV_X1 port map( A => A_s(41), ZN => n1134);
   U261 : INV_X1 port map( A => A_s(42), ZN => n1135);
   U262 : INV_X1 port map( A => A_s(43), ZN => n1136);
   U263 : INV_X1 port map( A => A_s(44), ZN => n1137);
   U264 : INV_X1 port map( A => A_s(45), ZN => n1138);
   U265 : INV_X1 port map( A => A_s(46), ZN => n1139);
   U266 : INV_X1 port map( A => A_s(47), ZN => n1140);
   U267 : INV_X1 port map( A => A_s(48), ZN => n1141);
   U268 : INV_X1 port map( A => A_s(49), ZN => n1142);
   U269 : INV_X1 port map( A => A_s(50), ZN => n1143);
   U270 : INV_X1 port map( A => A_s(51), ZN => n1144);
   U271 : INV_X1 port map( A => A_s(52), ZN => n1145);
   U272 : INV_X1 port map( A => A_s(53), ZN => n1146);
   U273 : INV_X1 port map( A => A_s(54), ZN => n1147);
   U274 : INV_X1 port map( A => A_s(55), ZN => n1148);
   U275 : INV_X1 port map( A => A_s(56), ZN => n1149);
   U276 : INV_X1 port map( A => A_s(57), ZN => n1150);
   U277 : INV_X1 port map( A => A_s(58), ZN => n1151);
   U278 : INV_X1 port map( A => A_s(59), ZN => n1152);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT60_i26 is

   port( A_s, A_ns, B : in std_logic_vector (59 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (59 downto 0));

end BOOTHENC_NBIT60_i26;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT60_i26 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, O_59_port, O_58_port, O_57_port, O_56_port, O_55_port,
      O_54_port, O_53_port, O_52_port, O_51_port, O_50_port, O_49_port, 
      O_48_port, O_47_port, O_46_port, O_45_port, O_44_port, O_43_port, 
      O_42_port, O_41_port, O_40_port, O_39_port, O_38_port, O_37_port, 
      O_36_port, O_35_port, O_34_port, O_33_port, O_32_port, O_31_port, 
      O_30_port, O_29_port, O_28_port, O_27_port, O_26_port, O_25_port, 
      O_24_port, O_23_port, O_22_port, O_21_port, O_20_port, O_19_port, 
      O_18_port, O_17_port, O_16_port, O_15_port, O_14_port, O_13_port, 
      O_12_port, O_11_port, O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, 
      O_5_port, O_4_port, O_3_port, O_2_port, O_1_port, n120, n121, n122, n123,
      n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, 
      n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, 
      n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, 
      n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n1027, 
      n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, 
      n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, 
      n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, 
      n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, 
      n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, 
      n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, 
      n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, 
      n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, 
      n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, 
      n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, 
      n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, 
      n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, 
      n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, 
      n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, 
      n1168, n1169, n1170, n1171, n1172, n1173 : std_logic;

begin
   O <= ( O_59_port, O_58_port, O_57_port, O_56_port, O_55_port, O_54_port, 
      O_53_port, O_52_port, O_51_port, O_50_port, O_49_port, O_48_port, 
      O_47_port, O_46_port, O_45_port, O_44_port, O_43_port, O_42_port, 
      O_41_port, O_40_port, O_39_port, O_38_port, O_37_port, O_36_port, 
      O_35_port, O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, 
      O_29_port, O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, 
      O_23_port, O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, 
      O_17_port, O_16_port, O_15_port, O_14_port, O_13_port, O_12_port, 
      O_11_port, O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, 
      O_4_port, O_3_port, O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(57), A_s(56), A_s(55), A_s(54), A_s(53), A_s(52), A_s(51), 
      A_s(50), A_s(49), A_s(48), A_s(47), A_s(46), A_s(45), A_s(44), A_s(43), 
      A_s(42), A_s(41), A_s(40), A_s(39), A_s(38), A_s(37), A_s(36), A_s(35), 
      A_s(34), A_s(33), A_s(32), A_s(31), A_s(30), A_s(29), A_s(28), A_s(27), 
      A_s(26), A_s(25), A_s(24), A_s(23), A_s(22), A_s(21), A_s(20), A_s(19), 
      A_s(18), A_s(17), A_s(16), A_s(15), A_s(14), A_s(13), A_s(12), A_s(11), 
      A_s(10), A_s(9), A_s(8), A_s(7), A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), 
      A_s(1), A_s(0), X_Logic0_port, X_Logic0_port );
   A_nso <= ( A_ns(57), A_ns(56), A_ns(55), A_ns(54), A_ns(53), A_ns(52), 
      A_ns(51), A_ns(50), A_ns(49), A_ns(48), A_ns(47), A_ns(46), A_ns(45), 
      A_ns(44), A_ns(43), A_ns(42), A_ns(41), A_ns(40), A_ns(39), A_ns(38), 
      A_ns(37), A_ns(36), A_ns(35), A_ns(34), A_ns(33), A_ns(32), A_ns(31), 
      A_ns(30), A_ns(29), A_ns(28), A_ns(27), A_ns(26), A_ns(25), A_ns(24), 
      A_ns(23), A_ns(22), A_ns(21), A_ns(20), A_ns(19), A_ns(18), A_ns(17), 
      A_ns(16), A_ns(15), A_ns(14), A_ns(13), A_ns(12), A_ns(11), A_ns(10), 
      A_ns(9), A_ns(8), A_ns(7), A_ns(6), A_ns(5), A_ns(4), A_ns(3), A_ns(2), 
      A_ns(1), A_ns(0), X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U241 : XOR2_X1 port map( A => B(25), B => B(26), Z => n182);
   U242 : NAND3_X1 port map( A1 => B(26), A2 => n1173, A3 => B(25), ZN => n120)
                           ;
   U2 : OAI221_X1 port map( B1 => n1053, B2 => n1090, C1 => n1042, C2 => n1056,
                           A => n160, ZN => O_29_port);
   U3 : OAI221_X1 port map( B1 => n1053, B2 => n1091, C1 => n1042, C2 => n1057,
                           A => n158, ZN => O_30_port);
   U4 : OAI221_X1 port map( B1 => n1052, B2 => n1099, C1 => n1043, C2 => n1065,
                           A => n150, ZN => O_38_port);
   U5 : OAI221_X1 port map( B1 => n1051, B2 => n1105, C1 => n1043, C2 => n1071,
                           A => n143, ZN => O_44_port);
   U6 : AOI22_X1 port map( A1 => A_ns(28), A2 => n1037, B1 => A_s(28), B2 => 
                           n1030, ZN => n160);
   U7 : AOI22_X1 port map( A1 => A_ns(58), A2 => n1040, B1 => A_s(58), B2 => 
                           n1033, ZN => n127);
   U8 : BUF_X1 port map( A => n1034, Z => n1037);
   U9 : BUF_X1 port map( A => n1027, Z => n1030);
   U10 : BUF_X1 port map( A => n1034, Z => n1038);
   U11 : BUF_X1 port map( A => n1027, Z => n1031);
   U12 : BUF_X1 port map( A => n1035, Z => n1039);
   U13 : BUF_X1 port map( A => n1028, Z => n1032);
   U14 : BUF_X1 port map( A => n1035, Z => n1040);
   U15 : BUF_X1 port map( A => n1028, Z => n1033);
   U16 : BUF_X1 port map( A => n1034, Z => n1036);
   U17 : BUF_X1 port map( A => n1027, Z => n1029);
   U18 : OAI221_X1 port map( B1 => n1050, B2 => n1120, C1 => n1045, C2 => n1086
                           , A => n127, ZN => O_59_port);
   U19 : AOI22_X1 port map( A1 => A_ns(29), A2 => n1037, B1 => A_s(29), B2 => 
                           n1030, ZN => n158);
   U20 : OAI221_X1 port map( B1 => n1052, B2 => n1096, C1 => n1043, C2 => n1062
                           , A => n153, ZN => O_35_port);
   U21 : AOI22_X1 port map( A1 => A_ns(34), A2 => n1038, B1 => A_s(34), B2 => 
                           n1031, ZN => n153);
   U22 : OAI221_X1 port map( B1 => n1052, B2 => n1095, C1 => n1042, C2 => n1061
                           , A => n154, ZN => O_34_port);
   U23 : AOI22_X1 port map( A1 => A_ns(33), A2 => n1038, B1 => A_s(33), B2 => 
                           n1031, ZN => n154);
   U24 : OAI221_X1 port map( B1 => n1053, B2 => n1088, C1 => n1042, C2 => n1087
                           , A => n162, ZN => O_27_port);
   U25 : AOI22_X1 port map( A1 => A_ns(26), A2 => n1037, B1 => A_s(26), B2 => 
                           n1030, ZN => n162);
   U26 : OAI221_X1 port map( B1 => n1052, B2 => n1093, C1 => n1042, C2 => n1059
                           , A => n156, ZN => O_32_port);
   U27 : AOI22_X1 port map( A1 => A_ns(31), A2 => n1037, B1 => A_s(31), B2 => 
                           n1030, ZN => n156);
   U28 : OAI221_X1 port map( B1 => n1052, B2 => n1097, C1 => n1043, C2 => n1063
                           , A => n152, ZN => O_36_port);
   U29 : AOI22_X1 port map( A1 => A_ns(35), A2 => n1038, B1 => A_s(35), B2 => 
                           n1031, ZN => n152);
   U30 : OAI221_X1 port map( B1 => n1052, B2 => n1092, C1 => n1042, C2 => n1058
                           , A => n157, ZN => O_31_port);
   U31 : AOI22_X1 port map( A1 => A_ns(30), A2 => n1037, B1 => A_s(30), B2 => 
                           n1030, ZN => n157);
   U32 : OAI221_X1 port map( B1 => n1052, B2 => n1094, C1 => n1042, C2 => n1060
                           , A => n155, ZN => O_33_port);
   U33 : AOI22_X1 port map( A1 => A_ns(32), A2 => n1038, B1 => A_s(32), B2 => 
                           n1031, ZN => n155);
   U34 : OAI221_X1 port map( B1 => n1053, B2 => n1089, C1 => n1042, C2 => n1055
                           , A => n161, ZN => O_28_port);
   U35 : AOI22_X1 port map( A1 => A_ns(27), A2 => n1037, B1 => A_s(27), B2 => 
                           n1030, ZN => n161);
   U36 : BUF_X1 port map( A => n1171, Z => n1027);
   U37 : BUF_X1 port map( A => n1172, Z => n1034);
   U38 : OAI221_X1 port map( B1 => n1051, B2 => n1112, C1 => n1044, C2 => n1078
                           , A => n135, ZN => O_51_port);
   U39 : AOI22_X1 port map( A1 => A_ns(50), A2 => n1039, B1 => A_s(50), B2 => 
                           n1032, ZN => n135);
   U40 : OAI221_X1 port map( B1 => n1052, B2 => n1102, C1 => n1043, C2 => n1068
                           , A => n146, ZN => O_41_port);
   U41 : AOI22_X1 port map( A1 => A_ns(40), A2 => n1038, B1 => A_s(40), B2 => 
                           n1031, ZN => n146);
   U42 : OAI221_X1 port map( B1 => n1051, B2 => n1104, C1 => n1043, C2 => n1070
                           , A => n144, ZN => O_43_port);
   U43 : AOI22_X1 port map( A1 => A_ns(42), A2 => n1038, B1 => A_s(42), B2 => 
                           n1031, ZN => n144);
   U44 : AOI22_X1 port map( A1 => A_ns(37), A2 => n1038, B1 => A_s(37), B2 => 
                           n1031, ZN => n150);
   U45 : AOI22_X1 port map( A1 => A_ns(43), A2 => n1039, B1 => A_s(43), B2 => 
                           n1032, ZN => n143);
   U46 : OAI221_X1 port map( B1 => n1051, B2 => n1108, C1 => n1044, C2 => n1074
                           , A => n140, ZN => O_47_port);
   U47 : AOI22_X1 port map( A1 => A_ns(46), A2 => n1039, B1 => A_s(46), B2 => 
                           n1032, ZN => n140);
   U48 : OAI221_X1 port map( B1 => n1051, B2 => n1110, C1 => n1044, C2 => n1076
                           , A => n138, ZN => O_49_port);
   U49 : AOI22_X1 port map( A1 => A_ns(48), A2 => n1039, B1 => A_s(48), B2 => 
                           n1032, ZN => n138);
   U50 : OAI221_X1 port map( B1 => n1051, B2 => n1103, C1 => n1043, C2 => n1069
                           , A => n145, ZN => O_42_port);
   U51 : AOI22_X1 port map( A1 => A_ns(41), A2 => n1038, B1 => A_s(41), B2 => 
                           n1031, ZN => n145);
   U52 : OAI221_X1 port map( B1 => n1052, B2 => n1101, C1 => n1043, C2 => n1067
                           , A => n147, ZN => O_40_port);
   U53 : AOI22_X1 port map( A1 => A_ns(39), A2 => n1038, B1 => A_s(39), B2 => 
                           n1031, ZN => n147);
   U54 : OAI221_X1 port map( B1 => n1051, B2 => n1107, C1 => n1043, C2 => n1073
                           , A => n141, ZN => O_46_port);
   U55 : AOI22_X1 port map( A1 => A_ns(45), A2 => n1039, B1 => A_s(45), B2 => 
                           n1032, ZN => n141);
   U56 : OAI221_X1 port map( B1 => n1051, B2 => n1109, C1 => n1044, C2 => n1075
                           , A => n139, ZN => O_48_port);
   U57 : AOI22_X1 port map( A1 => A_ns(47), A2 => n1039, B1 => A_s(47), B2 => 
                           n1032, ZN => n139);
   U58 : OAI221_X1 port map( B1 => n1051, B2 => n1111, C1 => n1044, C2 => n1077
                           , A => n136, ZN => O_50_port);
   U59 : AOI22_X1 port map( A1 => A_ns(49), A2 => n1039, B1 => A_s(49), B2 => 
                           n1032, ZN => n136);
   U60 : OAI221_X1 port map( B1 => n1052, B2 => n1098, C1 => n1043, C2 => n1064
                           , A => n151, ZN => O_37_port);
   U61 : AOI22_X1 port map( A1 => A_ns(36), A2 => n1038, B1 => A_s(36), B2 => 
                           n1031, ZN => n151);
   U62 : OAI221_X1 port map( B1 => n1052, B2 => n1100, C1 => n1043, C2 => n1066
                           , A => n149, ZN => O_39_port);
   U63 : AOI22_X1 port map( A1 => A_ns(38), A2 => n1038, B1 => A_s(38), B2 => 
                           n1031, ZN => n149);
   U64 : OAI221_X1 port map( B1 => n1051, B2 => n1106, C1 => n1043, C2 => n1072
                           , A => n142, ZN => O_45_port);
   U65 : AOI22_X1 port map( A1 => A_ns(44), A2 => n1039, B1 => A_s(44), B2 => 
                           n1032, ZN => n142);
   U66 : OAI221_X1 port map( B1 => n1050, B2 => n1117, C1 => n1044, C2 => n1083
                           , A => n130, ZN => O_56_port);
   U67 : AOI22_X1 port map( A1 => A_ns(55), A2 => n1040, B1 => A_s(55), B2 => 
                           n1033, ZN => n130);
   U68 : OAI221_X1 port map( B1 => n1050, B2 => n1118, C1 => n1044, C2 => n1084
                           , A => n129, ZN => O_57_port);
   U69 : AOI22_X1 port map( A1 => A_ns(56), A2 => n1040, B1 => A_s(56), B2 => 
                           n1033, ZN => n129);
   U70 : OAI221_X1 port map( B1 => n1051, B2 => n1113, C1 => n1044, C2 => n1079
                           , A => n134, ZN => O_52_port);
   U71 : AOI22_X1 port map( A1 => A_ns(51), A2 => n1039, B1 => A_s(51), B2 => 
                           n1032, ZN => n134);
   U72 : OAI221_X1 port map( B1 => n1050, B2 => n1114, C1 => n1044, C2 => n1080
                           , A => n133, ZN => O_53_port);
   U73 : AOI22_X1 port map( A1 => A_ns(52), A2 => n1039, B1 => A_s(52), B2 => 
                           n1032, ZN => n133);
   U74 : OAI221_X1 port map( B1 => n1050, B2 => n1115, C1 => n1044, C2 => n1081
                           , A => n132, ZN => O_54_port);
   U75 : AOI22_X1 port map( A1 => A_ns(53), A2 => n1039, B1 => A_s(53), B2 => 
                           n1032, ZN => n132);
   U76 : OAI221_X1 port map( B1 => n1050, B2 => n1116, C1 => n1044, C2 => n1082
                           , A => n131, ZN => O_55_port);
   U77 : AOI22_X1 port map( A1 => A_ns(54), A2 => n1040, B1 => A_s(54), B2 => 
                           n1033, ZN => n131);
   U78 : OAI221_X1 port map( B1 => n1050, B2 => n1119, C1 => n1044, C2 => n1085
                           , A => n128, ZN => O_58_port);
   U79 : AOI22_X1 port map( A1 => A_ns(57), A2 => n1040, B1 => A_s(57), B2 => 
                           n1033, ZN => n128);
   U80 : BUF_X1 port map( A => n1171, Z => n1028);
   U81 : BUF_X1 port map( A => n1172, Z => n1035);
   U82 : BUF_X1 port map( A => n1049, Z => n1053);
   U83 : BUF_X1 port map( A => n1047, Z => n1042);
   U84 : INV_X1 port map( A => n170, ZN => n1171);
   U85 : INV_X1 port map( A => n171, ZN => n1172);
   U86 : BUF_X1 port map( A => n1048, Z => n1052);
   U87 : BUF_X1 port map( A => n1046, Z => n1043);
   U88 : BUF_X1 port map( A => n1048, Z => n1051);
   U89 : BUF_X1 port map( A => n1048, Z => n1050);
   U90 : BUF_X1 port map( A => n1046, Z => n1044);
   U91 : BUF_X1 port map( A => n1046, Z => n1045);
   U92 : BUF_X1 port map( A => n1047, Z => n1041);
   U93 : BUF_X1 port map( A => n1049, Z => n1054);
   U94 : NAND2_X1 port map( A1 => n182, A2 => n1173, ZN => n170);
   U95 : NAND2_X1 port map( A1 => n182, A2 => n170, ZN => n171);
   U96 : BUF_X1 port map( A => n120, Z => n1049);
   U97 : BUF_X1 port map( A => n121, Z => n1047);
   U98 : BUF_X1 port map( A => n120, Z => n1048);
   U99 : BUF_X1 port map( A => n121, Z => n1046);
   U100 : OAI221_X1 port map( B1 => n1053, B2 => n1167, C1 => n1042, C2 => 
                           n1165, A => n165, ZN => O_24_port);
   U101 : INV_X1 port map( A => A_s(22), ZN => n1167);
   U102 : OAI221_X1 port map( B1 => n1053, B2 => n1170, C1 => n1042, C2 => 
                           n1169, A => n163, ZN => O_26_port);
   U103 : INV_X1 port map( A => A_s(24), ZN => n1170);
   U104 : INV_X1 port map( A => A_ns(24), ZN => n1169);
   U105 : AOI22_X1 port map( A1 => A_ns(25), A2 => n1037, B1 => A_s(25), B2 => 
                           n1030, ZN => n163);
   U106 : OAI221_X1 port map( B1 => n1053, B2 => n1160, C1 => n1041, C2 => 
                           n1158, A => n168, ZN => O_21_port);
   U107 : INV_X1 port map( A => A_s(19), ZN => n1160);
   U108 : INV_X1 port map( A => A_ns(19), ZN => n1158);
   U109 : OAI221_X1 port map( B1 => n1053, B2 => n1163, C1 => n1041, C2 => 
                           n1161, A => n167, ZN => O_22_port);
   U110 : INV_X1 port map( A => A_s(20), ZN => n1163);
   U111 : INV_X1 port map( A => A_ns(20), ZN => n1161);
   U112 : OAI221_X1 port map( B1 => n1053, B2 => n1164, C1 => n1042, C2 => 
                           n1162, A => n166, ZN => O_23_port);
   U113 : INV_X1 port map( A => A_s(21), ZN => n1164);
   U114 : INV_X1 port map( A => A_ns(21), ZN => n1162);
   U115 : OAI221_X1 port map( B1 => n1053, B2 => n1168, C1 => n1042, C2 => 
                           n1166, A => n164, ZN => O_25_port);
   U116 : INV_X1 port map( A => A_s(23), ZN => n1168);
   U117 : INV_X1 port map( A => B(27), ZN => n1173);
   U118 : OR3_X1 port map( A1 => B(25), A2 => B(26), A3 => n1173, ZN => n121);
   U119 : OAI221_X1 port map( B1 => n1054, B2 => n1148, C1 => n1041, C2 => 
                           n1146, A => n176, ZN => O_15_port);
   U120 : INV_X1 port map( A => A_s(13), ZN => n1148);
   U121 : INV_X1 port map( A => A_ns(13), ZN => n1146);
   U122 : OAI221_X1 port map( B1 => n1054, B2 => n1151, C1 => n1041, C2 => 
                           n1149, A => n175, ZN => O_16_port);
   U123 : INV_X1 port map( A => A_s(14), ZN => n1151);
   U124 : INV_X1 port map( A => A_ns(14), ZN => n1149);
   U125 : OAI221_X1 port map( B1 => n1054, B2 => n1152, C1 => n1041, C2 => 
                           n1150, A => n174, ZN => O_17_port);
   U126 : INV_X1 port map( A => A_s(15), ZN => n1152);
   U127 : INV_X1 port map( A => A_ns(15), ZN => n1150);
   U128 : OAI221_X1 port map( B1 => n1054, B2 => n1155, C1 => n1041, C2 => 
                           n1153, A => n173, ZN => O_18_port);
   U129 : INV_X1 port map( A => A_s(16), ZN => n1155);
   U130 : INV_X1 port map( A => A_ns(16), ZN => n1153);
   U131 : OAI221_X1 port map( B1 => n1054, B2 => n1156, C1 => n1041, C2 => 
                           n1154, A => n172, ZN => O_19_port);
   U132 : INV_X1 port map( A => A_s(17), ZN => n1156);
   U133 : INV_X1 port map( A => A_ns(17), ZN => n1154);
   U134 : OAI221_X1 port map( B1 => n1053, B2 => n1159, C1 => n1041, C2 => 
                           n1157, A => n169, ZN => O_20_port);
   U135 : INV_X1 port map( A => A_s(18), ZN => n1159);
   U136 : INV_X1 port map( A => A_ns(18), ZN => n1157);
   U137 : OAI221_X1 port map( B1 => n1050, B2 => n1132, C1 => n1045, C2 => 
                           n1130, A => n124, ZN => O_7_port);
   U138 : INV_X1 port map( A => A_s(5), ZN => n1132);
   U139 : INV_X1 port map( A => A_ns(5), ZN => n1130);
   U140 : OAI221_X1 port map( B1 => n1050, B2 => n1135, C1 => n1045, C2 => 
                           n1133, A => n123, ZN => O_8_port);
   U141 : INV_X1 port map( A => A_s(6), ZN => n1135);
   U142 : INV_X1 port map( A => A_ns(6), ZN => n1133);
   U143 : OAI221_X1 port map( B1 => n1050, B2 => n1136, C1 => n1045, C2 => 
                           n1134, A => n122, ZN => O_9_port);
   U144 : INV_X1 port map( A => A_s(7), ZN => n1136);
   U145 : INV_X1 port map( A => A_ns(7), ZN => n1134);
   U146 : OAI221_X1 port map( B1 => n1139, B2 => n1054, C1 => n1137, C2 => 
                           n1041, A => n181, ZN => O_10_port);
   U147 : INV_X1 port map( A => A_ns(8), ZN => n1137);
   U148 : INV_X1 port map( A => A_s(8), ZN => n1139);
   U149 : OAI221_X1 port map( B1 => n1054, B2 => n1140, C1 => n1041, C2 => 
                           n1138, A => n180, ZN => O_11_port);
   U150 : INV_X1 port map( A => A_s(9), ZN => n1140);
   U151 : INV_X1 port map( A => A_ns(9), ZN => n1138);
   U152 : OAI221_X1 port map( B1 => n1054, B2 => n1143, C1 => n1041, C2 => 
                           n1141, A => n179, ZN => O_12_port);
   U153 : INV_X1 port map( A => A_s(10), ZN => n1143);
   U154 : INV_X1 port map( A => A_ns(10), ZN => n1141);
   U155 : OAI221_X1 port map( B1 => n1054, B2 => n1144, C1 => n1041, C2 => 
                           n1142, A => n178, ZN => O_13_port);
   U156 : INV_X1 port map( A => A_s(11), ZN => n1144);
   U157 : INV_X1 port map( A => A_ns(11), ZN => n1142);
   U158 : OAI221_X1 port map( B1 => n1054, B2 => n1147, C1 => n1041, C2 => 
                           n1145, A => n177, ZN => O_14_port);
   U159 : INV_X1 port map( A => A_s(12), ZN => n1147);
   U160 : INV_X1 port map( A => A_ns(12), ZN => n1145);
   U161 : OAI22_X1 port map( A1 => n170, A2 => n1123, B1 => n171, B2 => n1121, 
                           ZN => O_1_port);
   U162 : OAI221_X1 port map( B1 => n1053, B2 => n1123, C1 => n1042, C2 => 
                           n1121, A => n159, ZN => O_2_port);
   U163 : AOI22_X1 port map( A1 => A_ns(1), A2 => n1037, B1 => A_s(1), B2 => 
                           n1030, ZN => n159);
   U164 : OAI221_X1 port map( B1 => n1052, B2 => n1124, C1 => n1043, C2 => 
                           n1122, A => n148, ZN => O_3_port);
   U165 : INV_X1 port map( A => A_s(1), ZN => n1124);
   U166 : INV_X1 port map( A => A_ns(1), ZN => n1122);
   U167 : OAI221_X1 port map( B1 => n1051, B2 => n1127, C1 => n1044, C2 => 
                           n1125, A => n137, ZN => O_4_port);
   U168 : INV_X1 port map( A => A_s(2), ZN => n1127);
   U169 : INV_X1 port map( A => A_ns(2), ZN => n1125);
   U170 : OAI221_X1 port map( B1 => n1050, B2 => n1128, C1 => n1045, C2 => 
                           n1126, A => n126, ZN => O_5_port);
   U171 : INV_X1 port map( A => A_s(3), ZN => n1128);
   U172 : INV_X1 port map( A => A_ns(3), ZN => n1126);
   U173 : OAI221_X1 port map( B1 => n1050, B2 => n1131, C1 => n1045, C2 => 
                           n1129, A => n125, ZN => O_6_port);
   U174 : INV_X1 port map( A => A_s(4), ZN => n1131);
   U175 : INV_X1 port map( A => A_ns(4), ZN => n1129);
   U176 : INV_X1 port map( A => A_ns(0), ZN => n1121);
   U177 : INV_X1 port map( A => A_s(0), ZN => n1123);
   U178 : AOI22_X1 port map( A1 => A_ns(2), A2 => n1038, B1 => A_s(2), B2 => 
                           n1031, ZN => n148);
   U179 : AOI22_X1 port map( A1 => A_ns(3), A2 => n1039, B1 => A_s(3), B2 => 
                           n1032, ZN => n137);
   U180 : AOI22_X1 port map( A1 => A_ns(4), A2 => n1040, B1 => A_s(4), B2 => 
                           n1033, ZN => n126);
   U181 : AOI22_X1 port map( A1 => A_ns(5), A2 => n1040, B1 => A_s(5), B2 => 
                           n1033, ZN => n125);
   U182 : AOI22_X1 port map( A1 => A_ns(6), A2 => n1040, B1 => A_s(6), B2 => 
                           n1033, ZN => n124);
   U183 : AOI22_X1 port map( A1 => A_ns(7), A2 => n1040, B1 => A_s(7), B2 => 
                           n1033, ZN => n123);
   U184 : AOI22_X1 port map( A1 => A_ns(8), A2 => n1040, B1 => A_s(8), B2 => 
                           n1033, ZN => n122);
   U185 : AOI22_X1 port map( A1 => A_ns(9), A2 => n1036, B1 => A_s(9), B2 => 
                           n1029, ZN => n181);
   U186 : AOI22_X1 port map( A1 => A_ns(10), A2 => n1036, B1 => A_s(10), B2 => 
                           n1029, ZN => n180);
   U187 : AOI22_X1 port map( A1 => A_ns(11), A2 => n1036, B1 => A_s(11), B2 => 
                           n1029, ZN => n179);
   U188 : AOI22_X1 port map( A1 => A_ns(12), A2 => n1036, B1 => A_s(12), B2 => 
                           n1029, ZN => n178);
   U189 : AOI22_X1 port map( A1 => A_ns(13), A2 => n1036, B1 => A_s(13), B2 => 
                           n1029, ZN => n177);
   U190 : AOI22_X1 port map( A1 => A_ns(14), A2 => n1036, B1 => A_s(14), B2 => 
                           n1029, ZN => n176);
   U191 : AOI22_X1 port map( A1 => A_ns(15), A2 => n1036, B1 => A_s(15), B2 => 
                           n1029, ZN => n175);
   U192 : AOI22_X1 port map( A1 => A_ns(16), A2 => n1036, B1 => A_s(16), B2 => 
                           n1029, ZN => n174);
   U193 : AOI22_X1 port map( A1 => A_ns(17), A2 => n1036, B1 => A_s(17), B2 => 
                           n1029, ZN => n173);
   U194 : AOI22_X1 port map( A1 => A_ns(18), A2 => n1036, B1 => A_s(18), B2 => 
                           n1029, ZN => n172);
   U195 : AOI22_X1 port map( A1 => A_ns(19), A2 => n1036, B1 => A_s(19), B2 => 
                           n1029, ZN => n169);
   U196 : AOI22_X1 port map( A1 => A_ns(20), A2 => n1036, B1 => A_s(20), B2 => 
                           n1029, ZN => n168);
   U197 : AOI22_X1 port map( A1 => A_ns(21), A2 => n1037, B1 => A_s(21), B2 => 
                           n1030, ZN => n167);
   U198 : AOI22_X1 port map( A1 => A_ns(22), A2 => n1037, B1 => A_s(22), B2 => 
                           n1030, ZN => n166);
   U199 : AOI22_X1 port map( A1 => A_ns(23), A2 => n1037, B1 => A_s(23), B2 => 
                           n1030, ZN => n165);
   U200 : AOI22_X1 port map( A1 => A_ns(24), A2 => n1037, B1 => A_s(24), B2 => 
                           n1030, ZN => n164);
   U201 : INV_X1 port map( A => A_ns(22), ZN => n1165);
   U202 : INV_X1 port map( A => A_ns(23), ZN => n1166);
   U203 : INV_X1 port map( A => A_ns(26), ZN => n1055);
   U204 : INV_X1 port map( A => A_ns(27), ZN => n1056);
   U205 : INV_X1 port map( A => A_ns(28), ZN => n1057);
   U206 : INV_X1 port map( A => A_ns(29), ZN => n1058);
   U207 : INV_X1 port map( A => A_ns(30), ZN => n1059);
   U208 : INV_X1 port map( A => A_ns(31), ZN => n1060);
   U209 : INV_X1 port map( A => A_ns(32), ZN => n1061);
   U210 : INV_X1 port map( A => A_ns(33), ZN => n1062);
   U211 : INV_X1 port map( A => A_ns(34), ZN => n1063);
   U212 : INV_X1 port map( A => A_ns(35), ZN => n1064);
   U213 : INV_X1 port map( A => A_ns(36), ZN => n1065);
   U214 : INV_X1 port map( A => A_ns(37), ZN => n1066);
   U215 : INV_X1 port map( A => A_ns(38), ZN => n1067);
   U216 : INV_X1 port map( A => A_ns(39), ZN => n1068);
   U217 : INV_X1 port map( A => A_ns(40), ZN => n1069);
   U218 : INV_X1 port map( A => A_ns(41), ZN => n1070);
   U219 : INV_X1 port map( A => A_ns(42), ZN => n1071);
   U220 : INV_X1 port map( A => A_ns(43), ZN => n1072);
   U221 : INV_X1 port map( A => A_ns(44), ZN => n1073);
   U222 : INV_X1 port map( A => A_ns(45), ZN => n1074);
   U223 : INV_X1 port map( A => A_ns(46), ZN => n1075);
   U224 : INV_X1 port map( A => A_ns(47), ZN => n1076);
   U225 : INV_X1 port map( A => A_ns(48), ZN => n1077);
   U226 : INV_X1 port map( A => A_ns(49), ZN => n1078);
   U227 : INV_X1 port map( A => A_ns(50), ZN => n1079);
   U228 : INV_X1 port map( A => A_ns(51), ZN => n1080);
   U229 : INV_X1 port map( A => A_ns(52), ZN => n1081);
   U230 : INV_X1 port map( A => A_ns(53), ZN => n1082);
   U231 : INV_X1 port map( A => A_ns(54), ZN => n1083);
   U232 : INV_X1 port map( A => A_ns(55), ZN => n1084);
   U233 : INV_X1 port map( A => A_ns(56), ZN => n1085);
   U234 : INV_X1 port map( A => A_ns(57), ZN => n1086);
   U235 : INV_X1 port map( A => A_ns(25), ZN => n1087);
   U236 : INV_X1 port map( A => A_s(25), ZN => n1088);
   U237 : INV_X1 port map( A => A_s(26), ZN => n1089);
   U238 : INV_X1 port map( A => A_s(27), ZN => n1090);
   U239 : INV_X1 port map( A => A_s(28), ZN => n1091);
   U240 : INV_X1 port map( A => A_s(29), ZN => n1092);
   U243 : INV_X1 port map( A => A_s(30), ZN => n1093);
   U244 : INV_X1 port map( A => A_s(31), ZN => n1094);
   U245 : INV_X1 port map( A => A_s(32), ZN => n1095);
   U246 : INV_X1 port map( A => A_s(33), ZN => n1096);
   U247 : INV_X1 port map( A => A_s(34), ZN => n1097);
   U248 : INV_X1 port map( A => A_s(35), ZN => n1098);
   U249 : INV_X1 port map( A => A_s(36), ZN => n1099);
   U250 : INV_X1 port map( A => A_s(37), ZN => n1100);
   U251 : INV_X1 port map( A => A_s(38), ZN => n1101);
   U252 : INV_X1 port map( A => A_s(39), ZN => n1102);
   U253 : INV_X1 port map( A => A_s(40), ZN => n1103);
   U254 : INV_X1 port map( A => A_s(41), ZN => n1104);
   U255 : INV_X1 port map( A => A_s(42), ZN => n1105);
   U256 : INV_X1 port map( A => A_s(43), ZN => n1106);
   U257 : INV_X1 port map( A => A_s(44), ZN => n1107);
   U258 : INV_X1 port map( A => A_s(45), ZN => n1108);
   U259 : INV_X1 port map( A => A_s(46), ZN => n1109);
   U260 : INV_X1 port map( A => A_s(47), ZN => n1110);
   U261 : INV_X1 port map( A => A_s(48), ZN => n1111);
   U262 : INV_X1 port map( A => A_s(49), ZN => n1112);
   U263 : INV_X1 port map( A => A_s(50), ZN => n1113);
   U264 : INV_X1 port map( A => A_s(51), ZN => n1114);
   U265 : INV_X1 port map( A => A_s(52), ZN => n1115);
   U266 : INV_X1 port map( A => A_s(53), ZN => n1116);
   U267 : INV_X1 port map( A => A_s(54), ZN => n1117);
   U268 : INV_X1 port map( A => A_s(55), ZN => n1118);
   U269 : INV_X1 port map( A => A_s(56), ZN => n1119);
   U270 : INV_X1 port map( A => A_s(57), ZN => n1120);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT58_i24 is

   port( A_s, A_ns, B : in std_logic_vector (57 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (57 downto 0));

end BOOTHENC_NBIT58_i24;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT58_i24 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, O_57_port, O_56_port, O_55_port, O_54_port, O_53_port,
      O_52_port, O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, 
      O_46_port, O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, 
      O_40_port, O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, 
      O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, 
      O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, 
      O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, 
      O_16_port, O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, 
      O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, 
      O_3_port, O_2_port, O_1_port, n116, n117, n118, n119, n120, n121, n122, 
      n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, 
      n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n1004, n1005, n1006, n1007, n1008, 
      n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, 
      n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, 
      n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, 
      n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, 
      n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, 
      n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, 
      n1069, n1070, n1071, n1072, n1073, n1074, n1075, A_so_36_port, n1077, 
      n1078, A_so_38_port, n1080, n1081, n1082, n1083, n1084, n1085, n1086, 
      n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, 
      n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, 
      n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, 
      n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, 
      n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, 
      n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, 
      n1147, n1148 : std_logic;

begin
   O <= ( O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, O_52_port, 
      O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, O_46_port, 
      O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, O_40_port, 
      O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, 
      O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, 
      O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, 
      O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, O_16_port, 
      O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, O_10_port, 
      O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, O_3_port, 
      O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(55), A_s(54), A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), 
      A_s(48), A_s(47), A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), 
      A_s(40), A_s(39), A_s(38), A_s(37), A_so_38_port, A_s(35), A_so_36_port, 
      A_s(33), A_s(32), A_s(31), A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), 
      A_s(25), A_s(24), A_s(23), A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), 
      A_s(17), A_s(16), A_s(15), A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), 
      A_s(9), A_s(8), A_s(7), A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), 
      A_s(0), X_Logic0_port, X_Logic0_port );
   A_nso <= ( A_ns(55), A_ns(54), A_ns(53), A_ns(52), A_ns(51), A_ns(50), 
      A_ns(49), A_ns(48), A_ns(47), A_ns(46), A_ns(45), A_ns(44), A_ns(43), 
      A_ns(42), A_ns(41), A_ns(40), A_ns(39), A_ns(38), A_ns(37), A_ns(36), 
      A_ns(35), A_ns(34), A_ns(33), A_ns(32), A_ns(31), A_ns(30), A_ns(29), 
      A_ns(28), A_ns(27), A_ns(26), A_ns(25), A_ns(24), A_ns(23), A_ns(22), 
      A_ns(21), A_ns(20), A_ns(19), A_ns(18), A_ns(17), A_ns(16), A_ns(15), 
      A_ns(14), A_ns(13), A_ns(12), A_ns(11), A_ns(10), A_ns(9), A_ns(8), 
      A_ns(7), A_ns(6), A_ns(5), A_ns(4), A_ns(3), A_ns(2), A_ns(1), A_ns(0), 
      X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U233 : XOR2_X1 port map( A => B(23), B => B(24), Z => n176);
   U234 : NAND3_X1 port map( A1 => B(24), A2 => n1148, A3 => B(23), ZN => n116)
                           ;
   U2 : OAI221_X1 port map( B1 => n1030, B2 => n1069, C1 => n1019, C2 => n1035,
                           A => n154, ZN => O_29_port);
   U3 : OAI221_X1 port map( B1 => n1028, B2 => n1082, C1 => n1020, C2 => n1046,
                           A => n141, ZN => O_40_port);
   U4 : OAI221_X1 port map( B1 => n1028, B2 => n1084, C1 => n1020, C2 => n1048,
                           A => n139, ZN => O_42_port);
   U5 : OAI221_X1 port map( B1 => n1029, B2 => n1074, C1 => n1019, C2 => n1040,
                           A => n148, ZN => O_34_port);
   U6 : OAI221_X1 port map( B1 => n1029, B2 => n1078, C1 => n1020, C2 => n1043,
                           A => n145, ZN => O_37_port);
   U7 : AOI22_X1 port map( A1 => A_ns(56), A2 => n1017, B1 => A_s(56), B2 => 
                           n1010, ZN => n123);
   U8 : BUF_X1 port map( A => n1011, Z => n1014);
   U9 : BUF_X1 port map( A => n1004, Z => n1007);
   U10 : BUF_X1 port map( A => n1011, Z => n1015);
   U11 : BUF_X1 port map( A => n1004, Z => n1008);
   U12 : BUF_X1 port map( A => n1012, Z => n1016);
   U13 : BUF_X1 port map( A => n1005, Z => n1009);
   U14 : BUF_X1 port map( A => n1012, Z => n1017);
   U15 : BUF_X1 port map( A => n1005, Z => n1010);
   U16 : BUF_X1 port map( A => n1011, Z => n1013);
   U17 : BUF_X1 port map( A => n1004, Z => n1006);
   U18 : AOI22_X1 port map( A1 => A_ns(36), A2 => n1015, B1 => A_so_38_port, B2
                           => n1008, ZN => n145);
   U19 : AOI22_X1 port map( A1 => A_ns(28), A2 => n1014, B1 => A_s(28), B2 => 
                           n1007, ZN => n154);
   U20 : OAI221_X1 port map( B1 => n1029, B2 => n1071, C1 => n1019, C2 => n1037
                           , A => n151, ZN => O_31_port);
   U21 : AOI22_X1 port map( A1 => A_ns(30), A2 => n1014, B1 => A_s(30), B2 => 
                           n1007, ZN => n151);
   U22 : OAI221_X1 port map( B1 => n1029, B2 => n1073, C1 => n1019, C2 => n1039
                           , A => n149, ZN => O_33_port);
   U23 : AOI22_X1 port map( A1 => A_ns(32), A2 => n1015, B1 => A_s(32), B2 => 
                           n1008, ZN => n149);
   U24 : OAI221_X1 port map( B1 => n1029, B2 => n1081, C1 => n1020, C2 => n1045
                           , A => n143, ZN => O_39_port);
   U25 : AOI22_X1 port map( A1 => A_ns(38), A2 => n1015, B1 => A_s(38), B2 => 
                           n1008, ZN => n143);
   U26 : OAI221_X1 port map( B1 => n1030, B2 => n1066, C1 => n1019, C2 => n1032
                           , A => n157, ZN => O_26_port);
   U27 : AOI22_X1 port map( A1 => A_ns(25), A2 => n1014, B1 => A_s(25), B2 => 
                           n1007, ZN => n157);
   U28 : OAI221_X1 port map( B1 => n1030, B2 => n1068, C1 => n1019, C2 => n1034
                           , A => n155, ZN => O_28_port);
   U29 : AOI22_X1 port map( A1 => A_ns(27), A2 => n1014, B1 => A_s(27), B2 => 
                           n1007, ZN => n155);
   U30 : OAI221_X1 port map( B1 => n1029, B2 => n1072, C1 => n1019, C2 => n1038
                           , A => n150, ZN => O_32_port);
   U31 : AOI22_X1 port map( A1 => A_ns(31), A2 => n1014, B1 => A_s(31), B2 => 
                           n1007, ZN => n150);
   U32 : AOI22_X1 port map( A1 => A_ns(33), A2 => n1015, B1 => A_s(33), B2 => 
                           n1008, ZN => n148);
   U33 : OAI221_X1 port map( B1 => n1029, B2 => n1077, C1 => n1020, C2 => n1042
                           , A => n146, ZN => O_36_port);
   U34 : AOI22_X1 port map( A1 => A_ns(35), A2 => n1015, B1 => A_s(35), B2 => 
                           n1008, ZN => n146);
   U35 : OAI221_X1 port map( B1 => n1029, B2 => n1080, C1 => n1020, C2 => n1044
                           , A => n144, ZN => O_38_port);
   U36 : AOI22_X1 port map( A1 => A_ns(37), A2 => n1015, B1 => A_s(37), B2 => 
                           n1008, ZN => n144);
   U37 : AOI22_X1 port map( A1 => A_ns(39), A2 => n1015, B1 => A_s(39), B2 => 
                           n1008, ZN => n141);
   U38 : OAI221_X1 port map( B1 => n1029, B2 => n1075, C1 => n1020, C2 => n1041
                           , A => n147, ZN => O_35_port);
   U39 : AOI22_X1 port map( A1 => A_ns(34), A2 => n1015, B1 => A_so_36_port, B2
                           => n1008, ZN => n147);
   U40 : OAI221_X1 port map( B1 => n1030, B2 => n1065, C1 => n1019, C2 => n1064
                           , A => n158, ZN => O_25_port);
   U41 : AOI22_X1 port map( A1 => A_ns(24), A2 => n1014, B1 => A_s(24), B2 => 
                           n1007, ZN => n158);
   U42 : OAI221_X1 port map( B1 => n1030, B2 => n1067, C1 => n1019, C2 => n1033
                           , A => n156, ZN => O_27_port);
   U43 : AOI22_X1 port map( A1 => A_ns(26), A2 => n1014, B1 => A_s(26), B2 => 
                           n1007, ZN => n156);
   U44 : OAI221_X1 port map( B1 => n1029, B2 => n1070, C1 => n1019, C2 => n1036
                           , A => n152, ZN => O_30_port);
   U45 : AOI22_X1 port map( A1 => A_ns(29), A2 => n1014, B1 => A_s(29), B2 => 
                           n1007, ZN => n152);
   U46 : BUF_X1 port map( A => n1146, Z => n1004);
   U47 : BUF_X1 port map( A => n1147, Z => n1011);
   U48 : OAI221_X1 port map( B1 => n1028, B2 => n1088, C1 => n1020, C2 => n1052
                           , A => n135, ZN => O_46_port);
   U49 : AOI22_X1 port map( A1 => A_ns(45), A2 => n1016, B1 => A_s(45), B2 => 
                           n1009, ZN => n135);
   U50 : OAI221_X1 port map( B1 => n1028, B2 => n1090, C1 => n1021, C2 => n1054
                           , A => n133, ZN => O_48_port);
   U51 : AOI22_X1 port map( A1 => A_ns(47), A2 => n1016, B1 => A_s(47), B2 => 
                           n1009, ZN => n133);
   U52 : OAI221_X1 port map( B1 => n1028, B2 => n1085, C1 => n1020, C2 => n1049
                           , A => n138, ZN => O_43_port);
   U53 : AOI22_X1 port map( A1 => A_ns(42), A2 => n1015, B1 => A_s(42), B2 => 
                           n1008, ZN => n138);
   U54 : AOI22_X1 port map( A1 => A_ns(41), A2 => n1015, B1 => A_s(41), B2 => 
                           n1008, ZN => n139);
   U55 : OAI221_X1 port map( B1 => n1028, B2 => n1086, C1 => n1020, C2 => n1050
                           , A => n137, ZN => O_44_port);
   U56 : AOI22_X1 port map( A1 => A_ns(43), A2 => n1016, B1 => A_s(43), B2 => 
                           n1009, ZN => n137);
   U57 : OAI221_X1 port map( B1 => n1028, B2 => n1087, C1 => n1020, C2 => n1051
                           , A => n136, ZN => O_45_port);
   U58 : AOI22_X1 port map( A1 => A_ns(44), A2 => n1016, B1 => A_s(44), B2 => 
                           n1009, ZN => n136);
   U59 : OAI221_X1 port map( B1 => n1028, B2 => n1089, C1 => n1021, C2 => n1053
                           , A => n134, ZN => O_47_port);
   U60 : AOI22_X1 port map( A1 => A_ns(46), A2 => n1016, B1 => A_s(46), B2 => 
                           n1009, ZN => n134);
   U61 : OAI221_X1 port map( B1 => n1028, B2 => n1091, C1 => n1021, C2 => n1055
                           , A => n132, ZN => O_49_port);
   U62 : AOI22_X1 port map( A1 => A_ns(48), A2 => n1016, B1 => A_s(48), B2 => 
                           n1009, ZN => n132);
   U63 : OAI221_X1 port map( B1 => n1027, B2 => n1093, C1 => n1021, C2 => n1057
                           , A => n129, ZN => O_51_port);
   U64 : AOI22_X1 port map( A1 => A_ns(50), A2 => n1016, B1 => A_s(50), B2 => 
                           n1009, ZN => n129);
   U65 : OAI221_X1 port map( B1 => n1028, B2 => n1083, C1 => n1020, C2 => n1047
                           , A => n140, ZN => O_41_port);
   U66 : AOI22_X1 port map( A1 => A_ns(40), A2 => n1015, B1 => A_s(40), B2 => 
                           n1008, ZN => n140);
   U67 : OAI221_X1 port map( B1 => n1027, B2 => n1097, C1 => n1021, C2 => n1061
                           , A => n125, ZN => O_55_port);
   U68 : AOI22_X1 port map( A1 => A_ns(54), A2 => n1017, B1 => A_s(54), B2 => 
                           n1010, ZN => n125);
   U69 : OAI221_X1 port map( B1 => n1027, B2 => n1098, C1 => n1021, C2 => n1062
                           , A => n124, ZN => O_56_port);
   U70 : AOI22_X1 port map( A1 => A_ns(55), A2 => n1017, B1 => A_s(55), B2 => 
                           n1010, ZN => n124);
   U71 : OAI221_X1 port map( B1 => n1028, B2 => n1092, C1 => n1021, C2 => n1056
                           , A => n130, ZN => O_50_port);
   U72 : AOI22_X1 port map( A1 => A_ns(49), A2 => n1016, B1 => A_s(49), B2 => 
                           n1009, ZN => n130);
   U73 : OAI221_X1 port map( B1 => n1027, B2 => n1094, C1 => n1021, C2 => n1058
                           , A => n128, ZN => O_52_port);
   U74 : AOI22_X1 port map( A1 => A_ns(51), A2 => n1016, B1 => A_s(51), B2 => 
                           n1009, ZN => n128);
   U75 : OAI221_X1 port map( B1 => n1027, B2 => n1095, C1 => n1021, C2 => n1059
                           , A => n127, ZN => O_53_port);
   U76 : AOI22_X1 port map( A1 => A_ns(52), A2 => n1016, B1 => A_s(52), B2 => 
                           n1009, ZN => n127);
   U77 : OAI221_X1 port map( B1 => n1027, B2 => n1096, C1 => n1021, C2 => n1060
                           , A => n126, ZN => O_54_port);
   U78 : AOI22_X1 port map( A1 => A_ns(53), A2 => n1016, B1 => A_s(53), B2 => 
                           n1009, ZN => n126);
   U79 : BUF_X1 port map( A => n1146, Z => n1005);
   U80 : BUF_X1 port map( A => n1147, Z => n1012);
   U81 : OAI221_X1 port map( B1 => n1027, B2 => n1099, C1 => n1021, C2 => n1063
                           , A => n123, ZN => O_57_port);
   U82 : BUF_X1 port map( A => n1026, Z => n1030);
   U83 : BUF_X1 port map( A => n1024, Z => n1019);
   U84 : INV_X1 port map( A => n164, ZN => n1146);
   U85 : INV_X1 port map( A => n165, ZN => n1147);
   U86 : BUF_X1 port map( A => n1025, Z => n1029);
   U87 : BUF_X1 port map( A => n1023, Z => n1020);
   U88 : BUF_X1 port map( A => n1025, Z => n1028);
   U89 : BUF_X1 port map( A => n1025, Z => n1027);
   U90 : BUF_X1 port map( A => n1023, Z => n1021);
   U91 : BUF_X1 port map( A => n1024, Z => n1018);
   U92 : BUF_X1 port map( A => n1026, Z => n1031);
   U93 : BUF_X1 port map( A => n1023, Z => n1022);
   U94 : NAND2_X1 port map( A1 => n176, A2 => n1148, ZN => n164);
   U95 : NAND2_X1 port map( A1 => n176, A2 => n164, ZN => n165);
   U96 : BUF_X1 port map( A => n117, Z => n1024);
   U97 : BUF_X1 port map( A => n116, Z => n1026);
   U98 : BUF_X1 port map( A => n116, Z => n1025);
   U99 : BUF_X1 port map( A => n117, Z => n1023);
   U100 : OAI221_X1 port map( B1 => n1030, B2 => n1145, C1 => n1019, C2 => 
                           n1144, A => n159, ZN => O_24_port);
   U101 : INV_X1 port map( A => A_s(22), ZN => n1145);
   U102 : INV_X1 port map( A => A_ns(22), ZN => n1144);
   U103 : AOI22_X1 port map( A1 => A_ns(23), A2 => n1014, B1 => A_s(23), B2 => 
                           n1007, ZN => n159);
   U104 : OAI221_X1 port map( B1 => n1030, B2 => n1142, C1 => n1018, C2 => 
                           n1140, A => n161, ZN => O_22_port);
   U105 : INV_X1 port map( A => A_s(20), ZN => n1142);
   U106 : OAI221_X1 port map( B1 => n1030, B2 => n1139, C1 => n1018, C2 => 
                           n1137, A => n162, ZN => O_21_port);
   U107 : INV_X1 port map( A => A_s(19), ZN => n1139);
   U108 : INV_X1 port map( A => A_ns(19), ZN => n1137);
   U109 : OAI221_X1 port map( B1 => n1030, B2 => n1143, C1 => n1019, C2 => 
                           n1141, A => n160, ZN => O_23_port);
   U110 : INV_X1 port map( A => A_s(21), ZN => n1143);
   U111 : INV_X1 port map( A => B(25), ZN => n1148);
   U112 : OR3_X1 port map( A1 => B(23), A2 => B(24), A3 => n1148, ZN => n117);
   U113 : OAI221_X1 port map( B1 => n1031, B2 => n1127, C1 => n1018, C2 => 
                           n1125, A => n170, ZN => O_15_port);
   U114 : INV_X1 port map( A => A_s(13), ZN => n1127);
   U115 : INV_X1 port map( A => A_ns(13), ZN => n1125);
   U116 : OAI221_X1 port map( B1 => n1031, B2 => n1130, C1 => n1018, C2 => 
                           n1128, A => n169, ZN => O_16_port);
   U117 : INV_X1 port map( A => A_s(14), ZN => n1130);
   U118 : INV_X1 port map( A => A_ns(14), ZN => n1128);
   U119 : OAI221_X1 port map( B1 => n1031, B2 => n1131, C1 => n1018, C2 => 
                           n1129, A => n168, ZN => O_17_port);
   U120 : INV_X1 port map( A => A_s(15), ZN => n1131);
   U121 : INV_X1 port map( A => A_ns(15), ZN => n1129);
   U122 : OAI221_X1 port map( B1 => n1030, B2 => n1134, C1 => n1018, C2 => 
                           n1132, A => n167, ZN => O_18_port);
   U123 : INV_X1 port map( A => A_s(16), ZN => n1134);
   U124 : INV_X1 port map( A => A_ns(16), ZN => n1132);
   U125 : OAI221_X1 port map( B1 => n1030, B2 => n1135, C1 => n1018, C2 => 
                           n1133, A => n166, ZN => O_19_port);
   U126 : INV_X1 port map( A => A_s(17), ZN => n1135);
   U127 : INV_X1 port map( A => A_ns(17), ZN => n1133);
   U128 : OAI221_X1 port map( B1 => n1030, B2 => n1138, C1 => n1018, C2 => 
                           n1136, A => n163, ZN => O_20_port);
   U129 : INV_X1 port map( A => A_s(18), ZN => n1138);
   U130 : INV_X1 port map( A => A_ns(18), ZN => n1136);
   U131 : OAI221_X1 port map( B1 => n1027, B2 => n1111, C1 => n1022, C2 => 
                           n1109, A => n120, ZN => O_7_port);
   U132 : INV_X1 port map( A => A_s(5), ZN => n1111);
   U133 : INV_X1 port map( A => A_ns(5), ZN => n1109);
   U134 : OAI221_X1 port map( B1 => n1027, B2 => n1114, C1 => n1022, C2 => 
                           n1112, A => n119, ZN => O_8_port);
   U135 : INV_X1 port map( A => A_s(6), ZN => n1114);
   U136 : INV_X1 port map( A => A_ns(6), ZN => n1112);
   U137 : OAI221_X1 port map( B1 => n1027, B2 => n1115, C1 => n1022, C2 => 
                           n1113, A => n118, ZN => O_9_port);
   U138 : INV_X1 port map( A => A_s(7), ZN => n1115);
   U139 : INV_X1 port map( A => A_ns(7), ZN => n1113);
   U140 : OAI221_X1 port map( B1 => n1118, B2 => n1031, C1 => n1116, C2 => 
                           n1018, A => n175, ZN => O_10_port);
   U141 : INV_X1 port map( A => A_ns(8), ZN => n1116);
   U142 : INV_X1 port map( A => A_s(8), ZN => n1118);
   U143 : OAI221_X1 port map( B1 => n1031, B2 => n1119, C1 => n1018, C2 => 
                           n1117, A => n174, ZN => O_11_port);
   U144 : INV_X1 port map( A => A_s(9), ZN => n1119);
   U145 : INV_X1 port map( A => A_ns(9), ZN => n1117);
   U146 : OAI221_X1 port map( B1 => n1031, B2 => n1122, C1 => n1018, C2 => 
                           n1120, A => n173, ZN => O_12_port);
   U147 : INV_X1 port map( A => A_s(10), ZN => n1122);
   U148 : INV_X1 port map( A => A_ns(10), ZN => n1120);
   U149 : OAI221_X1 port map( B1 => n1031, B2 => n1123, C1 => n1018, C2 => 
                           n1121, A => n172, ZN => O_13_port);
   U150 : INV_X1 port map( A => A_s(11), ZN => n1123);
   U151 : INV_X1 port map( A => A_ns(11), ZN => n1121);
   U152 : OAI221_X1 port map( B1 => n1031, B2 => n1126, C1 => n1018, C2 => 
                           n1124, A => n171, ZN => O_14_port);
   U153 : INV_X1 port map( A => A_s(12), ZN => n1126);
   U154 : INV_X1 port map( A => A_ns(12), ZN => n1124);
   U155 : OAI22_X1 port map( A1 => n164, A2 => n1102, B1 => n165, B2 => n1100, 
                           ZN => O_1_port);
   U156 : OAI221_X1 port map( B1 => n1029, B2 => n1102, C1 => n1019, C2 => 
                           n1100, A => n153, ZN => O_2_port);
   U157 : AOI22_X1 port map( A1 => A_ns(1), A2 => n1014, B1 => A_s(1), B2 => 
                           n1007, ZN => n153);
   U158 : OAI221_X1 port map( B1 => n1029, B2 => n1103, C1 => n1020, C2 => 
                           n1101, A => n142, ZN => O_3_port);
   U159 : INV_X1 port map( A => A_s(1), ZN => n1103);
   U160 : INV_X1 port map( A => A_ns(1), ZN => n1101);
   U161 : OAI221_X1 port map( B1 => n1028, B2 => n1106, C1 => n1021, C2 => 
                           n1104, A => n131, ZN => O_4_port);
   U162 : INV_X1 port map( A => A_s(2), ZN => n1106);
   U163 : INV_X1 port map( A => A_ns(2), ZN => n1104);
   U164 : OAI221_X1 port map( B1 => n1027, B2 => n1107, C1 => n1021, C2 => 
                           n1105, A => n122, ZN => O_5_port);
   U165 : INV_X1 port map( A => A_s(3), ZN => n1107);
   U166 : INV_X1 port map( A => A_ns(3), ZN => n1105);
   U167 : OAI221_X1 port map( B1 => n1027, B2 => n1110, C1 => n1022, C2 => 
                           n1108, A => n121, ZN => O_6_port);
   U168 : INV_X1 port map( A => A_s(4), ZN => n1110);
   U169 : INV_X1 port map( A => A_ns(4), ZN => n1108);
   U170 : INV_X1 port map( A => A_ns(0), ZN => n1100);
   U171 : INV_X1 port map( A => A_s(0), ZN => n1102);
   U172 : AOI22_X1 port map( A1 => A_ns(2), A2 => n1015, B1 => A_s(2), B2 => 
                           n1008, ZN => n142);
   U173 : AOI22_X1 port map( A1 => A_ns(3), A2 => n1016, B1 => A_s(3), B2 => 
                           n1009, ZN => n131);
   U174 : AOI22_X1 port map( A1 => A_ns(4), A2 => n1017, B1 => A_s(4), B2 => 
                           n1010, ZN => n122);
   U175 : AOI22_X1 port map( A1 => A_ns(5), A2 => n1017, B1 => A_s(5), B2 => 
                           n1010, ZN => n121);
   U176 : AOI22_X1 port map( A1 => A_ns(6), A2 => n1017, B1 => A_s(6), B2 => 
                           n1010, ZN => n120);
   U177 : AOI22_X1 port map( A1 => A_ns(7), A2 => n1017, B1 => A_s(7), B2 => 
                           n1010, ZN => n119);
   U178 : AOI22_X1 port map( A1 => A_ns(8), A2 => n1017, B1 => A_s(8), B2 => 
                           n1010, ZN => n118);
   U179 : AOI22_X1 port map( A1 => A_ns(9), A2 => n1013, B1 => A_s(9), B2 => 
                           n1006, ZN => n175);
   U180 : AOI22_X1 port map( A1 => A_ns(10), A2 => n1013, B1 => A_s(10), B2 => 
                           n1006, ZN => n174);
   U181 : AOI22_X1 port map( A1 => A_ns(11), A2 => n1013, B1 => A_s(11), B2 => 
                           n1006, ZN => n173);
   U182 : AOI22_X1 port map( A1 => A_ns(12), A2 => n1013, B1 => A_s(12), B2 => 
                           n1006, ZN => n172);
   U183 : AOI22_X1 port map( A1 => A_ns(13), A2 => n1013, B1 => A_s(13), B2 => 
                           n1006, ZN => n171);
   U184 : AOI22_X1 port map( A1 => A_ns(14), A2 => n1013, B1 => A_s(14), B2 => 
                           n1006, ZN => n170);
   U185 : AOI22_X1 port map( A1 => A_ns(15), A2 => n1013, B1 => A_s(15), B2 => 
                           n1006, ZN => n169);
   U186 : AOI22_X1 port map( A1 => A_ns(16), A2 => n1013, B1 => A_s(16), B2 => 
                           n1006, ZN => n168);
   U187 : AOI22_X1 port map( A1 => A_ns(17), A2 => n1013, B1 => A_s(17), B2 => 
                           n1006, ZN => n167);
   U188 : AOI22_X1 port map( A1 => A_ns(18), A2 => n1013, B1 => A_s(18), B2 => 
                           n1006, ZN => n166);
   U189 : AOI22_X1 port map( A1 => A_ns(19), A2 => n1013, B1 => A_s(19), B2 => 
                           n1006, ZN => n163);
   U190 : AOI22_X1 port map( A1 => A_ns(20), A2 => n1013, B1 => A_s(20), B2 => 
                           n1006, ZN => n162);
   U191 : AOI22_X1 port map( A1 => A_ns(21), A2 => n1014, B1 => A_s(21), B2 => 
                           n1007, ZN => n161);
   U192 : AOI22_X1 port map( A1 => A_ns(22), A2 => n1014, B1 => A_s(22), B2 => 
                           n1007, ZN => n160);
   U193 : INV_X1 port map( A => A_ns(20), ZN => n1140);
   U194 : INV_X1 port map( A => A_ns(21), ZN => n1141);
   U195 : INV_X1 port map( A => A_ns(24), ZN => n1032);
   U196 : INV_X1 port map( A => A_ns(25), ZN => n1033);
   U197 : INV_X1 port map( A => A_ns(26), ZN => n1034);
   U198 : INV_X1 port map( A => A_ns(27), ZN => n1035);
   U199 : INV_X1 port map( A => A_ns(28), ZN => n1036);
   U200 : INV_X1 port map( A => A_ns(29), ZN => n1037);
   U201 : INV_X1 port map( A => A_ns(30), ZN => n1038);
   U202 : INV_X1 port map( A => A_ns(31), ZN => n1039);
   U203 : INV_X1 port map( A => A_ns(32), ZN => n1040);
   U204 : INV_X1 port map( A => A_ns(33), ZN => n1041);
   U205 : INV_X1 port map( A => A_ns(34), ZN => n1042);
   U206 : INV_X1 port map( A => A_ns(35), ZN => n1043);
   U207 : INV_X1 port map( A => A_ns(36), ZN => n1044);
   U208 : INV_X1 port map( A => A_ns(37), ZN => n1045);
   U209 : INV_X1 port map( A => A_ns(38), ZN => n1046);
   U210 : INV_X1 port map( A => A_ns(39), ZN => n1047);
   U211 : INV_X1 port map( A => A_ns(40), ZN => n1048);
   U212 : INV_X1 port map( A => A_ns(41), ZN => n1049);
   U213 : INV_X1 port map( A => A_ns(42), ZN => n1050);
   U214 : INV_X1 port map( A => A_ns(43), ZN => n1051);
   U215 : INV_X1 port map( A => A_ns(44), ZN => n1052);
   U216 : INV_X1 port map( A => A_ns(45), ZN => n1053);
   U217 : INV_X1 port map( A => A_ns(46), ZN => n1054);
   U218 : INV_X1 port map( A => A_ns(47), ZN => n1055);
   U219 : INV_X1 port map( A => A_ns(48), ZN => n1056);
   U220 : INV_X1 port map( A => A_ns(49), ZN => n1057);
   U221 : INV_X1 port map( A => A_ns(50), ZN => n1058);
   U222 : INV_X1 port map( A => A_ns(51), ZN => n1059);
   U223 : INV_X1 port map( A => A_ns(52), ZN => n1060);
   U224 : INV_X1 port map( A => A_ns(53), ZN => n1061);
   U225 : INV_X1 port map( A => A_ns(54), ZN => n1062);
   U226 : INV_X1 port map( A => A_ns(55), ZN => n1063);
   U227 : INV_X1 port map( A => A_ns(23), ZN => n1064);
   U228 : INV_X1 port map( A => A_s(23), ZN => n1065);
   U229 : INV_X1 port map( A => A_s(24), ZN => n1066);
   U230 : INV_X1 port map( A => A_s(25), ZN => n1067);
   U231 : INV_X1 port map( A => A_s(26), ZN => n1068);
   U232 : INV_X1 port map( A => A_s(27), ZN => n1069);
   U235 : INV_X1 port map( A => A_s(28), ZN => n1070);
   U236 : INV_X1 port map( A => A_s(29), ZN => n1071);
   U237 : INV_X1 port map( A => A_s(30), ZN => n1072);
   U238 : INV_X1 port map( A => A_s(31), ZN => n1073);
   U239 : INV_X1 port map( A => A_s(32), ZN => n1074);
   U240 : INV_X1 port map( A => A_s(33), ZN => n1075);
   U241 : INV_X1 port map( A => n1077, ZN => A_so_36_port);
   U242 : INV_X1 port map( A => A_s(34), ZN => n1077);
   U243 : INV_X1 port map( A => A_s(35), ZN => n1078);
   U244 : INV_X1 port map( A => n1080, ZN => A_so_38_port);
   U245 : INV_X1 port map( A => A_s(36), ZN => n1080);
   U246 : INV_X1 port map( A => A_s(37), ZN => n1081);
   U247 : INV_X1 port map( A => A_s(38), ZN => n1082);
   U248 : INV_X1 port map( A => A_s(39), ZN => n1083);
   U249 : INV_X1 port map( A => A_s(40), ZN => n1084);
   U250 : INV_X1 port map( A => A_s(41), ZN => n1085);
   U251 : INV_X1 port map( A => A_s(42), ZN => n1086);
   U252 : INV_X1 port map( A => A_s(43), ZN => n1087);
   U253 : INV_X1 port map( A => A_s(44), ZN => n1088);
   U254 : INV_X1 port map( A => A_s(45), ZN => n1089);
   U255 : INV_X1 port map( A => A_s(46), ZN => n1090);
   U256 : INV_X1 port map( A => A_s(47), ZN => n1091);
   U257 : INV_X1 port map( A => A_s(48), ZN => n1092);
   U258 : INV_X1 port map( A => A_s(49), ZN => n1093);
   U259 : INV_X1 port map( A => A_s(50), ZN => n1094);
   U260 : INV_X1 port map( A => A_s(51), ZN => n1095);
   U261 : INV_X1 port map( A => A_s(52), ZN => n1096);
   U262 : INV_X1 port map( A => A_s(53), ZN => n1097);
   U263 : INV_X1 port map( A => A_s(54), ZN => n1098);
   U264 : INV_X1 port map( A => A_s(55), ZN => n1099);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT56_i22 is

   port( A_s, A_ns, B : in std_logic_vector (55 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (55 downto 0));

end BOOTHENC_NBIT56_i22;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT56_i22 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, O_55_port, O_54_port, O_53_port, O_52_port, O_51_port,
      O_50_port, O_49_port, O_48_port, O_47_port, O_46_port, O_45_port, 
      O_44_port, O_43_port, O_42_port, O_41_port, O_40_port, O_39_port, 
      O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, O_33_port, 
      O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, O_27_port, 
      O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, O_21_port, 
      O_20_port, O_19_port, O_18_port, O_17_port, O_16_port, O_15_port, 
      O_14_port, O_13_port, O_12_port, O_11_port, O_9_port, O_8_port, O_7_port,
      O_6_port, O_5_port, O_4_port, O_3_port, O_2_port, O_10_port, n111, n112, 
      n113, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n167, n168, n169, n170, n954, n955, n956, 
      n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, 
      n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, 
      n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, 
      n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, 
      n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, 
      n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, 
      n1024, n1025, n1026, n1027, n1028, n1029, A_so_50_port, n1031, n1032, 
      n1033, n1034, n1035, n1036, O_1_port, n1038, n1039, n1040, n1041, n1042, 
      n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, 
      n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, 
      n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, 
      n1073, n1074, n1075, n1076, n1077 : std_logic;

begin
   O <= ( O_55_port, O_54_port, O_53_port, O_52_port, O_51_port, O_50_port, 
      O_49_port, O_48_port, O_47_port, O_46_port, O_45_port, O_44_port, 
      O_43_port, O_42_port, O_41_port, O_40_port, O_39_port, O_38_port, 
      O_37_port, O_36_port, O_35_port, O_34_port, O_33_port, O_32_port, 
      O_31_port, O_30_port, O_29_port, O_28_port, O_27_port, O_26_port, 
      O_25_port, O_24_port, O_23_port, O_22_port, O_21_port, O_20_port, 
      O_19_port, O_18_port, O_17_port, O_16_port, O_15_port, O_14_port, 
      O_13_port, O_12_port, O_11_port, O_10_port, O_9_port, O_8_port, O_7_port,
      O_6_port, O_5_port, O_4_port, O_3_port, O_2_port, O_1_port, X_Logic0_port
      );
   A_so <= ( A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), A_so_50_port, A_s(47)
      , A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39),
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   A_nso <= ( A_ns(53), A_ns(52), A_ns(51), A_ns(50), A_ns(49), A_ns(48), 
      A_ns(47), A_ns(46), A_ns(45), A_ns(44), A_ns(43), A_ns(42), A_ns(41), 
      A_ns(40), A_ns(39), A_ns(38), A_ns(37), A_ns(36), A_ns(35), A_ns(34), 
      A_ns(33), A_ns(32), A_ns(31), A_ns(30), A_ns(29), A_ns(28), A_ns(27), 
      A_ns(26), A_ns(25), A_ns(24), A_ns(23), A_ns(22), A_ns(21), A_ns(20), 
      A_ns(19), A_ns(18), A_ns(17), A_ns(16), A_ns(15), A_ns(14), A_ns(13), 
      A_ns(12), A_ns(11), A_ns(10), A_ns(9), A_ns(8), A_ns(7), A_ns(6), A_ns(5)
      , A_ns(4), A_ns(3), A_ns(2), A_ns(1), A_ns(0), X_Logic0_port, 
      X_Logic0_port );
   
   X_Logic0_port <= '0';
   U224 : XOR2_X1 port map( A => B(21), B => B(22), Z => n170);
   U225 : NAND3_X1 port map( A1 => B(22), A2 => n1077, A3 => B(21), ZN => n119)
                           ;
   U2 : OAI221_X1 port map( B1 => n111, B2 => n972, C1 => n965, C2 => n1006, A 
                           => n153, ZN => O_25_port);
   U3 : INV_X1 port map( A => n969, ZN => n967);
   U4 : INV_X1 port map( A => n966, ZN => n964);
   U5 : INV_X1 port map( A => n966, ZN => n965);
   U6 : BUF_X1 port map( A => n955, Z => n958);
   U7 : INV_X1 port map( A => n969, ZN => n968);
   U8 : BUF_X1 port map( A => n955, Z => n959);
   U9 : AOI22_X1 port map( A1 => A_ns(54), A2 => n969, B1 => A_s(54), B2 => 
                           n966, ZN => n120);
   U10 : BUF_X1 port map( A => n956, Z => n960);
   U11 : BUF_X1 port map( A => n955, Z => n957);
   U12 : BUF_X1 port map( A => n956, Z => n961);
   U13 : OAI221_X1 port map( B1 => n111, B2 => n971, C1 => n965, C2 => n1005, A
                           => n154, ZN => O_24_port);
   U14 : OAI221_X1 port map( B1 => n111, B2 => n970, C1 => n965, C2 => n1004, A
                           => n155, ZN => O_23_port);
   U15 : AOI22_X1 port map( A1 => A_s(21), A2 => n958, B1 => A_ns(21), B2 => 
                           n962, ZN => n155);
   U16 : AOI22_X1 port map( A1 => A_s(23), A2 => n958, B1 => A_ns(23), B2 => 
                           n962, ZN => n153);
   U17 : OAI221_X1 port map( B1 => n111, B2 => n973, C1 => n965, C2 => n1007, A
                           => n152, ZN => O_26_port);
   U18 : AOI22_X1 port map( A1 => A_s(24), A2 => n958, B1 => A_ns(24), B2 => 
                           n962, ZN => n152);
   U19 : OAI221_X1 port map( B1 => n111, B2 => n974, C1 => n965, C2 => n1008, A
                           => n151, ZN => O_27_port);
   U20 : AOI22_X1 port map( A1 => A_s(25), A2 => n958, B1 => A_ns(25), B2 => 
                           n962, ZN => n151);
   U21 : AOI22_X1 port map( A1 => A_s(22), A2 => n958, B1 => A_ns(22), B2 => 
                           n962, ZN => n154);
   U22 : BUF_X1 port map( A => n1076, Z => n955);
   U23 : OAI221_X1 port map( B1 => n968, B2 => n989, C1 => n965, C2 => n1023, A
                           => n134, ZN => O_42_port);
   U24 : AOI22_X1 port map( A1 => A_s(40), A2 => n959, B1 => A_ns(40), B2 => 
                           n962, ZN => n134);
   U25 : OAI221_X1 port map( B1 => n111, B2 => n976, C1 => n965, C2 => n1010, A
                           => n149, ZN => O_29_port);
   U26 : AOI22_X1 port map( A1 => A_s(27), A2 => n958, B1 => A_ns(27), B2 => 
                           n962, ZN => n149);
   U27 : OAI221_X1 port map( B1 => n111, B2 => n978, C1 => n965, C2 => n1012, A
                           => n146, ZN => O_31_port);
   U28 : AOI22_X1 port map( A1 => A_s(29), A2 => n958, B1 => A_ns(29), B2 => 
                           n962, ZN => n146);
   U29 : OAI221_X1 port map( B1 => n968, B2 => n981, C1 => n965, C2 => n1015, A
                           => n143, ZN => O_34_port);
   U30 : AOI22_X1 port map( A1 => A_s(32), A2 => n959, B1 => A_ns(32), B2 => 
                           n962, ZN => n143);
   U31 : OAI221_X1 port map( B1 => n968, B2 => n983, C1 => n965, C2 => n1017, A
                           => n141, ZN => O_36_port);
   U32 : AOI22_X1 port map( A1 => A_s(34), A2 => n959, B1 => A_ns(34), B2 => 
                           n962, ZN => n141);
   U33 : OAI221_X1 port map( B1 => n968, B2 => n985, C1 => n965, C2 => n1019, A
                           => n139, ZN => O_38_port);
   U34 : AOI22_X1 port map( A1 => A_s(36), A2 => n959, B1 => A_ns(36), B2 => 
                           n962, ZN => n139);
   U35 : OAI221_X1 port map( B1 => n111, B2 => n980, C1 => n965, C2 => n1014, A
                           => n144, ZN => O_33_port);
   U36 : AOI22_X1 port map( A1 => A_s(31), A2 => n958, B1 => A_ns(31), B2 => 
                           n962, ZN => n144);
   U37 : OAI221_X1 port map( B1 => n968, B2 => n984, C1 => n965, C2 => n1018, A
                           => n140, ZN => O_37_port);
   U38 : AOI22_X1 port map( A1 => A_s(35), A2 => n959, B1 => A_ns(35), B2 => 
                           n962, ZN => n140);
   U39 : OAI221_X1 port map( B1 => n968, B2 => n986, C1 => n965, C2 => n1020, A
                           => n138, ZN => O_39_port);
   U40 : AOI22_X1 port map( A1 => A_s(37), A2 => n959, B1 => A_ns(37), B2 => 
                           n962, ZN => n138);
   U41 : OAI221_X1 port map( B1 => n968, B2 => n987, C1 => n965, C2 => n1021, A
                           => n136, ZN => O_40_port);
   U42 : AOI22_X1 port map( A1 => A_s(38), A2 => n959, B1 => A_ns(38), B2 => 
                           n962, ZN => n136);
   U43 : OAI221_X1 port map( B1 => n111, B2 => n977, C1 => n965, C2 => n1011, A
                           => n147, ZN => O_30_port);
   U44 : AOI22_X1 port map( A1 => A_s(28), A2 => n958, B1 => A_ns(28), B2 => 
                           n962, ZN => n147);
   U45 : OAI221_X1 port map( B1 => n111, B2 => n979, C1 => n965, C2 => n1013, A
                           => n145, ZN => O_32_port);
   U46 : AOI22_X1 port map( A1 => A_s(30), A2 => n958, B1 => A_ns(30), B2 => 
                           n962, ZN => n145);
   U47 : OAI221_X1 port map( B1 => n968, B2 => n988, C1 => n965, C2 => n1022, A
                           => n135, ZN => O_41_port);
   U48 : AOI22_X1 port map( A1 => A_s(39), A2 => n959, B1 => A_ns(39), B2 => 
                           n962, ZN => n135);
   U49 : OAI221_X1 port map( B1 => n968, B2 => n982, C1 => n965, C2 => n1016, A
                           => n142, ZN => O_35_port);
   U50 : AOI22_X1 port map( A1 => A_s(33), A2 => n959, B1 => A_ns(33), B2 => 
                           n962, ZN => n142);
   U51 : OAI221_X1 port map( B1 => n111, B2 => n975, C1 => n965, C2 => n1009, A
                           => n150, ZN => O_28_port);
   U52 : AOI22_X1 port map( A1 => A_s(26), A2 => n958, B1 => A_ns(26), B2 => 
                           n962, ZN => n150);
   U53 : OAI221_X1 port map( B1 => n968, B2 => n992, C1 => n965, C2 => n1026, A
                           => n131, ZN => O_45_port);
   U54 : AOI22_X1 port map( A1 => A_s(43), A2 => n960, B1 => A_ns(43), B2 => 
                           n963, ZN => n131);
   U55 : OAI221_X1 port map( B1 => n968, B2 => n998, C1 => n112, C2 => n1033, A
                           => n124, ZN => O_51_port);
   U56 : AOI22_X1 port map( A1 => A_s(49), A2 => n960, B1 => A_ns(49), B2 => 
                           n963, ZN => n124);
   U57 : OAI221_X1 port map( B1 => n968, B2 => n1001, C1 => n112, C2 => n1036, 
                           A => n121, ZN => O_54_port);
   U58 : AOI22_X1 port map( A1 => A_s(52), A2 => n960, B1 => A_ns(52), B2 => 
                           n963, ZN => n121);
   U59 : OAI221_X1 port map( B1 => n968, B2 => n991, C1 => n965, C2 => n1025, A
                           => n132, ZN => O_44_port);
   U60 : AOI22_X1 port map( A1 => A_s(42), A2 => n959, B1 => A_ns(42), B2 => 
                           n962, ZN => n132);
   U61 : OAI221_X1 port map( B1 => n968, B2 => n996, C1 => n112, C2 => n1031, A
                           => n127, ZN => O_49_port);
   U62 : AOI22_X1 port map( A1 => A_s(47), A2 => n960, B1 => A_ns(47), B2 => 
                           n963, ZN => n127);
   U63 : OAI221_X1 port map( B1 => n968, B2 => n1000, C1 => n112, C2 => n1035, 
                           A => n122, ZN => O_53_port);
   U64 : AOI22_X1 port map( A1 => A_s(51), A2 => n960, B1 => A_ns(51), B2 => 
                           n963, ZN => n122);
   U65 : OAI221_X1 port map( B1 => n968, B2 => n995, C1 => n112, C2 => n1029, A
                           => n128, ZN => O_48_port);
   U66 : AOI22_X1 port map( A1 => A_s(46), A2 => n960, B1 => A_ns(46), B2 => 
                           n963, ZN => n128);
   U67 : OAI221_X1 port map( B1 => n968, B2 => n990, C1 => n965, C2 => n1024, A
                           => n133, ZN => O_43_port);
   U68 : AOI22_X1 port map( A1 => A_s(41), A2 => n959, B1 => A_ns(41), B2 => 
                           n962, ZN => n133);
   U69 : OAI221_X1 port map( B1 => n968, B2 => n993, C1 => n965, C2 => n1027, A
                           => n130, ZN => O_46_port);
   U70 : AOI22_X1 port map( A1 => A_s(44), A2 => n960, B1 => A_ns(44), B2 => 
                           n963, ZN => n130);
   U71 : OAI221_X1 port map( B1 => n968, B2 => n994, C1 => n112, C2 => n1028, A
                           => n129, ZN => O_47_port);
   U72 : AOI22_X1 port map( A1 => A_s(45), A2 => n960, B1 => A_ns(45), B2 => 
                           n963, ZN => n129);
   U73 : OAI221_X1 port map( B1 => n968, B2 => n997, C1 => n112, C2 => n1032, A
                           => n125, ZN => O_50_port);
   U74 : AOI22_X1 port map( A1 => A_so_50_port, A2 => n960, B1 => A_ns(48), B2 
                           => n963, ZN => n125);
   U75 : OAI221_X1 port map( B1 => n968, B2 => n999, C1 => n112, C2 => n1034, A
                           => n123, ZN => O_52_port);
   U76 : AOI22_X1 port map( A1 => A_s(50), A2 => n960, B1 => A_ns(50), B2 => 
                           n963, ZN => n123);
   U77 : BUF_X1 port map( A => n1076, Z => n956);
   U78 : OAI221_X1 port map( B1 => n119, B2 => n1036, C1 => n954, C2 => n1001, 
                           A => n120, ZN => O_55_port);
   U79 : NAND2_X1 port map( A1 => n170, A2 => n964, ZN => n111);
   U80 : NAND2_X1 port map( A1 => n170, A2 => n1077, ZN => n112);
   U81 : INV_X1 port map( A => n119, ZN => n1076);
   U82 : INV_X1 port map( A => n954, ZN => n962);
   U83 : INV_X1 port map( A => n954, ZN => n963);
   U84 : OAI221_X1 port map( B1 => n967, B2 => n1002, C1 => n964, C2 => n1003, 
                           A => n156, ZN => O_22_port);
   U85 : AOI22_X1 port map( A1 => A_s(20), A2 => n957, B1 => A_ns(20), B2 => 
                           n963, ZN => n156);
   U86 : OR3_X1 port map( A1 => B(21), A2 => B(22), A3 => n1077, ZN => n954);
   U87 : INV_X1 port map( A => B(23), ZN => n1077);
   U88 : OAI221_X1 port map( B1 => n967, B2 => n1074, C1 => n964, C2 => n1075, 
                           A => n157, ZN => O_21_port);
   U89 : INV_X1 port map( A => A_ns(20), ZN => n1074);
   U90 : OAI221_X1 port map( B1 => n967, B2 => n1071, C1 => n964, C2 => n1073, 
                           A => n158, ZN => O_20_port);
   U91 : INV_X1 port map( A => A_ns(19), ZN => n1071);
   U92 : OAI221_X1 port map( B1 => n967, B2 => n1062, C1 => n964, C2 => n1064, 
                           A => n164, ZN => O_15_port);
   U93 : INV_X1 port map( A => A_ns(14), ZN => n1062);
   U94 : INV_X1 port map( A => A_s(14), ZN => n1064);
   U95 : OAI221_X1 port map( B1 => n967, B2 => n1063, C1 => n964, C2 => n1065, 
                           A => n163, ZN => O_16_port);
   U96 : INV_X1 port map( A => A_ns(15), ZN => n1063);
   U97 : OAI221_X1 port map( B1 => n967, B2 => n1066, C1 => n964, C2 => n1068, 
                           A => n162, ZN => O_17_port);
   U98 : INV_X1 port map( A => A_ns(16), ZN => n1066);
   U99 : OAI221_X1 port map( B1 => n967, B2 => n1067, C1 => n964, C2 => n1069, 
                           A => n161, ZN => O_18_port);
   U100 : INV_X1 port map( A => A_ns(17), ZN => n1067);
   U101 : OAI221_X1 port map( B1 => n967, B2 => n1070, C1 => n964, C2 => n1072,
                           A => n160, ZN => O_19_port);
   U102 : INV_X1 port map( A => A_ns(18), ZN => n1070);
   U103 : OAI221_X1 port map( B1 => n968, B2 => n1048, C1 => n112, C2 => n1050,
                           A => n116, ZN => O_7_port);
   U104 : INV_X1 port map( A => A_ns(6), ZN => n1048);
   U105 : INV_X1 port map( A => A_s(6), ZN => n1050);
   U106 : OAI221_X1 port map( B1 => n968, B2 => n1049, C1 => n112, C2 => n1051,
                           A => n115, ZN => O_8_port);
   U107 : INV_X1 port map( A => A_ns(7), ZN => n1049);
   U108 : INV_X1 port map( A => A_s(7), ZN => n1051);
   U109 : OAI221_X1 port map( B1 => n968, B2 => n1052, C1 => n112, C2 => n1053,
                           A => n113, ZN => O_9_port);
   U110 : AOI22_X1 port map( A1 => A_s(7), A2 => n961, B1 => A_ns(7), B2 => 
                           n963, ZN => n113);
   U111 : OAI221_X1 port map( B1 => n1053, B2 => n119, C1 => n1052, C2 => n954,
                           A => n169, ZN => O_10_port);
   U112 : AOI22_X1 port map( A1 => A_ns(9), A2 => n969, B1 => A_s(9), B2 => 
                           n966, ZN => n169);
   U113 : OAI221_X1 port map( B1 => n967, B2 => n1054, C1 => n964, C2 => n1056,
                           A => n168, ZN => O_11_port);
   U114 : INV_X1 port map( A => A_ns(10), ZN => n1054);
   U115 : INV_X1 port map( A => A_s(10), ZN => n1056);
   U116 : OAI221_X1 port map( B1 => n967, B2 => n1055, C1 => n964, C2 => n1057,
                           A => n167, ZN => O_12_port);
   U117 : INV_X1 port map( A => A_ns(11), ZN => n1055);
   U118 : INV_X1 port map( A => A_s(11), ZN => n1057);
   U119 : OAI221_X1 port map( B1 => n967, B2 => n1058, C1 => n964, C2 => n1060,
                           A => n166, ZN => O_13_port);
   U120 : INV_X1 port map( A => A_ns(12), ZN => n1058);
   U121 : INV_X1 port map( A => A_s(12), ZN => n1060);
   U122 : OAI221_X1 port map( B1 => n967, B2 => n1059, C1 => n964, C2 => n1061,
                           A => n165, ZN => O_14_port);
   U123 : INV_X1 port map( A => A_ns(13), ZN => n1059);
   U124 : INV_X1 port map( A => A_s(13), ZN => n1061);
   U125 : INV_X1 port map( A => n159, ZN => O_1_port);
   U126 : AOI22_X1 port map( A1 => n966, A2 => A_s(0), B1 => n969, B2 => 
                           A_ns(0), ZN => n159);
   U127 : OAI221_X1 port map( B1 => n111, B2 => n1038, C1 => n965, C2 => n1039,
                           A => n148, ZN => O_2_port);
   U128 : INV_X1 port map( A => A_ns(1), ZN => n1038);
   U129 : INV_X1 port map( A => A_s(1), ZN => n1039);
   U130 : OAI221_X1 port map( B1 => n968, B2 => n1040, C1 => n112, C2 => n1042,
                           A => n137, ZN => O_3_port);
   U131 : INV_X1 port map( A => A_ns(2), ZN => n1040);
   U132 : INV_X1 port map( A => A_s(2), ZN => n1042);
   U133 : OAI221_X1 port map( B1 => n967, B2 => n1041, C1 => n112, C2 => n1043,
                           A => n126, ZN => O_4_port);
   U134 : INV_X1 port map( A => A_ns(3), ZN => n1041);
   U135 : INV_X1 port map( A => A_s(3), ZN => n1043);
   U136 : OAI221_X1 port map( B1 => n967, B2 => n1044, C1 => n112, C2 => n1046,
                           A => n118, ZN => O_5_port);
   U137 : INV_X1 port map( A => A_ns(4), ZN => n1044);
   U138 : INV_X1 port map( A => A_s(4), ZN => n1046);
   U139 : OAI221_X1 port map( B1 => n967, B2 => n1045, C1 => n965, C2 => n1047,
                           A => n117, ZN => O_6_port);
   U140 : INV_X1 port map( A => A_ns(5), ZN => n1045);
   U141 : INV_X1 port map( A => A_s(5), ZN => n1047);
   U142 : INV_X1 port map( A => A_s(8), ZN => n1053);
   U143 : INV_X1 port map( A => A_ns(8), ZN => n1052);
   U144 : AOI22_X1 port map( A1 => A_s(0), A2 => n958, B1 => A_ns(0), B2 => 
                           n962, ZN => n148);
   U145 : AOI22_X1 port map( A1 => A_s(1), A2 => n959, B1 => A_ns(1), B2 => 
                           n962, ZN => n137);
   U146 : AOI22_X1 port map( A1 => A_s(2), A2 => n960, B1 => A_ns(2), B2 => 
                           n963, ZN => n126);
   U147 : AOI22_X1 port map( A1 => A_s(3), A2 => n960, B1 => A_ns(3), B2 => 
                           n963, ZN => n118);
   U148 : AOI22_X1 port map( A1 => A_s(4), A2 => n961, B1 => A_ns(4), B2 => 
                           n963, ZN => n117);
   U149 : AOI22_X1 port map( A1 => A_s(5), A2 => n961, B1 => A_ns(5), B2 => 
                           n963, ZN => n116);
   U150 : AOI22_X1 port map( A1 => A_s(6), A2 => n961, B1 => A_ns(6), B2 => 
                           n963, ZN => n115);
   U151 : AOI22_X1 port map( A1 => A_s(9), A2 => n957, B1 => A_ns(9), B2 => 
                           n963, ZN => n168);
   U152 : AOI22_X1 port map( A1 => A_s(10), A2 => n957, B1 => A_ns(10), B2 => 
                           n963, ZN => n167);
   U153 : AOI22_X1 port map( A1 => A_s(11), A2 => n957, B1 => A_ns(11), B2 => 
                           n963, ZN => n166);
   U154 : AOI22_X1 port map( A1 => A_s(12), A2 => n957, B1 => A_ns(12), B2 => 
                           n963, ZN => n165);
   U155 : AOI22_X1 port map( A1 => A_s(13), A2 => n957, B1 => A_ns(13), B2 => 
                           n963, ZN => n164);
   U156 : AOI22_X1 port map( A1 => A_s(14), A2 => n957, B1 => A_ns(14), B2 => 
                           n963, ZN => n163);
   U157 : AOI22_X1 port map( A1 => A_s(15), A2 => n957, B1 => A_ns(15), B2 => 
                           n963, ZN => n162);
   U158 : AOI22_X1 port map( A1 => A_s(16), A2 => n957, B1 => A_ns(16), B2 => 
                           n963, ZN => n161);
   U159 : AOI22_X1 port map( A1 => A_s(17), A2 => n957, B1 => A_ns(17), B2 => 
                           n963, ZN => n160);
   U160 : AOI22_X1 port map( A1 => A_s(18), A2 => n957, B1 => A_ns(18), B2 => 
                           n962, ZN => n158);
   U161 : AOI22_X1 port map( A1 => A_s(19), A2 => n957, B1 => A_ns(19), B2 => 
                           n962, ZN => n157);
   U162 : INV_X1 port map( A => A_s(15), ZN => n1065);
   U163 : INV_X1 port map( A => A_s(16), ZN => n1068);
   U164 : INV_X1 port map( A => A_s(17), ZN => n1069);
   U165 : INV_X1 port map( A => A_s(18), ZN => n1072);
   U166 : INV_X1 port map( A => A_s(19), ZN => n1073);
   U167 : INV_X1 port map( A => A_s(20), ZN => n1075);
   U168 : INV_X1 port map( A => n112, ZN => n966);
   U169 : INV_X1 port map( A => n111, ZN => n969);
   U170 : INV_X1 port map( A => A_ns(22), ZN => n970);
   U171 : INV_X1 port map( A => A_ns(23), ZN => n971);
   U172 : INV_X1 port map( A => A_ns(24), ZN => n972);
   U173 : INV_X1 port map( A => A_ns(25), ZN => n973);
   U174 : INV_X1 port map( A => A_ns(26), ZN => n974);
   U175 : INV_X1 port map( A => A_ns(27), ZN => n975);
   U176 : INV_X1 port map( A => A_ns(28), ZN => n976);
   U177 : INV_X1 port map( A => A_ns(29), ZN => n977);
   U178 : INV_X1 port map( A => A_ns(30), ZN => n978);
   U179 : INV_X1 port map( A => A_ns(31), ZN => n979);
   U180 : INV_X1 port map( A => A_ns(32), ZN => n980);
   U181 : INV_X1 port map( A => A_ns(33), ZN => n981);
   U182 : INV_X1 port map( A => A_ns(34), ZN => n982);
   U183 : INV_X1 port map( A => A_ns(35), ZN => n983);
   U184 : INV_X1 port map( A => A_ns(36), ZN => n984);
   U185 : INV_X1 port map( A => A_ns(37), ZN => n985);
   U186 : INV_X1 port map( A => A_ns(38), ZN => n986);
   U187 : INV_X1 port map( A => A_ns(39), ZN => n987);
   U188 : INV_X1 port map( A => A_ns(40), ZN => n988);
   U189 : INV_X1 port map( A => A_ns(41), ZN => n989);
   U190 : INV_X1 port map( A => A_ns(42), ZN => n990);
   U191 : INV_X1 port map( A => A_ns(43), ZN => n991);
   U192 : INV_X1 port map( A => A_ns(44), ZN => n992);
   U193 : INV_X1 port map( A => A_ns(45), ZN => n993);
   U194 : INV_X1 port map( A => A_ns(46), ZN => n994);
   U195 : INV_X1 port map( A => A_ns(47), ZN => n995);
   U196 : INV_X1 port map( A => A_ns(48), ZN => n996);
   U197 : INV_X1 port map( A => A_ns(49), ZN => n997);
   U198 : INV_X1 port map( A => A_ns(50), ZN => n998);
   U199 : INV_X1 port map( A => A_ns(51), ZN => n999);
   U200 : INV_X1 port map( A => A_ns(52), ZN => n1000);
   U201 : INV_X1 port map( A => A_ns(53), ZN => n1001);
   U202 : INV_X1 port map( A => A_ns(21), ZN => n1002);
   U203 : INV_X1 port map( A => A_s(21), ZN => n1003);
   U204 : INV_X1 port map( A => A_s(22), ZN => n1004);
   U205 : INV_X1 port map( A => A_s(23), ZN => n1005);
   U206 : INV_X1 port map( A => A_s(24), ZN => n1006);
   U207 : INV_X1 port map( A => A_s(25), ZN => n1007);
   U208 : INV_X1 port map( A => A_s(26), ZN => n1008);
   U209 : INV_X1 port map( A => A_s(27), ZN => n1009);
   U210 : INV_X1 port map( A => A_s(28), ZN => n1010);
   U211 : INV_X1 port map( A => A_s(29), ZN => n1011);
   U212 : INV_X1 port map( A => A_s(30), ZN => n1012);
   U213 : INV_X1 port map( A => A_s(31), ZN => n1013);
   U214 : INV_X1 port map( A => A_s(32), ZN => n1014);
   U215 : INV_X1 port map( A => A_s(33), ZN => n1015);
   U216 : INV_X1 port map( A => A_s(34), ZN => n1016);
   U217 : INV_X1 port map( A => A_s(35), ZN => n1017);
   U218 : INV_X1 port map( A => A_s(36), ZN => n1018);
   U219 : INV_X1 port map( A => A_s(37), ZN => n1019);
   U220 : INV_X1 port map( A => A_s(38), ZN => n1020);
   U221 : INV_X1 port map( A => A_s(39), ZN => n1021);
   U222 : INV_X1 port map( A => A_s(40), ZN => n1022);
   U223 : INV_X1 port map( A => A_s(41), ZN => n1023);
   U226 : INV_X1 port map( A => A_s(42), ZN => n1024);
   U227 : INV_X1 port map( A => A_s(43), ZN => n1025);
   U228 : INV_X1 port map( A => A_s(44), ZN => n1026);
   U229 : INV_X1 port map( A => A_s(45), ZN => n1027);
   U230 : INV_X1 port map( A => A_s(46), ZN => n1028);
   U231 : INV_X1 port map( A => A_s(47), ZN => n1029);
   U232 : INV_X1 port map( A => n1031, ZN => A_so_50_port);
   U233 : INV_X1 port map( A => A_s(48), ZN => n1031);
   U234 : INV_X1 port map( A => A_s(49), ZN => n1032);
   U235 : INV_X1 port map( A => A_s(50), ZN => n1033);
   U236 : INV_X1 port map( A => A_s(51), ZN => n1034);
   U237 : INV_X1 port map( A => A_s(52), ZN => n1035);
   U238 : INV_X1 port map( A => A_s(53), ZN => n1036);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT54_i20 is

   port( A_s, A_ns, B : in std_logic_vector (53 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (53 downto 0));

end BOOTHENC_NBIT54_i20;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT54_i20 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, O_53_port, O_52_port, O_51_port, O_50_port, O_49_port,
      O_48_port, O_47_port, O_46_port, O_45_port, O_44_port, O_43_port, 
      O_42_port, O_41_port, O_40_port, O_39_port, O_38_port, O_37_port, 
      O_36_port, O_35_port, O_34_port, O_33_port, O_32_port, O_31_port, 
      O_30_port, O_29_port, O_28_port, O_27_port, O_26_port, O_25_port, 
      O_24_port, O_23_port, O_22_port, O_21_port, O_20_port, O_19_port, 
      O_18_port, O_17_port, O_16_port, O_15_port, O_14_port, O_13_port, 
      O_12_port, O_11_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, 
      O_4_port, O_3_port, O_2_port, O_10_port, n107, n109, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n926, n927, n928, n929, n930, n931, n932, n933, n934, 
      n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, 
      n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, 
      n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, 
      n971, n972, n973, n974, A_so_21_port, n976, n977, n978, n979, n980, n981,
      n982, n983, n984, A_so_30_port, n986, n987, n988, n989, n990, n991, n992,
      n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, 
      n1004, n1005, n1006, n1007, n1008, A_so_53_port, n1010, O_1_port, n1012, 
      n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, 
      n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, 
      n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, 
      n1043, n1044, n1045, n1046, n1047 : std_logic;

begin
   O <= ( O_53_port, O_52_port, O_51_port, O_50_port, O_49_port, O_48_port, 
      O_47_port, O_46_port, O_45_port, O_44_port, O_43_port, O_42_port, 
      O_41_port, O_40_port, O_39_port, O_38_port, O_37_port, O_36_port, 
      O_35_port, O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, 
      O_29_port, O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, 
      O_23_port, O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, 
      O_17_port, O_16_port, O_15_port, O_14_port, O_13_port, O_12_port, 
      O_11_port, O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, 
      O_4_port, O_3_port, O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_so_53_port, A_s(50), A_s(49), A_s(48), A_s(47), A_s(46), A_s(45)
      , A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), A_s(38), A_s(37),
      A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), A_s(30), A_s(29), 
      A_so_30_port, A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), A_s(22), 
      A_s(21), A_s(20), A_so_21_port, A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   A_nso <= ( A_ns(51), A_ns(50), A_ns(49), A_ns(48), A_ns(47), A_ns(46), 
      A_ns(45), A_ns(44), A_ns(43), A_ns(42), A_ns(41), A_ns(40), A_ns(39), 
      A_ns(38), A_ns(37), A_ns(36), A_ns(35), A_ns(34), A_ns(33), A_ns(32), 
      A_ns(31), A_ns(30), A_ns(29), A_ns(28), A_ns(27), A_ns(26), A_ns(25), 
      A_ns(24), A_ns(23), A_ns(22), A_ns(21), A_ns(20), A_ns(19), A_ns(18), 
      A_ns(17), A_ns(16), A_ns(15), A_ns(14), A_ns(13), A_ns(12), A_ns(11), 
      A_ns(10), A_ns(9), A_ns(8), A_ns(7), A_ns(6), A_ns(5), A_ns(4), A_ns(3), 
      A_ns(2), A_ns(1), A_ns(0), X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U216 : XOR2_X1 port map( A => B(19), B => B(20), Z => n164);
   U217 : NAND3_X1 port map( A1 => B(20), A2 => n1047, A3 => B(19), ZN => n115)
                           ;
   U2 : OAI221_X1 port map( B1 => n940, B2 => n957, C1 => n938, C2 => n993, A 
                           => n135, ZN => O_36_port);
   U3 : OAI221_X1 port map( B1 => n107, B2 => n971, C1 => n937, C2 => n1007, A 
                           => n119, ZN => O_50_port);
   U4 : OAI221_X1 port map( B1 => n107, B2 => n972, C1 => n937, C2 => n1008, A 
                           => n118, ZN => O_51_port);
   U5 : OAI221_X1 port map( B1 => n940, B2 => n955, C1 => n938, C2 => n991, A 
                           => n137, ZN => O_34_port);
   U6 : OAI221_X1 port map( B1 => n939, B2 => n968, C1 => n938, C2 => n1004, A 
                           => n123, ZN => O_47_port);
   U7 : INV_X1 port map( A => A_ns(51), ZN => n973);
   U8 : INV_X1 port map( A => A_s(51), ZN => n1010);
   U9 : INV_X1 port map( A => n941, ZN => n939);
   U10 : INV_X1 port map( A => n941, ZN => n940);
   U11 : BUF_X1 port map( A => n928, Z => n930);
   U12 : BUF_X1 port map( A => n928, Z => n931);
   U13 : BUF_X1 port map( A => n928, Z => n932);
   U14 : BUF_X1 port map( A => n929, Z => n933);
   U15 : BUF_X1 port map( A => n929, Z => n934);
   U16 : OAI221_X1 port map( B1 => n107, B2 => n969, C1 => n937, C2 => n1005, A
                           => n122, ZN => O_48_port);
   U17 : AOI22_X1 port map( A1 => A_s(46), A2 => n933, B1 => A_ns(46), B2 => 
                           n936, ZN => n122);
   U18 : OAI221_X1 port map( B1 => n939, B2 => n942, C1 => n937, C2 => n977, A 
                           => n151, ZN => O_21_port);
   U19 : AOI22_X1 port map( A1 => A_so_21_port, A2 => n930, B1 => A_ns(19), B2 
                           => n935, ZN => n151);
   U20 : OAI221_X1 port map( B1 => n939, B2 => n943, C1 => n937, C2 => n978, A 
                           => n150, ZN => O_22_port);
   U21 : AOI22_X1 port map( A1 => A_s(20), A2 => n930, B1 => A_ns(20), B2 => 
                           n936, ZN => n150);
   U22 : OAI221_X1 port map( B1 => n940, B2 => n946, C1 => n938, C2 => n981, A 
                           => n147, ZN => O_25_port);
   U23 : AOI22_X1 port map( A1 => A_s(23), A2 => n931, B1 => A_ns(23), B2 => 
                           n936, ZN => n147);
   U24 : OAI221_X1 port map( B1 => n940, B2 => n945, C1 => n938, C2 => n980, A 
                           => n148, ZN => O_24_port);
   U25 : AOI22_X1 port map( A1 => A_s(22), A2 => n931, B1 => A_ns(22), B2 => 
                           n936, ZN => n148);
   U26 : OAI221_X1 port map( B1 => n940, B2 => n947, C1 => n938, C2 => n982, A 
                           => n146, ZN => O_26_port);
   U27 : AOI22_X1 port map( A1 => A_s(24), A2 => n931, B1 => A_ns(24), B2 => 
                           n936, ZN => n146);
   U28 : OAI221_X1 port map( B1 => n940, B2 => n948, C1 => n938, C2 => n983, A 
                           => n145, ZN => O_27_port);
   U29 : AOI22_X1 port map( A1 => A_s(25), A2 => n931, B1 => A_ns(25), B2 => 
                           n936, ZN => n145);
   U30 : OAI221_X1 port map( B1 => n940, B2 => n944, C1 => n938, C2 => n979, A 
                           => n149, ZN => O_23_port);
   U31 : AOI22_X1 port map( A1 => A_s(21), A2 => n931, B1 => A_ns(21), B2 => 
                           n935, ZN => n149);
   U32 : OAI221_X1 port map( B1 => n940, B2 => n949, C1 => n938, C2 => n984, A 
                           => n144, ZN => O_28_port);
   U33 : AOI22_X1 port map( A1 => A_s(26), A2 => n931, B1 => A_ns(26), B2 => 
                           n936, ZN => n144);
   U34 : OAI221_X1 port map( B1 => n940, B2 => n950, C1 => n938, C2 => n986, A 
                           => n143, ZN => O_29_port);
   U35 : AOI22_X1 port map( A1 => A_s(27), A2 => n931, B1 => A_ns(27), B2 => 
                           n936, ZN => n143);
   U36 : OAI221_X1 port map( B1 => n940, B2 => n951, C1 => n938, C2 => n987, A 
                           => n141, ZN => O_30_port);
   U37 : AOI22_X1 port map( A1 => A_so_30_port, A2 => n931, B1 => A_ns(28), B2 
                           => n936, ZN => n141);
   U38 : BUF_X1 port map( A => n1046, Z => n928);
   U39 : OAI221_X1 port map( B1 => n940, B2 => n961, C1 => n938, C2 => n997, A 
                           => n130, ZN => O_40_port);
   U40 : AOI22_X1 port map( A1 => A_s(38), A2 => n932, B1 => A_ns(38), B2 => 
                           n935, ZN => n130);
   U41 : OAI221_X1 port map( B1 => n940, B2 => n963, C1 => n938, C2 => n999, A 
                           => n128, ZN => O_42_port);
   U42 : AOI22_X1 port map( A1 => A_s(40), A2 => n932, B1 => A_ns(40), B2 => 
                           n935, ZN => n128);
   U43 : OAI221_X1 port map( B1 => n940, B2 => n953, C1 => n938, C2 => n989, A 
                           => n139, ZN => O_32_port);
   U44 : AOI22_X1 port map( A1 => A_s(30), A2 => n931, B1 => A_ns(30), B2 => 
                           n936, ZN => n139);
   U45 : OAI221_X1 port map( B1 => n940, B2 => n952, C1 => n938, C2 => n988, A 
                           => n140, ZN => O_31_port);
   U46 : AOI22_X1 port map( A1 => A_s(29), A2 => n931, B1 => A_ns(29), B2 => 
                           n936, ZN => n140);
   U47 : OAI221_X1 port map( B1 => n940, B2 => n954, C1 => n938, C2 => n990, A 
                           => n138, ZN => O_33_port);
   U48 : AOI22_X1 port map( A1 => A_s(31), A2 => n931, B1 => A_ns(31), B2 => 
                           n936, ZN => n138);
   U49 : OAI221_X1 port map( B1 => n940, B2 => n960, C1 => n938, C2 => n996, A 
                           => n132, ZN => O_39_port);
   U50 : AOI22_X1 port map( A1 => A_s(37), A2 => n932, B1 => A_ns(37), B2 => 
                           n935, ZN => n132);
   U51 : OAI221_X1 port map( B1 => n940, B2 => n958, C1 => n938, C2 => n994, A 
                           => n134, ZN => O_37_port);
   U52 : AOI22_X1 port map( A1 => A_s(35), A2 => n932, B1 => A_ns(35), B2 => 
                           n935, ZN => n134);
   U53 : OAI221_X1 port map( B1 => n940, B2 => n965, C1 => n938, C2 => n1001, A
                           => n126, ZN => O_44_port);
   U54 : AOI22_X1 port map( A1 => A_s(42), A2 => n932, B1 => A_ns(42), B2 => 
                           n935, ZN => n126);
   U55 : AOI22_X1 port map( A1 => A_s(32), A2 => n932, B1 => A_ns(32), B2 => 
                           n935, ZN => n137);
   U56 : AOI22_X1 port map( A1 => A_s(34), A2 => n932, B1 => A_ns(34), B2 => 
                           n935, ZN => n135);
   U57 : OAI221_X1 port map( B1 => n940, B2 => n962, C1 => n938, C2 => n998, A 
                           => n129, ZN => O_41_port);
   U58 : AOI22_X1 port map( A1 => A_s(39), A2 => n932, B1 => A_ns(39), B2 => 
                           n935, ZN => n129);
   U59 : OAI221_X1 port map( B1 => n940, B2 => n964, C1 => n938, C2 => n1000, A
                           => n127, ZN => O_43_port);
   U60 : AOI22_X1 port map( A1 => A_s(41), A2 => n932, B1 => A_ns(41), B2 => 
                           n935, ZN => n127);
   U61 : OAI221_X1 port map( B1 => n940, B2 => n959, C1 => n938, C2 => n995, A 
                           => n133, ZN => O_38_port);
   U62 : AOI22_X1 port map( A1 => A_s(36), A2 => n932, B1 => A_ns(36), B2 => 
                           n935, ZN => n133);
   U63 : OAI221_X1 port map( B1 => n940, B2 => n966, C1 => n938, C2 => n1002, A
                           => n125, ZN => O_45_port);
   U64 : AOI22_X1 port map( A1 => A_s(43), A2 => n933, B1 => A_ns(43), B2 => 
                           n936, ZN => n125);
   U65 : OAI221_X1 port map( B1 => n940, B2 => n956, C1 => n938, C2 => n992, A 
                           => n136, ZN => O_35_port);
   U66 : AOI22_X1 port map( A1 => A_s(33), A2 => n932, B1 => A_ns(33), B2 => 
                           n935, ZN => n136);
   U67 : OAI221_X1 port map( B1 => n107, B2 => n973, C1 => n937, C2 => n1010, A
                           => n117, ZN => O_52_port);
   U68 : AOI22_X1 port map( A1 => A_s(50), A2 => n933, B1 => A_ns(50), B2 => 
                           n936, ZN => n117);
   U69 : AOI22_X1 port map( A1 => A_s(49), A2 => n933, B1 => A_ns(49), B2 => 
                           n936, ZN => n118);
   U70 : OAI221_X1 port map( B1 => n939, B2 => n967, C1 => n938, C2 => n1003, A
                           => n124, ZN => O_46_port);
   U71 : AOI22_X1 port map( A1 => A_s(44), A2 => n933, B1 => A_ns(44), B2 => 
                           n936, ZN => n124);
   U72 : AOI22_X1 port map( A1 => A_s(45), A2 => n933, B1 => A_ns(45), B2 => 
                           n936, ZN => n123);
   U73 : OAI221_X1 port map( B1 => n107, B2 => n970, C1 => n937, C2 => n1006, A
                           => n121, ZN => O_49_port);
   U74 : AOI22_X1 port map( A1 => A_s(47), A2 => n933, B1 => A_ns(47), B2 => 
                           n936, ZN => n121);
   U75 : AOI22_X1 port map( A1 => A_s(48), A2 => n933, B1 => A_ns(48), B2 => 
                           n936, ZN => n119);
   U76 : AOI22_X1 port map( A1 => A_ns(52), A2 => n941, B1 => A_s(52), B2 => 
                           n926, ZN => n116);
   U77 : BUF_X1 port map( A => n1046, Z => n929);
   U78 : OAI221_X1 port map( B1 => n115, B2 => n1010, C1 => n927, C2 => n973, A
                           => n116, ZN => O_53_port);
   U79 : NAND2_X1 port map( A1 => n164, A2 => n937, ZN => n107);
   U80 : AND2_X1 port map( A1 => n164, A2 => n1047, ZN => n926);
   U81 : INV_X1 port map( A => n115, ZN => n1046);
   U82 : INV_X1 port map( A => n927, ZN => n935);
   U83 : INV_X1 port map( A => n927, ZN => n936);
   U84 : OAI221_X1 port map( B1 => n939, B2 => n974, C1 => n937, C2 => n976, A 
                           => n152, ZN => O_20_port);
   U85 : AOI22_X1 port map( A1 => A_s(18), A2 => n930, B1 => A_ns(18), B2 => 
                           n935, ZN => n152);
   U86 : OR3_X1 port map( A1 => B(19), A2 => B(20), A3 => n1047, ZN => n927);
   U87 : INV_X1 port map( A => B(21), ZN => n1047);
   U88 : OAI221_X1 port map( B1 => n939, B2 => n1036, C1 => n937, C2 => n1038, 
                           A => n158, ZN => O_15_port);
   U89 : INV_X1 port map( A => A_ns(14), ZN => n1036);
   U90 : INV_X1 port map( A => A_s(14), ZN => n1038);
   U91 : OAI221_X1 port map( B1 => n107, B2 => n1022, C1 => n937, C2 => n1024, 
                           A => n112, ZN => O_7_port);
   U92 : INV_X1 port map( A => A_ns(6), ZN => n1022);
   U93 : INV_X1 port map( A => A_s(6), ZN => n1024);
   U94 : OAI221_X1 port map( B1 => n107, B2 => n1023, C1 => n937, C2 => n1025, 
                           A => n111, ZN => O_8_port);
   U95 : INV_X1 port map( A => A_ns(7), ZN => n1023);
   U96 : INV_X1 port map( A => A_s(7), ZN => n1025);
   U97 : OAI221_X1 port map( B1 => n107, B2 => n1026, C1 => n937, C2 => n1027, 
                           A => n109, ZN => O_9_port);
   U98 : AOI22_X1 port map( A1 => A_s(7), A2 => n934, B1 => A_ns(7), B2 => n936
                           , ZN => n109);
   U99 : OAI221_X1 port map( B1 => n1027, B2 => n115, C1 => n1026, C2 => n927, 
                           A => n163, ZN => O_10_port);
   U100 : AOI22_X1 port map( A1 => A_ns(9), A2 => n941, B1 => A_s(9), B2 => 
                           n926, ZN => n163);
   U101 : OAI221_X1 port map( B1 => n939, B2 => n1028, C1 => n937, C2 => n1030,
                           A => n162, ZN => O_11_port);
   U102 : INV_X1 port map( A => A_ns(10), ZN => n1028);
   U103 : INV_X1 port map( A => A_s(10), ZN => n1030);
   U104 : OAI221_X1 port map( B1 => n939, B2 => n1029, C1 => n937, C2 => n1031,
                           A => n161, ZN => O_12_port);
   U105 : INV_X1 port map( A => A_ns(11), ZN => n1029);
   U106 : INV_X1 port map( A => A_s(11), ZN => n1031);
   U107 : OAI221_X1 port map( B1 => n939, B2 => n1032, C1 => n937, C2 => n1034,
                           A => n160, ZN => O_13_port);
   U108 : INV_X1 port map( A => A_ns(12), ZN => n1032);
   U109 : INV_X1 port map( A => A_s(12), ZN => n1034);
   U110 : OAI221_X1 port map( B1 => n939, B2 => n1033, C1 => n937, C2 => n1035,
                           A => n159, ZN => O_14_port);
   U111 : INV_X1 port map( A => A_ns(13), ZN => n1033);
   U112 : INV_X1 port map( A => A_s(13), ZN => n1035);
   U113 : INV_X1 port map( A => n153, ZN => O_1_port);
   U114 : AOI22_X1 port map( A1 => n926, A2 => A_s(0), B1 => n941, B2 => 
                           A_ns(0), ZN => n153);
   U115 : OAI221_X1 port map( B1 => n940, B2 => n1012, C1 => n938, C2 => n1013,
                           A => n142, ZN => O_2_port);
   U116 : INV_X1 port map( A => A_ns(1), ZN => n1012);
   U117 : INV_X1 port map( A => A_s(1), ZN => n1013);
   U118 : OAI221_X1 port map( B1 => n107, B2 => n1014, C1 => n937, C2 => n1016,
                           A => n131, ZN => O_3_port);
   U119 : INV_X1 port map( A => A_ns(2), ZN => n1014);
   U120 : INV_X1 port map( A => A_s(2), ZN => n1016);
   U121 : OAI221_X1 port map( B1 => n107, B2 => n1015, C1 => n937, C2 => n1017,
                           A => n120, ZN => O_4_port);
   U122 : INV_X1 port map( A => A_ns(3), ZN => n1015);
   U123 : INV_X1 port map( A => A_s(3), ZN => n1017);
   U124 : OAI221_X1 port map( B1 => n107, B2 => n1018, C1 => n937, C2 => n1020,
                           A => n114, ZN => O_5_port);
   U125 : INV_X1 port map( A => A_ns(4), ZN => n1018);
   U126 : INV_X1 port map( A => A_s(4), ZN => n1020);
   U127 : OAI221_X1 port map( B1 => n940, B2 => n1019, C1 => n937, C2 => n1021,
                           A => n113, ZN => O_6_port);
   U128 : INV_X1 port map( A => A_ns(5), ZN => n1019);
   U129 : INV_X1 port map( A => A_s(5), ZN => n1021);
   U130 : OAI221_X1 port map( B1 => n939, B2 => n1037, C1 => n937, C2 => n1039,
                           A => n157, ZN => O_16_port);
   U131 : INV_X1 port map( A => A_ns(15), ZN => n1037);
   U132 : INV_X1 port map( A => A_s(15), ZN => n1039);
   U133 : AOI22_X1 port map( A1 => A_s(14), A2 => n930, B1 => A_ns(14), B2 => 
                           n935, ZN => n157);
   U134 : OAI221_X1 port map( B1 => n939, B2 => n1044, C1 => n937, C2 => n1045,
                           A => n154, ZN => O_19_port);
   U135 : INV_X1 port map( A => A_ns(18), ZN => n1044);
   U136 : INV_X1 port map( A => A_s(18), ZN => n1045);
   U137 : AOI22_X1 port map( A1 => A_s(17), A2 => n930, B1 => A_ns(17), B2 => 
                           n935, ZN => n154);
   U138 : OAI221_X1 port map( B1 => n939, B2 => n1040, C1 => n937, C2 => n1042,
                           A => n156, ZN => O_17_port);
   U139 : INV_X1 port map( A => A_ns(16), ZN => n1040);
   U140 : INV_X1 port map( A => A_s(16), ZN => n1042);
   U141 : AOI22_X1 port map( A1 => A_s(15), A2 => n930, B1 => A_ns(15), B2 => 
                           n935, ZN => n156);
   U142 : OAI221_X1 port map( B1 => n939, B2 => n1041, C1 => n937, C2 => n1043,
                           A => n155, ZN => O_18_port);
   U143 : INV_X1 port map( A => A_ns(17), ZN => n1041);
   U144 : INV_X1 port map( A => A_s(17), ZN => n1043);
   U145 : AOI22_X1 port map( A1 => A_s(16), A2 => n930, B1 => A_ns(16), B2 => 
                           n935, ZN => n155);
   U146 : INV_X1 port map( A => A_s(8), ZN => n1027);
   U147 : INV_X1 port map( A => A_ns(8), ZN => n1026);
   U148 : AOI22_X1 port map( A1 => A_s(0), A2 => n931, B1 => A_ns(0), B2 => 
                           n936, ZN => n142);
   U149 : AOI22_X1 port map( A1 => A_s(1), A2 => n932, B1 => A_ns(1), B2 => 
                           n935, ZN => n131);
   U150 : AOI22_X1 port map( A1 => A_s(2), A2 => n933, B1 => A_ns(2), B2 => 
                           n936, ZN => n120);
   U151 : AOI22_X1 port map( A1 => A_s(3), A2 => n933, B1 => A_ns(3), B2 => 
                           n936, ZN => n114);
   U152 : AOI22_X1 port map( A1 => A_s(4), A2 => n933, B1 => A_ns(4), B2 => 
                           n936, ZN => n113);
   U153 : AOI22_X1 port map( A1 => A_s(5), A2 => n933, B1 => A_ns(5), B2 => 
                           n936, ZN => n112);
   U154 : AOI22_X1 port map( A1 => A_s(6), A2 => n934, B1 => A_ns(6), B2 => 
                           n936, ZN => n111);
   U155 : AOI22_X1 port map( A1 => A_s(9), A2 => n930, B1 => A_ns(9), B2 => 
                           n935, ZN => n162);
   U156 : AOI22_X1 port map( A1 => A_s(10), A2 => n930, B1 => A_ns(10), B2 => 
                           n935, ZN => n161);
   U157 : AOI22_X1 port map( A1 => A_s(11), A2 => n930, B1 => A_ns(11), B2 => 
                           n935, ZN => n160);
   U158 : AOI22_X1 port map( A1 => A_s(12), A2 => n930, B1 => A_ns(12), B2 => 
                           n935, ZN => n159);
   U159 : AOI22_X1 port map( A1 => A_s(13), A2 => n930, B1 => A_ns(13), B2 => 
                           n935, ZN => n158);
   U160 : INV_X1 port map( A => n926, ZN => n937);
   U161 : INV_X1 port map( A => n926, ZN => n938);
   U162 : INV_X1 port map( A => n107, ZN => n941);
   U163 : INV_X1 port map( A => A_ns(20), ZN => n942);
   U164 : INV_X1 port map( A => A_ns(21), ZN => n943);
   U165 : INV_X1 port map( A => A_ns(22), ZN => n944);
   U166 : INV_X1 port map( A => A_ns(23), ZN => n945);
   U167 : INV_X1 port map( A => A_ns(24), ZN => n946);
   U168 : INV_X1 port map( A => A_ns(25), ZN => n947);
   U169 : INV_X1 port map( A => A_ns(26), ZN => n948);
   U170 : INV_X1 port map( A => A_ns(27), ZN => n949);
   U171 : INV_X1 port map( A => A_ns(28), ZN => n950);
   U172 : INV_X1 port map( A => A_ns(29), ZN => n951);
   U173 : INV_X1 port map( A => A_ns(30), ZN => n952);
   U174 : INV_X1 port map( A => A_ns(31), ZN => n953);
   U175 : INV_X1 port map( A => A_ns(32), ZN => n954);
   U176 : INV_X1 port map( A => A_ns(33), ZN => n955);
   U177 : INV_X1 port map( A => A_ns(34), ZN => n956);
   U178 : INV_X1 port map( A => A_ns(35), ZN => n957);
   U179 : INV_X1 port map( A => A_ns(36), ZN => n958);
   U180 : INV_X1 port map( A => A_ns(37), ZN => n959);
   U181 : INV_X1 port map( A => A_ns(38), ZN => n960);
   U182 : INV_X1 port map( A => A_ns(39), ZN => n961);
   U183 : INV_X1 port map( A => A_ns(40), ZN => n962);
   U184 : INV_X1 port map( A => A_ns(41), ZN => n963);
   U185 : INV_X1 port map( A => A_ns(42), ZN => n964);
   U186 : INV_X1 port map( A => A_ns(43), ZN => n965);
   U187 : INV_X1 port map( A => A_ns(44), ZN => n966);
   U188 : INV_X1 port map( A => A_ns(45), ZN => n967);
   U189 : INV_X1 port map( A => A_ns(46), ZN => n968);
   U190 : INV_X1 port map( A => A_ns(47), ZN => n969);
   U191 : INV_X1 port map( A => A_ns(48), ZN => n970);
   U192 : INV_X1 port map( A => A_ns(49), ZN => n971);
   U193 : INV_X1 port map( A => A_ns(50), ZN => n972);
   U194 : INV_X1 port map( A => A_ns(19), ZN => n974);
   U195 : INV_X1 port map( A => n976, ZN => A_so_21_port);
   U196 : INV_X1 port map( A => A_s(19), ZN => n976);
   U197 : INV_X1 port map( A => A_s(20), ZN => n977);
   U198 : INV_X1 port map( A => A_s(21), ZN => n978);
   U199 : INV_X1 port map( A => A_s(22), ZN => n979);
   U200 : INV_X1 port map( A => A_s(23), ZN => n980);
   U201 : INV_X1 port map( A => A_s(24), ZN => n981);
   U202 : INV_X1 port map( A => A_s(25), ZN => n982);
   U203 : INV_X1 port map( A => A_s(26), ZN => n983);
   U204 : INV_X1 port map( A => A_s(27), ZN => n984);
   U205 : INV_X1 port map( A => n986, ZN => A_so_30_port);
   U206 : INV_X1 port map( A => A_s(28), ZN => n986);
   U207 : INV_X1 port map( A => A_s(29), ZN => n987);
   U208 : INV_X1 port map( A => A_s(30), ZN => n988);
   U209 : INV_X1 port map( A => A_s(31), ZN => n989);
   U210 : INV_X1 port map( A => A_s(32), ZN => n990);
   U211 : INV_X1 port map( A => A_s(33), ZN => n991);
   U212 : INV_X1 port map( A => A_s(34), ZN => n992);
   U213 : INV_X1 port map( A => A_s(35), ZN => n993);
   U214 : INV_X1 port map( A => A_s(36), ZN => n994);
   U215 : INV_X1 port map( A => A_s(37), ZN => n995);
   U218 : INV_X1 port map( A => A_s(38), ZN => n996);
   U219 : INV_X1 port map( A => A_s(39), ZN => n997);
   U220 : INV_X1 port map( A => A_s(40), ZN => n998);
   U221 : INV_X1 port map( A => A_s(41), ZN => n999);
   U222 : INV_X1 port map( A => A_s(42), ZN => n1000);
   U223 : INV_X1 port map( A => A_s(43), ZN => n1001);
   U224 : INV_X1 port map( A => A_s(44), ZN => n1002);
   U225 : INV_X1 port map( A => A_s(45), ZN => n1003);
   U226 : INV_X1 port map( A => A_s(46), ZN => n1004);
   U227 : INV_X1 port map( A => A_s(47), ZN => n1005);
   U228 : INV_X1 port map( A => A_s(48), ZN => n1006);
   U229 : INV_X1 port map( A => A_s(49), ZN => n1007);
   U230 : INV_X1 port map( A => A_s(50), ZN => n1008);
   U231 : INV_X1 port map( A => n1010, ZN => A_so_53_port);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT52_i18 is

   port( A_s, A_ns, B : in std_logic_vector (51 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (51 downto 0));

end BOOTHENC_NBIT52_i18;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT52_i18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI221_X4
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, O_49_port, O_50_port, O_51_port, O_48_port, O_47_port,
      O_46_port, O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, 
      O_40_port, O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, 
      O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, 
      O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, 
      O_22_port, O_21_port, O_20_port, O_19_port, O_2_port, O_3_port, O_4_port,
      O_5_port, O_6_port, O_7_port, O_8_port, O_9_port, O_10_port, O_11_port, 
      O_12_port, O_13_port, O_14_port, O_15_port, O_16_port, O_17_port, 
      O_18_port, n105, n107, n108, n109, n110, n111, n112, n113, n114, n115, 
      n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, 
      n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, 
      n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n949, n950, n951, n952, n953, 
      n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, 
      n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, 
      n978, n979, n980, n981, n982, n983, n984, A_nso_41_port, n986, n987, n988
      , n989, n990, n991, A_nso_47_port, n993, n994, n995, A_nso_50_port, n997,
      A_nso_51_port, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, 
      n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, 
      n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, 
      n1027, n1028, n1029, n1030, n1031, n1032, n1033, O_1_port, n1035, n1036, 
      n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, 
      n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, 
      n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066 : 
      std_logic;

begin
   O <= ( O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, O_46_port, 
      O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, O_40_port, 
      O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, 
      O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, 
      O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, 
      O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, O_16_port, 
      O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, O_10_port, 
      O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, O_3_port, 
      O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(49), A_s(48), A_s(47), A_s(46), A_s(45), A_s(44), A_s(43), 
      A_s(42), A_s(41), A_s(40), A_s(39), A_s(38), A_s(37), A_s(36), A_s(35), 
      A_s(34), A_s(33), A_s(32), A_s(31), A_s(30), A_s(29), A_s(28), A_s(27), 
      A_s(26), A_s(25), A_s(24), A_s(23), A_s(22), A_s(21), A_s(20), A_s(19), 
      A_s(18), A_s(17), A_s(16), A_s(15), A_s(14), A_s(13), A_s(12), A_s(11), 
      A_s(10), A_s(9), A_s(8), A_s(7), A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), 
      A_s(1), A_s(0), X_Logic0_port, X_Logic0_port );
   A_nso <= ( A_nso_51_port, A_nso_50_port, A_ns(47), A_ns(46), A_nso_47_port, 
      A_ns(44), A_ns(43), A_ns(42), A_ns(41), A_ns(40), A_nso_41_port, A_ns(38)
      , A_ns(37), A_ns(36), A_ns(35), A_ns(34), A_ns(33), A_ns(32), A_ns(31), 
      A_ns(30), A_ns(29), A_ns(28), A_ns(27), A_ns(26), A_ns(25), A_ns(24), 
      A_ns(23), A_ns(22), A_ns(21), A_ns(20), A_ns(19), A_ns(18), A_ns(17), 
      A_ns(16), A_ns(15), A_ns(14), A_ns(13), A_ns(12), A_ns(11), A_ns(10), 
      A_ns(9), A_ns(8), A_ns(7), A_ns(6), A_ns(5), A_ns(4), A_ns(3), A_ns(2), 
      A_ns(1), A_ns(0), X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U208 : XOR2_X1 port map( A => B(17), B => B(18), Z => n158);
   U209 : NAND3_X1 port map( A1 => B(18), A2 => n1066, A3 => B(17), ZN => n111)
                           ;
   U2 : OAI221_X1 port map( B1 => n962, B2 => n972, C1 => n961, C2 => n1010, A 
                           => n139, ZN => O_27_port);
   U3 : OAI221_X1 port map( B1 => n963, B2 => n993, C1 => n961, C2 => n1029, A 
                           => n118, ZN => O_46_port);
   U4 : OAI221_X4 port map( B1 => n963, B2 => n997, C1 => n961, C2 => n1032, A 
                           => n115, ZN => O_49_port);
   U5 : INV_X1 port map( A => A_ns(49), ZN => n999);
   U6 : BUF_X1 port map( A => n952, Z => n954);
   U7 : BUF_X1 port map( A => n952, Z => n955);
   U8 : BUF_X1 port map( A => n953, Z => n956);
   U9 : BUF_X1 port map( A => n953, Z => n957);
   U10 : INV_X1 port map( A => A_s(49), ZN => n1033);
   U11 : INV_X1 port map( A => n950, ZN => n961);
   U12 : OAI221_X1 port map( B1 => n962, B2 => n968, C1 => n961, C2 => n1006, A
                           => n143, ZN => O_23_port);
   U13 : AOI22_X1 port map( A1 => A_s(21), A2 => n955, B1 => A_ns(21), B2 => 
                           n958, ZN => n143);
   U14 : AOI22_X1 port map( A1 => A_s(25), A2 => n955, B1 => A_ns(25), B2 => 
                           n958, ZN => n139);
   U15 : OAI221_X1 port map( B1 => n962, B2 => n967, C1 => n960, C2 => n1005, A
                           => n144, ZN => O_22_port);
   U16 : AOI22_X1 port map( A1 => A_s(20), A2 => n954, B1 => A_ns(20), B2 => 
                           n959, ZN => n144);
   U17 : OAI221_X1 port map( B1 => n962, B2 => n966, C1 => n960, C2 => n1004, A
                           => n145, ZN => O_21_port);
   U18 : AOI22_X1 port map( A1 => A_s(19), A2 => n954, B1 => A_ns(19), B2 => 
                           n959, ZN => n145);
   U19 : OAI221_X1 port map( B1 => n963, B2 => n964, C1 => n960, C2 => n1002, A
                           => n148, ZN => O_19_port);
   U20 : AOI22_X1 port map( A1 => A_s(17), A2 => n954, B1 => A_ns(17), B2 => 
                           n958, ZN => n148);
   U21 : OAI221_X1 port map( B1 => n962, B2 => n971, C1 => n961, C2 => n1009, A
                           => n140, ZN => O_26_port);
   U22 : AOI22_X1 port map( A1 => A_s(24), A2 => n955, B1 => A_ns(24), B2 => 
                           n958, ZN => n140);
   U23 : OAI221_X1 port map( B1 => n962, B2 => n976, C1 => n961, C2 => n1014, A
                           => n134, ZN => O_31_port);
   U24 : AOI22_X1 port map( A1 => A_s(29), A2 => n955, B1 => A_ns(29), B2 => 
                           n958, ZN => n134);
   U25 : OAI221_X1 port map( B1 => n962, B2 => n975, C1 => n961, C2 => n1013, A
                           => n135, ZN => O_30_port);
   U26 : AOI22_X1 port map( A1 => A_s(28), A2 => n955, B1 => A_ns(28), B2 => 
                           n958, ZN => n135);
   U27 : OAI221_X1 port map( B1 => n962, B2 => n977, C1 => n961, C2 => n1015, A
                           => n133, ZN => O_32_port);
   U28 : AOI22_X1 port map( A1 => A_s(30), A2 => n955, B1 => A_ns(30), B2 => 
                           n958, ZN => n133);
   U29 : OAI221_X1 port map( B1 => n962, B2 => n965, C1 => n960, C2 => n1003, A
                           => n146, ZN => O_20_port);
   U30 : AOI22_X1 port map( A1 => A_s(18), A2 => n954, B1 => A_ns(18), B2 => 
                           n958, ZN => n146);
   U31 : OAI221_X1 port map( B1 => n962, B2 => n978, C1 => n961, C2 => n1016, A
                           => n132, ZN => O_33_port);
   U32 : AOI22_X1 port map( A1 => A_s(31), A2 => n955, B1 => A_ns(31), B2 => 
                           n958, ZN => n132);
   U33 : OAI221_X1 port map( B1 => n962, B2 => n969, C1 => n961, C2 => n1007, A
                           => n142, ZN => O_24_port);
   U34 : AOI22_X1 port map( A1 => A_s(22), A2 => n955, B1 => A_ns(22), B2 => 
                           n958, ZN => n142);
   U35 : OAI221_X1 port map( B1 => n962, B2 => n970, C1 => n961, C2 => n1008, A
                           => n141, ZN => O_25_port);
   U36 : AOI22_X1 port map( A1 => A_s(23), A2 => n955, B1 => A_ns(23), B2 => 
                           n958, ZN => n141);
   U37 : OAI221_X1 port map( B1 => n962, B2 => n973, C1 => n961, C2 => n1011, A
                           => n138, ZN => O_28_port);
   U38 : AOI22_X1 port map( A1 => A_s(26), A2 => n955, B1 => A_ns(26), B2 => 
                           n958, ZN => n138);
   U39 : OAI221_X1 port map( B1 => n962, B2 => n974, C1 => n961, C2 => n1012, A
                           => n137, ZN => O_29_port);
   U40 : AOI22_X1 port map( A1 => A_s(27), A2 => n955, B1 => A_ns(27), B2 => 
                           n958, ZN => n137);
   U41 : BUF_X1 port map( A => n1065, Z => n952);
   U42 : AOI22_X1 port map( A1 => A_s(44), A2 => n957, B1 => A_ns(44), B2 => 
                           n959, ZN => n118);
   U43 : OAI221_X1 port map( B1 => n963, B2 => n991, C1 => n961, C2 => n1028, A
                           => n119, ZN => O_45_port);
   U44 : AOI22_X1 port map( A1 => A_s(43), A2 => n957, B1 => A_ns(43), B2 => 
                           n959, ZN => n119);
   U45 : OAI221_X1 port map( B1 => n963, B2 => n983, C1 => n961, C2 => n1021, A
                           => n127, ZN => O_38_port);
   U46 : AOI22_X1 port map( A1 => A_s(36), A2 => n956, B1 => A_ns(36), B2 => 
                           n959, ZN => n127);
   U47 : OAI221_X1 port map( B1 => n963, B2 => n990, C1 => n961, C2 => n1027, A
                           => n120, ZN => O_44_port);
   U48 : AOI22_X1 port map( A1 => A_s(42), A2 => n956, B1 => A_ns(42), B2 => 
                           n959, ZN => n120);
   U49 : OAI221_X1 port map( B1 => n963, B2 => n995, C1 => n960, C2 => n1031, A
                           => n116, ZN => O_48_port);
   U50 : AOI22_X1 port map( A1 => A_s(46), A2 => n957, B1 => A_ns(46), B2 => 
                           n959, ZN => n116);
   U51 : AOI22_X1 port map( A1 => A_s(47), A2 => n957, B1 => A_ns(47), B2 => 
                           n959, ZN => n115);
   U52 : OAI221_X1 port map( B1 => n963, B2 => n986, C1 => n961, C2 => n1023, A
                           => n124, ZN => O_40_port);
   U53 : AOI22_X1 port map( A1 => A_s(38), A2 => n956, B1 => A_ns(38), B2 => 
                           n959, ZN => n124);
   U54 : OAI221_X1 port map( B1 => n963, B2 => n980, C1 => n961, C2 => n1018, A
                           => n130, ZN => O_35_port);
   U55 : AOI22_X1 port map( A1 => A_s(33), A2 => n956, B1 => A_ns(33), B2 => 
                           n959, ZN => n130);
   U56 : OAI221_X1 port map( B1 => n963, B2 => n984, C1 => n961, C2 => n1022, A
                           => n126, ZN => O_39_port);
   U57 : AOI22_X1 port map( A1 => A_s(37), A2 => n956, B1 => A_ns(37), B2 => 
                           n959, ZN => n126);
   U58 : OAI221_X1 port map( B1 => n963, B2 => n987, C1 => n961, C2 => n1024, A
                           => n123, ZN => O_41_port);
   U59 : AOI22_X1 port map( A1 => A_s(39), A2 => n956, B1 => A_nso_41_port, B2 
                           => n959, ZN => n123);
   U60 : OAI221_X1 port map( B1 => n963, B2 => n989, C1 => n961, C2 => n1026, A
                           => n121, ZN => O_43_port);
   U61 : AOI22_X1 port map( A1 => A_s(41), A2 => n956, B1 => A_ns(41), B2 => 
                           n959, ZN => n121);
   U62 : OAI221_X1 port map( B1 => n963, B2 => n994, C1 => n960, C2 => n1030, A
                           => n117, ZN => O_47_port);
   U63 : AOI22_X1 port map( A1 => A_s(45), A2 => n957, B1 => A_nso_47_port, B2 
                           => n959, ZN => n117);
   U64 : OAI221_X1 port map( B1 => n963, B2 => n979, C1 => n961, C2 => n1017, A
                           => n131, ZN => O_34_port);
   U65 : AOI22_X1 port map( A1 => A_s(32), A2 => n956, B1 => A_ns(32), B2 => 
                           n959, ZN => n131);
   U66 : OAI221_X1 port map( B1 => n963, B2 => n981, C1 => n961, C2 => n1019, A
                           => n129, ZN => O_36_port);
   U67 : AOI22_X1 port map( A1 => A_s(34), A2 => n956, B1 => A_ns(34), B2 => 
                           n959, ZN => n129);
   U68 : OAI221_X1 port map( B1 => n963, B2 => n988, C1 => n961, C2 => n1025, A
                           => n122, ZN => O_42_port);
   U69 : AOI22_X1 port map( A1 => A_s(40), A2 => n956, B1 => A_ns(40), B2 => 
                           n959, ZN => n122);
   U70 : OAI221_X1 port map( B1 => n963, B2 => n982, C1 => n961, C2 => n1020, A
                           => n128, ZN => O_37_port);
   U71 : AOI22_X1 port map( A1 => A_s(35), A2 => n956, B1 => A_ns(35), B2 => 
                           n959, ZN => n128);
   U72 : BUF_X1 port map( A => n1065, Z => n953);
   U73 : INV_X1 port map( A => n949, ZN => n963);
   U74 : OAI221_X1 port map( B1 => n963, B2 => n999, C1 => n960, C2 => n1033, A
                           => n113, ZN => O_50_port);
   U75 : AOI22_X1 port map( A1 => A_s(48), A2 => n957, B1 => A_nso_50_port, B2 
                           => n959, ZN => n113);
   U76 : AOI22_X1 port map( A1 => A_ns(50), A2 => n949, B1 => A_s(50), B2 => 
                           n950, ZN => n112);
   U77 : OAI221_X1 port map( B1 => n111, B2 => n1033, C1 => n951, C2 => n999, A
                           => n112, ZN => O_51_port);
   U78 : AND2_X1 port map( A1 => n158, A2 => n960, ZN => n949);
   U79 : AND2_X1 port map( A1 => n158, A2 => n1066, ZN => n950);
   U80 : INV_X1 port map( A => n111, ZN => n1065);
   U81 : INV_X1 port map( A => n951, ZN => n959);
   U82 : OAI221_X1 port map( B1 => n962, B2 => n1000, C1 => n960, C2 => n1001, 
                           A => n149, ZN => O_18_port);
   U83 : AOI22_X1 port map( A1 => A_s(16), A2 => n954, B1 => A_ns(16), B2 => 
                           n958, ZN => n149);
   U84 : OR3_X1 port map( A1 => B(17), A2 => B(18), A3 => n1066, ZN => n951);
   U85 : INV_X1 port map( A => B(19), ZN => n1066);
   U86 : OAI221_X1 port map( B1 => n962, B2 => n1060, C1 => n960, C2 => n1062, 
                           A => n151, ZN => O_16_port);
   U87 : INV_X1 port map( A => A_ns(15), ZN => n1060);
   U88 : OAI221_X1 port map( B1 => n962, B2 => n1063, C1 => n960, C2 => n1064, 
                           A => n150, ZN => O_17_port);
   U89 : INV_X1 port map( A => A_ns(16), ZN => n1063);
   U90 : OAI221_X1 port map( B1 => n962, B2 => n1059, C1 => n960, C2 => n1061, 
                           A => n152, ZN => O_15_port);
   U91 : INV_X1 port map( A => A_ns(14), ZN => n1059);
   U92 : INV_X1 port map( A => A_s(14), ZN => n1061);
   U93 : OAI221_X1 port map( B1 => n963, B2 => n1045, C1 => n960, C2 => n1047, 
                           A => n108, ZN => O_7_port);
   U94 : INV_X1 port map( A => A_ns(6), ZN => n1045);
   U95 : INV_X1 port map( A => A_s(6), ZN => n1047);
   U96 : OAI221_X1 port map( B1 => n963, B2 => n1046, C1 => n960, C2 => n1048, 
                           A => n107, ZN => O_8_port);
   U97 : INV_X1 port map( A => A_ns(7), ZN => n1046);
   U98 : INV_X1 port map( A => A_s(7), ZN => n1048);
   U99 : OAI221_X1 port map( B1 => n963, B2 => n1049, C1 => n960, C2 => n1050, 
                           A => n105, ZN => O_9_port);
   U100 : AOI22_X1 port map( A1 => A_s(7), A2 => n957, B1 => A_ns(7), B2 => 
                           n959, ZN => n105);
   U101 : OAI221_X1 port map( B1 => n1050, B2 => n111, C1 => n1049, C2 => n951,
                           A => n157, ZN => O_10_port);
   U102 : AOI22_X1 port map( A1 => A_ns(9), A2 => n949, B1 => A_s(9), B2 => 
                           n950, ZN => n157);
   U103 : OAI221_X1 port map( B1 => n962, B2 => n1051, C1 => n960, C2 => n1053,
                           A => n156, ZN => O_11_port);
   U104 : INV_X1 port map( A => A_ns(10), ZN => n1051);
   U105 : INV_X1 port map( A => A_s(10), ZN => n1053);
   U106 : OAI221_X1 port map( B1 => n962, B2 => n1052, C1 => n960, C2 => n1054,
                           A => n155, ZN => O_12_port);
   U107 : INV_X1 port map( A => A_ns(11), ZN => n1052);
   U108 : INV_X1 port map( A => A_s(11), ZN => n1054);
   U109 : OAI221_X1 port map( B1 => n962, B2 => n1055, C1 => n960, C2 => n1057,
                           A => n154, ZN => O_13_port);
   U110 : INV_X1 port map( A => A_ns(12), ZN => n1055);
   U111 : INV_X1 port map( A => A_s(12), ZN => n1057);
   U112 : OAI221_X1 port map( B1 => n962, B2 => n1056, C1 => n960, C2 => n1058,
                           A => n153, ZN => O_14_port);
   U113 : INV_X1 port map( A => A_ns(13), ZN => n1056);
   U114 : INV_X1 port map( A => A_s(13), ZN => n1058);
   U115 : INV_X1 port map( A => n147, ZN => O_1_port);
   U116 : AOI22_X1 port map( A1 => n950, A2 => A_s(0), B1 => n949, B2 => 
                           A_ns(0), ZN => n147);
   U117 : OAI221_X1 port map( B1 => n962, B2 => n1035, C1 => n961, C2 => n1036,
                           A => n136, ZN => O_2_port);
   U118 : INV_X1 port map( A => A_ns(1), ZN => n1035);
   U119 : INV_X1 port map( A => A_s(1), ZN => n1036);
   U120 : OAI221_X1 port map( B1 => n963, B2 => n1037, C1 => n960, C2 => n1039,
                           A => n125, ZN => O_3_port);
   U121 : INV_X1 port map( A => A_ns(2), ZN => n1037);
   U122 : INV_X1 port map( A => A_s(2), ZN => n1039);
   U123 : OAI221_X1 port map( B1 => n963, B2 => n1038, C1 => n960, C2 => n1040,
                           A => n114, ZN => O_4_port);
   U124 : INV_X1 port map( A => A_ns(3), ZN => n1038);
   U125 : INV_X1 port map( A => A_s(3), ZN => n1040);
   U126 : OAI221_X1 port map( B1 => n963, B2 => n1041, C1 => n960, C2 => n1043,
                           A => n110, ZN => O_5_port);
   U127 : INV_X1 port map( A => A_ns(4), ZN => n1041);
   U128 : INV_X1 port map( A => A_s(4), ZN => n1043);
   U129 : OAI221_X1 port map( B1 => n963, B2 => n1042, C1 => n960, C2 => n1044,
                           A => n109, ZN => O_6_port);
   U130 : INV_X1 port map( A => A_ns(5), ZN => n1042);
   U131 : INV_X1 port map( A => A_s(5), ZN => n1044);
   U132 : INV_X1 port map( A => A_s(8), ZN => n1050);
   U133 : INV_X1 port map( A => A_ns(8), ZN => n1049);
   U134 : AOI22_X1 port map( A1 => A_s(15), A2 => n954, B1 => A_ns(15), B2 => 
                           n958, ZN => n150);
   U135 : AOI22_X1 port map( A1 => A_s(0), A2 => n955, B1 => A_ns(0), B2 => 
                           n958, ZN => n136);
   U136 : AOI22_X1 port map( A1 => A_s(1), A2 => n956, B1 => A_ns(1), B2 => 
                           n959, ZN => n125);
   U137 : AOI22_X1 port map( A1 => A_s(2), A2 => n957, B1 => A_ns(2), B2 => 
                           n959, ZN => n114);
   U138 : AOI22_X1 port map( A1 => A_s(3), A2 => n957, B1 => A_ns(3), B2 => 
                           n959, ZN => n110);
   U139 : AOI22_X1 port map( A1 => A_s(4), A2 => n957, B1 => A_ns(4), B2 => 
                           n959, ZN => n109);
   U140 : AOI22_X1 port map( A1 => A_s(5), A2 => n957, B1 => A_ns(5), B2 => 
                           n959, ZN => n108);
   U141 : AOI22_X1 port map( A1 => A_s(6), A2 => n957, B1 => A_ns(6), B2 => 
                           n959, ZN => n107);
   U142 : AOI22_X1 port map( A1 => A_s(9), A2 => n954, B1 => A_ns(9), B2 => 
                           n958, ZN => n156);
   U143 : AOI22_X1 port map( A1 => A_s(10), A2 => n954, B1 => A_ns(10), B2 => 
                           n958, ZN => n155);
   U144 : AOI22_X1 port map( A1 => A_s(11), A2 => n954, B1 => A_ns(11), B2 => 
                           n958, ZN => n154);
   U145 : AOI22_X1 port map( A1 => A_s(12), A2 => n954, B1 => A_ns(12), B2 => 
                           n958, ZN => n153);
   U146 : AOI22_X1 port map( A1 => A_s(13), A2 => n954, B1 => A_ns(13), B2 => 
                           n958, ZN => n152);
   U147 : AOI22_X1 port map( A1 => A_s(14), A2 => n954, B1 => A_ns(14), B2 => 
                           n958, ZN => n151);
   U148 : INV_X1 port map( A => A_s(16), ZN => n1064);
   U149 : INV_X1 port map( A => A_s(15), ZN => n1062);
   U150 : INV_X1 port map( A => n951, ZN => n958);
   U151 : INV_X1 port map( A => n950, ZN => n960);
   U152 : INV_X1 port map( A => n949, ZN => n962);
   U153 : INV_X1 port map( A => A_ns(18), ZN => n964);
   U154 : INV_X1 port map( A => A_ns(19), ZN => n965);
   U155 : INV_X1 port map( A => A_ns(20), ZN => n966);
   U156 : INV_X1 port map( A => A_ns(21), ZN => n967);
   U157 : INV_X1 port map( A => A_ns(22), ZN => n968);
   U158 : INV_X1 port map( A => A_ns(23), ZN => n969);
   U159 : INV_X1 port map( A => A_ns(24), ZN => n970);
   U160 : INV_X1 port map( A => A_ns(25), ZN => n971);
   U161 : INV_X1 port map( A => A_ns(26), ZN => n972);
   U162 : INV_X1 port map( A => A_ns(27), ZN => n973);
   U163 : INV_X1 port map( A => A_ns(28), ZN => n974);
   U164 : INV_X1 port map( A => A_ns(29), ZN => n975);
   U165 : INV_X1 port map( A => A_ns(30), ZN => n976);
   U166 : INV_X1 port map( A => A_ns(31), ZN => n977);
   U167 : INV_X1 port map( A => A_ns(32), ZN => n978);
   U168 : INV_X1 port map( A => A_ns(33), ZN => n979);
   U169 : INV_X1 port map( A => A_ns(34), ZN => n980);
   U170 : INV_X1 port map( A => A_ns(35), ZN => n981);
   U171 : INV_X1 port map( A => A_ns(36), ZN => n982);
   U172 : INV_X1 port map( A => A_ns(37), ZN => n983);
   U173 : INV_X1 port map( A => A_ns(38), ZN => n984);
   U174 : INV_X1 port map( A => n986, ZN => A_nso_41_port);
   U175 : INV_X1 port map( A => A_ns(39), ZN => n986);
   U176 : INV_X1 port map( A => A_ns(40), ZN => n987);
   U177 : INV_X1 port map( A => A_ns(41), ZN => n988);
   U178 : INV_X1 port map( A => A_ns(42), ZN => n989);
   U179 : INV_X1 port map( A => A_ns(43), ZN => n990);
   U180 : INV_X1 port map( A => A_ns(44), ZN => n991);
   U181 : INV_X1 port map( A => n993, ZN => A_nso_47_port);
   U182 : INV_X1 port map( A => A_ns(45), ZN => n993);
   U183 : INV_X1 port map( A => A_ns(46), ZN => n994);
   U184 : INV_X1 port map( A => A_ns(47), ZN => n995);
   U185 : INV_X1 port map( A => n997, ZN => A_nso_50_port);
   U186 : INV_X1 port map( A => A_ns(48), ZN => n997);
   U187 : INV_X1 port map( A => n999, ZN => A_nso_51_port);
   U188 : INV_X1 port map( A => A_ns(17), ZN => n1000);
   U189 : INV_X1 port map( A => A_s(17), ZN => n1001);
   U190 : INV_X1 port map( A => A_s(18), ZN => n1002);
   U191 : INV_X1 port map( A => A_s(19), ZN => n1003);
   U192 : INV_X1 port map( A => A_s(20), ZN => n1004);
   U193 : INV_X1 port map( A => A_s(21), ZN => n1005);
   U194 : INV_X1 port map( A => A_s(22), ZN => n1006);
   U195 : INV_X1 port map( A => A_s(23), ZN => n1007);
   U196 : INV_X1 port map( A => A_s(24), ZN => n1008);
   U197 : INV_X1 port map( A => A_s(25), ZN => n1009);
   U198 : INV_X1 port map( A => A_s(26), ZN => n1010);
   U199 : INV_X1 port map( A => A_s(27), ZN => n1011);
   U200 : INV_X1 port map( A => A_s(28), ZN => n1012);
   U201 : INV_X1 port map( A => A_s(29), ZN => n1013);
   U202 : INV_X1 port map( A => A_s(30), ZN => n1014);
   U203 : INV_X1 port map( A => A_s(31), ZN => n1015);
   U204 : INV_X1 port map( A => A_s(32), ZN => n1016);
   U205 : INV_X1 port map( A => A_s(33), ZN => n1017);
   U206 : INV_X1 port map( A => A_s(34), ZN => n1018);
   U207 : INV_X1 port map( A => A_s(35), ZN => n1019);
   U210 : INV_X1 port map( A => A_s(36), ZN => n1020);
   U211 : INV_X1 port map( A => A_s(37), ZN => n1021);
   U212 : INV_X1 port map( A => A_s(38), ZN => n1022);
   U213 : INV_X1 port map( A => A_s(39), ZN => n1023);
   U214 : INV_X1 port map( A => A_s(40), ZN => n1024);
   U215 : INV_X1 port map( A => A_s(41), ZN => n1025);
   U216 : INV_X1 port map( A => A_s(42), ZN => n1026);
   U217 : INV_X1 port map( A => A_s(43), ZN => n1027);
   U218 : INV_X1 port map( A => A_s(44), ZN => n1028);
   U219 : INV_X1 port map( A => A_s(45), ZN => n1029);
   U220 : INV_X1 port map( A => A_s(46), ZN => n1030);
   U221 : INV_X1 port map( A => A_s(47), ZN => n1031);
   U222 : INV_X1 port map( A => A_s(48), ZN => n1032);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT50_i16 is

   port( A_s, A_ns, B : in std_logic_vector (49 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (49 downto 0));

end BOOTHENC_NBIT50_i16;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT50_i16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, O_47_port, O_48_port, O_49_port, O_46_port, O_45_port,
      O_44_port, O_43_port, O_42_port, O_41_port, O_40_port, O_39_port, 
      O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, O_33_port, 
      O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, O_27_port, 
      O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, O_21_port, 
      O_20_port, O_19_port, O_18_port, O_17_port, O_2_port, O_3_port, O_4_port,
      O_5_port, O_6_port, O_7_port, O_8_port, O_9_port, O_10_port, O_11_port, 
      O_12_port, O_13_port, O_14_port, O_15_port, O_16_port, n101, n103, n104, 
      n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, 
      n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, 
      n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, 
      n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, 
      n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, 
      n970, n971, n972, A_nso_18_port, n974, A_nso_19_port, n976, A_nso_20_port
      , n978, A_nso_21_port, n980, A_nso_22_port, n982, A_nso_23_port, n984, 
      A_nso_24_port, n986, A_nso_25_port, n988, A_nso_26_port, n990, 
      A_nso_27_port, n992, A_nso_28_port, n994, A_nso_29_port, n996, 
      A_nso_30_port, n998, A_nso_31_port, n1000, A_nso_32_port, n1002, 
      A_nso_33_port, n1004, A_nso_34_port, n1006, A_nso_35_port, n1008, 
      A_nso_36_port, n1010, A_nso_37_port, n1012, A_nso_38_port, n1014, n1015, 
      A_nso_40_port, n1017, A_nso_41_port, n1019, A_nso_42_port, n1021, 
      A_nso_43_port, n1023, A_nso_44_port, n1025, n1026, A_nso_46_port, n1028, 
      A_nso_47_port, n1030, n1031, n1032, A_nso_17_port, n1034, A_so_17_port, 
      n1036, A_so_18_port, n1038, A_so_19_port, n1040, A_so_20_port, n1042, 
      A_so_21_port, n1044, A_so_22_port, n1046, A_so_23_port, n1048, 
      A_so_24_port, n1050, A_so_25_port, n1052, n1053, A_so_27_port, n1055, 
      n1056, A_so_29_port, n1058, n1059, n1060, A_so_32_port, n1062, 
      A_so_33_port, n1064, n1065, n1066, n1067, n1068, n1069, n1070, 
      A_so_40_port, n1072, n1073, n1074, n1075, n1076, A_so_45_port, n1078, 
      n1079, n1080, n1081, n1082, O_1_port, n1084, n1085, n1086, n1087, n1088, 
      n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, 
      n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, 
      n1109, n1110, n1111 : std_logic;

begin
   O <= ( O_49_port, O_48_port, O_47_port, O_46_port, O_45_port, O_44_port, 
      O_43_port, O_42_port, O_41_port, O_40_port, O_39_port, O_38_port, 
      O_37_port, O_36_port, O_35_port, O_34_port, O_33_port, O_32_port, 
      O_31_port, O_30_port, O_29_port, O_28_port, O_27_port, O_26_port, 
      O_25_port, O_24_port, O_23_port, O_22_port, O_21_port, O_20_port, 
      O_19_port, O_18_port, O_17_port, O_16_port, O_15_port, O_14_port, 
      O_13_port, O_12_port, O_11_port, O_10_port, O_9_port, O_8_port, O_7_port,
      O_6_port, O_5_port, O_4_port, O_3_port, O_2_port, O_1_port, X_Logic0_port
      );
   A_so <= ( A_s(47), A_s(46), A_s(45), A_s(44), A_so_45_port, A_s(42), A_s(41)
      , A_s(40), A_s(39), A_so_40_port, A_s(37), A_s(36), A_s(35), A_s(34), 
      A_s(33), A_s(32), A_so_33_port, A_so_32_port, A_s(29), A_s(28), 
      A_so_29_port, A_s(26), A_so_27_port, A_s(24), A_so_25_port, A_so_24_port,
      A_so_23_port, A_so_22_port, A_so_21_port, A_so_20_port, A_so_19_port, 
      A_so_18_port, A_so_17_port, A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), 
      A_s(9), A_s(8), A_s(7), A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), 
      A_s(0), X_Logic0_port, X_Logic0_port );
   A_nso <= ( A_ns(47), A_ns(46), A_nso_47_port, A_nso_46_port, A_ns(43), 
      A_nso_44_port, A_nso_43_port, A_nso_42_port, A_nso_41_port, A_nso_40_port
      , A_ns(37), A_nso_38_port, A_nso_37_port, A_nso_36_port, A_nso_35_port, 
      A_nso_34_port, A_nso_33_port, A_nso_32_port, A_nso_31_port, A_nso_30_port
      , A_nso_29_port, A_nso_28_port, A_nso_27_port, A_nso_26_port, 
      A_nso_25_port, A_nso_24_port, A_nso_23_port, A_nso_22_port, A_nso_21_port
      , A_nso_20_port, A_nso_19_port, A_nso_18_port, A_nso_17_port, A_ns(14), 
      A_ns(13), A_ns(12), A_ns(11), A_ns(10), A_ns(9), A_ns(8), A_ns(7), 
      A_ns(6), A_ns(5), A_ns(4), A_ns(3), A_ns(2), A_ns(1), A_ns(0), 
      X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U200 : XOR2_X1 port map( A => B(15), B => B(16), Z => n152);
   U201 : NAND3_X1 port map( A1 => B(16), A2 => n1111, A3 => B(15), ZN => n108)
                           ;
   U2 : OAI221_X1 port map( B1 => n972, B2 => n1028, C1 => n970, C2 => n1079, A
                           => n113, ZN => O_45_port);
   U3 : OAI221_X1 port map( B1 => n971, B2 => n976, C1 => n969, C2 => n1040, A 
                           => n143, ZN => O_18_port);
   U4 : OAI221_X1 port map( B1 => n971, B2 => n992, C1 => n970, C2 => n1055, A 
                           => n134, ZN => O_26_port);
   U5 : OAI221_X1 port map( B1 => n971, B2 => n1002, C1 => n970, C2 => n1062, A
                           => n128, ZN => O_31_port);
   U6 : CLKBUF_X1 port map( A => n961, Z => n964);
   U7 : CLKBUF_X1 port map( A => n1110, Z => n962);
   U8 : AND2_X1 port map( A1 => n152, A2 => n1111, ZN => n959);
   U9 : INV_X1 port map( A => A_ns(47), ZN => n1032);
   U10 : BUF_X1 port map( A => n961, Z => n963);
   U11 : BUF_X1 port map( A => n962, Z => n965);
   U12 : BUF_X1 port map( A => n962, Z => n966);
   U13 : OAI221_X1 port map( B1 => n972, B2 => n1021, C1 => n970, C2 => n1074, 
                           A => n117, ZN => O_41_port);
   U14 : OAI221_X1 port map( B1 => n972, B2 => n1025, C1 => n970, C2 => n1076, 
                           A => n115, ZN => O_43_port);
   U15 : AOI22_X1 port map( A1 => A_s(41), A2 => n965, B1 => A_nso_43_port, B2 
                           => n968, ZN => n115);
   U16 : INV_X1 port map( A => n959, ZN => n970);
   U17 : OAI221_X1 port map( B1 => n972, B2 => n986, C1 => n970, C2 => n1050, A
                           => n137, ZN => O_23_port);
   U18 : AOI22_X1 port map( A1 => A_so_23_port, A2 => n964, B1 => A_nso_23_port
                           , B2 => n967, ZN => n137);
   U19 : OAI221_X1 port map( B1 => n971, B2 => n978, C1 => n969, C2 => n1042, A
                           => n142, ZN => O_19_port);
   U20 : AOI22_X1 port map( A1 => A_so_19_port, A2 => n963, B1 => A_nso_19_port
                           , B2 => n968, ZN => n142);
   U21 : AOI22_X1 port map( A1 => A_so_18_port, A2 => n963, B1 => A_nso_18_port
                           , B2 => n967, ZN => n143);
   U22 : AOI22_X1 port map( A1 => A_s(29), A2 => n964, B1 => A_nso_31_port, B2 
                           => n967, ZN => n128);
   U23 : OAI221_X1 port map( B1 => n971, B2 => n982, C1 => n969, C2 => n1046, A
                           => n139, ZN => O_21_port);
   U24 : AOI22_X1 port map( A1 => A_so_21_port, A2 => n963, B1 => A_nso_21_port
                           , B2 => n968, ZN => n139);
   U25 : OAI221_X1 port map( B1 => n971, B2 => n1006, C1 => n970, C2 => n1065, 
                           A => n126, ZN => O_33_port);
   U26 : AOI22_X1 port map( A1 => A_so_33_port, A2 => n964, B1 => A_nso_33_port
                           , B2 => n967, ZN => n126);
   U27 : OAI221_X1 port map( B1 => n971, B2 => n994, C1 => n970, C2 => n1056, A
                           => n133, ZN => O_27_port);
   U28 : AOI22_X1 port map( A1 => A_so_27_port, A2 => n964, B1 => A_nso_27_port
                           , B2 => n967, ZN => n133);
   U29 : OAI221_X1 port map( B1 => n972, B2 => n990, C1 => n970, C2 => n1053, A
                           => n135, ZN => O_25_port);
   U30 : AOI22_X1 port map( A1 => A_so_25_port, A2 => n964, B1 => A_nso_25_port
                           , B2 => n967, ZN => n135);
   U31 : OAI221_X1 port map( B1 => n972, B2 => n1010, C1 => n970, C2 => n1067, 
                           A => n124, ZN => O_35_port);
   U32 : AOI22_X1 port map( A1 => A_s(33), A2 => n965, B1 => A_nso_35_port, B2 
                           => n968, ZN => n124);
   U33 : OAI221_X1 port map( B1 => n972, B2 => n1014, C1 => n970, C2 => n1069, 
                           A => n122, ZN => O_37_port);
   U34 : AOI22_X1 port map( A1 => A_s(35), A2 => n965, B1 => A_nso_37_port, B2 
                           => n968, ZN => n122);
   U35 : OAI221_X1 port map( B1 => n971, B2 => n998, C1 => n970, C2 => n1059, A
                           => n131, ZN => O_29_port);
   U36 : AOI22_X1 port map( A1 => A_so_29_port, A2 => n964, B1 => A_nso_29_port
                           , B2 => n967, ZN => n131);
   U37 : BUF_X1 port map( A => n1110, Z => n961);
   U38 : AOI22_X1 port map( A1 => A_so_45_port, A2 => n966, B1 => A_ns(43), B2 
                           => n968, ZN => n113);
   U39 : OAI221_X1 port map( B1 => n972, B2 => n1032, C1 => n969, C2 => n1082, 
                           A => n110, ZN => O_48_port);
   U40 : AOI22_X1 port map( A1 => A_s(46), A2 => n966, B1 => A_ns(46), B2 => 
                           n968, ZN => n110);
   U41 : OAI221_X1 port map( B1 => n972, B2 => n1031, C1 => n970, C2 => n1081, 
                           A => n111, ZN => O_47_port);
   U42 : AOI22_X1 port map( A1 => A_s(45), A2 => n966, B1 => A_nso_47_port, B2 
                           => n968, ZN => n111);
   U43 : OAI221_X1 port map( B1 => n972, B2 => n1017, C1 => n970, C2 => n1072, 
                           A => n120, ZN => O_39_port);
   U44 : AOI22_X1 port map( A1 => A_s(37), A2 => n965, B1 => A_ns(37), B2 => 
                           n968, ZN => n120);
   U45 : AOI22_X1 port map( A1 => A_s(39), A2 => n965, B1 => A_nso_41_port, B2 
                           => n968, ZN => n117);
   U46 : INV_X1 port map( A => n958, ZN => n972);
   U47 : OAI221_X1 port map( B1 => n108, B2 => n1082, C1 => n960, C2 => n1032, 
                           A => n109, ZN => O_49_port);
   U48 : OAI221_X1 port map( B1 => n972, B2 => n1026, C1 => n970, C2 => n1078, 
                           A => n114, ZN => O_44_port);
   U49 : AOI22_X1 port map( A1 => A_s(42), A2 => n965, B1 => A_nso_44_port, B2 
                           => n968, ZN => n114);
   U50 : OAI221_X1 port map( B1 => n972, B2 => n1023, C1 => n970, C2 => n1075, 
                           A => n116, ZN => O_42_port);
   U51 : AOI22_X1 port map( A1 => A_s(40), A2 => n965, B1 => A_nso_42_port, B2 
                           => n968, ZN => n116);
   U52 : OAI221_X1 port map( B1 => n971, B2 => n984, C1 => n969, C2 => n1048, A
                           => n138, ZN => O_22_port);
   U53 : AOI22_X1 port map( A1 => A_so_22_port, A2 => n963, B1 => A_nso_22_port
                           , B2 => n968, ZN => n138);
   U54 : OAI221_X1 port map( B1 => n971, B2 => n974, C1 => n969, C2 => n1038, A
                           => n144, ZN => O_17_port);
   U55 : AOI22_X1 port map( A1 => A_so_17_port, A2 => n963, B1 => A_nso_17_port
                           , B2 => n967, ZN => n144);
   U56 : OAI221_X1 port map( B1 => n972, B2 => n988, C1 => n970, C2 => n1052, A
                           => n136, ZN => O_24_port);
   U57 : AOI22_X1 port map( A1 => A_so_24_port, A2 => n964, B1 => A_nso_24_port
                           , B2 => n967, ZN => n136);
   U58 : AOI22_X1 port map( A1 => A_s(24), A2 => n964, B1 => A_nso_26_port, B2 
                           => n967, ZN => n134);
   U59 : OAI221_X1 port map( B1 => n971, B2 => n996, C1 => n970, C2 => n1058, A
                           => n132, ZN => O_28_port);
   U60 : AOI22_X1 port map( A1 => A_s(26), A2 => n964, B1 => A_nso_28_port, B2 
                           => n967, ZN => n132);
   U61 : OAI221_X1 port map( B1 => n971, B2 => n1000, C1 => n970, C2 => n1060, 
                           A => n129, ZN => O_30_port);
   U62 : AOI22_X1 port map( A1 => A_s(28), A2 => n964, B1 => A_nso_30_port, B2 
                           => n967, ZN => n129);
   U63 : OAI221_X1 port map( B1 => n971, B2 => n980, C1 => n969, C2 => n1044, A
                           => n140, ZN => O_20_port);
   U64 : AOI22_X1 port map( A1 => A_so_20_port, A2 => n963, B1 => A_nso_20_port
                           , B2 => n968, ZN => n140);
   U65 : OAI221_X1 port map( B1 => n971, B2 => n1004, C1 => n970, C2 => n1064, 
                           A => n127, ZN => O_32_port);
   U66 : AOI22_X1 port map( A1 => A_so_32_port, A2 => n964, B1 => A_nso_32_port
                           , B2 => n967, ZN => n127);
   U67 : OAI221_X1 port map( B1 => n972, B2 => n1008, C1 => n970, C2 => n1066, 
                           A => n125, ZN => O_34_port);
   U68 : AOI22_X1 port map( A1 => A_s(32), A2 => n965, B1 => A_nso_34_port, B2 
                           => n968, ZN => n125);
   U69 : OAI221_X1 port map( B1 => n972, B2 => n1012, C1 => n970, C2 => n1068, 
                           A => n123, ZN => O_36_port);
   U70 : AOI22_X1 port map( A1 => A_s(34), A2 => n965, B1 => A_nso_36_port, B2 
                           => n968, ZN => n123);
   U71 : INV_X1 port map( A => n960, ZN => n967);
   U72 : AND2_X1 port map( A1 => n152, A2 => n969, ZN => n958);
   U73 : INV_X1 port map( A => n108, ZN => n1110);
   U74 : OAI221_X1 port map( B1 => n972, B2 => n1015, C1 => n970, C2 => n1070, 
                           A => n121, ZN => O_38_port);
   U75 : AOI22_X1 port map( A1 => A_s(36), A2 => n965, B1 => A_nso_38_port, B2 
                           => n968, ZN => n121);
   U76 : OAI221_X1 port map( B1 => n972, B2 => n1019, C1 => n970, C2 => n1073, 
                           A => n118, ZN => O_40_port);
   U77 : AOI22_X1 port map( A1 => A_so_40_port, A2 => n965, B1 => A_nso_40_port
                           , B2 => n968, ZN => n118);
   U78 : OAI221_X1 port map( B1 => n972, B2 => n1030, C1 => n970, C2 => n1080, 
                           A => n112, ZN => O_46_port);
   U79 : AOI22_X1 port map( A1 => A_s(44), A2 => n966, B1 => A_nso_46_port, B2 
                           => n968, ZN => n112);
   U80 : INV_X1 port map( A => n960, ZN => n968);
   U81 : AOI22_X1 port map( A1 => A_ns(48), A2 => n958, B1 => A_s(48), B2 => 
                           n959, ZN => n109);
   U82 : INV_X1 port map( A => A_s(47), ZN => n1082);
   U83 : OAI221_X1 port map( B1 => n971, B2 => n1034, C1 => n969, C2 => n1036, 
                           A => n145, ZN => O_16_port);
   U84 : AOI22_X1 port map( A1 => A_s(14), A2 => n963, B1 => A_ns(14), B2 => 
                           n968, ZN => n145);
   U85 : OR3_X1 port map( A1 => B(15), A2 => B(16), A3 => n1111, ZN => n960);
   U86 : INV_X1 port map( A => B(17), ZN => n1111);
   U87 : OAI221_X1 port map( B1 => n971, B2 => n1108, C1 => n969, C2 => n1109, 
                           A => n146, ZN => O_15_port);
   U88 : INV_X1 port map( A => A_ns(14), ZN => n1108);
   U89 : OAI221_X1 port map( B1 => n972, B2 => n1094, C1 => n969, C2 => n1096, 
                           A => n104, ZN => O_7_port);
   U90 : INV_X1 port map( A => A_ns(6), ZN => n1094);
   U91 : INV_X1 port map( A => A_s(6), ZN => n1096);
   U92 : OAI221_X1 port map( B1 => n972, B2 => n1095, C1 => n969, C2 => n1097, 
                           A => n103, ZN => O_8_port);
   U93 : INV_X1 port map( A => A_ns(7), ZN => n1095);
   U94 : INV_X1 port map( A => A_s(7), ZN => n1097);
   U95 : OAI221_X1 port map( B1 => n972, B2 => n1098, C1 => n969, C2 => n1099, 
                           A => n101, ZN => O_9_port);
   U96 : AOI22_X1 port map( A1 => A_s(7), A2 => n966, B1 => A_ns(7), B2 => n967
                           , ZN => n101);
   U97 : OAI221_X1 port map( B1 => n1099, B2 => n108, C1 => n1098, C2 => n960, 
                           A => n151, ZN => O_10_port);
   U98 : AOI22_X1 port map( A1 => A_ns(9), A2 => n958, B1 => A_s(9), B2 => n959
                           , ZN => n151);
   U99 : OAI221_X1 port map( B1 => n971, B2 => n1100, C1 => n969, C2 => n1102, 
                           A => n150, ZN => O_11_port);
   U100 : INV_X1 port map( A => A_ns(10), ZN => n1100);
   U101 : INV_X1 port map( A => A_s(10), ZN => n1102);
   U102 : OAI221_X1 port map( B1 => n971, B2 => n1101, C1 => n969, C2 => n1103,
                           A => n149, ZN => O_12_port);
   U103 : INV_X1 port map( A => A_ns(11), ZN => n1101);
   U104 : INV_X1 port map( A => A_s(11), ZN => n1103);
   U105 : OAI221_X1 port map( B1 => n971, B2 => n1104, C1 => n969, C2 => n1106,
                           A => n148, ZN => O_13_port);
   U106 : INV_X1 port map( A => A_ns(12), ZN => n1104);
   U107 : INV_X1 port map( A => A_s(12), ZN => n1106);
   U108 : OAI221_X1 port map( B1 => n971, B2 => n1105, C1 => n969, C2 => n1107,
                           A => n147, ZN => O_14_port);
   U109 : INV_X1 port map( A => A_ns(13), ZN => n1105);
   U110 : INV_X1 port map( A => n141, ZN => O_1_port);
   U111 : AOI22_X1 port map( A1 => n959, A2 => A_s(0), B1 => n958, B2 => 
                           A_ns(0), ZN => n141);
   U112 : OAI221_X1 port map( B1 => n971, B2 => n1084, C1 => n970, C2 => n1085,
                           A => n130, ZN => O_2_port);
   U113 : INV_X1 port map( A => A_ns(1), ZN => n1084);
   U114 : INV_X1 port map( A => A_s(1), ZN => n1085);
   U115 : OAI221_X1 port map( B1 => n972, B2 => n1086, C1 => n969, C2 => n1088,
                           A => n119, ZN => O_3_port);
   U116 : INV_X1 port map( A => A_ns(2), ZN => n1086);
   U117 : INV_X1 port map( A => A_s(2), ZN => n1088);
   U118 : OAI221_X1 port map( B1 => n972, B2 => n1087, C1 => n969, C2 => n1089,
                           A => n107, ZN => O_4_port);
   U119 : INV_X1 port map( A => A_ns(3), ZN => n1087);
   U120 : INV_X1 port map( A => A_s(3), ZN => n1089);
   U121 : OAI221_X1 port map( B1 => n972, B2 => n1090, C1 => n969, C2 => n1092,
                           A => n106, ZN => O_5_port);
   U122 : INV_X1 port map( A => A_ns(4), ZN => n1090);
   U123 : INV_X1 port map( A => A_s(4), ZN => n1092);
   U124 : OAI221_X1 port map( B1 => n972, B2 => n1091, C1 => n969, C2 => n1093,
                           A => n105, ZN => O_6_port);
   U125 : INV_X1 port map( A => A_ns(5), ZN => n1091);
   U126 : INV_X1 port map( A => A_s(5), ZN => n1093);
   U127 : INV_X1 port map( A => A_s(8), ZN => n1099);
   U128 : INV_X1 port map( A => A_ns(8), ZN => n1098);
   U129 : AOI22_X1 port map( A1 => A_s(0), A2 => n964, B1 => A_ns(0), B2 => 
                           n967, ZN => n130);
   U130 : AOI22_X1 port map( A1 => A_s(1), A2 => n965, B1 => A_ns(1), B2 => 
                           n968, ZN => n119);
   U131 : AOI22_X1 port map( A1 => A_s(2), A2 => n966, B1 => A_ns(2), B2 => 
                           n967, ZN => n107);
   U132 : AOI22_X1 port map( A1 => A_s(3), A2 => n966, B1 => A_ns(3), B2 => 
                           n967, ZN => n106);
   U133 : AOI22_X1 port map( A1 => A_s(4), A2 => n966, B1 => A_ns(4), B2 => 
                           n967, ZN => n105);
   U134 : AOI22_X1 port map( A1 => A_s(5), A2 => n966, B1 => A_ns(5), B2 => 
                           n967, ZN => n104);
   U135 : AOI22_X1 port map( A1 => A_s(6), A2 => n966, B1 => A_ns(6), B2 => 
                           n967, ZN => n103);
   U136 : AOI22_X1 port map( A1 => A_s(9), A2 => n963, B1 => A_ns(9), B2 => 
                           n968, ZN => n150);
   U137 : AOI22_X1 port map( A1 => A_s(10), A2 => n963, B1 => A_ns(10), B2 => 
                           n968, ZN => n149);
   U138 : AOI22_X1 port map( A1 => A_s(11), A2 => n963, B1 => A_ns(11), B2 => 
                           n968, ZN => n148);
   U139 : AOI22_X1 port map( A1 => A_s(12), A2 => n963, B1 => A_ns(12), B2 => 
                           n968, ZN => n147);
   U140 : AOI22_X1 port map( A1 => A_s(13), A2 => n963, B1 => A_ns(13), B2 => 
                           n968, ZN => n146);
   U141 : INV_X1 port map( A => A_s(13), ZN => n1107);
   U142 : INV_X1 port map( A => A_s(14), ZN => n1109);
   U143 : INV_X1 port map( A => n959, ZN => n969);
   U144 : INV_X1 port map( A => n958, ZN => n971);
   U145 : INV_X1 port map( A => n974, ZN => A_nso_18_port);
   U146 : INV_X1 port map( A => A_ns(16), ZN => n974);
   U147 : INV_X1 port map( A => n976, ZN => A_nso_19_port);
   U148 : INV_X1 port map( A => A_ns(17), ZN => n976);
   U149 : INV_X1 port map( A => n978, ZN => A_nso_20_port);
   U150 : INV_X1 port map( A => A_ns(18), ZN => n978);
   U151 : INV_X1 port map( A => n980, ZN => A_nso_21_port);
   U152 : INV_X1 port map( A => A_ns(19), ZN => n980);
   U153 : INV_X1 port map( A => n982, ZN => A_nso_22_port);
   U154 : INV_X1 port map( A => A_ns(20), ZN => n982);
   U155 : INV_X1 port map( A => n984, ZN => A_nso_23_port);
   U156 : INV_X1 port map( A => A_ns(21), ZN => n984);
   U157 : INV_X1 port map( A => n986, ZN => A_nso_24_port);
   U158 : INV_X1 port map( A => A_ns(22), ZN => n986);
   U159 : INV_X1 port map( A => n988, ZN => A_nso_25_port);
   U160 : INV_X1 port map( A => A_ns(23), ZN => n988);
   U161 : INV_X1 port map( A => n990, ZN => A_nso_26_port);
   U162 : INV_X1 port map( A => A_ns(24), ZN => n990);
   U163 : INV_X1 port map( A => n992, ZN => A_nso_27_port);
   U164 : INV_X1 port map( A => A_ns(25), ZN => n992);
   U165 : INV_X1 port map( A => n994, ZN => A_nso_28_port);
   U166 : INV_X1 port map( A => A_ns(26), ZN => n994);
   U167 : INV_X1 port map( A => n996, ZN => A_nso_29_port);
   U168 : INV_X1 port map( A => A_ns(27), ZN => n996);
   U169 : INV_X1 port map( A => n998, ZN => A_nso_30_port);
   U170 : INV_X1 port map( A => A_ns(28), ZN => n998);
   U171 : INV_X1 port map( A => n1000, ZN => A_nso_31_port);
   U172 : INV_X1 port map( A => A_ns(29), ZN => n1000);
   U173 : INV_X1 port map( A => n1002, ZN => A_nso_32_port);
   U174 : INV_X1 port map( A => A_ns(30), ZN => n1002);
   U175 : INV_X1 port map( A => n1004, ZN => A_nso_33_port);
   U176 : INV_X1 port map( A => A_ns(31), ZN => n1004);
   U177 : INV_X1 port map( A => n1006, ZN => A_nso_34_port);
   U178 : INV_X1 port map( A => A_ns(32), ZN => n1006);
   U179 : INV_X1 port map( A => n1008, ZN => A_nso_35_port);
   U180 : INV_X1 port map( A => A_ns(33), ZN => n1008);
   U181 : INV_X1 port map( A => n1010, ZN => A_nso_36_port);
   U182 : INV_X1 port map( A => A_ns(34), ZN => n1010);
   U183 : INV_X1 port map( A => n1012, ZN => A_nso_37_port);
   U184 : INV_X1 port map( A => A_ns(35), ZN => n1012);
   U185 : INV_X1 port map( A => n1014, ZN => A_nso_38_port);
   U186 : INV_X1 port map( A => A_ns(36), ZN => n1014);
   U187 : INV_X1 port map( A => A_ns(37), ZN => n1015);
   U188 : INV_X1 port map( A => n1017, ZN => A_nso_40_port);
   U189 : INV_X1 port map( A => A_ns(38), ZN => n1017);
   U190 : INV_X1 port map( A => n1019, ZN => A_nso_41_port);
   U191 : INV_X1 port map( A => A_ns(39), ZN => n1019);
   U192 : INV_X1 port map( A => n1021, ZN => A_nso_42_port);
   U193 : INV_X1 port map( A => A_ns(40), ZN => n1021);
   U194 : INV_X1 port map( A => n1023, ZN => A_nso_43_port);
   U195 : INV_X1 port map( A => A_ns(41), ZN => n1023);
   U196 : INV_X1 port map( A => n1025, ZN => A_nso_44_port);
   U197 : INV_X1 port map( A => A_ns(42), ZN => n1025);
   U198 : INV_X1 port map( A => A_ns(43), ZN => n1026);
   U199 : INV_X1 port map( A => n1028, ZN => A_nso_46_port);
   U202 : INV_X1 port map( A => A_ns(44), ZN => n1028);
   U203 : INV_X1 port map( A => n1030, ZN => A_nso_47_port);
   U204 : INV_X1 port map( A => A_ns(45), ZN => n1030);
   U205 : INV_X1 port map( A => A_ns(46), ZN => n1031);
   U206 : INV_X1 port map( A => n1034, ZN => A_nso_17_port);
   U207 : INV_X1 port map( A => A_ns(15), ZN => n1034);
   U208 : INV_X1 port map( A => n1036, ZN => A_so_17_port);
   U209 : INV_X1 port map( A => A_s(15), ZN => n1036);
   U210 : INV_X1 port map( A => n1038, ZN => A_so_18_port);
   U211 : INV_X1 port map( A => A_s(16), ZN => n1038);
   U212 : INV_X1 port map( A => n1040, ZN => A_so_19_port);
   U213 : INV_X1 port map( A => A_s(17), ZN => n1040);
   U214 : INV_X1 port map( A => n1042, ZN => A_so_20_port);
   U215 : INV_X1 port map( A => A_s(18), ZN => n1042);
   U216 : INV_X1 port map( A => n1044, ZN => A_so_21_port);
   U217 : INV_X1 port map( A => A_s(19), ZN => n1044);
   U218 : INV_X1 port map( A => n1046, ZN => A_so_22_port);
   U219 : INV_X1 port map( A => A_s(20), ZN => n1046);
   U220 : INV_X1 port map( A => n1048, ZN => A_so_23_port);
   U221 : INV_X1 port map( A => A_s(21), ZN => n1048);
   U222 : INV_X1 port map( A => n1050, ZN => A_so_24_port);
   U223 : INV_X1 port map( A => A_s(22), ZN => n1050);
   U224 : INV_X1 port map( A => n1052, ZN => A_so_25_port);
   U225 : INV_X1 port map( A => A_s(23), ZN => n1052);
   U226 : INV_X1 port map( A => A_s(24), ZN => n1053);
   U227 : INV_X1 port map( A => n1055, ZN => A_so_27_port);
   U228 : INV_X1 port map( A => A_s(25), ZN => n1055);
   U229 : INV_X1 port map( A => A_s(26), ZN => n1056);
   U230 : INV_X1 port map( A => n1058, ZN => A_so_29_port);
   U231 : INV_X1 port map( A => A_s(27), ZN => n1058);
   U232 : INV_X1 port map( A => A_s(28), ZN => n1059);
   U233 : INV_X1 port map( A => A_s(29), ZN => n1060);
   U234 : INV_X1 port map( A => n1062, ZN => A_so_32_port);
   U235 : INV_X1 port map( A => A_s(30), ZN => n1062);
   U236 : INV_X1 port map( A => n1064, ZN => A_so_33_port);
   U237 : INV_X1 port map( A => A_s(31), ZN => n1064);
   U238 : INV_X1 port map( A => A_s(32), ZN => n1065);
   U239 : INV_X1 port map( A => A_s(33), ZN => n1066);
   U240 : INV_X1 port map( A => A_s(34), ZN => n1067);
   U241 : INV_X1 port map( A => A_s(35), ZN => n1068);
   U242 : INV_X1 port map( A => A_s(36), ZN => n1069);
   U243 : INV_X1 port map( A => A_s(37), ZN => n1070);
   U244 : INV_X1 port map( A => n1072, ZN => A_so_40_port);
   U245 : INV_X1 port map( A => A_s(38), ZN => n1072);
   U246 : INV_X1 port map( A => A_s(39), ZN => n1073);
   U247 : INV_X1 port map( A => A_s(40), ZN => n1074);
   U248 : INV_X1 port map( A => A_s(41), ZN => n1075);
   U249 : INV_X1 port map( A => A_s(42), ZN => n1076);
   U250 : INV_X1 port map( A => n1078, ZN => A_so_45_port);
   U251 : INV_X1 port map( A => A_s(43), ZN => n1078);
   U252 : INV_X1 port map( A => A_s(44), ZN => n1079);
   U253 : INV_X1 port map( A => A_s(45), ZN => n1080);
   U254 : INV_X1 port map( A => A_s(46), ZN => n1081);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT48_i14 is

   port( A_s, A_ns, B : in std_logic_vector (47 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (47 downto 0));

end BOOTHENC_NBIT48_i14;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT48_i14 is

   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105
      , n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
      n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, 
      n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, 
      n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
      n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, 
      n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, 
      n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, 
      n190, n191, n192, n193, n999, n1000, n1001, n1002, n1003, n1004, n1005, 
      n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, 
      n1016, n1017, n1018, n1019, n1020, n1021, n1022, O_2_port, n1024, 
      O_1_port, O_3_port, n1027, O_4_port, n1029, O_5_port, n1031, O_6_port, 
      n1033, O_7_port, n1035, O_8_port, n1037, O_9_port, n1039, O_10_port, 
      n1041, O_11_port, n1043, O_12_port, n1045, O_13_port, n1047, O_14_port, 
      n1049, O_45_port, O_46_port, n1052, O_47_port, n1054, O_44_port, n1056, 
      O_43_port, n1058, O_42_port, n1060, O_41_port, n1062, O_40_port, n1064, 
      O_39_port, n1066, O_38_port, n1068, O_37_port, n1070, O_36_port, n1072, 
      O_35_port, n1074, O_34_port, n1076, O_33_port, n1078, O_32_port, n1080, 
      O_31_port, n1082, O_30_port, n1084, O_29_port, n1086, O_28_port, n1088, 
      O_27_port, n1090, O_26_port, n1092, O_25_port, n1094, O_24_port, n1096, 
      O_23_port, n1098, O_22_port, n1100, O_21_port, n1102, O_20_port, n1104, 
      O_19_port, n1106, O_18_port, n1108, O_17_port, n1110, O_16_port, n1112, 
      O_15_port, n1114, n1115, n1116, n1117 : std_logic;

begin
   O <= ( O_47_port, O_46_port, O_45_port, O_44_port, O_43_port, O_42_port, 
      O_41_port, O_40_port, O_39_port, O_38_port, O_37_port, O_36_port, 
      O_35_port, O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, 
      O_29_port, O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, 
      O_23_port, O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, 
      O_17_port, O_16_port, O_15_port, O_14_port, O_13_port, O_12_port, 
      O_11_port, O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, 
      O_4_port, O_3_port, O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), 
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   A_nso <= ( A_ns(45), A_ns(44), A_ns(43), A_ns(42), A_ns(41), A_ns(40), 
      A_ns(39), A_ns(38), A_ns(37), A_ns(36), A_ns(35), A_ns(34), A_ns(33), 
      A_ns(32), A_ns(31), A_ns(30), A_ns(29), A_ns(28), A_ns(27), A_ns(26), 
      A_ns(25), A_ns(24), A_ns(23), A_ns(22), A_ns(21), A_ns(20), A_ns(19), 
      A_ns(18), A_ns(17), A_ns(16), A_ns(15), A_ns(14), A_ns(13), A_ns(12), 
      A_ns(11), A_ns(10), A_ns(9), A_ns(8), A_ns(7), A_ns(6), A_ns(5), A_ns(4),
      A_ns(3), A_ns(2), A_ns(1), A_ns(0), X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U194 : XOR2_X1 port map( A => B(13), B => B(14), Z => n193);
   U2 : CLKBUF_X1 port map( A => n1116, Z => n999);
   U3 : CLKBUF_X1 port map( A => n97, Z => n1017);
   U4 : CLKBUF_X1 port map( A => n100, Z => n1005);
   U5 : CLKBUF_X1 port map( A => n99, Z => n1011);
   U6 : CLKBUF_X1 port map( A => n1000, Z => n1003);
   U7 : CLKBUF_X1 port map( A => n1018, Z => n1021);
   U8 : CLKBUF_X1 port map( A => n1012, Z => n1015);
   U9 : CLKBUF_X1 port map( A => n1006, Z => n1009);
   U10 : BUF_X1 port map( A => n1000, Z => n1004);
   U11 : BUF_X1 port map( A => n999, Z => n1002);
   U12 : BUF_X1 port map( A => n999, Z => n1001);
   U13 : BUF_X1 port map( A => n1018, Z => n1022);
   U14 : BUF_X1 port map( A => n1116, Z => n1000);
   U15 : BUF_X1 port map( A => n1017, Z => n1020);
   U16 : BUF_X1 port map( A => n1017, Z => n1019);
   U17 : INV_X1 port map( A => n118, ZN => O_47_port);
   U18 : BUF_X1 port map( A => n1012, Z => n1016);
   U19 : BUF_X1 port map( A => n1006, Z => n1010);
   U20 : INV_X1 port map( A => n180, ZN => O_17_port);
   U21 : AOI221_X1 port map( B1 => n1022, B2 => A_ns(16), C1 => n1004, C2 => 
                           A_s(16), A => n1112, ZN => n180);
   U22 : INV_X1 port map( A => n181, ZN => n1112);
   U23 : AOI22_X1 port map( A1 => A_s(15), A2 => n1016, B1 => A_ns(15), B2 => 
                           n1010, ZN => n181);
   U24 : BUF_X1 port map( A => n97, Z => n1018);
   U25 : INV_X1 port map( A => n192, ZN => n1116);
   U26 : BUF_X1 port map( A => n1011, Z => n1014);
   U27 : BUF_X1 port map( A => n1005, Z => n1008);
   U28 : BUF_X1 port map( A => n1011, Z => n1013);
   U29 : BUF_X1 port map( A => n1005, Z => n1007);
   U30 : NAND2_X1 port map( A1 => n193, A2 => n1117, ZN => n192);
   U31 : BUF_X1 port map( A => n100, Z => n1006);
   U32 : BUF_X1 port map( A => n99, Z => n1012);
   U33 : AND2_X1 port map( A1 => n193, A2 => n192, ZN => n97);
   U34 : AOI221_X1 port map( B1 => n1016, B2 => A_s(45), C1 => n1010, C2 => 
                           A_ns(45), A => n1054, ZN => n118);
   U35 : INV_X1 port map( A => n119, ZN => n1054);
   U36 : AOI22_X1 port map( A1 => A_ns(46), A2 => n1019, B1 => A_s(46), B2 => 
                           n1001, ZN => n119);
   U37 : INV_X1 port map( A => n120, ZN => O_46_port);
   U38 : AOI221_X1 port map( B1 => n1019, B2 => A_ns(45), C1 => n1001, C2 => 
                           A_s(45), A => n1052, ZN => n120);
   U39 : INV_X1 port map( A => n121, ZN => n1052);
   U40 : AOI22_X1 port map( A1 => A_s(44), A2 => n1013, B1 => A_ns(44), B2 => 
                           n1007, ZN => n121);
   U41 : INV_X1 port map( A => n172, ZN => O_21_port);
   U42 : AOI221_X1 port map( B1 => n1021, B2 => A_ns(20), C1 => n1004, C2 => 
                           A_s(20), A => n1104, ZN => n172);
   U43 : INV_X1 port map( A => n173, ZN => n1104);
   U44 : AOI22_X1 port map( A1 => A_s(19), A2 => n1016, B1 => A_ns(19), B2 => 
                           n1010, ZN => n173);
   U45 : INV_X1 port map( A => n174, ZN => O_20_port);
   U46 : AOI221_X1 port map( B1 => n1021, B2 => A_ns(19), C1 => n1004, C2 => 
                           A_s(19), A => n1106, ZN => n174);
   U47 : INV_X1 port map( A => n175, ZN => n1106);
   U48 : AOI22_X1 port map( A1 => A_s(18), A2 => n1016, B1 => A_ns(18), B2 => 
                           n1010, ZN => n175);
   U49 : NOR3_X1 port map( A1 => B(13), A2 => B(14), A3 => n1117, ZN => n100);
   U50 : INV_X1 port map( A => n186, ZN => O_14_port);
   U51 : INV_X1 port map( A => n187, ZN => n1049);
   U52 : AOI22_X1 port map( A1 => A_s(12), A2 => n1016, B1 => A_ns(12), B2 => 
                           n1010, ZN => n187);
   U53 : INV_X1 port map( A => n138, ZN => O_37_port);
   U54 : AOI221_X1 port map( B1 => n1020, B2 => A_ns(36), C1 => n1002, C2 => 
                           A_s(36), A => n1072, ZN => n138);
   U55 : INV_X1 port map( A => n139, ZN => n1072);
   U56 : AOI22_X1 port map( A1 => A_s(35), A2 => n1014, B1 => A_ns(35), B2 => 
                           n1008, ZN => n139);
   U57 : INV_X1 port map( A => n134, ZN => O_39_port);
   U58 : AOI221_X1 port map( B1 => n1020, B2 => A_ns(38), C1 => n1002, C2 => 
                           A_s(38), A => n1068, ZN => n134);
   U59 : INV_X1 port map( A => n135, ZN => n1068);
   U60 : AOI22_X1 port map( A1 => A_s(37), A2 => n1014, B1 => A_ns(37), B2 => 
                           n1008, ZN => n135);
   U61 : INV_X1 port map( A => n136, ZN => O_38_port);
   U62 : AOI221_X1 port map( B1 => n1020, B2 => A_ns(37), C1 => n1002, C2 => 
                           A_s(37), A => n1070, ZN => n136);
   U63 : INV_X1 port map( A => n137, ZN => n1070);
   U64 : AOI22_X1 port map( A1 => A_s(36), A2 => n1014, B1 => A_ns(36), B2 => 
                           n1008, ZN => n137);
   U65 : INV_X1 port map( A => n140, ZN => O_36_port);
   U66 : AOI221_X1 port map( B1 => n1020, B2 => A_ns(35), C1 => n1002, C2 => 
                           A_s(35), A => n1074, ZN => n140);
   U67 : INV_X1 port map( A => n141, ZN => n1074);
   U68 : AOI22_X1 port map( A1 => A_s(34), A2 => n1014, B1 => A_ns(34), B2 => 
                           n1008, ZN => n141);
   U69 : INV_X1 port map( A => B(15), ZN => n1117);
   U70 : INV_X1 port map( A => n176, ZN => O_19_port);
   U71 : AOI221_X1 port map( B1 => n1022, B2 => A_ns(18), C1 => n1004, C2 => 
                           A_s(18), A => n1108, ZN => n176);
   U72 : INV_X1 port map( A => n177, ZN => n1108);
   U73 : AOI22_X1 port map( A1 => A_s(17), A2 => n1016, B1 => A_ns(17), B2 => 
                           n1010, ZN => n177);
   U74 : INV_X1 port map( A => n160, ZN => O_27_port);
   U75 : AOI221_X1 port map( B1 => n1021, B2 => A_ns(26), C1 => n1003, C2 => 
                           A_s(26), A => n1092, ZN => n160);
   U76 : INV_X1 port map( A => n161, ZN => n1092);
   U77 : AOI22_X1 port map( A1 => A_s(25), A2 => n1015, B1 => A_ns(25), B2 => 
                           n1009, ZN => n161);
   U78 : INV_X1 port map( A => n164, ZN => O_25_port);
   U79 : AOI221_X1 port map( B1 => n1021, B2 => A_ns(24), C1 => n1003, C2 => 
                           A_s(24), A => n1096, ZN => n164);
   U80 : INV_X1 port map( A => n165, ZN => n1096);
   U81 : AOI22_X1 port map( A1 => A_s(23), A2 => n1015, B1 => A_ns(23), B2 => 
                           n1009, ZN => n165);
   U82 : INV_X1 port map( A => n156, ZN => O_29_port);
   U83 : AOI221_X1 port map( B1 => n1021, B2 => A_ns(28), C1 => n1003, C2 => 
                           A_s(28), A => n1088, ZN => n156);
   U84 : INV_X1 port map( A => n157, ZN => n1088);
   U85 : AOI22_X1 port map( A1 => A_s(27), A2 => n1015, B1 => A_ns(27), B2 => 
                           n1009, ZN => n157);
   U86 : INV_X1 port map( A => n146, ZN => O_33_port);
   U87 : AOI221_X1 port map( B1 => n1020, B2 => A_ns(32), C1 => n1003, C2 => 
                           A_s(32), A => n1080, ZN => n146);
   U88 : INV_X1 port map( A => n147, ZN => n1080);
   U89 : AOI22_X1 port map( A1 => A_s(31), A2 => n1014, B1 => A_ns(31), B2 => 
                           n1008, ZN => n147);
   U90 : INV_X1 port map( A => n142, ZN => O_35_port);
   U91 : AOI221_X1 port map( B1 => n1020, B2 => A_ns(34), C1 => n1002, C2 => 
                           A_s(34), A => n1076, ZN => n142);
   U92 : INV_X1 port map( A => n143, ZN => n1076);
   U93 : AOI22_X1 port map( A1 => A_s(33), A2 => n1014, B1 => A_ns(33), B2 => 
                           n1008, ZN => n143);
   U94 : INV_X1 port map( A => n168, ZN => O_23_port);
   U95 : AOI221_X1 port map( B1 => n1021, B2 => A_ns(22), C1 => n1003, C2 => 
                           A_s(22), A => n1100, ZN => n168);
   U96 : INV_X1 port map( A => n169, ZN => n1100);
   U97 : AOI22_X1 port map( A1 => A_s(21), A2 => n1015, B1 => A_ns(21), B2 => 
                           n1009, ZN => n169);
   U98 : INV_X1 port map( A => n150, ZN => O_31_port);
   U99 : AOI221_X1 port map( B1 => n1021, B2 => A_ns(30), C1 => n1003, C2 => 
                           A_s(30), A => n1084, ZN => n150);
   U100 : INV_X1 port map( A => n151, ZN => n1084);
   U101 : AOI22_X1 port map( A1 => A_s(29), A2 => n1015, B1 => A_ns(29), B2 => 
                           n1009, ZN => n151);
   U102 : INV_X1 port map( A => n182, ZN => O_16_port);
   U103 : AOI221_X1 port map( B1 => n1022, B2 => A_ns(15), C1 => n1004, C2 => 
                           A_s(15), A => n1114, ZN => n182);
   U104 : INV_X1 port map( A => n183, ZN => n1114);
   U105 : AOI22_X1 port map( A1 => A_s(14), A2 => n1016, B1 => A_ns(14), B2 => 
                           n1010, ZN => n183);
   U106 : INV_X1 port map( A => n144, ZN => O_34_port);
   U107 : AOI221_X1 port map( B1 => n1020, B2 => A_ns(33), C1 => n1002, C2 => 
                           A_s(33), A => n1078, ZN => n144);
   U108 : INV_X1 port map( A => n145, ZN => n1078);
   U109 : AOI22_X1 port map( A1 => A_s(32), A2 => n1014, B1 => A_ns(32), B2 => 
                           n1008, ZN => n145);
   U110 : INV_X1 port map( A => n132, ZN => O_40_port);
   U111 : AOI221_X1 port map( B1 => n1020, B2 => A_ns(39), C1 => n1002, C2 => 
                           A_s(39), A => n1066, ZN => n132);
   U112 : INV_X1 port map( A => n133, ZN => n1066);
   U113 : AOI22_X1 port map( A1 => A_s(38), A2 => n1014, B1 => A_ns(38), B2 => 
                           n1008, ZN => n133);
   U114 : INV_X1 port map( A => n178, ZN => O_18_port);
   U115 : AOI221_X1 port map( B1 => n1022, B2 => A_ns(17), C1 => n1004, C2 => 
                           A_s(17), A => n1110, ZN => n178);
   U116 : INV_X1 port map( A => n179, ZN => n1110);
   U117 : AOI22_X1 port map( A1 => A_s(16), A2 => n1016, B1 => A_ns(16), B2 => 
                           n1010, ZN => n179);
   U118 : INV_X1 port map( A => n184, ZN => O_15_port);
   U119 : AOI221_X1 port map( B1 => n1022, B2 => A_ns(14), C1 => n1004, C2 => 
                           A_s(14), A => n1115, ZN => n184);
   U120 : INV_X1 port map( A => n185, ZN => n1115);
   U121 : INV_X1 port map( A => n158, ZN => O_28_port);
   U122 : AOI221_X1 port map( B1 => n1021, B2 => A_ns(27), C1 => n1003, C2 => 
                           A_s(27), A => n1090, ZN => n158);
   U123 : INV_X1 port map( A => n159, ZN => n1090);
   U124 : AOI22_X1 port map( A1 => A_s(26), A2 => n1015, B1 => A_ns(26), B2 => 
                           n1009, ZN => n159);
   U125 : INV_X1 port map( A => n170, ZN => O_22_port);
   U126 : AOI221_X1 port map( B1 => n1021, B2 => A_ns(21), C1 => n1003, C2 => 
                           A_s(21), A => n1102, ZN => n170);
   U127 : INV_X1 port map( A => n171, ZN => n1102);
   U128 : AOI22_X1 port map( A1 => A_s(20), A2 => n1015, B1 => A_ns(20), B2 => 
                           n1009, ZN => n171);
   U129 : INV_X1 port map( A => n166, ZN => O_24_port);
   U130 : AOI221_X1 port map( B1 => n1021, B2 => A_ns(23), C1 => n1003, C2 => 
                           A_s(23), A => n1098, ZN => n166);
   U131 : INV_X1 port map( A => n167, ZN => n1098);
   U132 : AOI22_X1 port map( A1 => A_s(22), A2 => n1015, B1 => A_ns(22), B2 => 
                           n1009, ZN => n167);
   U133 : INV_X1 port map( A => n162, ZN => O_26_port);
   U134 : AOI221_X1 port map( B1 => n1021, B2 => A_ns(25), C1 => n1003, C2 => 
                           A_s(25), A => n1094, ZN => n162);
   U135 : INV_X1 port map( A => n163, ZN => n1094);
   U136 : AOI22_X1 port map( A1 => A_s(24), A2 => n1015, B1 => A_ns(24), B2 => 
                           n1009, ZN => n163);
   U137 : INV_X1 port map( A => n152, ZN => O_30_port);
   U138 : AOI221_X1 port map( B1 => n1021, B2 => A_ns(29), C1 => n1003, C2 => 
                           A_s(29), A => n1086, ZN => n152);
   U139 : INV_X1 port map( A => n153, ZN => n1086);
   U140 : AOI22_X1 port map( A1 => A_s(28), A2 => n1015, B1 => A_ns(28), B2 => 
                           n1009, ZN => n153);
   U141 : INV_X1 port map( A => n148, ZN => O_32_port);
   U142 : AOI221_X1 port map( B1 => n1020, B2 => A_ns(31), C1 => n1003, C2 => 
                           A_s(31), A => n1082, ZN => n148);
   U143 : INV_X1 port map( A => n149, ZN => n1082);
   U144 : AOI22_X1 port map( A1 => A_s(30), A2 => n1015, B1 => A_ns(30), B2 => 
                           n1009, ZN => n149);
   U145 : AND3_X1 port map( A1 => B(13), A2 => n1117, A3 => B(14), ZN => n99);
   U146 : INV_X1 port map( A => n124, ZN => O_44_port);
   U147 : AOI221_X1 port map( B1 => n1019, B2 => A_ns(43), C1 => n1002, C2 => 
                           A_s(43), A => n1058, ZN => n124);
   U148 : INV_X1 port map( A => n125, ZN => n1058);
   U149 : AOI22_X1 port map( A1 => A_s(42), A2 => n1013, B1 => A_ns(42), B2 => 
                           n1007, ZN => n125);
   U150 : INV_X1 port map( A => n122, ZN => O_45_port);
   U151 : AOI221_X1 port map( B1 => n1019, B2 => A_ns(44), C1 => n1002, C2 => 
                           A_s(44), A => n1056, ZN => n122);
   U152 : INV_X1 port map( A => n123, ZN => n1056);
   U153 : AOI22_X1 port map( A1 => A_s(43), A2 => n1013, B1 => A_ns(43), B2 => 
                           n1007, ZN => n123);
   U154 : INV_X1 port map( A => n130, ZN => O_41_port);
   U155 : AOI221_X1 port map( B1 => n1020, B2 => A_ns(40), C1 => n1002, C2 => 
                           A_s(40), A => n1064, ZN => n130);
   U156 : INV_X1 port map( A => n131, ZN => n1064);
   U157 : AOI22_X1 port map( A1 => A_s(39), A2 => n1014, B1 => A_ns(39), B2 => 
                           n1008, ZN => n131);
   U158 : INV_X1 port map( A => n126, ZN => O_43_port);
   U159 : AOI221_X1 port map( B1 => n1020, B2 => A_ns(42), C1 => n1002, C2 => 
                           A_s(42), A => n1060, ZN => n126);
   U160 : INV_X1 port map( A => n127, ZN => n1060);
   U161 : AOI22_X1 port map( A1 => A_s(41), A2 => n1014, B1 => A_ns(41), B2 => 
                           n1008, ZN => n127);
   U162 : INV_X1 port map( A => n128, ZN => O_42_port);
   U163 : AOI221_X1 port map( B1 => n1020, B2 => A_ns(41), C1 => n1002, C2 => 
                           A_s(41), A => n1062, ZN => n128);
   U164 : INV_X1 port map( A => n129, ZN => n1062);
   U165 : AOI22_X1 port map( A1 => A_s(40), A2 => n1014, B1 => A_ns(40), B2 => 
                           n1008, ZN => n129);
   U166 : INV_X1 port map( A => n188, ZN => O_12_port);
   U167 : AOI221_X1 port map( B1 => A_ns(11), B2 => n1022, C1 => A_s(11), C2 =>
                           n1001, A => n1045, ZN => n188);
   U168 : INV_X1 port map( A => n105, ZN => O_7_port);
   U169 : AOI221_X1 port map( B1 => n1019, B2 => A_ns(6), C1 => n1001, C2 => 
                           A_s(6), A => n1035, ZN => n105);
   U170 : INV_X1 port map( A => n106, ZN => n1035);
   U171 : INV_X1 port map( A => n112, ZN => O_8_port);
   U172 : AOI221_X1 port map( B1 => n1019, B2 => A_ns(7), C1 => n1001, C2 => 
                           A_s(7), A => n1037, ZN => n112);
   U173 : INV_X1 port map( A => n113, ZN => n1037);
   U174 : INV_X1 port map( A => n103, ZN => O_9_port);
   U175 : AOI221_X1 port map( B1 => n1019, B2 => A_ns(8), C1 => n1001, C2 => 
                           A_s(8), A => n1039, ZN => n103);
   U176 : INV_X1 port map( A => n104, ZN => n1039);
   U177 : INV_X1 port map( A => n190, ZN => O_10_port);
   U178 : AOI221_X1 port map( B1 => n1019, B2 => A_ns(9), C1 => n1001, C2 => 
                           A_s(9), A => n1041, ZN => n190);
   U179 : INV_X1 port map( A => n191, ZN => n1041);
   U180 : INV_X1 port map( A => n101, ZN => O_11_port);
   U181 : AOI221_X1 port map( B1 => n1019, B2 => A_ns(10), C1 => n1001, C2 => 
                           A_s(10), A => n1043, ZN => n101);
   U182 : INV_X1 port map( A => n102, ZN => n1043);
   U183 : INV_X1 port map( A => n96, ZN => O_13_port);
   U184 : AOI221_X1 port map( B1 => n1020, B2 => A_ns(12), C1 => n1002, C2 => 
                           A_s(12), A => n1047, ZN => n96);
   U185 : INV_X1 port map( A => n111, ZN => O_1_port);
   U186 : AOI22_X1 port map( A1 => n1001, A2 => A_s(0), B1 => n1022, B2 => 
                           A_ns(0), ZN => n111);
   U187 : INV_X1 port map( A => n154, ZN => O_2_port);
   U188 : AOI221_X1 port map( B1 => n1021, B2 => A_ns(1), C1 => n1003, C2 => 
                           A_s(1), A => n1024, ZN => n154);
   U189 : INV_X1 port map( A => n155, ZN => n1024);
   U190 : INV_X1 port map( A => n109, ZN => O_3_port);
   U191 : AOI221_X1 port map( B1 => n1019, B2 => A_ns(2), C1 => n1001, C2 => 
                           A_s(2), A => n1027, ZN => n109);
   U192 : INV_X1 port map( A => n110, ZN => n1027);
   U193 : INV_X1 port map( A => n116, ZN => O_4_port);
   U195 : AOI221_X1 port map( B1 => n1019, B2 => A_ns(3), C1 => n1001, C2 => 
                           A_s(3), A => n1029, ZN => n116);
   U196 : INV_X1 port map( A => n117, ZN => n1029);
   U197 : INV_X1 port map( A => n107, ZN => O_5_port);
   U198 : AOI221_X1 port map( B1 => n1019, B2 => A_ns(4), C1 => n1001, C2 => 
                           A_s(4), A => n1031, ZN => n107);
   U199 : INV_X1 port map( A => n108, ZN => n1031);
   U200 : INV_X1 port map( A => n114, ZN => O_6_port);
   U201 : AOI221_X1 port map( B1 => n1019, B2 => A_ns(5), C1 => n1001, C2 => 
                           A_s(5), A => n1033, ZN => n114);
   U202 : INV_X1 port map( A => n115, ZN => n1033);
   U203 : INV_X1 port map( A => n189, ZN => n1045);
   U204 : AOI22_X1 port map( A1 => A_s(10), A2 => n1016, B1 => A_ns(10), B2 => 
                           n1010, ZN => n189);
   U205 : INV_X1 port map( A => n98, ZN => n1047);
   U206 : AOI22_X1 port map( A1 => A_s(11), A2 => n1014, B1 => A_ns(11), B2 => 
                           n1008, ZN => n98);
   U207 : AOI22_X1 port map( A1 => A_s(0), A2 => n1015, B1 => A_ns(0), B2 => 
                           n1009, ZN => n155);
   U208 : AOI22_X1 port map( A1 => A_s(1), A2 => n1013, B1 => A_ns(1), B2 => 
                           n1007, ZN => n110);
   U209 : AOI22_X1 port map( A1 => A_s(2), A2 => n1013, B1 => A_ns(2), B2 => 
                           n1007, ZN => n117);
   U210 : AOI22_X1 port map( A1 => A_s(3), A2 => n1013, B1 => A_ns(3), B2 => 
                           n1007, ZN => n108);
   U211 : AOI22_X1 port map( A1 => A_s(4), A2 => n1013, B1 => A_ns(4), B2 => 
                           n1007, ZN => n115);
   U212 : AOI22_X1 port map( A1 => A_s(5), A2 => n1013, B1 => A_ns(5), B2 => 
                           n1007, ZN => n106);
   U213 : AOI22_X1 port map( A1 => A_s(6), A2 => n1013, B1 => A_ns(6), B2 => 
                           n1007, ZN => n113);
   U214 : AOI22_X1 port map( A1 => A_s(7), A2 => n1013, B1 => A_ns(7), B2 => 
                           n1007, ZN => n104);
   U215 : AOI22_X1 port map( A1 => A_s(8), A2 => n1013, B1 => A_ns(8), B2 => 
                           n1007, ZN => n191);
   U216 : AOI22_X1 port map( A1 => A_s(9), A2 => n1013, B1 => A_ns(9), B2 => 
                           n1007, ZN => n102);
   U217 : AOI22_X1 port map( A1 => A_s(13), A2 => n1016, B1 => A_ns(13), B2 => 
                           n1010, ZN => n185);
   U218 : AOI221_X1 port map( B1 => n1022, B2 => A_ns(13), C1 => n1004, C2 => 
                           A_s(13), A => n1049, ZN => n186);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT46_i12 is

   port( A_s, A_ns, B : in std_logic_vector (45 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (45 downto 0));

end BOOTHENC_NBIT46_i12;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT46_i12 is

   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, 
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, 
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, 
      n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, 
      O_2_port, n985, O_1_port, O_3_port, n988, O_4_port, n990, O_5_port, n992,
      O_6_port, n994, O_7_port, n996, O_8_port, n998, O_9_port, n1000, 
      O_10_port, n1002, O_11_port, n1004, O_12_port, n1006, O_43_port, 
      O_44_port, n1009, O_45_port, n1011, O_42_port, n1013, O_41_port, n1015, 
      O_40_port, n1017, O_39_port, n1019, O_38_port, n1021, O_37_port, n1023, 
      O_36_port, n1025, O_35_port, n1027, O_34_port, n1029, O_33_port, n1031, 
      O_32_port, n1033, O_31_port, n1035, O_30_port, n1037, O_29_port, n1039, 
      O_28_port, n1041, O_27_port, n1043, O_26_port, n1045, O_25_port, n1047, 
      O_24_port, n1049, O_23_port, n1051, O_22_port, n1053, O_21_port, n1055, 
      O_20_port, n1057, O_19_port, n1059, O_18_port, n1061, O_17_port, n1063, 
      O_16_port, n1065, O_15_port, n1067, O_14_port, n1069, O_13_port, n1071, 
      n1072, n1073, n1074 : std_logic;

begin
   O <= ( O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, O_40_port, 
      O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, 
      O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, 
      O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, 
      O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, O_16_port, 
      O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, O_10_port, 
      O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, O_3_port, 
      O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), A_s(38), A_s(37), 
      A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), A_s(30), A_s(29), 
      A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), A_s(22), A_s(21), 
      A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), A_s(14), A_s(13), 
      A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), A_s(6), A_s(5), A_s(4)
      , A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, X_Logic0_port );
   A_nso <= ( A_ns(43), A_ns(42), A_ns(41), A_ns(40), A_ns(39), A_ns(38), 
      A_ns(37), A_ns(36), A_ns(35), A_ns(34), A_ns(33), A_ns(32), A_ns(31), 
      A_ns(30), A_ns(29), A_ns(28), A_ns(27), A_ns(26), A_ns(25), A_ns(24), 
      A_ns(23), A_ns(22), A_ns(21), A_ns(20), A_ns(19), A_ns(18), A_ns(17), 
      A_ns(16), A_ns(15), A_ns(14), A_ns(13), A_ns(12), A_ns(11), A_ns(10), 
      A_ns(9), A_ns(8), A_ns(7), A_ns(6), A_ns(5), A_ns(4), A_ns(3), A_ns(2), 
      A_ns(1), A_ns(0), X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U186 : XOR2_X1 port map( A => B(11), B => B(12), Z => n185);
   U2 : CLKBUF_X1 port map( A => n960, Z => n963);
   U3 : CLKBUF_X1 port map( A => n979, Z => n982);
   U4 : CLKBUF_X1 port map( A => n1073, Z => n961);
   U5 : CLKBUF_X1 port map( A => n973, Z => n976);
   U6 : CLKBUF_X1 port map( A => n967, Z => n970);
   U7 : CLKBUF_X1 port map( A => n93, Z => n978);
   U8 : CLKBUF_X1 port map( A => n96, Z => n966);
   U9 : CLKBUF_X1 port map( A => n95, Z => n972);
   U10 : BUF_X1 port map( A => n960, Z => n962);
   U11 : BUF_X1 port map( A => n961, Z => n965);
   U12 : BUF_X1 port map( A => n961, Z => n964);
   U13 : BUF_X1 port map( A => n979, Z => n983);
   U14 : BUF_X1 port map( A => n1073, Z => n960);
   U15 : BUF_X1 port map( A => n978, Z => n981);
   U16 : BUF_X1 port map( A => n978, Z => n980);
   U17 : INV_X1 port map( A => n112, ZN => O_45_port);
   U18 : BUF_X1 port map( A => n973, Z => n977);
   U19 : BUF_X1 port map( A => n967, Z => n971);
   U20 : BUF_X1 port map( A => n93, Z => n979);
   U21 : INV_X1 port map( A => n184, ZN => n1073);
   U22 : INV_X1 port map( A => n174, ZN => O_15_port);
   U23 : AOI221_X1 port map( B1 => n983, B2 => A_ns(14), C1 => n965, C2 => 
                           A_s(14), A => n1069, ZN => n174);
   U24 : INV_X1 port map( A => n175, ZN => n1069);
   U25 : AOI22_X1 port map( A1 => A_s(13), A2 => n977, B1 => A_ns(13), B2 => 
                           n971, ZN => n175);
   U26 : BUF_X1 port map( A => n972, Z => n975);
   U27 : BUF_X1 port map( A => n966, Z => n969);
   U28 : BUF_X1 port map( A => n972, Z => n974);
   U29 : BUF_X1 port map( A => n966, Z => n968);
   U30 : NAND2_X1 port map( A1 => n185, A2 => n1074, ZN => n184);
   U31 : BUF_X1 port map( A => n96, Z => n967);
   U32 : BUF_X1 port map( A => n95, Z => n973);
   U33 : AND2_X1 port map( A1 => n185, A2 => n184, ZN => n93);
   U34 : AOI221_X1 port map( B1 => n977, B2 => A_s(43), C1 => n971, C2 => 
                           A_ns(43), A => n1011, ZN => n112);
   U35 : INV_X1 port map( A => n113, ZN => n1011);
   U36 : AOI22_X1 port map( A1 => A_ns(44), A2 => n980, B1 => A_s(44), B2 => 
                           n962, ZN => n113);
   U37 : INV_X1 port map( A => n114, ZN => O_44_port);
   U38 : AOI221_X1 port map( B1 => n980, B2 => A_ns(43), C1 => n962, C2 => 
                           A_s(43), A => n1009, ZN => n114);
   U39 : INV_X1 port map( A => n115, ZN => n1009);
   U40 : AOI22_X1 port map( A1 => A_s(42), A2 => n974, B1 => A_ns(42), B2 => 
                           n968, ZN => n115);
   U41 : INV_X1 port map( A => n176, ZN => O_14_port);
   U42 : AOI221_X1 port map( B1 => n983, B2 => A_ns(13), C1 => n965, C2 => 
                           A_s(13), A => n1071, ZN => n176);
   U43 : INV_X1 port map( A => n177, ZN => n1071);
   U44 : AOI22_X1 port map( A1 => A_s(12), A2 => n977, B1 => A_ns(12), B2 => 
                           n971, ZN => n177);
   U45 : NOR3_X1 port map( A1 => B(11), A2 => B(12), A3 => n1074, ZN => n96);
   U46 : INV_X1 port map( A => n180, ZN => O_12_port);
   U47 : INV_X1 port map( A => n181, ZN => n1006);
   U48 : AOI22_X1 port map( A1 => A_s(10), A2 => n977, B1 => A_ns(10), B2 => 
                           n971, ZN => n181);
   U49 : INV_X1 port map( A => B(13), ZN => n1074);
   U50 : INV_X1 port map( A => n178, ZN => O_13_port);
   U51 : AOI221_X1 port map( B1 => n983, B2 => A_ns(12), C1 => n965, C2 => 
                           A_s(12), A => n1072, ZN => n178);
   U52 : INV_X1 port map( A => n179, ZN => n1072);
   U53 : AND3_X1 port map( A1 => B(11), A2 => n1074, A3 => B(12), ZN => n95);
   U54 : INV_X1 port map( A => n154, ZN => O_25_port);
   U55 : AOI221_X1 port map( B1 => n982, B2 => A_ns(24), C1 => n964, C2 => 
                           A_s(24), A => n1049, ZN => n154);
   U56 : INV_X1 port map( A => n155, ZN => n1049);
   U57 : AOI22_X1 port map( A1 => A_s(23), A2 => n976, B1 => A_ns(23), B2 => 
                           n970, ZN => n155);
   U58 : INV_X1 port map( A => n148, ZN => O_28_port);
   U59 : AOI221_X1 port map( B1 => n982, B2 => A_ns(27), C1 => n964, C2 => 
                           A_s(27), A => n1043, ZN => n148);
   U60 : INV_X1 port map( A => n149, ZN => n1043);
   U61 : AOI22_X1 port map( A1 => A_s(26), A2 => n976, B1 => A_ns(26), B2 => 
                           n970, ZN => n149);
   U62 : INV_X1 port map( A => n162, ZN => O_21_port);
   U63 : AOI221_X1 port map( B1 => n982, B2 => A_ns(20), C1 => n964, C2 => 
                           A_s(20), A => n1057, ZN => n162);
   U64 : INV_X1 port map( A => n163, ZN => n1057);
   U65 : AOI22_X1 port map( A1 => A_s(19), A2 => n976, B1 => A_ns(19), B2 => 
                           n970, ZN => n163);
   U66 : INV_X1 port map( A => n146, ZN => O_29_port);
   U67 : AOI221_X1 port map( B1 => n981, B2 => A_ns(28), C1 => n964, C2 => 
                           A_s(28), A => n1041, ZN => n146);
   U68 : INV_X1 port map( A => n147, ZN => n1041);
   U69 : AOI22_X1 port map( A1 => A_s(27), A2 => n976, B1 => A_ns(27), B2 => 
                           n970, ZN => n147);
   U70 : INV_X1 port map( A => n156, ZN => O_24_port);
   U71 : AOI221_X1 port map( B1 => n982, B2 => A_ns(23), C1 => n964, C2 => 
                           A_s(23), A => n1051, ZN => n156);
   U72 : INV_X1 port map( A => n157, ZN => n1051);
   U73 : AOI22_X1 port map( A1 => A_s(22), A2 => n976, B1 => A_ns(22), B2 => 
                           n970, ZN => n157);
   U74 : INV_X1 port map( A => n124, ZN => O_39_port);
   U75 : AOI221_X1 port map( B1 => n981, B2 => A_ns(38), C1 => n963, C2 => 
                           A_s(38), A => n1021, ZN => n124);
   U76 : INV_X1 port map( A => n125, ZN => n1021);
   U77 : AOI22_X1 port map( A1 => A_s(37), A2 => n975, B1 => A_ns(37), B2 => 
                           n969, ZN => n125);
   U78 : INV_X1 port map( A => n116, ZN => O_43_port);
   U79 : AOI221_X1 port map( B1 => n980, B2 => A_ns(42), C1 => n962, C2 => 
                           A_s(42), A => n1013, ZN => n116);
   U80 : INV_X1 port map( A => n117, ZN => n1013);
   U81 : AOI22_X1 port map( A1 => A_s(41), A2 => n974, B1 => A_ns(41), B2 => 
                           n968, ZN => n117);
   U82 : INV_X1 port map( A => n166, ZN => O_19_port);
   U83 : AOI221_X1 port map( B1 => n982, B2 => A_ns(18), C1 => n964, C2 => 
                           A_s(18), A => n1061, ZN => n166);
   U84 : INV_X1 port map( A => n167, ZN => n1061);
   U85 : AOI22_X1 port map( A1 => A_s(17), A2 => n977, B1 => A_ns(17), B2 => 
                           n971, ZN => n167);
   U86 : INV_X1 port map( A => n128, ZN => O_37_port);
   U87 : AOI221_X1 port map( B1 => n981, B2 => A_ns(36), C1 => n963, C2 => 
                           A_s(36), A => n1025, ZN => n128);
   U88 : INV_X1 port map( A => n129, ZN => n1025);
   U89 : AOI22_X1 port map( A1 => A_s(35), A2 => n975, B1 => A_ns(35), B2 => 
                           n969, ZN => n129);
   U90 : INV_X1 port map( A => n118, ZN => O_42_port);
   U91 : AOI221_X1 port map( B1 => n980, B2 => A_ns(41), C1 => n963, C2 => 
                           A_s(41), A => n1015, ZN => n118);
   U92 : INV_X1 port map( A => n119, ZN => n1015);
   U93 : AOI22_X1 port map( A1 => A_s(40), A2 => n974, B1 => A_ns(40), B2 => 
                           n968, ZN => n119);
   U94 : INV_X1 port map( A => n152, ZN => O_26_port);
   U95 : AOI221_X1 port map( B1 => n982, B2 => A_ns(25), C1 => n964, C2 => 
                           A_s(25), A => n1047, ZN => n152);
   U96 : INV_X1 port map( A => n153, ZN => n1047);
   U97 : AOI22_X1 port map( A1 => A_s(24), A2 => n976, B1 => A_ns(24), B2 => 
                           n970, ZN => n153);
   U98 : INV_X1 port map( A => n172, ZN => O_16_port);
   U99 : AOI221_X1 port map( B1 => n982, B2 => A_ns(15), C1 => n965, C2 => 
                           A_s(15), A => n1067, ZN => n172);
   U100 : INV_X1 port map( A => n173, ZN => n1067);
   U101 : AOI22_X1 port map( A1 => A_s(14), A2 => n976, B1 => A_ns(14), B2 => 
                           n970, ZN => n173);
   U102 : INV_X1 port map( A => n140, ZN => O_31_port);
   U103 : AOI221_X1 port map( B1 => n981, B2 => A_ns(30), C1 => n963, C2 => 
                           A_s(30), A => n1037, ZN => n140);
   U104 : INV_X1 port map( A => n141, ZN => n1037);
   U105 : AOI22_X1 port map( A1 => A_s(29), A2 => n975, B1 => A_ns(29), B2 => 
                           n969, ZN => n141);
   U106 : INV_X1 port map( A => n150, ZN => O_27_port);
   U107 : AOI221_X1 port map( B1 => n982, B2 => A_ns(26), C1 => n964, C2 => 
                           A_s(26), A => n1045, ZN => n150);
   U108 : INV_X1 port map( A => n151, ZN => n1045);
   U109 : AOI22_X1 port map( A1 => A_s(25), A2 => n976, B1 => A_ns(25), B2 => 
                           n970, ZN => n151);
   U110 : INV_X1 port map( A => n136, ZN => O_33_port);
   U111 : AOI221_X1 port map( B1 => n981, B2 => A_ns(32), C1 => n963, C2 => 
                           A_s(32), A => n1033, ZN => n136);
   U112 : INV_X1 port map( A => n137, ZN => n1033);
   U113 : AOI22_X1 port map( A1 => A_s(31), A2 => n975, B1 => A_ns(31), B2 => 
                           n969, ZN => n137);
   U114 : INV_X1 port map( A => n132, ZN => O_35_port);
   U115 : AOI221_X1 port map( B1 => n981, B2 => A_ns(34), C1 => n963, C2 => 
                           A_s(34), A => n1029, ZN => n132);
   U116 : INV_X1 port map( A => n133, ZN => n1029);
   U117 : AOI22_X1 port map( A1 => A_s(33), A2 => n975, B1 => A_ns(33), B2 => 
                           n969, ZN => n133);
   U118 : INV_X1 port map( A => n158, ZN => O_23_port);
   U119 : AOI221_X1 port map( B1 => n982, B2 => A_ns(22), C1 => n964, C2 => 
                           A_s(22), A => n1053, ZN => n158);
   U120 : INV_X1 port map( A => n159, ZN => n1053);
   U121 : AOI22_X1 port map( A1 => A_s(21), A2 => n976, B1 => A_ns(21), B2 => 
                           n970, ZN => n159);
   U122 : INV_X1 port map( A => n170, ZN => O_17_port);
   U123 : AOI221_X1 port map( B1 => n982, B2 => A_ns(16), C1 => n965, C2 => 
                           A_s(16), A => n1065, ZN => n170);
   U124 : INV_X1 port map( A => n171, ZN => n1065);
   U125 : AOI22_X1 port map( A1 => A_s(15), A2 => n977, B1 => A_ns(15), B2 => 
                           n971, ZN => n171);
   U126 : INV_X1 port map( A => n120, ZN => O_41_port);
   U127 : AOI221_X1 port map( B1 => n980, B2 => A_ns(40), C1 => n963, C2 => 
                           A_s(40), A => n1017, ZN => n120);
   U128 : INV_X1 port map( A => n121, ZN => n1017);
   U129 : AOI22_X1 port map( A1 => A_s(39), A2 => n974, B1 => A_ns(39), B2 => 
                           n968, ZN => n121);
   U130 : INV_X1 port map( A => n160, ZN => O_22_port);
   U131 : AOI221_X1 port map( B1 => n982, B2 => A_ns(21), C1 => n964, C2 => 
                           A_s(21), A => n1055, ZN => n160);
   U132 : INV_X1 port map( A => n161, ZN => n1055);
   U133 : AOI22_X1 port map( A1 => A_s(20), A2 => n976, B1 => A_ns(20), B2 => 
                           n970, ZN => n161);
   U134 : INV_X1 port map( A => n164, ZN => O_20_port);
   U135 : AOI221_X1 port map( B1 => n982, B2 => A_ns(19), C1 => n964, C2 => 
                           A_s(19), A => n1059, ZN => n164);
   U136 : INV_X1 port map( A => n165, ZN => n1059);
   U137 : AOI22_X1 port map( A1 => A_s(18), A2 => n976, B1 => A_ns(18), B2 => 
                           n970, ZN => n165);
   U138 : INV_X1 port map( A => n138, ZN => O_32_port);
   U139 : AOI221_X1 port map( B1 => n981, B2 => A_ns(31), C1 => n963, C2 => 
                           A_s(31), A => n1035, ZN => n138);
   U140 : INV_X1 port map( A => n139, ZN => n1035);
   U141 : AOI22_X1 port map( A1 => A_s(30), A2 => n975, B1 => A_ns(30), B2 => 
                           n969, ZN => n139);
   U142 : INV_X1 port map( A => n168, ZN => O_18_port);
   U143 : AOI221_X1 port map( B1 => n982, B2 => A_ns(17), C1 => n965, C2 => 
                           A_s(17), A => n1063, ZN => n168);
   U144 : INV_X1 port map( A => n169, ZN => n1063);
   U145 : AOI22_X1 port map( A1 => A_s(16), A2 => n977, B1 => A_ns(16), B2 => 
                           n971, ZN => n169);
   U146 : INV_X1 port map( A => n142, ZN => O_30_port);
   U147 : AOI221_X1 port map( B1 => n981, B2 => A_ns(29), C1 => n964, C2 => 
                           A_s(29), A => n1039, ZN => n142);
   U148 : INV_X1 port map( A => n143, ZN => n1039);
   U149 : AOI22_X1 port map( A1 => A_s(28), A2 => n975, B1 => A_ns(28), B2 => 
                           n969, ZN => n143);
   U150 : INV_X1 port map( A => n134, ZN => O_34_port);
   U151 : AOI221_X1 port map( B1 => n981, B2 => A_ns(33), C1 => n963, C2 => 
                           A_s(33), A => n1031, ZN => n134);
   U152 : INV_X1 port map( A => n135, ZN => n1031);
   U153 : AOI22_X1 port map( A1 => A_s(32), A2 => n975, B1 => A_ns(32), B2 => 
                           n969, ZN => n135);
   U154 : INV_X1 port map( A => n130, ZN => O_36_port);
   U155 : AOI221_X1 port map( B1 => n981, B2 => A_ns(35), C1 => n963, C2 => 
                           A_s(35), A => n1027, ZN => n130);
   U156 : INV_X1 port map( A => n131, ZN => n1027);
   U157 : AOI22_X1 port map( A1 => A_s(34), A2 => n975, B1 => A_ns(34), B2 => 
                           n969, ZN => n131);
   U158 : INV_X1 port map( A => n126, ZN => O_38_port);
   U159 : AOI221_X1 port map( B1 => n981, B2 => A_ns(37), C1 => n963, C2 => 
                           A_s(37), A => n1023, ZN => n126);
   U160 : INV_X1 port map( A => n127, ZN => n1023);
   U161 : AOI22_X1 port map( A1 => A_s(36), A2 => n975, B1 => A_ns(36), B2 => 
                           n969, ZN => n127);
   U162 : INV_X1 port map( A => n122, ZN => O_40_port);
   U163 : AOI221_X1 port map( B1 => n980, B2 => A_ns(39), C1 => n963, C2 => 
                           A_s(39), A => n1019, ZN => n122);
   U164 : INV_X1 port map( A => n123, ZN => n1019);
   U165 : AOI22_X1 port map( A1 => A_s(38), A2 => n975, B1 => A_ns(38), B2 => 
                           n969, ZN => n123);
   U166 : INV_X1 port map( A => n92, ZN => O_11_port);
   U167 : AOI221_X1 port map( B1 => n981, B2 => A_ns(10), C1 => n963, C2 => 
                           A_s(10), A => n1004, ZN => n92);
   U168 : INV_X1 port map( A => n99, ZN => O_7_port);
   U169 : AOI221_X1 port map( B1 => n980, B2 => A_ns(6), C1 => n962, C2 => 
                           A_s(6), A => n996, ZN => n99);
   U170 : INV_X1 port map( A => n100, ZN => n996);
   U171 : INV_X1 port map( A => n106, ZN => O_8_port);
   U172 : AOI221_X1 port map( B1 => n980, B2 => A_ns(7), C1 => n962, C2 => 
                           A_s(7), A => n998, ZN => n106);
   U173 : INV_X1 port map( A => n107, ZN => n998);
   U174 : INV_X1 port map( A => n97, ZN => O_9_port);
   U175 : AOI221_X1 port map( B1 => n980, B2 => A_ns(8), C1 => n962, C2 => 
                           A_s(8), A => n1000, ZN => n97);
   U176 : INV_X1 port map( A => n98, ZN => n1000);
   U177 : INV_X1 port map( A => n182, ZN => O_10_port);
   U178 : AOI221_X1 port map( B1 => A_ns(9), B2 => n983, C1 => A_s(9), C2 => 
                           n962, A => n1002, ZN => n182);
   U179 : INV_X1 port map( A => n105, ZN => O_1_port);
   U180 : AOI22_X1 port map( A1 => n962, A2 => A_s(0), B1 => n983, B2 => 
                           A_ns(0), ZN => n105);
   U181 : INV_X1 port map( A => n144, ZN => O_2_port);
   U182 : AOI221_X1 port map( B1 => n981, B2 => A_ns(1), C1 => n964, C2 => 
                           A_s(1), A => n985, ZN => n144);
   U183 : INV_X1 port map( A => n145, ZN => n985);
   U184 : INV_X1 port map( A => n103, ZN => O_3_port);
   U185 : AOI221_X1 port map( B1 => n980, B2 => A_ns(2), C1 => n962, C2 => 
                           A_s(2), A => n988, ZN => n103);
   U187 : INV_X1 port map( A => n104, ZN => n988);
   U188 : INV_X1 port map( A => n110, ZN => O_4_port);
   U189 : AOI221_X1 port map( B1 => n980, B2 => A_ns(3), C1 => n962, C2 => 
                           A_s(3), A => n990, ZN => n110);
   U190 : INV_X1 port map( A => n111, ZN => n990);
   U191 : INV_X1 port map( A => n101, ZN => O_5_port);
   U192 : AOI221_X1 port map( B1 => n980, B2 => A_ns(4), C1 => n962, C2 => 
                           A_s(4), A => n992, ZN => n101);
   U193 : INV_X1 port map( A => n102, ZN => n992);
   U194 : INV_X1 port map( A => n108, ZN => O_6_port);
   U195 : AOI221_X1 port map( B1 => n980, B2 => A_ns(5), C1 => n962, C2 => 
                           A_s(5), A => n994, ZN => n108);
   U196 : INV_X1 port map( A => n109, ZN => n994);
   U197 : INV_X1 port map( A => n183, ZN => n1002);
   U198 : AOI22_X1 port map( A1 => A_s(8), A2 => n974, B1 => A_ns(8), B2 => 
                           n968, ZN => n183);
   U199 : INV_X1 port map( A => n94, ZN => n1004);
   U200 : AOI22_X1 port map( A1 => A_s(9), A2 => n975, B1 => A_ns(9), B2 => 
                           n969, ZN => n94);
   U201 : AOI22_X1 port map( A1 => A_s(0), A2 => n976, B1 => A_ns(0), B2 => 
                           n970, ZN => n145);
   U202 : AOI22_X1 port map( A1 => A_s(1), A2 => n974, B1 => A_ns(1), B2 => 
                           n968, ZN => n104);
   U203 : AOI22_X1 port map( A1 => A_s(2), A2 => n974, B1 => A_ns(2), B2 => 
                           n968, ZN => n111);
   U204 : AOI22_X1 port map( A1 => A_s(3), A2 => n974, B1 => A_ns(3), B2 => 
                           n968, ZN => n102);
   U205 : AOI22_X1 port map( A1 => A_s(4), A2 => n974, B1 => A_ns(4), B2 => 
                           n968, ZN => n109);
   U206 : AOI22_X1 port map( A1 => A_s(5), A2 => n974, B1 => A_ns(5), B2 => 
                           n968, ZN => n100);
   U207 : AOI22_X1 port map( A1 => A_s(6), A2 => n974, B1 => A_ns(6), B2 => 
                           n968, ZN => n107);
   U208 : AOI22_X1 port map( A1 => A_s(7), A2 => n974, B1 => A_ns(7), B2 => 
                           n968, ZN => n98);
   U209 : AOI22_X1 port map( A1 => A_s(11), A2 => n977, B1 => A_ns(11), B2 => 
                           n971, ZN => n179);
   U210 : AOI221_X1 port map( B1 => n983, B2 => A_ns(11), C1 => n962, C2 => 
                           A_s(11), A => n1006, ZN => n180);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT44_i10 is

   port( A_s, A_ns, B : in std_logic_vector (43 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (43 downto 0));

end BOOTHENC_NBIT44_i10;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT44_i10 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
      n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, 
      n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, 
      n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, 
      n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n924, n925, n926, n927, n928, 
      n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, 
      n941, n942, n943, n944, n945, n946, n947, O_2_port, n949, O_1_port, 
      O_3_port, n952, O_4_port, n954, O_5_port, n956, O_6_port, n958, O_7_port,
      n960, O_8_port, n962, O_9_port, n964, O_10_port, n966, O_41_port, 
      O_42_port, n969, O_43_port, n971, O_40_port, n973, O_39_port, n975, 
      O_38_port, n977, O_37_port, n979, O_36_port, n981, O_35_port, n983, 
      O_34_port, n985, O_33_port, n987, O_32_port, n989, O_31_port, n991, 
      O_30_port, n993, O_29_port, n995, O_28_port, n997, O_27_port, n999, 
      O_26_port, n1001, O_25_port, n1003, O_24_port, n1005, O_23_port, n1007, 
      O_22_port, n1009, O_21_port, n1011, O_20_port, n1013, O_19_port, n1015, 
      O_18_port, n1017, O_17_port, n1019, O_16_port, n1021, O_15_port, n1023, 
      O_14_port, n1025, O_13_port, n1027, O_12_port, n1029, O_11_port, n1031, 
      n1032, n1033, n1034 : std_logic;

begin
   O <= ( O_43_port, O_42_port, O_41_port, O_40_port, O_39_port, O_38_port, 
      O_37_port, O_36_port, O_35_port, O_34_port, O_33_port, O_32_port, 
      O_31_port, O_30_port, O_29_port, O_28_port, O_27_port, O_26_port, 
      O_25_port, O_24_port, O_23_port, O_22_port, O_21_port, O_20_port, 
      O_19_port, O_18_port, O_17_port, O_16_port, O_15_port, O_14_port, 
      O_13_port, O_12_port, O_11_port, O_10_port, O_9_port, O_8_port, O_7_port,
      O_6_port, O_5_port, O_4_port, O_3_port, O_2_port, O_1_port, X_Logic0_port
      );
   A_so <= ( A_s(41), A_s(40), A_s(39), A_s(38), A_s(37), A_s(36), A_s(35), 
      A_s(34), A_s(33), A_s(32), A_s(31), A_s(30), A_s(29), A_s(28), A_s(27), 
      A_s(26), A_s(25), A_s(24), A_s(23), A_s(22), A_s(21), A_s(20), A_s(19), 
      A_s(18), A_s(17), A_s(16), A_s(15), A_s(14), A_s(13), A_s(12), A_s(11), 
      A_s(10), A_s(9), A_s(8), A_s(7), A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), 
      A_s(1), A_s(0), X_Logic0_port, X_Logic0_port );
   A_nso <= ( A_ns(41), A_ns(40), A_ns(39), A_ns(38), A_ns(37), A_ns(36), 
      A_ns(35), A_ns(34), A_ns(33), A_ns(32), A_ns(31), A_ns(30), A_ns(29), 
      A_ns(28), A_ns(27), A_ns(26), A_ns(25), A_ns(24), A_ns(23), A_ns(22), 
      A_ns(21), A_ns(20), A_ns(19), A_ns(18), A_ns(17), A_ns(16), A_ns(15), 
      A_ns(14), A_ns(13), A_ns(12), A_ns(11), A_ns(10), A_ns(9), A_ns(8), 
      A_ns(7), A_ns(6), A_ns(5), A_ns(4), A_ns(3), A_ns(2), A_ns(1), A_ns(0), 
      X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U178 : XOR2_X1 port map( A => B(10), B => B(9), Z => n177);
   U2 : CLKBUF_X1 port map( A => n924, Z => n927);
   U3 : CLKBUF_X1 port map( A => n942, Z => n945);
   U4 : CLKBUF_X1 port map( A => n92, Z => n930);
   U5 : CLKBUF_X1 port map( A => n91, Z => n936);
   U6 : CLKBUF_X1 port map( A => n925, Z => n928);
   U7 : BUF_X2 port map( A => n943, Z => n946);
   U8 : CLKBUF_X1 port map( A => n943, Z => n947);
   U9 : CLKBUF_X1 port map( A => n89, Z => n942);
   U10 : CLKBUF_X1 port map( A => n937, Z => n940);
   U11 : CLKBUF_X1 port map( A => n931, Z => n934);
   U12 : BUF_X1 port map( A => n924, Z => n926);
   U13 : BUF_X1 port map( A => n925, Z => n929);
   U14 : BUF_X1 port map( A => n942, Z => n944);
   U15 : BUF_X1 port map( A => n1033, Z => n924);
   U16 : BUF_X1 port map( A => n1033, Z => n925);
   U17 : INV_X1 port map( A => n168, ZN => O_13_port);
   U18 : AOI221_X1 port map( B1 => n947, B2 => A_ns(12), C1 => n929, C2 => 
                           A_s(12), A => n1029, ZN => n168);
   U19 : INV_X1 port map( A => n106, ZN => O_43_port);
   U20 : INV_X1 port map( A => n169, ZN => n1029);
   U21 : AOI22_X1 port map( A1 => A_s(11), A2 => n941, B1 => A_ns(11), B2 => 
                           n935, ZN => n169);
   U22 : BUF_X1 port map( A => n937, Z => n941);
   U23 : BUF_X1 port map( A => n931, Z => n935);
   U24 : BUF_X1 port map( A => n89, Z => n943);
   U25 : INV_X1 port map( A => n176, ZN => n1033);
   U26 : BUF_X1 port map( A => n936, Z => n939);
   U27 : BUF_X1 port map( A => n930, Z => n933);
   U28 : BUF_X1 port map( A => n936, Z => n938);
   U29 : BUF_X1 port map( A => n930, Z => n932);
   U30 : INV_X1 port map( A => n170, ZN => O_12_port);
   U31 : NAND2_X1 port map( A1 => n177, A2 => n1034, ZN => n176);
   U32 : BUF_X1 port map( A => n92, Z => n931);
   U33 : BUF_X1 port map( A => n91, Z => n937);
   U34 : AND2_X1 port map( A1 => n177, A2 => n176, ZN => n89);
   U35 : AOI221_X1 port map( B1 => n941, B2 => A_s(41), C1 => n935, C2 => 
                           A_ns(41), A => n971, ZN => n106);
   U36 : INV_X1 port map( A => n107, ZN => n971);
   U37 : AOI22_X1 port map( A1 => A_ns(42), A2 => n944, B1 => A_s(42), B2 => 
                           n926, ZN => n107);
   U38 : INV_X1 port map( A => n108, ZN => O_42_port);
   U39 : AOI221_X1 port map( B1 => n944, B2 => A_ns(41), C1 => n926, C2 => 
                           A_s(41), A => n969, ZN => n108);
   U40 : INV_X1 port map( A => n109, ZN => n969);
   U41 : AOI22_X1 port map( A1 => A_s(40), A2 => n938, B1 => A_ns(40), B2 => 
                           n932, ZN => n109);
   U42 : INV_X1 port map( A => n174, ZN => O_10_port);
   U43 : INV_X1 port map( A => n175, ZN => n966);
   U44 : AOI22_X1 port map( A1 => A_s(8), A2 => n938, B1 => A_ns(8), B2 => n932
                           , ZN => n175);
   U45 : AOI221_X1 port map( B1 => n947, B2 => A_ns(11), C1 => n929, C2 => 
                           A_s(11), A => n1031, ZN => n170);
   U46 : INV_X1 port map( A => n171, ZN => n1031);
   U47 : AOI22_X1 port map( A1 => A_s(10), A2 => n941, B1 => A_ns(10), B2 => 
                           n935, ZN => n171);
   U48 : NOR3_X1 port map( A1 => B(10), A2 => B(9), A3 => n1034, ZN => n92);
   U49 : INV_X1 port map( A => n164, ZN => O_15_port);
   U50 : AOI221_X1 port map( B1 => n946, B2 => A_ns(14), C1 => n928, C2 => 
                           A_s(14), A => n1025, ZN => n164);
   U51 : INV_X1 port map( A => n165, ZN => n1025);
   U52 : AOI22_X1 port map( A1 => A_s(13), A2 => n941, B1 => A_ns(13), B2 => 
                           n935, ZN => n165);
   U53 : INV_X1 port map( A => n166, ZN => O_14_port);
   U54 : AOI221_X1 port map( B1 => n946, B2 => A_ns(13), C1 => n929, C2 => 
                           A_s(13), A => n1027, ZN => n166);
   U55 : INV_X1 port map( A => n167, ZN => n1027);
   U56 : AOI22_X1 port map( A1 => A_s(12), A2 => n941, B1 => A_ns(12), B2 => 
                           n935, ZN => n167);
   U57 : INV_X1 port map( A => B(11), ZN => n1034);
   U58 : INV_X1 port map( A => n172, ZN => O_11_port);
   U59 : AOI221_X1 port map( B1 => n946, B2 => A_ns(10), C1 => n929, C2 => 
                           A_s(10), A => n1032, ZN => n172);
   U60 : INV_X1 port map( A => n173, ZN => n1032);
   U61 : INV_X1 port map( A => n162, ZN => O_16_port);
   U62 : AOI221_X1 port map( B1 => n946, B2 => A_ns(15), C1 => n928, C2 => 
                           A_s(15), A => n1023, ZN => n162);
   U63 : INV_X1 port map( A => n163, ZN => n1023);
   U64 : AOI22_X1 port map( A1 => A_s(14), A2 => n940, B1 => A_ns(14), B2 => 
                           n934, ZN => n163);
   U65 : INV_X1 port map( A => n156, ZN => O_19_port);
   U66 : AOI221_X1 port map( B1 => n946, B2 => A_ns(18), C1 => n928, C2 => 
                           A_s(18), A => n1017, ZN => n156);
   U67 : INV_X1 port map( A => n157, ZN => n1017);
   U68 : AOI22_X1 port map( A1 => A_s(17), A2 => n940, B1 => A_ns(17), B2 => 
                           n934, ZN => n157);
   U69 : INV_X1 port map( A => n160, ZN => O_17_port);
   U70 : AOI221_X1 port map( B1 => n946, B2 => A_ns(16), C1 => n928, C2 => 
                           A_s(16), A => n1021, ZN => n160);
   U71 : INV_X1 port map( A => n161, ZN => n1021);
   U72 : AOI22_X1 port map( A1 => A_s(15), A2 => n940, B1 => A_ns(15), B2 => 
                           n934, ZN => n161);
   U73 : INV_X1 port map( A => n158, ZN => O_18_port);
   U74 : AOI221_X1 port map( B1 => n946, B2 => A_ns(17), C1 => n928, C2 => 
                           A_s(17), A => n1019, ZN => n158);
   U75 : INV_X1 port map( A => n159, ZN => n1019);
   U76 : AOI22_X1 port map( A1 => A_s(16), A2 => n940, B1 => A_ns(16), B2 => 
                           n934, ZN => n159);
   U77 : AND3_X1 port map( A1 => B(10), A2 => n1034, A3 => B(9), ZN => n91);
   U78 : INV_X1 port map( A => n144, ZN => O_25_port);
   U79 : AOI221_X1 port map( B1 => n946, B2 => A_ns(24), C1 => n928, C2 => 
                           A_s(24), A => n1005, ZN => n144);
   U80 : INV_X1 port map( A => n145, ZN => n1005);
   U81 : AOI22_X1 port map( A1 => A_s(23), A2 => n940, B1 => A_ns(23), B2 => 
                           n934, ZN => n145);
   U82 : INV_X1 port map( A => n140, ZN => O_27_port);
   U83 : AOI221_X1 port map( B1 => n945, B2 => A_ns(26), C1 => n928, C2 => 
                           A_s(26), A => n1001, ZN => n140);
   U84 : INV_X1 port map( A => n141, ZN => n1001);
   U85 : AOI22_X1 port map( A1 => A_s(25), A2 => n940, B1 => A_ns(25), B2 => 
                           n934, ZN => n141);
   U86 : INV_X1 port map( A => n154, ZN => O_20_port);
   U87 : AOI221_X1 port map( B1 => n946, B2 => A_ns(19), C1 => n928, C2 => 
                           A_s(19), A => n1015, ZN => n154);
   U88 : INV_X1 port map( A => n155, ZN => n1015);
   U89 : AOI22_X1 port map( A1 => A_s(18), A2 => n940, B1 => A_ns(18), B2 => 
                           n934, ZN => n155);
   U90 : INV_X1 port map( A => n138, ZN => O_28_port);
   U91 : AOI221_X1 port map( B1 => n945, B2 => A_ns(27), C1 => n927, C2 => 
                           A_s(27), A => n999, ZN => n138);
   U92 : INV_X1 port map( A => n139, ZN => n999);
   U93 : AOI22_X1 port map( A1 => A_s(26), A2 => n939, B1 => A_ns(26), B2 => 
                           n933, ZN => n139);
   U94 : INV_X1 port map( A => n142, ZN => O_26_port);
   U95 : AOI221_X1 port map( B1 => n945, B2 => A_ns(25), C1 => n928, C2 => 
                           A_s(25), A => n1003, ZN => n142);
   U96 : INV_X1 port map( A => n143, ZN => n1003);
   U97 : AOI22_X1 port map( A1 => A_s(24), A2 => n940, B1 => A_ns(24), B2 => 
                           n934, ZN => n143);
   U98 : INV_X1 port map( A => n132, ZN => O_30_port);
   U99 : AOI221_X1 port map( B1 => n945, B2 => A_ns(29), C1 => n927, C2 => 
                           A_s(29), A => n995, ZN => n132);
   U100 : INV_X1 port map( A => n133, ZN => n995);
   U101 : AOI22_X1 port map( A1 => A_s(28), A2 => n939, B1 => A_ns(28), B2 => 
                           n933, ZN => n133);
   U102 : INV_X1 port map( A => n118, ZN => O_37_port);
   U103 : AOI221_X1 port map( B1 => n944, B2 => A_ns(36), C1 => n927, C2 => 
                           A_s(36), A => n981, ZN => n118);
   U104 : INV_X1 port map( A => n119, ZN => n981);
   U105 : AOI22_X1 port map( A1 => A_s(35), A2 => n939, B1 => A_ns(35), B2 => 
                           n933, ZN => n119);
   U106 : INV_X1 port map( A => n114, ZN => O_39_port);
   U107 : AOI221_X1 port map( B1 => n944, B2 => A_ns(38), C1 => n926, C2 => 
                           A_s(38), A => n977, ZN => n114);
   U108 : INV_X1 port map( A => n115, ZN => n977);
   U109 : AOI22_X1 port map( A1 => A_s(37), A2 => n938, B1 => A_ns(37), B2 => 
                           n932, ZN => n115);
   U110 : INV_X1 port map( A => n110, ZN => O_41_port);
   U111 : AOI221_X1 port map( B1 => n944, B2 => A_ns(40), C1 => n926, C2 => 
                           A_s(40), A => n973, ZN => n110);
   U112 : INV_X1 port map( A => n111, ZN => n973);
   U113 : AOI22_X1 port map( A1 => A_s(39), A2 => n938, B1 => A_ns(39), B2 => 
                           n932, ZN => n111);
   U114 : INV_X1 port map( A => n116, ZN => O_38_port);
   U115 : AOI221_X1 port map( B1 => n944, B2 => A_ns(37), C1 => n927, C2 => 
                           A_s(37), A => n979, ZN => n116);
   U116 : INV_X1 port map( A => n117, ZN => n979);
   U117 : AOI22_X1 port map( A1 => A_s(36), A2 => n938, B1 => A_ns(36), B2 => 
                           n932, ZN => n117);
   U118 : INV_X1 port map( A => n112, ZN => O_40_port);
   U119 : AOI221_X1 port map( B1 => n944, B2 => A_ns(39), C1 => n926, C2 => 
                           A_s(39), A => n975, ZN => n112);
   U120 : INV_X1 port map( A => n113, ZN => n975);
   U121 : AOI22_X1 port map( A1 => A_s(38), A2 => n938, B1 => A_ns(38), B2 => 
                           n932, ZN => n113);
   U122 : INV_X1 port map( A => n146, ZN => O_24_port);
   U123 : AOI221_X1 port map( B1 => n946, B2 => A_ns(23), C1 => n928, C2 => 
                           A_s(23), A => n1007, ZN => n146);
   U124 : INV_X1 port map( A => n147, ZN => n1007);
   U125 : AOI22_X1 port map( A1 => A_s(22), A2 => n940, B1 => A_ns(22), B2 => 
                           n934, ZN => n147);
   U126 : INV_X1 port map( A => n136, ZN => O_29_port);
   U127 : AOI221_X1 port map( B1 => n945, B2 => A_ns(28), C1 => n927, C2 => 
                           A_s(28), A => n997, ZN => n136);
   U128 : INV_X1 port map( A => n137, ZN => n997);
   U129 : AOI22_X1 port map( A1 => A_s(27), A2 => n939, B1 => A_ns(27), B2 => 
                           n933, ZN => n137);
   U130 : INV_X1 port map( A => n152, ZN => O_21_port);
   U131 : AOI221_X1 port map( B1 => n946, B2 => A_ns(20), C1 => n928, C2 => 
                           A_s(20), A => n1013, ZN => n152);
   U132 : INV_X1 port map( A => n153, ZN => n1013);
   U133 : AOI22_X1 port map( A1 => A_s(19), A2 => n940, B1 => A_ns(19), B2 => 
                           n934, ZN => n153);
   U134 : INV_X1 port map( A => n126, ZN => O_33_port);
   U135 : AOI221_X1 port map( B1 => n945, B2 => A_ns(32), C1 => n927, C2 => 
                           A_s(32), A => n989, ZN => n126);
   U136 : INV_X1 port map( A => n127, ZN => n989);
   U137 : AOI22_X1 port map( A1 => A_s(31), A2 => n939, B1 => A_ns(31), B2 => 
                           n933, ZN => n127);
   U138 : INV_X1 port map( A => n122, ZN => O_35_port);
   U139 : AOI221_X1 port map( B1 => n945, B2 => A_ns(34), C1 => n927, C2 => 
                           A_s(34), A => n985, ZN => n122);
   U140 : INV_X1 port map( A => n123, ZN => n985);
   U141 : AOI22_X1 port map( A1 => A_s(33), A2 => n939, B1 => A_ns(33), B2 => 
                           n933, ZN => n123);
   U142 : INV_X1 port map( A => n130, ZN => O_31_port);
   U143 : AOI221_X1 port map( B1 => n945, B2 => A_ns(30), C1 => n927, C2 => 
                           A_s(30), A => n993, ZN => n130);
   U144 : INV_X1 port map( A => n131, ZN => n993);
   U145 : AOI22_X1 port map( A1 => A_s(29), A2 => n939, B1 => A_ns(29), B2 => 
                           n933, ZN => n131);
   U146 : INV_X1 port map( A => n148, ZN => O_23_port);
   U147 : AOI221_X1 port map( B1 => n946, B2 => A_ns(22), C1 => n928, C2 => 
                           A_s(22), A => n1009, ZN => n148);
   U148 : INV_X1 port map( A => n149, ZN => n1009);
   U149 : AOI22_X1 port map( A1 => A_s(21), A2 => n940, B1 => A_ns(21), B2 => 
                           n934, ZN => n149);
   U150 : INV_X1 port map( A => n128, ZN => O_32_port);
   U151 : AOI221_X1 port map( B1 => n945, B2 => A_ns(31), C1 => n927, C2 => 
                           A_s(31), A => n991, ZN => n128);
   U152 : INV_X1 port map( A => n129, ZN => n991);
   U153 : AOI22_X1 port map( A1 => A_s(30), A2 => n939, B1 => A_ns(30), B2 => 
                           n933, ZN => n129);
   U154 : INV_X1 port map( A => n150, ZN => O_22_port);
   U155 : AOI221_X1 port map( B1 => n946, B2 => A_ns(21), C1 => n928, C2 => 
                           A_s(21), A => n1011, ZN => n150);
   U156 : INV_X1 port map( A => n151, ZN => n1011);
   U157 : AOI22_X1 port map( A1 => A_s(20), A2 => n940, B1 => A_ns(20), B2 => 
                           n934, ZN => n151);
   U158 : INV_X1 port map( A => n120, ZN => O_36_port);
   U159 : AOI221_X1 port map( B1 => n945, B2 => A_ns(35), C1 => n927, C2 => 
                           A_s(35), A => n983, ZN => n120);
   U160 : INV_X1 port map( A => n121, ZN => n983);
   U161 : AOI22_X1 port map( A1 => A_s(34), A2 => n939, B1 => A_ns(34), B2 => 
                           n933, ZN => n121);
   U162 : INV_X1 port map( A => n124, ZN => O_34_port);
   U163 : AOI221_X1 port map( B1 => n945, B2 => A_ns(33), C1 => n927, C2 => 
                           A_s(33), A => n987, ZN => n124);
   U164 : INV_X1 port map( A => n125, ZN => n987);
   U165 : AOI22_X1 port map( A1 => A_s(32), A2 => n939, B1 => A_ns(32), B2 => 
                           n933, ZN => n125);
   U166 : INV_X1 port map( A => n93, ZN => O_7_port);
   U167 : AOI221_X1 port map( B1 => n944, B2 => A_ns(6), C1 => n926, C2 => 
                           A_s(6), A => n960, ZN => n93);
   U168 : INV_X1 port map( A => n88, ZN => O_9_port);
   U169 : AOI221_X1 port map( B1 => n945, B2 => A_ns(8), C1 => n927, C2 => 
                           A_s(8), A => n964, ZN => n88);
   U170 : INV_X1 port map( A => n100, ZN => O_8_port);
   U171 : AOI221_X1 port map( B1 => A_ns(7), B2 => n947, C1 => A_s(7), C2 => 
                           n926, A => n962, ZN => n100);
   U172 : INV_X1 port map( A => n99, ZN => O_1_port);
   U173 : INV_X1 port map( A => n97, ZN => O_3_port);
   U174 : AOI221_X1 port map( B1 => n944, B2 => A_ns(2), C1 => n926, C2 => 
                           A_s(2), A => n952, ZN => n97);
   U175 : INV_X1 port map( A => n102, ZN => O_6_port);
   U176 : AOI221_X1 port map( B1 => n944, B2 => A_ns(5), C1 => n926, C2 => 
                           A_s(5), A => n958, ZN => n102);
   U177 : INV_X1 port map( A => n134, ZN => O_2_port);
   U179 : AOI221_X1 port map( B1 => n945, B2 => A_ns(1), C1 => n927, C2 => 
                           A_s(1), A => n949, ZN => n134);
   U180 : INV_X1 port map( A => n104, ZN => O_4_port);
   U181 : AOI221_X1 port map( B1 => n944, B2 => A_ns(3), C1 => n926, C2 => 
                           A_s(3), A => n954, ZN => n104);
   U182 : INV_X1 port map( A => n95, ZN => O_5_port);
   U183 : AOI221_X1 port map( B1 => n944, B2 => A_ns(4), C1 => n926, C2 => 
                           A_s(4), A => n956, ZN => n95);
   U184 : INV_X1 port map( A => n135, ZN => n949);
   U185 : AOI22_X1 port map( A1 => A_s(0), A2 => n939, B1 => A_ns(0), B2 => 
                           n933, ZN => n135);
   U186 : INV_X1 port map( A => n98, ZN => n952);
   U187 : AOI22_X1 port map( A1 => A_s(1), A2 => n938, B1 => A_ns(1), B2 => 
                           n932, ZN => n98);
   U188 : INV_X1 port map( A => n105, ZN => n954);
   U189 : AOI22_X1 port map( A1 => A_s(2), A2 => n938, B1 => A_ns(2), B2 => 
                           n932, ZN => n105);
   U190 : INV_X1 port map( A => n96, ZN => n956);
   U191 : AOI22_X1 port map( A1 => A_s(3), A2 => n938, B1 => A_ns(3), B2 => 
                           n932, ZN => n96);
   U192 : INV_X1 port map( A => n103, ZN => n958);
   U193 : AOI22_X1 port map( A1 => A_s(4), A2 => n938, B1 => A_ns(4), B2 => 
                           n932, ZN => n103);
   U194 : INV_X1 port map( A => n94, ZN => n960);
   U195 : AOI22_X1 port map( A1 => A_s(5), A2 => n938, B1 => A_ns(5), B2 => 
                           n932, ZN => n94);
   U196 : INV_X1 port map( A => n101, ZN => n962);
   U197 : AOI22_X1 port map( A1 => A_s(6), A2 => n938, B1 => A_ns(6), B2 => 
                           n932, ZN => n101);
   U198 : INV_X1 port map( A => n90, ZN => n964);
   U199 : AOI22_X1 port map( A1 => A_s(7), A2 => n939, B1 => A_ns(7), B2 => 
                           n933, ZN => n90);
   U200 : AOI22_X1 port map( A1 => n926, A2 => A_s(0), B1 => n947, B2 => 
                           A_ns(0), ZN => n99);
   U201 : AOI221_X1 port map( B1 => n944, B2 => A_ns(9), C1 => n926, C2 => 
                           A_s(9), A => n966, ZN => n174);
   U202 : AOI22_X1 port map( A1 => A_s(9), A2 => n941, B1 => A_ns(9), B2 => 
                           n935, ZN => n173);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT42_i8 is

   port( A_s, A_ns, B : in std_logic_vector (41 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (41 downto 0));

end BOOTHENC_NBIT42_i8;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT42_i8 is

   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
      n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, 
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, 
      n168, n169, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, 
      n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, 
      n901, n902, O_2_port, n904, O_1_port, O_3_port, n907, O_4_port, n909, 
      O_5_port, n911, O_6_port, n913, O_7_port, n915, O_8_port, n917, O_39_port
      , O_40_port, n920, O_41_port, n922, O_38_port, n924, O_37_port, n926, 
      O_36_port, n928, O_35_port, n930, O_34_port, n932, O_33_port, n934, 
      O_32_port, n936, O_31_port, n938, O_30_port, n940, O_29_port, n942, 
      O_28_port, n944, O_27_port, n946, O_26_port, n948, O_25_port, n950, 
      O_24_port, n952, O_23_port, n954, O_22_port, n956, O_21_port, n958, 
      O_20_port, n960, O_19_port, n962, O_18_port, n964, O_17_port, n966, 
      O_16_port, n968, O_15_port, n970, O_14_port, n972, O_13_port, n974, 
      O_12_port, n976, O_11_port, n978, O_10_port, n980, n981, O_9_port, n983, 
      n984, n985 : std_logic;

begin
   O <= ( O_41_port, O_40_port, O_39_port, O_38_port, O_37_port, O_36_port, 
      O_35_port, O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, 
      O_29_port, O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, 
      O_23_port, O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, 
      O_17_port, O_16_port, O_15_port, O_14_port, O_13_port, O_12_port, 
      O_11_port, O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, 
      O_4_port, O_3_port, O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(39), A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), 
      A_s(32), A_s(31), A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), 
      A_s(24), A_s(23), A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), 
      A_s(16), A_s(15), A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), 
      A_s(8), A_s(7), A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), 
      X_Logic0_port, X_Logic0_port );
   A_nso <= ( A_ns(39), A_ns(38), A_ns(37), A_ns(36), A_ns(35), A_ns(34), 
      A_ns(33), A_ns(32), A_ns(31), A_ns(30), A_ns(29), A_ns(28), A_ns(27), 
      A_ns(26), A_ns(25), A_ns(24), A_ns(23), A_ns(22), A_ns(21), A_ns(20), 
      A_ns(19), A_ns(18), A_ns(17), A_ns(16), A_ns(15), A_ns(14), A_ns(13), 
      A_ns(12), A_ns(11), A_ns(10), A_ns(9), A_ns(8), A_ns(7), A_ns(6), A_ns(5)
      , A_ns(4), A_ns(3), A_ns(2), A_ns(1), A_ns(0), X_Logic0_port, 
      X_Logic0_port );
   
   X_Logic0_port <= '0';
   U170 : XOR2_X1 port map( A => B(7), B => B(8), Z => n169);
   U2 : CLKBUF_X1 port map( A => n898, Z => n902);
   U3 : BUF_X2 port map( A => n879, Z => n881);
   U4 : CLKBUF_X1 port map( A => n879, Z => n882);
   U5 : BUF_X2 port map( A => n897, Z => n899);
   U6 : CLKBUF_X1 port map( A => n984, Z => n880);
   U7 : CLKBUF_X1 port map( A => n897, Z => n900);
   U8 : BUF_X2 port map( A => n891, Z => n893);
   U9 : BUF_X2 port map( A => n885, Z => n887);
   U10 : CLKBUF_X1 port map( A => n85, Z => n898);
   U11 : CLKBUF_X1 port map( A => n891, Z => n894);
   U12 : CLKBUF_X1 port map( A => n885, Z => n888);
   U13 : CLKBUF_X1 port map( A => n88, Z => n886);
   U14 : CLKBUF_X1 port map( A => n87, Z => n892);
   U15 : BUF_X1 port map( A => n880, Z => n883);
   U16 : BUF_X1 port map( A => n880, Z => n884);
   U17 : BUF_X1 port map( A => n984, Z => n879);
   U18 : BUF_X1 port map( A => n898, Z => n901);
   U19 : INV_X1 port map( A => n102, ZN => O_41_port);
   U20 : BUF_X1 port map( A => n85, Z => n897);
   U21 : INV_X1 port map( A => n168, ZN => n984);
   U22 : BUF_X1 port map( A => n892, Z => n895);
   U23 : BUF_X1 port map( A => n886, Z => n889);
   U24 : BUF_X1 port map( A => n892, Z => n896);
   U25 : BUF_X1 port map( A => n886, Z => n890);
   U26 : INV_X1 port map( A => n143, ZN => n958);
   U27 : AOI22_X1 port map( A1 => A_s(20), A2 => n895, B1 => A_ns(20), B2 => 
                           n889, ZN => n143);
   U28 : INV_X1 port map( A => n164, ZN => O_11_port);
   U29 : AOI221_X1 port map( B1 => n901, B2 => A_ns(10), C1 => n884, C2 => 
                           A_s(10), A => n980, ZN => n164);
   U30 : INV_X1 port map( A => n165, ZN => n980);
   U31 : AOI22_X1 port map( A1 => A_s(9), A2 => n896, B1 => A_ns(9), B2 => n890
                           , ZN => n165);
   U32 : AOI22_X1 port map( A1 => A_s(26), A2 => n894, B1 => A_ns(26), B2 => 
                           n888, ZN => n131);
   U33 : INV_X1 port map( A => n125, ZN => n942);
   U34 : AOI22_X1 port map( A1 => A_s(28), A2 => n894, B1 => A_ns(28), B2 => 
                           n888, ZN => n125);
   U35 : AOI22_X1 port map( A1 => A_s(34), A2 => n893, B1 => A_ns(34), B2 => 
                           n887, ZN => n113);
   U36 : AOI22_X1 port map( A1 => A_s(36), A2 => n893, B1 => A_ns(36), B2 => 
                           n887, ZN => n109);
   U37 : INV_X1 port map( A => n122, ZN => O_31_port);
   U38 : AOI221_X1 port map( B1 => n900, B2 => A_ns(30), C1 => n882, C2 => 
                           A_s(30), A => n940, ZN => n122);
   U39 : INV_X1 port map( A => n136, ZN => O_25_port);
   U40 : INV_X1 port map( A => n144, ZN => O_21_port);
   U41 : INV_X1 port map( A => n114, ZN => O_35_port);
   U42 : AOI221_X1 port map( B1 => n899, B2 => A_ns(34), C1 => n882, C2 => 
                           A_s(34), A => n932, ZN => n114);
   U43 : INV_X1 port map( A => n132, ZN => O_27_port);
   U44 : AOI221_X1 port map( B1 => n900, B2 => A_ns(26), C1 => n882, C2 => 
                           A_s(26), A => n948, ZN => n132);
   U45 : INV_X1 port map( A => n110, ZN => O_37_port);
   U46 : AOI221_X1 port map( B1 => n899, B2 => A_ns(36), C1 => n881, C2 => 
                           A_s(36), A => n928, ZN => n110);
   U47 : INV_X1 port map( A => n111, ZN => n928);
   U48 : INV_X1 port map( A => n128, ZN => O_29_port);
   U49 : AOI221_X1 port map( B1 => n900, B2 => A_ns(28), C1 => n882, C2 => 
                           A_s(28), A => n944, ZN => n128);
   U50 : INV_X1 port map( A => n129, ZN => n944);
   U51 : NAND2_X1 port map( A1 => n169, A2 => n985, ZN => n168);
   U52 : AND2_X1 port map( A1 => n169, A2 => n168, ZN => n85);
   U53 : BUF_X1 port map( A => n88, Z => n885);
   U54 : BUF_X1 port map( A => n87, Z => n891);
   U55 : AOI221_X1 port map( B1 => n896, B2 => A_s(39), C1 => n890, C2 => 
                           A_ns(39), A => n922, ZN => n102);
   U56 : INV_X1 port map( A => n103, ZN => n922);
   U57 : AOI22_X1 port map( A1 => A_ns(40), A2 => n899, B1 => A_s(40), B2 => 
                           n881, ZN => n103);
   U58 : INV_X1 port map( A => n104, ZN => O_40_port);
   U59 : AOI221_X1 port map( B1 => n899, B2 => A_ns(39), C1 => n881, C2 => 
                           A_s(39), A => n920, ZN => n104);
   U60 : INV_X1 port map( A => n105, ZN => n920);
   U61 : AOI22_X1 port map( A1 => A_s(38), A2 => n893, B1 => A_ns(38), B2 => 
                           n887, ZN => n105);
   U62 : INV_X1 port map( A => n112, ZN => O_36_port);
   U63 : AOI221_X1 port map( B1 => n899, B2 => A_ns(35), C1 => n882, C2 => 
                           A_s(35), A => n930, ZN => n112);
   U64 : INV_X1 port map( A => n113, ZN => n930);
   U65 : INV_X1 port map( A => n130, ZN => O_28_port);
   U66 : AOI221_X1 port map( B1 => n900, B2 => A_ns(27), C1 => n882, C2 => 
                           A_s(27), A => n946, ZN => n130);
   U67 : INV_X1 port map( A => n131, ZN => n946);
   U68 : INV_X1 port map( A => n142, ZN => O_22_port);
   U69 : AOI221_X1 port map( B1 => n901, B2 => A_ns(21), C1 => n883, C2 => 
                           A_s(21), A => n958, ZN => n142);
   U70 : INV_X1 port map( A => n108, ZN => O_38_port);
   U71 : AOI221_X1 port map( B1 => n899, B2 => A_ns(37), C1 => n881, C2 => 
                           A_s(37), A => n926, ZN => n108);
   U72 : INV_X1 port map( A => n109, ZN => n926);
   U73 : INV_X1 port map( A => n124, ZN => O_30_port);
   U74 : AOI221_X1 port map( B1 => n900, B2 => A_ns(29), C1 => n882, C2 => 
                           A_s(29), A => n942, ZN => n124);
   U75 : INV_X1 port map( A => n96, ZN => O_8_port);
   U76 : INV_X1 port map( A => n97, ZN => n917);
   U77 : AOI22_X1 port map( A1 => A_s(6), A2 => n893, B1 => A_ns(6), B2 => n887
                           , ZN => n97);
   U78 : INV_X1 port map( A => B(9), ZN => n985);
   U79 : AOI221_X1 port map( B1 => n901, B2 => A_ns(20), C1 => n883, C2 => 
                           A_s(20), A => n960, ZN => n144);
   U80 : INV_X1 port map( A => n145, ZN => n960);
   U81 : AOI22_X1 port map( A1 => A_s(19), A2 => n895, B1 => A_ns(19), B2 => 
                           n889, ZN => n145);
   U82 : INV_X1 port map( A => n162, ZN => O_12_port);
   U83 : AOI221_X1 port map( B1 => n901, B2 => A_ns(11), C1 => n884, C2 => 
                           A_s(11), A => n978, ZN => n162);
   U84 : INV_X1 port map( A => n163, ZN => n978);
   U85 : AOI22_X1 port map( A1 => A_s(10), A2 => n896, B1 => A_ns(10), B2 => 
                           n890, ZN => n163);
   U86 : INV_X1 port map( A => n94, ZN => O_9_port);
   U87 : AOI221_X1 port map( B1 => n899, B2 => A_ns(8), C1 => n881, C2 => 
                           A_s(8), A => n983, ZN => n94);
   U88 : INV_X1 port map( A => n95, ZN => n983);
   U89 : INV_X1 port map( A => n160, ZN => O_13_port);
   U90 : AOI221_X1 port map( B1 => n901, B2 => A_ns(12), C1 => n883, C2 => 
                           A_s(12), A => n976, ZN => n160);
   U91 : INV_X1 port map( A => n161, ZN => n976);
   U92 : AOI22_X1 port map( A1 => A_s(11), A2 => n896, B1 => A_ns(11), B2 => 
                           n890, ZN => n161);
   U93 : NOR3_X1 port map( A1 => B(7), A2 => B(8), A3 => n985, ZN => n88);
   U94 : INV_X1 port map( A => n166, ZN => O_10_port);
   U95 : AOI221_X1 port map( B1 => n899, B2 => A_ns(9), C1 => n881, C2 => 
                           A_s(9), A => n981, ZN => n166);
   U96 : INV_X1 port map( A => n167, ZN => n981);
   U97 : AOI22_X1 port map( A1 => A_s(8), A2 => n893, B1 => A_ns(8), B2 => n887
                           , ZN => n167);
   U98 : INV_X1 port map( A => n158, ZN => O_14_port);
   U99 : AOI221_X1 port map( B1 => n901, B2 => A_ns(13), C1 => n883, C2 => 
                           A_s(13), A => n974, ZN => n158);
   U100 : INV_X1 port map( A => n159, ZN => n974);
   U101 : AOI22_X1 port map( A1 => A_s(12), A2 => n895, B1 => A_ns(12), B2 => 
                           n889, ZN => n159);
   U102 : INV_X1 port map( A => n154, ZN => O_16_port);
   U103 : AOI221_X1 port map( B1 => n901, B2 => A_ns(15), C1 => n883, C2 => 
                           A_s(15), A => n970, ZN => n154);
   U104 : INV_X1 port map( A => n155, ZN => n970);
   U105 : AOI22_X1 port map( A1 => A_s(14), A2 => n895, B1 => A_ns(14), B2 => 
                           n889, ZN => n155);
   U106 : INV_X1 port map( A => n140, ZN => O_23_port);
   U107 : AOI221_X1 port map( B1 => n901, B2 => A_ns(22), C1 => n883, C2 => 
                           A_s(22), A => n956, ZN => n140);
   U108 : INV_X1 port map( A => n141, ZN => n956);
   U109 : AOI22_X1 port map( A1 => A_s(21), A2 => n895, B1 => A_ns(21), B2 => 
                           n889, ZN => n141);
   U110 : INV_X1 port map( A => n148, ZN => O_19_port);
   U111 : AOI221_X1 port map( B1 => n901, B2 => A_ns(18), C1 => n883, C2 => 
                           A_s(18), A => n964, ZN => n148);
   U112 : INV_X1 port map( A => n149, ZN => n964);
   U113 : AOI22_X1 port map( A1 => A_s(17), A2 => n895, B1 => A_ns(17), B2 => 
                           n889, ZN => n149);
   U114 : INV_X1 port map( A => n152, ZN => O_17_port);
   U115 : AOI221_X1 port map( B1 => n901, B2 => A_ns(16), C1 => n883, C2 => 
                           A_s(16), A => n968, ZN => n152);
   U116 : INV_X1 port map( A => n153, ZN => n968);
   U117 : AOI22_X1 port map( A1 => A_s(15), A2 => n895, B1 => A_ns(15), B2 => 
                           n889, ZN => n153);
   U118 : INV_X1 port map( A => n156, ZN => O_15_port);
   U119 : AOI221_X1 port map( B1 => n901, B2 => A_ns(14), C1 => n883, C2 => 
                           A_s(14), A => n972, ZN => n156);
   U120 : INV_X1 port map( A => n157, ZN => n972);
   U121 : AOI22_X1 port map( A1 => A_s(13), A2 => n895, B1 => A_ns(13), B2 => 
                           n889, ZN => n157);
   U122 : INV_X1 port map( A => n150, ZN => O_18_port);
   U123 : AOI221_X1 port map( B1 => n901, B2 => A_ns(17), C1 => n883, C2 => 
                           A_s(17), A => n966, ZN => n150);
   U124 : INV_X1 port map( A => n151, ZN => n966);
   U125 : AOI22_X1 port map( A1 => A_s(16), A2 => n895, B1 => A_ns(16), B2 => 
                           n889, ZN => n151);
   U126 : INV_X1 port map( A => n146, ZN => O_20_port);
   U127 : AOI221_X1 port map( B1 => n901, B2 => A_ns(19), C1 => n883, C2 => 
                           A_s(19), A => n962, ZN => n146);
   U128 : INV_X1 port map( A => n147, ZN => n962);
   U129 : AOI22_X1 port map( A1 => A_s(18), A2 => n895, B1 => A_ns(18), B2 => 
                           n889, ZN => n147);
   U130 : AND3_X1 port map( A1 => B(7), A2 => n985, A3 => B(8), ZN => n87);
   U131 : AOI221_X1 port map( B1 => n900, B2 => A_ns(24), C1 => n883, C2 => 
                           A_s(24), A => n952, ZN => n136);
   U132 : INV_X1 port map( A => n137, ZN => n952);
   U133 : AOI22_X1 port map( A1 => A_s(23), A2 => n895, B1 => A_ns(23), B2 => 
                           n889, ZN => n137);
   U134 : INV_X1 port map( A => n138, ZN => O_24_port);
   U135 : AOI221_X1 port map( B1 => n900, B2 => A_ns(23), C1 => n883, C2 => 
                           A_s(23), A => n954, ZN => n138);
   U136 : INV_X1 port map( A => n139, ZN => n954);
   U137 : AOI22_X1 port map( A1 => A_s(22), A2 => n895, B1 => A_ns(22), B2 => 
                           n889, ZN => n139);
   U138 : INV_X1 port map( A => n134, ZN => O_26_port);
   U139 : AOI221_X1 port map( B1 => n900, B2 => A_ns(25), C1 => n882, C2 => 
                           A_s(25), A => n950, ZN => n134);
   U140 : INV_X1 port map( A => n135, ZN => n950);
   U141 : AOI22_X1 port map( A1 => A_s(24), A2 => n894, B1 => A_ns(24), B2 => 
                           n888, ZN => n135);
   U142 : AOI22_X1 port map( A1 => A_s(27), A2 => n894, B1 => A_ns(27), B2 => 
                           n888, ZN => n129);
   U143 : AOI22_X1 port map( A1 => A_s(35), A2 => n893, B1 => A_ns(35), B2 => 
                           n887, ZN => n111);
   U144 : INV_X1 port map( A => n106, ZN => O_39_port);
   U145 : AOI221_X1 port map( B1 => n899, B2 => A_ns(38), C1 => n881, C2 => 
                           A_s(38), A => n924, ZN => n106);
   U146 : INV_X1 port map( A => n107, ZN => n924);
   U147 : AOI22_X1 port map( A1 => A_s(37), A2 => n893, B1 => A_ns(37), B2 => 
                           n887, ZN => n107);
   U148 : INV_X1 port map( A => n120, ZN => O_32_port);
   U149 : AOI221_X1 port map( B1 => n900, B2 => A_ns(31), C1 => n882, C2 => 
                           A_s(31), A => n938, ZN => n120);
   U150 : INV_X1 port map( A => n121, ZN => n938);
   U151 : AOI22_X1 port map( A1 => A_s(30), A2 => n894, B1 => A_ns(30), B2 => 
                           n888, ZN => n121);
   U152 : INV_X1 port map( A => n133, ZN => n948);
   U153 : AOI22_X1 port map( A1 => A_s(25), A2 => n894, B1 => A_ns(25), B2 => 
                           n888, ZN => n133);
   U154 : INV_X1 port map( A => n123, ZN => n940);
   U155 : AOI22_X1 port map( A1 => A_s(29), A2 => n894, B1 => A_ns(29), B2 => 
                           n888, ZN => n123);
   U156 : INV_X1 port map( A => n115, ZN => n932);
   U157 : AOI22_X1 port map( A1 => A_s(33), A2 => n894, B1 => A_ns(33), B2 => 
                           n888, ZN => n115);
   U158 : INV_X1 port map( A => n118, ZN => O_33_port);
   U159 : AOI221_X1 port map( B1 => n900, B2 => A_ns(32), C1 => n882, C2 => 
                           A_s(32), A => n936, ZN => n118);
   U160 : INV_X1 port map( A => n119, ZN => n936);
   U161 : AOI22_X1 port map( A1 => A_s(31), A2 => n894, B1 => A_ns(31), B2 => 
                           n888, ZN => n119);
   U162 : INV_X1 port map( A => n116, ZN => O_34_port);
   U163 : AOI221_X1 port map( B1 => n900, B2 => A_ns(33), C1 => n882, C2 => 
                           A_s(33), A => n934, ZN => n116);
   U164 : INV_X1 port map( A => n117, ZN => n934);
   U165 : AOI22_X1 port map( A1 => A_s(32), A2 => n894, B1 => A_ns(32), B2 => 
                           n888, ZN => n117);
   U166 : INV_X1 port map( A => n93, ZN => O_1_port);
   U167 : AOI22_X1 port map( A1 => n881, A2 => A_s(0), B1 => n902, B2 => 
                           A_ns(0), ZN => n93);
   U168 : INV_X1 port map( A => n89, ZN => O_5_port);
   U169 : AOI221_X1 port map( B1 => n899, B2 => A_ns(4), C1 => n881, C2 => 
                           A_s(4), A => n911, ZN => n89);
   U171 : INV_X1 port map( A => n90, ZN => n911);
   U172 : AOI22_X1 port map( A1 => A_s(3), A2 => n893, B1 => A_ns(3), B2 => 
                           n887, ZN => n90);
   U173 : INV_X1 port map( A => n126, ZN => O_2_port);
   U174 : AOI221_X1 port map( B1 => n900, B2 => A_ns(1), C1 => n882, C2 => 
                           A_s(1), A => n904, ZN => n126);
   U175 : INV_X1 port map( A => n127, ZN => n904);
   U176 : AOI22_X1 port map( A1 => A_s(0), A2 => n894, B1 => A_ns(0), B2 => 
                           n888, ZN => n127);
   U177 : INV_X1 port map( A => n100, ZN => O_4_port);
   U178 : AOI221_X1 port map( B1 => n899, B2 => A_ns(3), C1 => n881, C2 => 
                           A_s(3), A => n909, ZN => n100);
   U179 : INV_X1 port map( A => n101, ZN => n909);
   U180 : AOI22_X1 port map( A1 => A_s(2), A2 => n893, B1 => A_ns(2), B2 => 
                           n887, ZN => n101);
   U181 : INV_X1 port map( A => n91, ZN => O_3_port);
   U182 : AOI221_X1 port map( B1 => n899, B2 => A_ns(2), C1 => n881, C2 => 
                           A_s(2), A => n907, ZN => n91);
   U183 : INV_X1 port map( A => n92, ZN => n907);
   U184 : AOI22_X1 port map( A1 => A_s(1), A2 => n893, B1 => A_ns(1), B2 => 
                           n887, ZN => n92);
   U185 : INV_X1 port map( A => n84, ZN => O_7_port);
   U186 : AOI221_X1 port map( B1 => n900, B2 => A_ns(6), C1 => n882, C2 => 
                           A_s(6), A => n915, ZN => n84);
   U187 : INV_X1 port map( A => n86, ZN => n915);
   U188 : AOI22_X1 port map( A1 => A_s(5), A2 => n894, B1 => A_ns(5), B2 => 
                           n888, ZN => n86);
   U189 : INV_X1 port map( A => n98, ZN => O_6_port);
   U190 : AOI221_X1 port map( B1 => A_ns(5), B2 => n902, C1 => A_s(5), C2 => 
                           n881, A => n913, ZN => n98);
   U191 : INV_X1 port map( A => n99, ZN => n913);
   U192 : AOI22_X1 port map( A1 => A_s(4), A2 => n893, B1 => A_ns(4), B2 => 
                           n887, ZN => n99);
   U193 : AOI22_X1 port map( A1 => A_s(7), A2 => n893, B1 => A_ns(7), B2 => 
                           n887, ZN => n95);
   U194 : AOI221_X1 port map( B1 => n899, B2 => A_ns(7), C1 => n881, C2 => 
                           A_s(7), A => n917, ZN => n96);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT40_i6 is

   port( A_s, A_ns, B : in std_logic_vector (39 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (39 downto 0));

end BOOTHENC_NBIT40_i6;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT40_i6 is

   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
      n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104
      , n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
      n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, 
      n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, 
      n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, 
      n153, n154, n155, n156, n157, n158, n159, n160, n161, n832, n833, n834, 
      n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, 
      n847, n848, n849, O_2_port, n851, O_1_port, O_3_port, n854, O_4_port, 
      n856, O_5_port, n858, O_6_port, n860, O_37_port, O_38_port, n863, 
      O_39_port, n865, O_36_port, n867, O_35_port, n869, O_34_port, n871, 
      O_33_port, n873, O_32_port, n875, O_31_port, n877, O_30_port, n879, 
      O_29_port, n881, O_28_port, n883, O_27_port, n885, O_26_port, n887, 
      O_25_port, n889, O_24_port, n891, O_23_port, n893, O_22_port, n895, 
      O_21_port, n897, O_20_port, n899, O_19_port, n901, O_18_port, n903, 
      O_17_port, n905, O_16_port, n907, O_15_port, n909, O_14_port, n911, 
      O_13_port, n913, O_12_port, n915, O_11_port, n917, O_10_port, n919, n920,
      O_9_port, O_8_port, n923, O_7_port, n925, n926, n927, n928 : std_logic;

begin
   O <= ( O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, 
      O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, 
      O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, 
      O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, O_16_port, 
      O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, O_10_port, 
      O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, O_3_port, 
      O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   A_nso <= ( A_ns(37), A_ns(36), A_ns(35), A_ns(34), A_ns(33), A_ns(32), 
      A_ns(31), A_ns(30), A_ns(29), A_ns(28), A_ns(27), A_ns(26), A_ns(25), 
      A_ns(24), A_ns(23), A_ns(22), A_ns(21), A_ns(20), A_ns(19), A_ns(18), 
      A_ns(17), A_ns(16), A_ns(15), A_ns(14), A_ns(13), A_ns(12), A_ns(11), 
      A_ns(10), A_ns(9), A_ns(8), A_ns(7), A_ns(6), A_ns(5), A_ns(4), A_ns(3), 
      A_ns(2), A_ns(1), A_ns(0), X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U162 : XOR2_X1 port map( A => B(5), B => B(6), Z => n161);
   U2 : AND2_X1 port map( A1 => n161, A2 => n160, ZN => n81);
   U3 : INV_X1 port map( A => n98, ZN => O_39_port);
   U4 : AOI221_X1 port map( B1 => n846, B2 => A_s(37), C1 => n840, C2 => 
                           A_ns(37), A => n865, ZN => n98);
   U5 : INV_X1 port map( A => n124, ZN => O_27_port);
   U6 : BUF_X2 port map( A => n927, Z => n832);
   U7 : CLKBUF_X1 port map( A => n927, Z => n834);
   U8 : CLKBUF_X1 port map( A => n927, Z => n833);
   U9 : BUF_X2 port map( A => n841, Z => n843);
   U10 : BUF_X2 port map( A => n835, Z => n837);
   U11 : CLKBUF_X1 port map( A => n841, Z => n844);
   U12 : CLKBUF_X1 port map( A => n835, Z => n838);
   U13 : CLKBUF_X1 port map( A => n84, Z => n836);
   U14 : CLKBUF_X1 port map( A => n83, Z => n842);
   U15 : BUF_X2 port map( A => n81, Z => n847);
   U16 : INV_X1 port map( A => n160, ZN => n927);
   U17 : INV_X1 port map( A => n88, ZN => O_9_port);
   U18 : AOI221_X1 port map( B1 => n847, B2 => A_ns(8), C1 => n832, C2 => 
                           A_s(8), A => n923, ZN => n88);
   U19 : INV_X1 port map( A => n89, ZN => n923);
   U20 : AOI22_X1 port map( A1 => A_s(7), A2 => n843, B1 => A_ns(7), B2 => n837
                           , ZN => n89);
   U21 : CLKBUF_X1 port map( A => n81, Z => n849);
   U22 : BUF_X1 port map( A => n842, Z => n845);
   U23 : BUF_X1 port map( A => n836, Z => n839);
   U24 : BUF_X1 port map( A => n842, Z => n846);
   U25 : BUF_X1 port map( A => n836, Z => n840);
   U26 : AOI22_X1 port map( A1 => A_s(36), A2 => n843, B1 => A_ns(36), B2 => 
                           n837, ZN => n101);
   U27 : INV_X1 port map( A => n113, ZN => n877);
   U28 : AOI22_X1 port map( A1 => A_s(30), A2 => n844, B1 => A_ns(30), B2 => 
                           n838, ZN => n113);
   U29 : INV_X1 port map( A => n123, ZN => n885);
   U30 : AOI22_X1 port map( A1 => A_s(26), A2 => n844, B1 => A_ns(26), B2 => 
                           n838, ZN => n123);
   U31 : CLKBUF_X1 port map( A => n81, Z => n848);
   U32 : INV_X1 port map( A => n105, ZN => n869);
   U33 : AOI22_X1 port map( A1 => A_s(34), A2 => n843, B1 => A_ns(34), B2 => 
                           n837, ZN => n105);
   U34 : INV_X1 port map( A => n110, ZN => O_33_port);
   U35 : AOI221_X1 port map( B1 => n847, B2 => A_ns(32), C1 => n833, C2 => 
                           A_s(32), A => n875, ZN => n110);
   U36 : INV_X1 port map( A => n111, ZN => n875);
   U37 : INV_X1 port map( A => n106, ZN => O_35_port);
   U38 : AOI221_X1 port map( B1 => n847, B2 => A_ns(34), C1 => n832, C2 => 
                           A_s(34), A => n871, ZN => n106);
   U39 : INV_X1 port map( A => n120, ZN => O_29_port);
   U40 : AOI221_X1 port map( B1 => n848, B2 => A_ns(28), C1 => n833, C2 => 
                           A_s(28), A => n883, ZN => n120);
   U41 : INV_X1 port map( A => n102, ZN => O_37_port);
   U42 : AOI221_X1 port map( B1 => n847, B2 => A_ns(36), C1 => n832, C2 => 
                           A_s(36), A => n867, ZN => n102);
   U43 : INV_X1 port map( A => n103, ZN => n867);
   U44 : NAND2_X1 port map( A1 => n161, A2 => n928, ZN => n160);
   U45 : INV_X1 port map( A => n100, ZN => O_38_port);
   U46 : AOI221_X1 port map( B1 => n847, B2 => A_ns(37), C1 => n832, C2 => 
                           A_s(37), A => n863, ZN => n100);
   U47 : INV_X1 port map( A => n101, ZN => n863);
   U48 : BUF_X1 port map( A => n84, Z => n835);
   U49 : BUF_X1 port map( A => n83, Z => n841);
   U50 : INV_X1 port map( A => n99, ZN => n865);
   U51 : AOI22_X1 port map( A1 => A_ns(38), A2 => n847, B1 => A_s(38), B2 => 
                           n832, ZN => n99);
   U52 : INV_X1 port map( A => n112, ZN => O_32_port);
   U53 : AOI221_X1 port map( B1 => n848, B2 => A_ns(31), C1 => n833, C2 => 
                           A_s(31), A => n877, ZN => n112);
   U54 : INV_X1 port map( A => n154, ZN => O_12_port);
   U55 : AOI221_X1 port map( B1 => n849, B2 => A_ns(11), C1 => n834, C2 => 
                           A_s(11), A => n917, ZN => n154);
   U56 : INV_X1 port map( A => n155, ZN => n917);
   U57 : AOI22_X1 port map( A1 => A_s(10), A2 => n845, B1 => A_ns(10), B2 => 
                           n839, ZN => n155);
   U58 : NOR3_X1 port map( A1 => B(5), A2 => B(6), A3 => n928, ZN => n84);
   U59 : INV_X1 port map( A => n122, ZN => O_28_port);
   U60 : AOI221_X1 port map( B1 => n848, B2 => A_ns(27), C1 => n833, C2 => 
                           A_s(27), A => n885, ZN => n122);
   U61 : INV_X1 port map( A => n94, ZN => O_6_port);
   U62 : INV_X1 port map( A => n95, ZN => n860);
   U63 : AOI22_X1 port map( A1 => A_s(4), A2 => n843, B1 => A_ns(4), B2 => n837
                           , ZN => n95);
   U64 : INV_X1 port map( A => n158, ZN => O_10_port);
   U65 : AOI221_X1 port map( B1 => n847, B2 => A_ns(9), C1 => n832, C2 => 
                           A_s(9), A => n920, ZN => n158);
   U66 : INV_X1 port map( A => n159, ZN => n920);
   U67 : AOI22_X1 port map( A1 => A_s(8), A2 => n843, B1 => A_ns(8), B2 => n837
                           , ZN => n159);
   U68 : INV_X1 port map( A => n104, ZN => O_36_port);
   U69 : AOI221_X1 port map( B1 => n847, B2 => A_ns(35), C1 => n832, C2 => 
                           A_s(35), A => n869, ZN => n104);
   U70 : INV_X1 port map( A => B(7), ZN => n928);
   U71 : INV_X1 port map( A => n92, ZN => O_7_port);
   U72 : AOI221_X1 port map( B1 => n847, B2 => A_ns(6), C1 => n832, C2 => 
                           A_s(6), A => n926, ZN => n92);
   U73 : INV_X1 port map( A => n93, ZN => n926);
   U74 : INV_X1 port map( A => n156, ZN => O_11_port);
   U75 : AOI221_X1 port map( B1 => n849, B2 => A_ns(10), C1 => n834, C2 => 
                           A_s(10), A => n919, ZN => n156);
   U76 : INV_X1 port map( A => n157, ZN => n919);
   U77 : AOI22_X1 port map( A1 => A_s(9), A2 => n846, B1 => A_ns(9), B2 => n840
                           , ZN => n157);
   U78 : INV_X1 port map( A => n90, ZN => O_8_port);
   U79 : AOI221_X1 port map( B1 => n847, B2 => A_ns(7), C1 => n832, C2 => 
                           A_s(7), A => n925, ZN => n90);
   U80 : INV_X1 port map( A => n91, ZN => n925);
   U81 : AOI22_X1 port map( A1 => A_s(6), A2 => n843, B1 => A_ns(6), B2 => n837
                           , ZN => n91);
   U82 : AND3_X1 port map( A1 => B(5), A2 => n928, A3 => B(6), ZN => n83);
   U83 : INV_X1 port map( A => n130, ZN => O_24_port);
   U84 : AOI221_X1 port map( B1 => n848, B2 => A_ns(23), C1 => n833, C2 => 
                           A_s(23), A => n893, ZN => n130);
   U85 : INV_X1 port map( A => n131, ZN => n893);
   U86 : AOI22_X1 port map( A1 => A_s(22), A2 => n844, B1 => A_ns(22), B2 => 
                           n838, ZN => n131);
   U87 : INV_X1 port map( A => n134, ZN => O_22_port);
   U88 : AOI221_X1 port map( B1 => n848, B2 => A_ns(21), C1 => n834, C2 => 
                           A_s(21), A => n897, ZN => n134);
   U89 : INV_X1 port map( A => n135, ZN => n897);
   U90 : AOI22_X1 port map( A1 => A_s(20), A2 => n845, B1 => A_ns(20), B2 => 
                           n839, ZN => n135);
   U91 : INV_X1 port map( A => n126, ZN => O_26_port);
   U92 : AOI221_X1 port map( B1 => n848, B2 => A_ns(25), C1 => n833, C2 => 
                           A_s(25), A => n889, ZN => n126);
   U93 : INV_X1 port map( A => n127, ZN => n889);
   U94 : AOI22_X1 port map( A1 => A_s(24), A2 => n844, B1 => A_ns(24), B2 => 
                           n838, ZN => n127);
   U95 : INV_X1 port map( A => n136, ZN => O_21_port);
   U96 : AOI221_X1 port map( B1 => n849, B2 => A_ns(20), C1 => n834, C2 => 
                           A_s(20), A => n899, ZN => n136);
   U97 : INV_X1 port map( A => n137, ZN => n899);
   U98 : AOI22_X1 port map( A1 => A_s(19), A2 => n845, B1 => A_ns(19), B2 => 
                           n839, ZN => n137);
   U99 : INV_X1 port map( A => n138, ZN => O_20_port);
   U100 : AOI221_X1 port map( B1 => n849, B2 => A_ns(19), C1 => n834, C2 => 
                           A_s(19), A => n901, ZN => n138);
   U101 : INV_X1 port map( A => n139, ZN => n901);
   U102 : AOI22_X1 port map( A1 => A_s(18), A2 => n845, B1 => A_ns(18), B2 => 
                           n839, ZN => n139);
   U103 : INV_X1 port map( A => n150, ZN => O_14_port);
   U104 : AOI221_X1 port map( B1 => n849, B2 => A_ns(13), C1 => n834, C2 => 
                           A_s(13), A => n913, ZN => n150);
   U105 : INV_X1 port map( A => n151, ZN => n913);
   U106 : AOI22_X1 port map( A1 => A_s(12), A2 => n845, B1 => A_ns(12), B2 => 
                           n839, ZN => n151);
   U107 : INV_X1 port map( A => n146, ZN => O_16_port);
   U108 : AOI221_X1 port map( B1 => n849, B2 => A_ns(15), C1 => n834, C2 => 
                           A_s(15), A => n909, ZN => n146);
   U109 : INV_X1 port map( A => n147, ZN => n909);
   U110 : AOI22_X1 port map( A1 => A_s(14), A2 => n845, B1 => A_ns(14), B2 => 
                           n839, ZN => n147);
   U111 : INV_X1 port map( A => n132, ZN => O_23_port);
   U112 : AOI221_X1 port map( B1 => n848, B2 => A_ns(22), C1 => n834, C2 => 
                           A_s(22), A => n895, ZN => n132);
   U113 : INV_X1 port map( A => n133, ZN => n895);
   U114 : AOI22_X1 port map( A1 => A_s(21), A2 => n845, B1 => A_ns(21), B2 => 
                           n839, ZN => n133);
   U115 : INV_X1 port map( A => n140, ZN => O_19_port);
   U116 : AOI221_X1 port map( B1 => n849, B2 => A_ns(18), C1 => n834, C2 => 
                           A_s(18), A => n903, ZN => n140);
   U117 : INV_X1 port map( A => n141, ZN => n903);
   U118 : AOI22_X1 port map( A1 => A_s(17), A2 => n845, B1 => A_ns(17), B2 => 
                           n839, ZN => n141);
   U119 : INV_X1 port map( A => n128, ZN => O_25_port);
   U120 : AOI221_X1 port map( B1 => n848, B2 => A_ns(24), C1 => n833, C2 => 
                           A_s(24), A => n891, ZN => n128);
   U121 : INV_X1 port map( A => n129, ZN => n891);
   U122 : AOI22_X1 port map( A1 => A_s(23), A2 => n844, B1 => A_ns(23), B2 => 
                           n838, ZN => n129);
   U123 : INV_X1 port map( A => n152, ZN => O_13_port);
   U124 : AOI221_X1 port map( B1 => n849, B2 => A_ns(12), C1 => n834, C2 => 
                           A_s(12), A => n915, ZN => n152);
   U125 : INV_X1 port map( A => n153, ZN => n915);
   U126 : AOI22_X1 port map( A1 => A_s(11), A2 => n845, B1 => A_ns(11), B2 => 
                           n839, ZN => n153);
   U127 : INV_X1 port map( A => n148, ZN => O_15_port);
   U128 : AOI221_X1 port map( B1 => n849, B2 => A_ns(14), C1 => n834, C2 => 
                           A_s(14), A => n911, ZN => n148);
   U129 : INV_X1 port map( A => n149, ZN => n911);
   U130 : AOI22_X1 port map( A1 => A_s(13), A2 => n845, B1 => A_ns(13), B2 => 
                           n839, ZN => n149);
   U131 : INV_X1 port map( A => n144, ZN => O_17_port);
   U132 : AOI221_X1 port map( B1 => n849, B2 => A_ns(16), C1 => n834, C2 => 
                           A_s(16), A => n907, ZN => n144);
   U133 : INV_X1 port map( A => n145, ZN => n907);
   U134 : AOI22_X1 port map( A1 => A_s(15), A2 => n845, B1 => A_ns(15), B2 => 
                           n839, ZN => n145);
   U135 : INV_X1 port map( A => n142, ZN => O_18_port);
   U136 : AOI221_X1 port map( B1 => n849, B2 => A_ns(17), C1 => n834, C2 => 
                           A_s(17), A => n905, ZN => n142);
   U137 : INV_X1 port map( A => n143, ZN => n905);
   U138 : AOI22_X1 port map( A1 => A_s(16), A2 => n845, B1 => A_ns(16), B2 => 
                           n839, ZN => n143);
   U139 : INV_X1 port map( A => n116, ZN => O_30_port);
   U140 : AOI221_X1 port map( B1 => n848, B2 => A_ns(29), C1 => n833, C2 => 
                           A_s(29), A => n881, ZN => n116);
   U141 : INV_X1 port map( A => n117, ZN => n881);
   U142 : AOI22_X1 port map( A1 => A_s(28), A2 => n844, B1 => A_ns(28), B2 => 
                           n838, ZN => n117);
   U143 : AOI22_X1 port map( A1 => A_s(31), A2 => n844, B1 => A_ns(31), B2 => 
                           n838, ZN => n111);
   U144 : AOI22_X1 port map( A1 => A_s(35), A2 => n843, B1 => A_ns(35), B2 => 
                           n837, ZN => n103);
   U145 : INV_X1 port map( A => n108, ZN => O_34_port);
   U146 : AOI221_X1 port map( B1 => n847, B2 => A_ns(33), C1 => n833, C2 => 
                           A_s(33), A => n873, ZN => n108);
   U147 : INV_X1 port map( A => n109, ZN => n873);
   U148 : AOI22_X1 port map( A1 => A_s(32), A2 => n843, B1 => A_ns(32), B2 => 
                           n837, ZN => n109);
   U149 : INV_X1 port map( A => n114, ZN => O_31_port);
   U150 : AOI221_X1 port map( B1 => n848, B2 => A_ns(30), C1 => n833, C2 => 
                           A_s(30), A => n879, ZN => n114);
   U151 : INV_X1 port map( A => n115, ZN => n879);
   U152 : AOI22_X1 port map( A1 => A_s(29), A2 => n844, B1 => A_ns(29), B2 => 
                           n838, ZN => n115);
   U153 : INV_X1 port map( A => n121, ZN => n883);
   U154 : AOI22_X1 port map( A1 => A_s(27), A2 => n844, B1 => A_ns(27), B2 => 
                           n838, ZN => n121);
   U155 : AOI221_X1 port map( B1 => n848, B2 => A_ns(26), C1 => n833, C2 => 
                           A_s(26), A => n887, ZN => n124);
   U156 : INV_X1 port map( A => n125, ZN => n887);
   U157 : AOI22_X1 port map( A1 => A_s(25), A2 => n844, B1 => A_ns(25), B2 => 
                           n838, ZN => n125);
   U158 : INV_X1 port map( A => n107, ZN => n871);
   U159 : AOI22_X1 port map( A1 => A_s(33), A2 => n843, B1 => A_ns(33), B2 => 
                           n837, ZN => n107);
   U160 : INV_X1 port map( A => n96, ZN => O_4_port);
   U161 : AOI221_X1 port map( B1 => A_ns(3), B2 => n849, C1 => A_s(3), C2 => 
                           n832, A => n856, ZN => n96);
   U163 : INV_X1 port map( A => n80, ZN => O_5_port);
   U164 : AOI221_X1 port map( B1 => n848, B2 => A_ns(4), C1 => n833, C2 => 
                           A_s(4), A => n858, ZN => n80);
   U165 : INV_X1 port map( A => n85, ZN => O_3_port);
   U166 : AOI221_X1 port map( B1 => n847, B2 => A_ns(2), C1 => n832, C2 => 
                           A_s(2), A => n854, ZN => n85);
   U167 : INV_X1 port map( A => n86, ZN => n854);
   U168 : INV_X1 port map( A => n87, ZN => O_1_port);
   U169 : AOI22_X1 port map( A1 => n832, A2 => A_s(0), B1 => n849, B2 => 
                           A_ns(0), ZN => n87);
   U170 : INV_X1 port map( A => n118, ZN => O_2_port);
   U171 : AOI221_X1 port map( B1 => n848, B2 => A_ns(1), C1 => n833, C2 => 
                           A_s(1), A => n851, ZN => n118);
   U172 : INV_X1 port map( A => n119, ZN => n851);
   U173 : INV_X1 port map( A => n97, ZN => n856);
   U174 : AOI22_X1 port map( A1 => A_s(2), A2 => n843, B1 => A_ns(2), B2 => 
                           n837, ZN => n97);
   U175 : INV_X1 port map( A => n82, ZN => n858);
   U176 : AOI22_X1 port map( A1 => A_s(3), A2 => n844, B1 => A_ns(3), B2 => 
                           n838, ZN => n82);
   U177 : AOI22_X1 port map( A1 => A_s(0), A2 => n844, B1 => A_ns(0), B2 => 
                           n838, ZN => n119);
   U178 : AOI22_X1 port map( A1 => A_s(1), A2 => n843, B1 => A_ns(1), B2 => 
                           n837, ZN => n86);
   U179 : AOI22_X1 port map( A1 => A_s(5), A2 => n843, B1 => A_ns(5), B2 => 
                           n837, ZN => n93);
   U180 : AOI221_X1 port map( B1 => n847, B2 => A_ns(5), C1 => n832, C2 => 
                           A_s(5), A => n860, ZN => n94);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT38_i4 is

   port( A_s, A_ns, B : in std_logic_vector (37 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (37 downto 0));

end BOOTHENC_NBIT38_i4;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT38_i4 is

   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
      n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, 
      n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, 
      n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, 
      n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, 
      n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, 
      n149, n150, n151, n152, n153, n787, n788, n789, n790, n791, n792, n793, 
      n794, n795, n796, n797, n798, O_2_port, n800, O_1_port, O_3_port, n803, 
      O_4_port, n805, O_35_port, O_36_port, n808, O_37_port, n810, O_34_port, 
      n812, O_33_port, n814, O_32_port, n816, O_31_port, n818, O_30_port, n820,
      O_29_port, n822, O_28_port, n824, O_27_port, n826, O_26_port, n828, 
      O_25_port, n830, O_24_port, n832, O_23_port, n834, O_22_port, n836, 
      O_21_port, n838, O_20_port, n840, O_19_port, n842, O_18_port, n844, 
      O_17_port, n846, O_16_port, n848, O_15_port, n850, O_14_port, n852, 
      O_13_port, n854, O_12_port, n856, O_11_port, n858, O_10_port, n860, n861,
      O_9_port, O_8_port, n864, O_7_port, n866, O_6_port, n868, O_5_port, n870,
      n871, n872, n873 : std_logic;

begin
   O <= ( O_37_port, O_36_port, O_35_port, O_34_port, O_33_port, O_32_port, 
      O_31_port, O_30_port, O_29_port, O_28_port, O_27_port, O_26_port, 
      O_25_port, O_24_port, O_23_port, O_22_port, O_21_port, O_20_port, 
      O_19_port, O_18_port, O_17_port, O_16_port, O_15_port, O_14_port, 
      O_13_port, O_12_port, O_11_port, O_10_port, O_9_port, O_8_port, O_7_port,
      O_6_port, O_5_port, O_4_port, O_3_port, O_2_port, O_1_port, X_Logic0_port
      );
   A_so <= ( A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), A_s(30), A_s(29), 
      A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), A_s(22), A_s(21), 
      A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), A_s(14), A_s(13), 
      A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), A_s(6), A_s(5), A_s(4)
      , A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, X_Logic0_port );
   A_nso <= ( A_ns(35), A_ns(34), A_ns(33), A_ns(32), A_ns(31), A_ns(30), 
      A_ns(29), A_ns(28), A_ns(27), A_ns(26), A_ns(25), A_ns(24), A_ns(23), 
      A_ns(22), A_ns(21), A_ns(20), A_ns(19), A_ns(18), A_ns(17), A_ns(16), 
      A_ns(15), A_ns(14), A_ns(13), A_ns(12), A_ns(11), A_ns(10), A_ns(9), 
      A_ns(8), A_ns(7), A_ns(6), A_ns(5), A_ns(4), A_ns(3), A_ns(2), A_ns(1), 
      A_ns(0), X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U154 : XOR2_X1 port map( A => B(3), B => B(4), Z => n153);
   U2 : INV_X1 port map( A => n84, ZN => O_8_port);
   U3 : AND2_X1 port map( A1 => n153, A2 => n152, ZN => n77);
   U4 : BUF_X2 port map( A => n872, Z => n787);
   U5 : CLKBUF_X1 port map( A => n872, Z => n789);
   U6 : CLKBUF_X1 port map( A => n872, Z => n788);
   U7 : BUF_X2 port map( A => n79, Z => n793);
   U8 : BUF_X2 port map( A => n80, Z => n790);
   U9 : CLKBUF_X1 port map( A => n79, Z => n795);
   U10 : CLKBUF_X1 port map( A => n80, Z => n792);
   U11 : CLKBUF_X1 port map( A => n79, Z => n794);
   U12 : CLKBUF_X1 port map( A => n80, Z => n791);
   U13 : BUF_X2 port map( A => n77, Z => n796);
   U14 : CLKBUF_X1 port map( A => n77, Z => n798);
   U15 : INV_X1 port map( A => n152, ZN => n872);
   U16 : INV_X1 port map( A => n86, ZN => O_7_port);
   U17 : AOI221_X1 port map( B1 => n796, B2 => A_ns(6), C1 => n787, C2 => 
                           A_s(6), A => n868, ZN => n86);
   U18 : INV_X1 port map( A => n87, ZN => n868);
   U19 : AOI22_X1 port map( A1 => A_s(5), A2 => n793, B1 => A_ns(5), B2 => n790
                           , ZN => n87);
   U20 : CLKBUF_X1 port map( A => n77, Z => n797);
   U21 : INV_X1 port map( A => n105, ZN => n818);
   U22 : AOI22_X1 port map( A1 => A_s(30), A2 => n793, B1 => A_ns(30), B2 => 
                           n790, ZN => n105);
   U23 : INV_X1 port map( A => n102, ZN => O_33_port);
   U24 : AOI221_X1 port map( B1 => n796, B2 => A_ns(32), C1 => n788, C2 => 
                           A_s(32), A => n816, ZN => n102);
   U25 : INV_X1 port map( A => n94, ZN => O_37_port);
   U26 : INV_X1 port map( A => n98, ZN => O_35_port);
   U27 : AOI221_X1 port map( B1 => n796, B2 => A_ns(34), C1 => n787, C2 => 
                           A_s(34), A => n812, ZN => n98);
   U28 : NAND2_X1 port map( A1 => n153, A2 => n873, ZN => n152);
   U29 : INV_X1 port map( A => n104, ZN => O_32_port);
   U30 : AOI221_X1 port map( B1 => n796, B2 => A_ns(31), C1 => n788, C2 => 
                           A_s(31), A => n818, ZN => n104);
   U31 : NOR3_X1 port map( A1 => B(3), A2 => B(4), A3 => n873, ZN => n80);
   U32 : AND3_X1 port map( A1 => B(3), A2 => n873, A3 => B(4), ZN => n79);
   U33 : INV_X1 port map( A => n92, ZN => O_4_port);
   U34 : INV_X1 port map( A => n93, ZN => n805);
   U35 : AOI22_X1 port map( A1 => A_s(2), A2 => n793, B1 => A_ns(2), B2 => n790
                           , ZN => n93);
   U36 : INV_X1 port map( A => n90, ZN => O_5_port);
   U37 : AOI221_X1 port map( B1 => n796, B2 => A_ns(4), C1 => n787, C2 => 
                           A_s(4), A => n871, ZN => n90);
   U38 : INV_X1 port map( A => n91, ZN => n871);
   U39 : INV_X1 port map( A => n142, ZN => O_14_port);
   U40 : AOI221_X1 port map( B1 => n798, B2 => A_ns(13), C1 => n789, C2 => 
                           A_s(13), A => n854, ZN => n142);
   U41 : INV_X1 port map( A => n143, ZN => n854);
   U42 : AOI22_X1 port map( A1 => A_s(12), A2 => n795, B1 => A_ns(12), B2 => 
                           n792, ZN => n143);
   U43 : INV_X1 port map( A => B(5), ZN => n873);
   U44 : INV_X1 port map( A => n144, ZN => O_13_port);
   U45 : AOI221_X1 port map( B1 => n798, B2 => A_ns(12), C1 => n789, C2 => 
                           A_s(12), A => n856, ZN => n144);
   U46 : INV_X1 port map( A => n145, ZN => n856);
   U47 : AOI22_X1 port map( A1 => A_s(11), A2 => n795, B1 => A_ns(11), B2 => 
                           n792, ZN => n145);
   U48 : AOI221_X1 port map( B1 => n796, B2 => A_ns(7), C1 => n787, C2 => 
                           A_s(7), A => n866, ZN => n84);
   U49 : INV_X1 port map( A => n85, ZN => n866);
   U50 : AOI22_X1 port map( A1 => A_s(6), A2 => n793, B1 => A_ns(6), B2 => n790
                           , ZN => n85);
   U51 : INV_X1 port map( A => n140, ZN => O_15_port);
   U52 : AOI221_X1 port map( B1 => n798, B2 => A_ns(14), C1 => n789, C2 => 
                           A_s(14), A => n852, ZN => n140);
   U53 : INV_X1 port map( A => n141, ZN => n852);
   U54 : AOI22_X1 port map( A1 => A_s(13), A2 => n795, B1 => A_ns(13), B2 => 
                           n792, ZN => n141);
   U55 : INV_X1 port map( A => n82, ZN => O_9_port);
   U56 : AOI221_X1 port map( B1 => n796, B2 => A_ns(8), C1 => n787, C2 => 
                           A_s(8), A => n864, ZN => n82);
   U57 : INV_X1 port map( A => n83, ZN => n864);
   U58 : AOI22_X1 port map( A1 => A_s(7), A2 => n793, B1 => A_ns(7), B2 => n790
                           , ZN => n83);
   U59 : INV_X1 port map( A => n148, ZN => O_11_port);
   U60 : AOI221_X1 port map( B1 => n798, B2 => A_ns(10), C1 => n789, C2 => 
                           A_s(10), A => n860, ZN => n148);
   U61 : INV_X1 port map( A => n149, ZN => n860);
   U62 : AOI22_X1 port map( A1 => A_s(9), A2 => n795, B1 => A_ns(9), B2 => n792
                           , ZN => n149);
   U63 : INV_X1 port map( A => n138, ZN => O_16_port);
   U64 : AOI221_X1 port map( B1 => n798, B2 => A_ns(15), C1 => n789, C2 => 
                           A_s(15), A => n850, ZN => n138);
   U65 : INV_X1 port map( A => n139, ZN => n850);
   U66 : AOI22_X1 port map( A1 => A_s(14), A2 => n795, B1 => A_ns(14), B2 => 
                           n792, ZN => n139);
   U67 : INV_X1 port map( A => n88, ZN => O_6_port);
   U68 : AOI221_X1 port map( B1 => n796, B2 => A_ns(5), C1 => n787, C2 => 
                           A_s(5), A => n870, ZN => n88);
   U69 : INV_X1 port map( A => n89, ZN => n870);
   U70 : AOI22_X1 port map( A1 => A_s(4), A2 => n793, B1 => A_ns(4), B2 => n790
                           , ZN => n89);
   U71 : INV_X1 port map( A => n150, ZN => O_10_port);
   U72 : AOI221_X1 port map( B1 => n796, B2 => A_ns(9), C1 => n787, C2 => 
                           A_s(9), A => n861, ZN => n150);
   U73 : INV_X1 port map( A => n151, ZN => n861);
   U74 : AOI22_X1 port map( A1 => A_s(8), A2 => n793, B1 => A_ns(8), B2 => n790
                           , ZN => n151);
   U75 : INV_X1 port map( A => n146, ZN => O_12_port);
   U76 : AOI221_X1 port map( B1 => n798, B2 => A_ns(11), C1 => n789, C2 => 
                           A_s(11), A => n858, ZN => n146);
   U77 : INV_X1 port map( A => n147, ZN => n858);
   U78 : AOI22_X1 port map( A1 => A_s(10), A2 => n795, B1 => A_ns(10), B2 => 
                           n792, ZN => n147);
   U79 : INV_X1 port map( A => n106, ZN => O_31_port);
   U80 : AOI221_X1 port map( B1 => n797, B2 => A_ns(30), C1 => n788, C2 => 
                           A_s(30), A => n820, ZN => n106);
   U81 : INV_X1 port map( A => n107, ZN => n820);
   U82 : AOI22_X1 port map( A1 => A_s(29), A2 => n794, B1 => A_ns(29), B2 => 
                           n791, ZN => n107);
   U83 : INV_X1 port map( A => n132, ZN => O_19_port);
   U84 : AOI221_X1 port map( B1 => n798, B2 => A_ns(18), C1 => n789, C2 => 
                           A_s(18), A => n844, ZN => n132);
   U85 : INV_X1 port map( A => n133, ZN => n844);
   U86 : AOI22_X1 port map( A1 => A_s(17), A2 => n795, B1 => A_ns(17), B2 => 
                           n792, ZN => n133);
   U87 : INV_X1 port map( A => n120, ZN => O_25_port);
   U88 : AOI221_X1 port map( B1 => n797, B2 => A_ns(24), C1 => n788, C2 => 
                           A_s(24), A => n832, ZN => n120);
   U89 : INV_X1 port map( A => n121, ZN => n832);
   U90 : AOI22_X1 port map( A1 => A_s(23), A2 => n794, B1 => A_ns(23), B2 => 
                           n791, ZN => n121);
   U91 : INV_X1 port map( A => n114, ZN => O_28_port);
   U92 : AOI221_X1 port map( B1 => n797, B2 => A_ns(27), C1 => n788, C2 => 
                           A_s(27), A => n826, ZN => n114);
   U93 : INV_X1 port map( A => n115, ZN => n826);
   U94 : AOI22_X1 port map( A1 => A_s(26), A2 => n794, B1 => A_ns(26), B2 => 
                           n791, ZN => n115);
   U95 : INV_X1 port map( A => n108, ZN => O_30_port);
   U96 : AOI221_X1 port map( B1 => n797, B2 => A_ns(29), C1 => n788, C2 => 
                           A_s(29), A => n822, ZN => n108);
   U97 : INV_X1 port map( A => n109, ZN => n822);
   U98 : AOI22_X1 port map( A1 => A_s(28), A2 => n794, B1 => A_ns(28), B2 => 
                           n791, ZN => n109);
   U99 : INV_X1 port map( A => n126, ZN => O_22_port);
   U100 : AOI221_X1 port map( B1 => n797, B2 => A_ns(21), C1 => n788, C2 => 
                           A_s(21), A => n838, ZN => n126);
   U101 : INV_X1 port map( A => n127, ZN => n838);
   U102 : AOI22_X1 port map( A1 => A_s(20), A2 => n794, B1 => A_ns(20), B2 => 
                           n791, ZN => n127);
   U103 : INV_X1 port map( A => n128, ZN => O_21_port);
   U104 : AOI221_X1 port map( B1 => n797, B2 => A_ns(20), C1 => n789, C2 => 
                           A_s(20), A => n840, ZN => n128);
   U105 : INV_X1 port map( A => n129, ZN => n840);
   U106 : AOI22_X1 port map( A1 => A_s(19), A2 => n795, B1 => A_ns(19), B2 => 
                           n792, ZN => n129);
   U107 : INV_X1 port map( A => n124, ZN => O_23_port);
   U108 : AOI221_X1 port map( B1 => n797, B2 => A_ns(22), C1 => n788, C2 => 
                           A_s(22), A => n836, ZN => n124);
   U109 : INV_X1 port map( A => n125, ZN => n836);
   U110 : AOI22_X1 port map( A1 => A_s(21), A2 => n794, B1 => A_ns(21), B2 => 
                           n791, ZN => n125);
   U111 : INV_X1 port map( A => n112, ZN => O_29_port);
   U112 : AOI221_X1 port map( B1 => n797, B2 => A_ns(28), C1 => n788, C2 => 
                           A_s(28), A => n824, ZN => n112);
   U113 : INV_X1 port map( A => n113, ZN => n824);
   U114 : AOI22_X1 port map( A1 => A_s(27), A2 => n794, B1 => A_ns(27), B2 => 
                           n791, ZN => n113);
   U115 : INV_X1 port map( A => n116, ZN => O_27_port);
   U116 : AOI221_X1 port map( B1 => n797, B2 => A_ns(26), C1 => n788, C2 => 
                           A_s(26), A => n828, ZN => n116);
   U117 : INV_X1 port map( A => n117, ZN => n828);
   U118 : AOI22_X1 port map( A1 => A_s(25), A2 => n794, B1 => A_ns(25), B2 => 
                           n791, ZN => n117);
   U119 : INV_X1 port map( A => n118, ZN => O_26_port);
   U120 : AOI221_X1 port map( B1 => n797, B2 => A_ns(25), C1 => n788, C2 => 
                           A_s(25), A => n830, ZN => n118);
   U121 : INV_X1 port map( A => n119, ZN => n830);
   U122 : AOI22_X1 port map( A1 => A_s(24), A2 => n794, B1 => A_ns(24), B2 => 
                           n791, ZN => n119);
   U123 : INV_X1 port map( A => n134, ZN => O_18_port);
   U124 : AOI221_X1 port map( B1 => n797, B2 => A_ns(17), C1 => n789, C2 => 
                           A_s(17), A => n846, ZN => n134);
   U125 : INV_X1 port map( A => n135, ZN => n846);
   U126 : AOI22_X1 port map( A1 => A_s(16), A2 => n795, B1 => A_ns(16), B2 => 
                           n792, ZN => n135);
   U127 : INV_X1 port map( A => n136, ZN => O_17_port);
   U128 : AOI221_X1 port map( B1 => n798, B2 => A_ns(16), C1 => n789, C2 => 
                           A_s(16), A => n848, ZN => n136);
   U129 : INV_X1 port map( A => n137, ZN => n848);
   U130 : AOI22_X1 port map( A1 => A_s(15), A2 => n795, B1 => A_ns(15), B2 => 
                           n792, ZN => n137);
   U131 : INV_X1 port map( A => n122, ZN => O_24_port);
   U132 : AOI221_X1 port map( B1 => n797, B2 => A_ns(23), C1 => n788, C2 => 
                           A_s(23), A => n834, ZN => n122);
   U133 : INV_X1 port map( A => n123, ZN => n834);
   U134 : AOI22_X1 port map( A1 => A_s(22), A2 => n794, B1 => A_ns(22), B2 => 
                           n791, ZN => n123);
   U135 : INV_X1 port map( A => n130, ZN => O_20_port);
   U136 : AOI221_X1 port map( B1 => n798, B2 => A_ns(19), C1 => n789, C2 => 
                           A_s(19), A => n842, ZN => n130);
   U137 : INV_X1 port map( A => n131, ZN => n842);
   U138 : AOI22_X1 port map( A1 => A_s(18), A2 => n795, B1 => A_ns(18), B2 => 
                           n792, ZN => n131);
   U139 : INV_X1 port map( A => n96, ZN => O_36_port);
   U140 : AOI221_X1 port map( B1 => n796, B2 => A_ns(35), C1 => n787, C2 => 
                           A_s(35), A => n808, ZN => n96);
   U141 : INV_X1 port map( A => n97, ZN => n808);
   U142 : AOI22_X1 port map( A1 => A_s(34), A2 => n793, B1 => A_ns(34), B2 => 
                           n790, ZN => n97);
   U143 : INV_X1 port map( A => n100, ZN => O_34_port);
   U144 : AOI221_X1 port map( B1 => n796, B2 => A_ns(33), C1 => n787, C2 => 
                           A_s(33), A => n814, ZN => n100);
   U145 : INV_X1 port map( A => n101, ZN => n814);
   U146 : AOI22_X1 port map( A1 => A_s(32), A2 => n793, B1 => A_ns(32), B2 => 
                           n790, ZN => n101);
   U147 : INV_X1 port map( A => n99, ZN => n812);
   U148 : AOI22_X1 port map( A1 => A_s(33), A2 => n793, B1 => A_ns(33), B2 => 
                           n790, ZN => n99);
   U149 : INV_X1 port map( A => n103, ZN => n816);
   U150 : AOI22_X1 port map( A1 => A_s(31), A2 => n793, B1 => A_ns(31), B2 => 
                           n790, ZN => n103);
   U151 : AOI221_X1 port map( B1 => n795, B2 => A_s(35), C1 => n792, C2 => 
                           A_ns(35), A => n810, ZN => n94);
   U152 : INV_X1 port map( A => n95, ZN => n810);
   U153 : AOI22_X1 port map( A1 => A_ns(36), A2 => n796, B1 => A_s(36), B2 => 
                           n787, ZN => n95);
   U155 : INV_X1 port map( A => n81, ZN => O_1_port);
   U156 : AOI22_X1 port map( A1 => n787, A2 => A_s(0), B1 => n798, B2 => 
                           A_ns(0), ZN => n81);
   U157 : INV_X1 port map( A => n110, ZN => O_2_port);
   U158 : AOI221_X1 port map( B1 => A_ns(1), B2 => n798, C1 => A_s(1), C2 => 
                           n787, A => n800, ZN => n110);
   U159 : INV_X1 port map( A => n76, ZN => O_3_port);
   U160 : AOI221_X1 port map( B1 => n797, B2 => A_ns(2), C1 => n788, C2 => 
                           A_s(2), A => n803, ZN => n76);
   U161 : INV_X1 port map( A => n111, ZN => n800);
   U162 : AOI22_X1 port map( A1 => A_s(0), A2 => n794, B1 => A_ns(0), B2 => 
                           n791, ZN => n111);
   U163 : INV_X1 port map( A => n78, ZN => n803);
   U164 : AOI22_X1 port map( A1 => A_s(1), A2 => n794, B1 => A_ns(1), B2 => 
                           n791, ZN => n78);
   U165 : AOI22_X1 port map( A1 => A_s(3), A2 => n793, B1 => A_ns(3), B2 => 
                           n790, ZN => n91);
   U166 : AOI221_X1 port map( B1 => n796, B2 => A_ns(3), C1 => n787, C2 => 
                           A_s(3), A => n805, ZN => n92);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT36_i2 is

   port( A_s, A_ns, B : in std_logic_vector (35 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (35 downto 0));

end BOOTHENC_NBIT36_i2;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT36_i2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X4
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X4
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, O_7_port, O_4_port, O_2_port, O_35_port, O_33_port, 
      O_31_port, O_29_port, O_27_port, O_25_port, O_23_port, O_21_port, 
      O_19_port, O_17_port, O_15_port, O_13_port, O_11_port, O_10_port, 
      O_9_port, O_5_port, n59, n60, n62, n63, n64, n65, n66, n67, n68, n69, n71
      , n72, n73, n74, n75, n76, n77, n78, n79, n80, n82, n83, n84, n85, n86, 
      n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n98, n99, n100, n101, 
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, net262743, 
      net265977, net267111, net267109, net268509, net272336, net273081, 
      net273334, net273346, net273374, n698, O_1_port, n700, n701, n702, n703, 
      n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, 
      n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, 
      n728, n729, n730, n731, n732, n733, n734, A_nso_3_port, O_3_port, n737, 
      A_nso_5_port, n739, A_nso_7_port, n741, A_nso_9_port, n743, A_nso_11_port
      , n745, A_nso_13_port, n747, A_nso_15_port, n749, A_nso_17_port, n751, 
      A_nso_19_port, n753, A_nso_21_port, n755, A_nso_23_port, n757, 
      A_nso_25_port, n759, A_nso_27_port, n761, A_nso_29_port, n763, 
      A_nso_31_port, n765, A_nso_33_port, n767, A_nso_35_port, n769, 
      A_so_5_port, n771, A_so_6_port, n773, A_so_8_port, n775, A_so_10_port, 
      n777, A_so_12_port, n779, A_so_14_port, n781, A_so_16_port, n783, n784, 
      n785, n786, n787, n788, n789, n790, n791, n792, n793, O_34_port, 
      O_32_port, O_30_port, O_28_port, O_26_port, O_24_port, O_22_port, 
      O_20_port, O_18_port, O_16_port, O_14_port, O_12_port, O_8_port, O_6_port
      : std_logic;

begin
   O <= ( O_35_port, O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, 
      O_29_port, O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, 
      O_23_port, O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, 
      O_17_port, O_16_port, O_15_port, O_14_port, O_13_port, O_12_port, 
      O_11_port, O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, 
      O_4_port, O_3_port, O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(33), A_s(32), A_s(31), A_s(30), A_s(29), A_s(28), A_s(27), 
      A_s(26), A_s(25), A_s(24), A_s(23), A_s(22), A_s(21), A_s(20), A_s(19), 
      A_s(18), A_s(17), A_s(16), A_s(15), A_so_16_port, A_s(13), A_so_14_port, 
      A_s(11), A_so_12_port, A_s(9), A_so_10_port, A_s(7), A_so_8_port, A_s(5),
      A_so_6_port, A_so_5_port, A_s(2), net265977, A_s(0), X_Logic0_port, 
      X_Logic0_port );
   A_nso <= ( A_nso_35_port, A_ns(32), A_nso_33_port, A_ns(30), A_nso_31_port, 
      A_ns(28), A_nso_29_port, A_ns(26), A_nso_27_port, A_ns(24), A_nso_25_port
      , A_ns(22), A_nso_23_port, A_ns(20), A_nso_21_port, A_ns(18), 
      A_nso_19_port, A_ns(16), A_nso_17_port, A_ns(14), A_nso_15_port, A_ns(12)
      , A_nso_13_port, A_ns(10), A_nso_11_port, A_ns(8), A_nso_9_port, A_ns(6),
      A_nso_7_port, A_ns(4), A_nso_5_port, net267109, A_nso_3_port, A_ns(0), 
      X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : OR3_X2 port map( A1 => n71, A2 => net272336, A3 => n737, ZN => O_3_port
                           );
   U3 : INV_X1 port map( A => n741, ZN => A_nso_7_port);
   U4 : INV_X1 port map( A => A_ns(0), ZN => n724);
   U5 : NOR2_X1 port map( A1 => net273081, A2 => n723, ZN => n716);
   U6 : INV_X1 port map( A => A_s(0), ZN => n723);
   U7 : NAND2_X1 port map( A1 => n727, A2 => A_ns(0), ZN => n728);
   U8 : NOR2_X1 port map( A1 => B(3), A2 => n722, ZN => n718);
   U9 : INV_X1 port map( A => n739, ZN => A_nso_5_port);
   U10 : AND3_X1 port map( A1 => A_s(1), A2 => B(1), A3 => B(2), ZN => n698);
   U11 : OR2_X1 port map( A1 => n716, A2 => n717, ZN => O_1_port);
   U12 : AOI221_X1 port map( B1 => n710, B2 => A_s(5), C1 => net273346, C2 => 
                           A_ns(4), A => n67, ZN => n66);
   U13 : OAI221_X4 port map( B1 => net273081, B2 => n783, C1 => net262743, C2 
                           => n749, A => n104, ZN => O_15_port);
   U14 : OAI221_X4 port map( B1 => net273081, B2 => n786, C1 => net262743, C2 
                           => n755, A => n94, ZN => O_21_port);
   U15 : OAI221_X4 port map( B1 => net273081, B2 => n784, C1 => net262743, C2 
                           => n751, A => n101, ZN => O_17_port);
   U16 : OAI21_X1 port map( B1 => n730, B2 => n732, A => B(3), ZN => n706);
   U17 : AND2_X1 port map( A1 => A_ns(2), A2 => n700, ZN => n726);
   U18 : XOR2_X1 port map( A => B(2), B => B(1), Z => n700);
   U19 : INV_X1 port map( A => n722, ZN => n701);
   U20 : INV_X1 port map( A => n64, ZN => net268509);
   U21 : BUF_X2 port map( A => net268509, Z => n715);
   U22 : OR2_X1 port map( A1 => net273081, A2 => n773, ZN => n702);
   U23 : OR2_X1 port map( A1 => net262743, A2 => n739, ZN => n703);
   U24 : NAND3_X1 port map( A1 => n702, A2 => n703, A3 => n68, ZN => O_5_port);
   U25 : NAND2_X1 port map( A1 => n733, A2 => n704, ZN => n705);
   U26 : NAND2_X1 port map( A1 => n705, A2 => n706, ZN => n734);
   U27 : INV_X1 port map( A => B(3), ZN => n704);
   U28 : NOR2_X1 port map( A1 => B(3), A2 => n719, ZN => net273374);
   U29 : INV_X1 port map( A => n739, ZN => n707);
   U30 : CLKBUF_X1 port map( A => n725, Z => n708);
   U31 : INV_X1 port map( A => net273374, ZN => n709);
   U32 : INV_X2 port map( A => n709, ZN => n710);
   U33 : XOR2_X1 port map( A => B(2), B => B(1), Z => n711);
   U34 : XNOR2_X1 port map( A => B(2), B => B(1), ZN => n712);
   U35 : AND2_X4 port map( A1 => n718, A2 => B(2), ZN => n713);
   U36 : INV_X2 port map( A => n713, ZN => n63);
   U37 : CLKBUF_X1 port map( A => A_ns(2), Z => n714);
   U38 : NOR2_X1 port map( A1 => B(2), A2 => n701, ZN => n727);
   U39 : NOR2_X1 port map( A1 => B(2), A2 => B(1), ZN => n720);
   U40 : INV_X1 port map( A => B(1), ZN => n722);
   U41 : NAND2_X1 port map( A1 => n711, A2 => B(3), ZN => n64);
   U42 : NOR2_X1 port map( A1 => n724, A2 => net273334, ZN => n717);
   U43 : OR2_X2 port map( A1 => B(3), A2 => n712, ZN => net273081);
   U44 : NAND2_X2 port map( A1 => n720, A2 => B(3), ZN => net262743);
   U45 : MUX2_X1 port map( A => n698, B => n726, S => B(3), Z => n71);
   U46 : INV_X2 port map( A => net262743, ZN => net273346);
   U47 : NAND3_X1 port map( A1 => B(2), A2 => n701, A3 => A_s(0), ZN => n729);
   U48 : MUX2_X1 port map( A => n729, B => n728, S => B(3), Z => n721);
   U49 : INV_X1 port map( A => n730, ZN => A_nso_3_port);
   U50 : INV_X1 port map( A => A_s(1), ZN => n725);
   U51 : INV_X1 port map( A => n708, ZN => net265977);
   U52 : XNOR2_X1 port map( A => B(2), B => B(1), ZN => n719);
   U53 : NOR2_X1 port map( A1 => net262743, A2 => n730, ZN => net272336);
   U54 : INV_X1 port map( A => A_ns(1), ZN => n730);
   U55 : XNOR2_X1 port map( A => B(2), B => B(1), ZN => n731);
   U56 : XNOR2_X1 port map( A => B(2), B => B(1), ZN => n732);
   U57 : NAND2_X1 port map( A1 => n734, A2 => n721, ZN => O_2_port);
   U58 : OR2_X1 port map( A1 => n731, A2 => n725, ZN => n733);
   U59 : OAI221_X1 port map( B1 => net273081, B2 => n792, C1 => net262743, C2 
                           => n767, A => n75, ZN => O_33_port);
   U60 : OAI221_X1 port map( B1 => net273081, B2 => n790, C1 => net262743, C2 
                           => n763, A => n82, ZN => O_29_port);
   U61 : OAI221_X1 port map( B1 => net273081, B2 => n789, C1 => net262743, C2 
                           => n761, A => n85, ZN => O_27_port);
   U62 : OAI221_X1 port map( B1 => net273081, B2 => n791, C1 => net262743, C2 
                           => n765, A => n78, ZN => O_31_port);
   U63 : OAI221_X1 port map( B1 => net273081, B2 => n788, C1 => net262743, C2 
                           => n759, A => n88, ZN => O_25_port);
   U64 : OAI221_X1 port map( B1 => net273081, B2 => n793, C1 => net262743, C2 
                           => n769, A => n72, ZN => O_35_port);
   U65 : CLKBUF_X3 port map( A => n64, Z => net273334);
   U66 : AOI221_X4 port map( B1 => n710, B2 => A_s(11), C1 => net273346, C2 => 
                           A_ns(10), A => n109, ZN => n108);
   U67 : AND2_X1 port map( A1 => net273374, A2 => A_s(2), ZN => n737);
   U68 : AOI221_X4 port map( B1 => n710, B2 => A_s(7), C1 => net273346, C2 => 
                           A_ns(6), A => n62, ZN => n60);
   U69 : AOI221_X4 port map( B1 => n710, B2 => A_s(19), C1 => net273346, C2 => 
                           A_ns(18), A => n96, ZN => n95);
   U70 : AOI221_X4 port map( B1 => n710, B2 => A_s(17), C1 => net273346, C2 => 
                           A_ns(16), A => n100, ZN => n99);
   U71 : AOI221_X4 port map( B1 => n710, B2 => A_s(15), C1 => net273346, C2 => 
                           A_ns(14), A => n103, ZN => n102);
   U72 : AOI221_X4 port map( B1 => n710, B2 => A_s(13), C1 => net273346, C2 => 
                           A_ns(12), A => n106, ZN => n105);
   U73 : AOI221_X4 port map( B1 => n710, B2 => A_s(33), C1 => net273346, C2 => 
                           A_ns(32), A => n74, ZN => n73);
   U74 : AOI221_X4 port map( B1 => n710, B2 => A_s(31), C1 => net273346, C2 => 
                           A_ns(30), A => n77, ZN => n76);
   U75 : AOI221_X4 port map( B1 => n710, B2 => A_s(29), C1 => net273346, C2 => 
                           A_ns(28), A => n80, ZN => n79);
   U76 : AOI221_X4 port map( B1 => n710, B2 => A_s(27), C1 => net273346, C2 => 
                           A_ns(26), A => n84, ZN => n83);
   U77 : AOI221_X4 port map( B1 => n710, B2 => A_s(23), C1 => net273346, C2 => 
                           A_ns(22), A => n90, ZN => n89);
   U78 : AOI221_X4 port map( B1 => n710, B2 => A_s(21), C1 => net273346, C2 => 
                           A_ns(20), A => n93, ZN => n92);
   U79 : AOI221_X4 port map( B1 => n710, B2 => A_s(25), C1 => net273346, C2 => 
                           A_ns(24), A => n87, ZN => n86);
   U80 : INV_X1 port map( A => A_ns(33), ZN => n769);
   U81 : INV_X1 port map( A => n76, ZN => O_32_port);
   U82 : INV_X1 port map( A => n714, ZN => net267111);
   U83 : INV_X1 port map( A => A_ns(15), ZN => n751);
   U84 : INV_X1 port map( A => A_ns(11), ZN => n747);
   U85 : INV_X1 port map( A => A_ns(7), ZN => n743);
   U86 : INV_X1 port map( A => A_ns(5), ZN => n741);
   U87 : INV_X1 port map( A => A_ns(13), ZN => n749);
   U88 : INV_X1 port map( A => A_ns(17), ZN => n753);
   U89 : INV_X1 port map( A => A_ns(9), ZN => n745);
   U90 : INV_X1 port map( A => A_ns(31), ZN => n767);
   U91 : INV_X1 port map( A => A_ns(23), ZN => n759);
   U92 : INV_X1 port map( A => A_ns(27), ZN => n763);
   U93 : INV_X1 port map( A => A_ns(19), ZN => n755);
   U94 : INV_X1 port map( A => A_ns(21), ZN => n757);
   U95 : INV_X1 port map( A => A_ns(25), ZN => n761);
   U96 : INV_X1 port map( A => A_ns(29), ZN => n765);
   U97 : OAI221_X1 port map( B1 => net273081, B2 => n771, C1 => net262743, C2 
                           => net267111, A => n69, ZN => O_4_port);
   U98 : OAI221_X1 port map( B1 => net273081, B2 => n777, C1 => net262743, C2 
                           => n743, A => n59, ZN => O_9_port);
   U99 : INV_X1 port map( A => n108, ZN => O_12_port);
   U100 : INV_X1 port map( A => n105, ZN => O_14_port);
   U101 : INV_X1 port map( A => n102, ZN => O_16_port);
   U102 : INV_X1 port map( A => n99, ZN => O_18_port);
   U103 : INV_X1 port map( A => n60, ZN => O_8_port);
   U104 : INV_X1 port map( A => n66, ZN => O_6_port);
   U105 : INV_X1 port map( A => A_s(8), ZN => n777);
   U106 : INV_X1 port map( A => A_s(4), ZN => n773);
   U107 : INV_X1 port map( A => A_s(6), ZN => n775);
   U108 : OAI221_X1 port map( B1 => n777, B2 => n63, C1 => net273334, C2 => 
                           n745, A => n111, ZN => O_10_port);
   U109 : OAI221_X1 port map( B1 => net273081, B2 => n775, C1 => net262743, C2 
                           => n741, A => n65, ZN => O_7_port);
   U110 : OAI221_X1 port map( B1 => net273081, B2 => n779, C1 => net262743, C2 
                           => n745, A => n110, ZN => O_11_port);
   U111 : INV_X1 port map( A => n73, ZN => O_34_port);
   U112 : INV_X1 port map( A => n79, ZN => O_30_port);
   U113 : INV_X1 port map( A => n89, ZN => O_24_port);
   U114 : INV_X1 port map( A => n86, ZN => O_26_port);
   U115 : INV_X1 port map( A => n95, ZN => O_20_port);
   U116 : INV_X1 port map( A => n83, ZN => O_28_port);
   U117 : INV_X1 port map( A => n92, ZN => O_22_port);
   U118 : INV_X1 port map( A => A_s(10), ZN => n779);
   U119 : INV_X1 port map( A => A_s(12), ZN => n781);
   U120 : INV_X1 port map( A => A_s(14), ZN => n783);
   U121 : INV_X1 port map( A => A_s(16), ZN => n784);
   U122 : INV_X1 port map( A => A_s(20), ZN => n786);
   U123 : INV_X1 port map( A => A_s(24), ZN => n788);
   U124 : INV_X1 port map( A => A_s(18), ZN => n785);
   U125 : INV_X1 port map( A => A_s(22), ZN => n787);
   U126 : INV_X1 port map( A => A_s(26), ZN => n789);
   U127 : INV_X1 port map( A => A_s(28), ZN => n790);
   U128 : INV_X1 port map( A => A_s(30), ZN => n791);
   U129 : INV_X1 port map( A => A_s(32), ZN => n792);
   U130 : OAI221_X1 port map( B1 => net273081, B2 => n787, C1 => net262743, C2 
                           => n757, A => n91, ZN => O_23_port);
   U131 : OAI221_X1 port map( B1 => net273081, B2 => n785, C1 => net262743, C2 
                           => n753, A => n98, ZN => O_19_port);
   U132 : OAI221_X1 port map( B1 => net273081, B2 => n781, C1 => net262743, C2 
                           => n747, A => n107, ZN => O_13_port);
   U133 : AOI22_X1 port map( A1 => A_s(9), A2 => n710, B1 => A_ns(8), B2 => 
                           net273346, ZN => n111);
   U134 : OAI22_X1 port map( A1 => n792, A2 => n63, B1 => n769, B2 => net273334
                           , ZN => n74);
   U135 : OAI22_X1 port map( A1 => n791, A2 => n63, B1 => n767, B2 => net273334
                           , ZN => n77);
   U136 : OAI22_X1 port map( A1 => n790, A2 => n63, B1 => n765, B2 => net273334
                           , ZN => n80);
   U137 : OAI22_X1 port map( A1 => n789, A2 => n63, B1 => n763, B2 => net273334
                           , ZN => n84);
   U138 : OAI22_X1 port map( A1 => n788, A2 => n63, B1 => n761, B2 => net273334
                           , ZN => n87);
   U139 : OAI22_X1 port map( A1 => n787, A2 => n63, B1 => n759, B2 => net273334
                           , ZN => n90);
   U140 : OAI22_X1 port map( A1 => n786, A2 => n63, B1 => n757, B2 => net273334
                           , ZN => n93);
   U141 : OAI22_X1 port map( A1 => n785, A2 => n63, B1 => n755, B2 => net273334
                           , ZN => n96);
   U142 : OAI22_X1 port map( A1 => n784, A2 => n63, B1 => n753, B2 => net273334
                           , ZN => n100);
   U143 : OAI22_X1 port map( A1 => n783, A2 => n63, B1 => n751, B2 => net273334
                           , ZN => n103);
   U144 : OAI22_X1 port map( A1 => n781, A2 => n63, B1 => n749, B2 => net273334
                           , ZN => n106);
   U145 : OAI22_X1 port map( A1 => n779, A2 => n63, B1 => n747, B2 => net273334
                           , ZN => n109);
   U146 : OAI22_X1 port map( A1 => n775, A2 => n63, B1 => net273334, B2 => n743
                           , ZN => n62);
   U147 : OAI22_X1 port map( A1 => n773, A2 => n63, B1 => n741, B2 => n64, ZN 
                           => n67);
   U148 : AOI22_X1 port map( A1 => A_s(33), A2 => n713, B1 => A_ns(34), B2 => 
                           net268509, ZN => n72);
   U149 : AOI22_X1 port map( A1 => A_s(31), A2 => n713, B1 => A_ns(32), B2 => 
                           net268509, ZN => n75);
   U150 : AOI22_X1 port map( A1 => A_s(29), A2 => n713, B1 => A_ns(30), B2 => 
                           n715, ZN => n78);
   U151 : AOI22_X1 port map( A1 => A_s(27), A2 => n713, B1 => A_ns(28), B2 => 
                           net268509, ZN => n82);
   U152 : AOI22_X1 port map( A1 => A_s(25), A2 => n713, B1 => A_ns(26), B2 => 
                           net268509, ZN => n85);
   U153 : AOI22_X1 port map( A1 => A_s(23), A2 => n713, B1 => A_ns(24), B2 => 
                           n715, ZN => n88);
   U154 : AOI22_X1 port map( A1 => A_s(21), A2 => n713, B1 => A_ns(22), B2 => 
                           n715, ZN => n91);
   U155 : AOI22_X1 port map( A1 => A_s(19), A2 => n713, B1 => A_ns(20), B2 => 
                           n715, ZN => n94);
   U156 : AOI22_X1 port map( A1 => A_s(17), A2 => n713, B1 => A_ns(18), B2 => 
                           n715, ZN => n98);
   U157 : AOI22_X1 port map( A1 => A_s(15), A2 => n713, B1 => A_ns(16), B2 => 
                           n715, ZN => n101);
   U158 : AOI22_X1 port map( A1 => A_s(13), A2 => n713, B1 => A_ns(14), B2 => 
                           n715, ZN => n104);
   U159 : AOI22_X1 port map( A1 => A_s(11), A2 => n713, B1 => A_ns(12), B2 => 
                           n715, ZN => n107);
   U160 : AOI22_X1 port map( A1 => A_s(9), A2 => n713, B1 => A_ns(10), B2 => 
                           n715, ZN => n110);
   U161 : AOI22_X1 port map( A1 => A_s(7), A2 => n713, B1 => A_ns(8), B2 => 
                           n715, ZN => n59);
   U162 : AOI22_X1 port map( A1 => A_s(5), A2 => n713, B1 => A_ns(6), B2 => 
                           n715, ZN => n65);
   U163 : AOI22_X1 port map( A1 => A_so_5_port, A2 => n713, B1 => A_ns(4), B2 
                           => n715, ZN => n68);
   U164 : AOI22_X1 port map( A1 => A_s(2), A2 => n713, B1 => n707, B2 => 
                           net268509, ZN => n69);
   U165 : INV_X1 port map( A => net267111, ZN => net267109);
   U166 : INV_X1 port map( A => A_ns(3), ZN => n739);
   U167 : INV_X1 port map( A => n743, ZN => A_nso_9_port);
   U168 : INV_X1 port map( A => n745, ZN => A_nso_11_port);
   U169 : INV_X1 port map( A => n747, ZN => A_nso_13_port);
   U170 : INV_X1 port map( A => n749, ZN => A_nso_15_port);
   U171 : INV_X1 port map( A => n751, ZN => A_nso_17_port);
   U172 : INV_X1 port map( A => n753, ZN => A_nso_19_port);
   U173 : INV_X1 port map( A => n755, ZN => A_nso_21_port);
   U174 : INV_X1 port map( A => n757, ZN => A_nso_23_port);
   U175 : INV_X1 port map( A => n759, ZN => A_nso_25_port);
   U176 : INV_X1 port map( A => n761, ZN => A_nso_27_port);
   U177 : INV_X1 port map( A => n763, ZN => A_nso_29_port);
   U178 : INV_X1 port map( A => n765, ZN => A_nso_31_port);
   U179 : INV_X1 port map( A => n767, ZN => A_nso_33_port);
   U180 : INV_X1 port map( A => n769, ZN => A_nso_35_port);
   U181 : INV_X1 port map( A => n771, ZN => A_so_5_port);
   U182 : INV_X1 port map( A => A_s(3), ZN => n771);
   U183 : INV_X1 port map( A => n773, ZN => A_so_6_port);
   U184 : INV_X1 port map( A => n775, ZN => A_so_8_port);
   U185 : INV_X1 port map( A => n777, ZN => A_so_10_port);
   U186 : INV_X1 port map( A => n779, ZN => A_so_12_port);
   U187 : INV_X1 port map( A => n781, ZN => A_so_14_port);
   U188 : INV_X1 port map( A => n783, ZN => A_so_16_port);
   U189 : INV_X1 port map( A => A_s(34), ZN => n793);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT34_i0 is

   port( A_s, A_ns, B : in std_logic_vector (33 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (33 downto 0));

end BOOTHENC_NBIT34_i0;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT34_i0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X4
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, n41, n42, n43, n44, n45, n46, n47, n49, n50, n51, n53,
      n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68
      , n69, n70, n71, n72, n73, net267007, net267041, net267119, net267125, 
      net267123, net267121, net267131, net267129, net267127, net268556, 
      net278130, net278161, n52, n40, n429, n430, n431, n432, n433, n434, n435,
      A_nso_6_port, n437, n438, A_nso_8_port, n440, n441, A_nso_10_port, n443, 
      n444, A_nso_12_port, n446, n447, A_nso_14_port, n449, n450, A_nso_16_port
      , n452, n453, A_nso_18_port, n455, n456, A_nso_20_port, n458, n459, 
      A_nso_22_port, n461, n462, A_nso_24_port, n464, n465, A_nso_26_port, n467
      , n468, A_nso_28_port, n470, n471, A_nso_30_port, n473, n474, 
      A_nso_32_port, n476, n477, n478, n479, n480, n481 : std_logic;

begin
   A_so <= ( A_s(32), A_s(31), A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), 
      A_s(25), A_s(24), A_s(23), A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), 
      A_s(17), A_s(16), A_s(15), A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), 
      A_s(9), A_s(8), A_s(7), A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), 
      A_s(0), X_Logic0_port );
   A_nso <= ( A_ns(32), A_nso_32_port, A_ns(30), A_nso_30_port, A_ns(28), 
      A_nso_28_port, A_ns(26), A_nso_26_port, A_ns(24), A_nso_24_port, A_ns(22)
      , A_nso_22_port, A_ns(20), A_nso_20_port, A_ns(18), A_nso_18_port, 
      A_ns(16), A_nso_16_port, A_ns(14), A_nso_14_port, A_ns(12), A_nso_12_port
      , A_ns(10), A_nso_10_port, A_ns(8), A_nso_8_port, A_ns(6), A_nso_6_port, 
      A_ns(4), net278130, A_ns(2), A_ns(1), A_ns(0), X_Logic0_port );
   
   X_Logic0_port <= '0';
   U3 : OAI221_X1 port map( B1 => net267119, B2 => n459, C1 => net267123, C2 =>
                           n461, A => n61, ZN => O(21));
   U4 : OAI221_X1 port map( B1 => net267119, B2 => n461, C1 => net267123, C2 =>
                           n462, A => n60, ZN => O(22));
   U5 : OAI221_X1 port map( B1 => net267119, B2 => n449, C1 => net267125, C2 =>
                           n450, A => n69, ZN => O(14));
   U6 : OAI221_X1 port map( B1 => net267119, B2 => n467, C1 => net267123, C2 =>
                           n468, A => n56, ZN => O(26));
   U7 : OAI221_X1 port map( B1 => net267119, B2 => n470, C1 => net267123, C2 =>
                           n471, A => n54, ZN => O(28));
   U8 : INV_X1 port map( A => A_ns(29), ZN => n473);
   U9 : OR2_X1 port map( A1 => n431, A2 => B(0), ZN => n429);
   U10 : INV_X1 port map( A => A_ns(3), ZN => n430);
   U11 : CLKBUF_X3 port map( A => A_ns(3), Z => net278130);
   U12 : OAI221_X4 port map( B1 => net267119, B2 => n443, C1 => net267121, C2 
                           => n444, A => n73, ZN => O(10));
   U13 : BUF_X4 port map( A => n429, Z => net267119);
   U14 : OAI221_X1 port map( B1 => n433, B2 => n429, C1 => n432, C2 => 
                           net267121, A => n52, ZN => O(2));
   U15 : NAND2_X1 port map( A1 => A_s(2), A2 => n435, ZN => n52);
   U16 : CLKBUF_X3 port map( A => n40, Z => net267121);
   U17 : INV_X1 port map( A => A_ns(2), ZN => n432);
   U18 : CLKBUF_X1 port map( A => n432, Z => n434);
   U19 : OAI221_X1 port map( B1 => n429, B2 => net267041, C1 => net267121, C2 
                           => net267007, A => n46, ZN => O(4));
   U20 : OAI221_X1 port map( B1 => n429, B2 => n434, C1 => n430, C2 => 
                           net267121, A => n47, ZN => O(3));
   U21 : INV_X1 port map( A => B(1), ZN => n431);
   U22 : AND2_X1 port map( A1 => B(0), A2 => n431, ZN => n435);
   U23 : INV_X1 port map( A => A_ns(1), ZN => n433);
   U24 : CLKBUF_X1 port map( A => n433, Z => net278161);
   U25 : CLKBUF_X1 port map( A => n435, Z => net267129);
   U26 : CLKBUF_X1 port map( A => n435, Z => net267131);
   U27 : CLKBUF_X3 port map( A => n435, Z => net267127);
   U28 : NAND2_X1 port map( A1 => B(1), A2 => B(0), ZN => n40);
   U29 : CLKBUF_X1 port map( A => n40, Z => net267123);
   U30 : CLKBUF_X1 port map( A => n40, Z => net267125);
   U31 : OAI221_X4 port map( B1 => net267119, B2 => n464, C1 => net267123, C2 
                           => n465, A => n58, ZN => O(24));
   U32 : OAI221_X1 port map( B1 => net267119, B2 => n476, C1 => net267121, C2 
                           => n477, A => n49, ZN => O(32));
   U33 : INV_X1 port map( A => A_ns(32), ZN => n477);
   U34 : INV_X1 port map( A => A_ns(31), ZN => n476);
   U35 : OAI22_X1 port map( A1 => net268556, A2 => n480, B1 => net267121, B2 =>
                           n479, ZN => O(0));
   U36 : INV_X1 port map( A => A_ns(0), ZN => n479);
   U37 : OAI221_X1 port map( B1 => net267119, B2 => n446, C1 => net267125, C2 
                           => n447, A => n71, ZN => O(12));
   U38 : NAND2_X1 port map( A1 => A_s(12), A2 => net267127, ZN => n71);
   U39 : OAI221_X1 port map( B1 => net267119, B2 => n444, C1 => net267125, C2 
                           => n446, A => n72, ZN => O(11));
   U40 : NAND2_X1 port map( A1 => A_s(11), A2 => net267127, ZN => n72);
   U41 : NAND2_X1 port map( A1 => A_s(14), A2 => net267127, ZN => n69);
   U42 : OAI221_X1 port map( B1 => net267119, B2 => n441, C1 => net267123, C2 
                           => n443, A => n41, ZN => O(9));
   U43 : NAND2_X1 port map( A1 => A_s(9), A2 => net267127, ZN => n41);
   U44 : OAI221_X1 port map( B1 => net267119, B2 => n438, C1 => net267121, C2 
                           => n440, A => n43, ZN => O(7));
   U45 : NAND2_X1 port map( A1 => A_s(7), A2 => net267127, ZN => n43);
   U46 : OAI221_X1 port map( B1 => net267119, B2 => n455, C1 => net267125, C2 
                           => n456, A => n65, ZN => O(18));
   U47 : NAND2_X1 port map( A1 => A_s(18), A2 => net267127, ZN => n65);
   U48 : OAI221_X1 port map( B1 => net267119, B2 => net267007, C1 => net267121,
                           C2 => n437, A => n45, ZN => O(5));
   U49 : NAND2_X1 port map( A1 => A_s(5), A2 => net267129, ZN => n45);
   U50 : OAI221_X1 port map( B1 => net267119, B2 => n440, C1 => n441, C2 => 
                           net267121, A => n42, ZN => O(8));
   U51 : NAND2_X1 port map( A1 => A_s(8), A2 => net267127, ZN => n42);
   U52 : NAND2_X1 port map( A1 => A_s(10), A2 => net267127, ZN => n73);
   U53 : OAI221_X1 port map( B1 => net267119, B2 => n437, C1 => net267121, C2 
                           => n438, A => n44, ZN => O(6));
   U54 : NAND2_X1 port map( A1 => A_s(6), A2 => net267127, ZN => n44);
   U55 : OAI221_X1 port map( B1 => net267119, B2 => n456, C1 => net267123, C2 
                           => n458, A => n64, ZN => O(19));
   U56 : NAND2_X1 port map( A1 => A_s(19), A2 => net267127, ZN => n64);
   U57 : OAI221_X1 port map( B1 => net267119, B2 => n453, C1 => net267125, C2 
                           => n455, A => n66, ZN => O(17));
   U58 : NAND2_X1 port map( A1 => A_s(17), A2 => net267127, ZN => n66);
   U59 : NAND2_X1 port map( A1 => A_s(4), A2 => net267131, ZN => n46);
   U60 : OAI221_X1 port map( B1 => net267119, B2 => n447, C1 => net267125, C2 
                           => n449, A => n70, ZN => O(13));
   U61 : NAND2_X1 port map( A1 => A_s(13), A2 => net267127, ZN => n70);
   U62 : OAI221_X1 port map( B1 => net267119, B2 => n450, C1 => net267125, C2 
                           => n452, A => n68, ZN => O(15));
   U63 : NAND2_X1 port map( A1 => A_s(15), A2 => net267127, ZN => n68);
   U64 : OAI221_X1 port map( B1 => net267119, B2 => n452, C1 => net267125, C2 
                           => n453, A => n67, ZN => O(16));
   U65 : NAND2_X1 port map( A1 => A_s(16), A2 => net267127, ZN => n67);
   U66 : NAND2_X1 port map( A1 => A_s(3), A2 => net267131, ZN => n47);
   U67 : INV_X1 port map( A => A_ns(19), ZN => n458);
   U68 : INV_X1 port map( A => A_ns(5), ZN => n437);
   U69 : INV_X1 port map( A => A_ns(7), ZN => n440);
   U70 : INV_X1 port map( A => A_ns(3), ZN => net267041);
   U71 : INV_X1 port map( A => A_ns(9), ZN => n443);
   U72 : INV_X1 port map( A => A_ns(11), ZN => n446);
   U73 : INV_X1 port map( A => A_ns(13), ZN => n449);
   U74 : INV_X1 port map( A => A_ns(17), ZN => n455);
   U75 : INV_X1 port map( A => A_ns(15), ZN => n452);
   U76 : OAI222_X1 port map( A1 => n481, A2 => net268556, B1 => n477, B2 => 
                           net267119, C1 => n478, C2 => net267121, ZN => O(33))
                           ;
   U77 : OAI221_X1 port map( B1 => net267119, B2 => n473, C1 => net267121, C2 
                           => n474, A => n51, ZN => O(30));
   U78 : NAND2_X1 port map( A1 => A_s(30), A2 => net267127, ZN => n51);
   U79 : OAI221_X1 port map( B1 => net267119, B2 => n465, C1 => net267123, C2 
                           => n467, A => n57, ZN => O(25));
   U80 : NAND2_X1 port map( A1 => A_s(25), A2 => net267127, ZN => n57);
   U81 : OAI221_X1 port map( B1 => net267119, B2 => n462, C1 => net267123, C2 
                           => n464, A => n59, ZN => O(23));
   U82 : NAND2_X1 port map( A1 => A_s(23), A2 => net267127, ZN => n59);
   U83 : OAI221_X1 port map( B1 => net267119, B2 => n468, C1 => net267123, C2 
                           => n470, A => n55, ZN => O(27));
   U84 : NAND2_X1 port map( A1 => A_s(27), A2 => net267127, ZN => n55);
   U85 : OAI221_X1 port map( B1 => net267119, B2 => n458, C1 => net267123, C2 
                           => n459, A => n62, ZN => O(20));
   U86 : NAND2_X1 port map( A1 => A_s(20), A2 => net267127, ZN => n62);
   U87 : NAND2_X1 port map( A1 => A_s(28), A2 => net267127, ZN => n54);
   U88 : NAND2_X1 port map( A1 => A_s(21), A2 => net267127, ZN => n61);
   U89 : NAND2_X1 port map( A1 => A_s(24), A2 => net267127, ZN => n58);
   U90 : NAND2_X1 port map( A1 => A_s(26), A2 => net267127, ZN => n56);
   U91 : NAND2_X1 port map( A1 => A_s(22), A2 => net267127, ZN => n60);
   U92 : OAI221_X1 port map( B1 => net267119, B2 => n471, C1 => net267123, C2 
                           => n473, A => n53, ZN => O(29));
   U93 : NAND2_X1 port map( A1 => A_s(29), A2 => net267127, ZN => n53);
   U94 : OAI221_X1 port map( B1 => net267119, B2 => n474, C1 => net267121, C2 
                           => n476, A => n50, ZN => O(31));
   U95 : NAND2_X1 port map( A1 => A_s(31), A2 => net267127, ZN => n50);
   U96 : INV_X1 port map( A => A_ns(23), ZN => n464);
   U97 : INV_X1 port map( A => A_ns(21), ZN => n461);
   U98 : INV_X1 port map( A => A_ns(27), ZN => n470);
   U99 : INV_X1 port map( A => A_ns(25), ZN => n467);
   U100 : NAND2_X1 port map( A1 => A_s(32), A2 => net267127, ZN => n49);
   U101 : OAI221_X1 port map( B1 => net267119, B2 => n479, C1 => net267123, C2 
                           => net278161, A => n63, ZN => O(1));
   U102 : NAND2_X1 port map( A1 => A_s(1), A2 => net267127, ZN => n63);
   U103 : INV_X1 port map( A => net267129, ZN => net268556);
   U104 : INV_X1 port map( A => A_ns(4), ZN => net267007);
   U105 : INV_X1 port map( A => n437, ZN => A_nso_6_port);
   U106 : INV_X1 port map( A => A_ns(6), ZN => n438);
   U107 : INV_X1 port map( A => n440, ZN => A_nso_8_port);
   U108 : INV_X1 port map( A => A_ns(8), ZN => n441);
   U109 : INV_X1 port map( A => n443, ZN => A_nso_10_port);
   U110 : INV_X1 port map( A => A_ns(10), ZN => n444);
   U111 : INV_X1 port map( A => n446, ZN => A_nso_12_port);
   U112 : INV_X1 port map( A => A_ns(12), ZN => n447);
   U113 : INV_X1 port map( A => n449, ZN => A_nso_14_port);
   U114 : INV_X1 port map( A => A_ns(14), ZN => n450);
   U115 : INV_X1 port map( A => n452, ZN => A_nso_16_port);
   U116 : INV_X1 port map( A => A_ns(16), ZN => n453);
   U117 : INV_X1 port map( A => n455, ZN => A_nso_18_port);
   U118 : INV_X1 port map( A => A_ns(18), ZN => n456);
   U119 : INV_X1 port map( A => n458, ZN => A_nso_20_port);
   U120 : INV_X1 port map( A => A_ns(20), ZN => n459);
   U121 : INV_X1 port map( A => n461, ZN => A_nso_22_port);
   U122 : INV_X1 port map( A => A_ns(22), ZN => n462);
   U123 : INV_X1 port map( A => n464, ZN => A_nso_24_port);
   U124 : INV_X1 port map( A => A_ns(24), ZN => n465);
   U125 : INV_X1 port map( A => n467, ZN => A_nso_26_port);
   U126 : INV_X1 port map( A => A_ns(26), ZN => n468);
   U127 : INV_X1 port map( A => n470, ZN => A_nso_28_port);
   U128 : INV_X1 port map( A => A_ns(28), ZN => n471);
   U129 : INV_X1 port map( A => n473, ZN => A_nso_30_port);
   U130 : INV_X1 port map( A => A_ns(30), ZN => n474);
   U131 : INV_X1 port map( A => n476, ZN => A_nso_32_port);
   U132 : INV_X1 port map( A => A_ns(33), ZN => n478);
   U133 : INV_X1 port map( A => A_s(0), ZN => n480);
   U134 : INV_X1 port map( A => A_s(33), ZN => n481);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHMUL_NBIT32 is

   port( A, B : in std_logic_vector (31 downto 0);  S : out std_logic_vector 
         (63 downto 0));

end BOOTHMUL_NBIT32;

architecture SYN_BEHAVIOURAL of BOOTHMUL_NBIT32 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BOOTHMUL_NBIT32_DW01_sub_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component RCA_NBIT64
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT62
      port( A, B : in std_logic_vector (61 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (61 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT60
      port( A, B : in std_logic_vector (59 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (59 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT58
      port( A, B : in std_logic_vector (57 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (57 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT56
      port( A, B : in std_logic_vector (55 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (55 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT54
      port( A, B : in std_logic_vector (53 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (53 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT52
      port( A, B : in std_logic_vector (51 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (51 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT50
      port( A, B : in std_logic_vector (49 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (49 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT48
      port( A, B : in std_logic_vector (47 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (47 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT46
      port( A, B : in std_logic_vector (45 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (45 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT44
      port( A, B : in std_logic_vector (43 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (43 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT42
      port( A, B : in std_logic_vector (41 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (41 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT40
      port( A, B : in std_logic_vector (39 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (39 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT38
      port( A, B : in std_logic_vector (37 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (37 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT36
      port( A, B : in std_logic_vector (35 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (35 downto 0);  Co : out std_logic);
   end component;
   
   component BOOTHENC_NBIT64_i30
      port( A_s, A_ns, B : in std_logic_vector (63 downto 0);  O, A_so, A_nso :
            out std_logic_vector (63 downto 0));
   end component;
   
   component BOOTHENC_NBIT62_i28
      port( A_s, A_ns, B : in std_logic_vector (61 downto 0);  O, A_so, A_nso :
            out std_logic_vector (61 downto 0));
   end component;
   
   component BOOTHENC_NBIT60_i26
      port( A_s, A_ns, B : in std_logic_vector (59 downto 0);  O, A_so, A_nso :
            out std_logic_vector (59 downto 0));
   end component;
   
   component BOOTHENC_NBIT58_i24
      port( A_s, A_ns, B : in std_logic_vector (57 downto 0);  O, A_so, A_nso :
            out std_logic_vector (57 downto 0));
   end component;
   
   component BOOTHENC_NBIT56_i22
      port( A_s, A_ns, B : in std_logic_vector (55 downto 0);  O, A_so, A_nso :
            out std_logic_vector (55 downto 0));
   end component;
   
   component BOOTHENC_NBIT54_i20
      port( A_s, A_ns, B : in std_logic_vector (53 downto 0);  O, A_so, A_nso :
            out std_logic_vector (53 downto 0));
   end component;
   
   component BOOTHENC_NBIT52_i18
      port( A_s, A_ns, B : in std_logic_vector (51 downto 0);  O, A_so, A_nso :
            out std_logic_vector (51 downto 0));
   end component;
   
   component BOOTHENC_NBIT50_i16
      port( A_s, A_ns, B : in std_logic_vector (49 downto 0);  O, A_so, A_nso :
            out std_logic_vector (49 downto 0));
   end component;
   
   component BOOTHENC_NBIT48_i14
      port( A_s, A_ns, B : in std_logic_vector (47 downto 0);  O, A_so, A_nso :
            out std_logic_vector (47 downto 0));
   end component;
   
   component BOOTHENC_NBIT46_i12
      port( A_s, A_ns, B : in std_logic_vector (45 downto 0);  O, A_so, A_nso :
            out std_logic_vector (45 downto 0));
   end component;
   
   component BOOTHENC_NBIT44_i10
      port( A_s, A_ns, B : in std_logic_vector (43 downto 0);  O, A_so, A_nso :
            out std_logic_vector (43 downto 0));
   end component;
   
   component BOOTHENC_NBIT42_i8
      port( A_s, A_ns, B : in std_logic_vector (41 downto 0);  O, A_so, A_nso :
            out std_logic_vector (41 downto 0));
   end component;
   
   component BOOTHENC_NBIT40_i6
      port( A_s, A_ns, B : in std_logic_vector (39 downto 0);  O, A_so, A_nso :
            out std_logic_vector (39 downto 0));
   end component;
   
   component BOOTHENC_NBIT38_i4
      port( A_s, A_ns, B : in std_logic_vector (37 downto 0);  O, A_so, A_nso :
            out std_logic_vector (37 downto 0));
   end component;
   
   component BOOTHENC_NBIT36_i2
      port( A_s, A_ns, B : in std_logic_vector (35 downto 0);  O, A_so, A_nso :
            out std_logic_vector (35 downto 0));
   end component;
   
   component BOOTHENC_NBIT34_i0
      port( A_s, A_ns, B : in std_logic_vector (33 downto 0);  O, A_so, A_nso :
            out std_logic_vector (33 downto 0));
   end component;
   
   signal X_Logic0_port, A_n_65, A_n_30_port, A_n_29_port, A_n_28_port, 
      A_n_27_port, A_n_26_port, A_n_25_port, A_n_24_port, A_n_23_port, 
      A_n_22_port, A_n_21_port, A_n_20_port, A_n_19_port, A_n_18_port, 
      A_n_17_port, A_n_16_port, A_n_15_port, A_n_14_port, A_n_13_port, 
      A_n_12_port, A_n_11_port, A_n_10_port, A_n_9_port, A_n_8_port, A_n_7_port
      , A_n_6_port, A_n_5_port, A_n_4_port, A_n_3_port, A_n_2_port, A_n_1_port,
      A_n_0_port, SHIFT_1_31_port, SHIFT_1_30_port, SHIFT_1_29_port, 
      SHIFT_1_28_port, SHIFT_1_27_port, SHIFT_1_26_port, SHIFT_1_25_port, 
      SHIFT_1_24_port, SHIFT_1_23_port, SHIFT_1_22_port, SHIFT_1_21_port, 
      SHIFT_1_20_port, SHIFT_1_19_port, SHIFT_1_18_port, SHIFT_1_17_port, 
      SHIFT_1_16_port, SHIFT_1_15_port, SHIFT_1_14_port, SHIFT_1_13_port, 
      SHIFT_1_12_port, SHIFT_1_11_port, SHIFT_1_10_port, SHIFT_1_9_port, 
      SHIFT_1_8_port, SHIFT_1_7_port, SHIFT_1_6_port, SHIFT_1_5_port, 
      SHIFT_1_4_port, SHIFT_1_3_port, SHIFT_1_2_port, SHIFT_1_1_port, 
      SHIFT_1_0_port, SHIFT_15_61_port, SHIFT_15_60_port, SHIFT_15_59_port, 
      SHIFT_15_58_port, SHIFT_15_57_port, SHIFT_15_56_port, SHIFT_15_55_port, 
      SHIFT_15_54_port, SHIFT_15_53_port, SHIFT_15_52_port, SHIFT_15_51_port, 
      SHIFT_15_50_port, SHIFT_15_49_port, SHIFT_15_48_port, SHIFT_15_47_port, 
      SHIFT_15_46_port, SHIFT_15_45_port, SHIFT_15_44_port, SHIFT_15_43_port, 
      SHIFT_15_42_port, SHIFT_15_41_port, SHIFT_15_40_port, SHIFT_15_39_port, 
      SHIFT_15_38_port, SHIFT_15_37_port, SHIFT_15_36_port, SHIFT_15_35_port, 
      SHIFT_15_34_port, SHIFT_15_33_port, SHIFT_15_32_port, SHIFT_15_31_port, 
      SHIFT_15_30_port, SHIFT_15_29_port, SHIFT_15_28_port, SHIFT_15_27_port, 
      SHIFT_15_26_port, SHIFT_15_25_port, SHIFT_15_24_port, SHIFT_15_23_port, 
      SHIFT_15_22_port, SHIFT_15_21_port, SHIFT_15_20_port, SHIFT_15_19_port, 
      SHIFT_15_18_port, SHIFT_15_17_port, SHIFT_15_16_port, SHIFT_15_15_port, 
      SHIFT_15_14_port, SHIFT_15_13_port, SHIFT_15_12_port, SHIFT_15_11_port, 
      SHIFT_15_10_port, SHIFT_15_9_port, SHIFT_15_8_port, SHIFT_15_7_port, 
      SHIFT_15_6_port, SHIFT_15_5_port, SHIFT_15_4_port, SHIFT_15_3_port, 
      SHIFT_15_2_port, SHIFT_15_1_port, SHIFT_15_0_port, SHIFT_14_59_port, 
      SHIFT_14_58_port, SHIFT_14_57_port, SHIFT_14_56_port, SHIFT_14_55_port, 
      SHIFT_14_54_port, SHIFT_14_53_port, SHIFT_14_52_port, SHIFT_14_51_port, 
      SHIFT_14_50_port, SHIFT_14_49_port, SHIFT_14_48_port, SHIFT_14_47_port, 
      SHIFT_14_46_port, SHIFT_14_45_port, SHIFT_14_44_port, SHIFT_14_43_port, 
      SHIFT_14_42_port, SHIFT_14_41_port, SHIFT_14_40_port, SHIFT_14_39_port, 
      SHIFT_14_38_port, SHIFT_14_37_port, SHIFT_14_36_port, SHIFT_14_35_port, 
      SHIFT_14_34_port, SHIFT_14_33_port, SHIFT_14_32_port, SHIFT_14_31_port, 
      SHIFT_14_30_port, SHIFT_14_29_port, SHIFT_14_28_port, SHIFT_14_27_port, 
      SHIFT_14_26_port, SHIFT_14_25_port, SHIFT_14_24_port, SHIFT_14_23_port, 
      SHIFT_14_22_port, SHIFT_14_21_port, SHIFT_14_20_port, SHIFT_14_19_port, 
      SHIFT_14_18_port, SHIFT_14_17_port, SHIFT_14_16_port, SHIFT_14_15_port, 
      SHIFT_14_14_port, SHIFT_14_13_port, SHIFT_14_12_port, SHIFT_14_11_port, 
      SHIFT_14_10_port, SHIFT_14_9_port, SHIFT_14_8_port, SHIFT_14_7_port, 
      SHIFT_14_6_port, SHIFT_14_5_port, SHIFT_14_4_port, SHIFT_14_3_port, 
      SHIFT_14_2_port, SHIFT_14_1_port, SHIFT_14_0_port, SHIFT_13_57_port, 
      SHIFT_13_56_port, SHIFT_13_55_port, SHIFT_13_54_port, SHIFT_13_53_port, 
      SHIFT_13_52_port, SHIFT_13_51_port, SHIFT_13_50_port, SHIFT_13_49_port, 
      SHIFT_13_48_port, SHIFT_13_47_port, SHIFT_13_46_port, SHIFT_13_45_port, 
      SHIFT_13_44_port, SHIFT_13_43_port, SHIFT_13_42_port, SHIFT_13_41_port, 
      SHIFT_13_40_port, SHIFT_13_39_port, SHIFT_13_38_port, SHIFT_13_37_port, 
      SHIFT_13_36_port, SHIFT_13_35_port, SHIFT_13_34_port, SHIFT_13_33_port, 
      SHIFT_13_32_port, SHIFT_13_31_port, SHIFT_13_30_port, SHIFT_13_29_port, 
      SHIFT_13_28_port, SHIFT_13_27_port, SHIFT_13_26_port, SHIFT_13_25_port, 
      SHIFT_13_24_port, SHIFT_13_23_port, SHIFT_13_22_port, SHIFT_13_21_port, 
      SHIFT_13_20_port, SHIFT_13_19_port, SHIFT_13_18_port, SHIFT_13_17_port, 
      SHIFT_13_16_port, SHIFT_13_15_port, SHIFT_13_14_port, SHIFT_13_13_port, 
      SHIFT_13_12_port, SHIFT_13_11_port, SHIFT_13_10_port, SHIFT_13_9_port, 
      SHIFT_13_8_port, SHIFT_13_7_port, SHIFT_13_6_port, SHIFT_13_5_port, 
      SHIFT_13_4_port, SHIFT_13_3_port, SHIFT_13_2_port, SHIFT_13_1_port, 
      SHIFT_13_0_port, SHIFT_12_55_port, SHIFT_12_54_port, SHIFT_12_53_port, 
      SHIFT_12_52_port, SHIFT_12_51_port, SHIFT_12_50_port, SHIFT_12_49_port, 
      SHIFT_12_48_port, SHIFT_12_47_port, SHIFT_12_46_port, SHIFT_12_45_port, 
      SHIFT_12_44_port, SHIFT_12_43_port, SHIFT_12_42_port, SHIFT_12_41_port, 
      SHIFT_12_40_port, SHIFT_12_39_port, SHIFT_12_38_port, SHIFT_12_37_port, 
      SHIFT_12_36_port, SHIFT_12_35_port, SHIFT_12_34_port, SHIFT_12_33_port, 
      SHIFT_12_32_port, SHIFT_12_31_port, SHIFT_12_30_port, SHIFT_12_29_port, 
      SHIFT_12_28_port, SHIFT_12_27_port, SHIFT_12_26_port, SHIFT_12_25_port, 
      SHIFT_12_24_port, SHIFT_12_23_port, SHIFT_12_22_port, SHIFT_12_21_port, 
      SHIFT_12_20_port, SHIFT_12_19_port, SHIFT_12_18_port, SHIFT_12_17_port, 
      SHIFT_12_16_port, SHIFT_12_15_port, SHIFT_12_14_port, SHIFT_12_13_port, 
      SHIFT_12_12_port, SHIFT_12_11_port, SHIFT_12_10_port, SHIFT_12_9_port, 
      SHIFT_12_8_port, SHIFT_12_7_port, SHIFT_12_6_port, SHIFT_12_5_port, 
      SHIFT_12_4_port, SHIFT_12_3_port, SHIFT_12_2_port, SHIFT_12_1_port, 
      SHIFT_12_0_port, SHIFT_11_53_port, SHIFT_11_52_port, SHIFT_11_51_port, 
      SHIFT_11_50_port, SHIFT_11_49_port, SHIFT_11_48_port, SHIFT_11_47_port, 
      SHIFT_11_46_port, SHIFT_11_45_port, SHIFT_11_44_port, SHIFT_11_43_port, 
      SHIFT_11_42_port, SHIFT_11_41_port, SHIFT_11_40_port, SHIFT_11_39_port, 
      SHIFT_11_38_port, SHIFT_11_37_port, SHIFT_11_36_port, SHIFT_11_35_port, 
      SHIFT_11_34_port, SHIFT_11_33_port, SHIFT_11_32_port, SHIFT_11_31_port, 
      SHIFT_11_30_port, SHIFT_11_29_port, SHIFT_11_28_port, SHIFT_11_27_port, 
      SHIFT_11_26_port, SHIFT_11_25_port, SHIFT_11_24_port, SHIFT_11_23_port, 
      SHIFT_11_22_port, SHIFT_11_21_port, SHIFT_11_20_port, SHIFT_11_19_port, 
      SHIFT_11_18_port, SHIFT_11_17_port, SHIFT_11_16_port, SHIFT_11_15_port, 
      SHIFT_11_14_port, SHIFT_11_13_port, SHIFT_11_12_port, SHIFT_11_11_port, 
      SHIFT_11_10_port, SHIFT_11_9_port, SHIFT_11_8_port, SHIFT_11_7_port, 
      SHIFT_11_6_port, SHIFT_11_5_port, SHIFT_11_4_port, SHIFT_11_3_port, 
      SHIFT_11_2_port, SHIFT_11_1_port, SHIFT_11_0_port, SHIFT_10_51_port, 
      SHIFT_10_50_port, SHIFT_10_49_port, SHIFT_10_48_port, SHIFT_10_47_port, 
      SHIFT_10_46_port, SHIFT_10_45_port, SHIFT_10_44_port, SHIFT_10_43_port, 
      SHIFT_10_42_port, SHIFT_10_41_port, SHIFT_10_40_port, SHIFT_10_39_port, 
      SHIFT_10_38_port, SHIFT_10_37_port, SHIFT_10_36_port, SHIFT_10_35_port, 
      SHIFT_10_34_port, SHIFT_10_33_port, SHIFT_10_32_port, SHIFT_10_31_port, 
      SHIFT_10_30_port, SHIFT_10_29_port, SHIFT_10_28_port, SHIFT_10_27_port, 
      SHIFT_10_26_port, SHIFT_10_25_port, SHIFT_10_24_port, SHIFT_10_23_port, 
      SHIFT_10_22_port, SHIFT_10_21_port, SHIFT_10_20_port, SHIFT_10_19_port, 
      SHIFT_10_18_port, SHIFT_10_17_port, SHIFT_10_16_port, SHIFT_10_15_port, 
      SHIFT_10_14_port, SHIFT_10_13_port, SHIFT_10_12_port, SHIFT_10_11_port, 
      SHIFT_10_10_port, SHIFT_10_9_port, SHIFT_10_8_port, SHIFT_10_7_port, 
      SHIFT_10_6_port, SHIFT_10_5_port, SHIFT_10_4_port, SHIFT_10_3_port, 
      SHIFT_10_2_port, SHIFT_10_1_port, SHIFT_10_0_port, SHIFT_9_49_port, 
      SHIFT_9_48_port, SHIFT_9_47_port, SHIFT_9_46_port, SHIFT_9_45_port, 
      SHIFT_9_44_port, SHIFT_9_43_port, SHIFT_9_42_port, SHIFT_9_41_port, 
      SHIFT_9_40_port, SHIFT_9_39_port, SHIFT_9_38_port, SHIFT_9_37_port, 
      SHIFT_9_36_port, SHIFT_9_35_port, SHIFT_9_34_port, SHIFT_9_33_port, 
      SHIFT_9_32_port, SHIFT_9_31_port, SHIFT_9_30_port, SHIFT_9_29_port, 
      SHIFT_9_28_port, SHIFT_9_27_port, SHIFT_9_26_port, SHIFT_9_25_port, 
      SHIFT_9_24_port, SHIFT_9_23_port, SHIFT_9_22_port, SHIFT_9_21_port, 
      SHIFT_9_20_port, SHIFT_9_19_port, SHIFT_9_18_port, SHIFT_9_17_port, 
      SHIFT_9_16_port, SHIFT_9_15_port, SHIFT_9_14_port, SHIFT_9_13_port, 
      SHIFT_9_12_port, SHIFT_9_11_port, SHIFT_9_10_port, SHIFT_9_9_port, 
      SHIFT_9_8_port, SHIFT_9_7_port, SHIFT_9_6_port, SHIFT_9_5_port, 
      SHIFT_9_4_port, SHIFT_9_3_port, SHIFT_9_2_port, SHIFT_9_1_port, 
      SHIFT_9_0_port, SHIFT_8_47_port, SHIFT_8_46_port, SHIFT_8_45_port, 
      SHIFT_8_44_port, SHIFT_8_43_port, SHIFT_8_42_port, SHIFT_8_41_port, 
      SHIFT_8_40_port, SHIFT_8_39_port, SHIFT_8_38_port, SHIFT_8_37_port, 
      SHIFT_8_36_port, SHIFT_8_35_port, SHIFT_8_34_port, SHIFT_8_33_port, 
      SHIFT_8_32_port, SHIFT_8_31_port, SHIFT_8_30_port, SHIFT_8_29_port, 
      SHIFT_8_28_port, SHIFT_8_27_port, SHIFT_8_26_port, SHIFT_8_25_port, 
      SHIFT_8_24_port, SHIFT_8_23_port, SHIFT_8_22_port, SHIFT_8_21_port, 
      SHIFT_8_20_port, SHIFT_8_19_port, SHIFT_8_18_port, SHIFT_8_17_port, 
      SHIFT_8_16_port, SHIFT_8_15_port, SHIFT_8_14_port, SHIFT_8_13_port, 
      SHIFT_8_12_port, SHIFT_8_11_port, SHIFT_8_10_port, SHIFT_8_9_port, 
      SHIFT_8_8_port, SHIFT_8_7_port, SHIFT_8_6_port, SHIFT_8_5_port, 
      SHIFT_8_4_port, SHIFT_8_3_port, SHIFT_8_2_port, SHIFT_8_1_port, 
      SHIFT_8_0_port, SHIFT_7_45_port, SHIFT_7_44_port, SHIFT_7_43_port, 
      SHIFT_7_42_port, SHIFT_7_41_port, SHIFT_7_40_port, SHIFT_7_39_port, 
      SHIFT_7_38_port, SHIFT_7_37_port, SHIFT_7_36_port, SHIFT_7_35_port, 
      SHIFT_7_34_port, SHIFT_7_33_port, SHIFT_7_32_port, SHIFT_7_31_port, 
      SHIFT_7_30_port, SHIFT_7_29_port, SHIFT_7_28_port, SHIFT_7_27_port, 
      SHIFT_7_26_port, SHIFT_7_25_port, SHIFT_7_24_port, SHIFT_7_23_port, 
      SHIFT_7_22_port, SHIFT_7_21_port, SHIFT_7_20_port, SHIFT_7_19_port, 
      SHIFT_7_18_port, SHIFT_7_17_port, SHIFT_7_16_port, SHIFT_7_15_port, 
      SHIFT_7_14_port, SHIFT_7_13_port, SHIFT_7_12_port, SHIFT_7_11_port, 
      SHIFT_7_10_port, SHIFT_7_9_port, SHIFT_7_8_port, SHIFT_7_7_port, 
      SHIFT_7_6_port, SHIFT_7_5_port, SHIFT_7_4_port, SHIFT_7_3_port, 
      SHIFT_7_2_port, SHIFT_7_1_port, SHIFT_7_0_port, SHIFT_6_43_port, 
      SHIFT_6_42_port, SHIFT_6_41_port, SHIFT_6_40_port, SHIFT_6_39_port, 
      SHIFT_6_38_port, SHIFT_6_37_port, SHIFT_6_36_port, SHIFT_6_35_port, 
      SHIFT_6_34_port, SHIFT_6_33_port, SHIFT_6_32_port, SHIFT_6_31_port, 
      SHIFT_6_30_port, SHIFT_6_29_port, SHIFT_6_28_port, SHIFT_6_27_port, 
      SHIFT_6_26_port, SHIFT_6_25_port, SHIFT_6_24_port, SHIFT_6_23_port, 
      SHIFT_6_22_port, SHIFT_6_21_port, SHIFT_6_20_port, SHIFT_6_19_port, 
      SHIFT_6_18_port, SHIFT_6_17_port, SHIFT_6_16_port, SHIFT_6_15_port, 
      SHIFT_6_14_port, SHIFT_6_13_port, SHIFT_6_12_port, SHIFT_6_11_port, 
      SHIFT_6_10_port, SHIFT_6_9_port, SHIFT_6_8_port, SHIFT_6_7_port, 
      SHIFT_6_6_port, SHIFT_6_5_port, SHIFT_6_4_port, SHIFT_6_3_port, 
      SHIFT_6_2_port, SHIFT_6_1_port, SHIFT_6_0_port, SHIFT_5_41_port, 
      SHIFT_5_40_port, SHIFT_5_39_port, SHIFT_5_38_port, SHIFT_5_37_port, 
      SHIFT_5_36_port, SHIFT_5_35_port, SHIFT_5_34_port, SHIFT_5_33_port, 
      SHIFT_5_32_port, SHIFT_5_31_port, SHIFT_5_30_port, SHIFT_5_29_port, 
      SHIFT_5_28_port, SHIFT_5_27_port, SHIFT_5_26_port, SHIFT_5_25_port, 
      SHIFT_5_24_port, SHIFT_5_23_port, SHIFT_5_22_port, SHIFT_5_21_port, 
      SHIFT_5_20_port, SHIFT_5_19_port, SHIFT_5_18_port, SHIFT_5_17_port, 
      SHIFT_5_16_port, SHIFT_5_15_port, SHIFT_5_14_port, SHIFT_5_13_port, 
      SHIFT_5_12_port, SHIFT_5_11_port, SHIFT_5_10_port, SHIFT_5_9_port, 
      SHIFT_5_8_port, SHIFT_5_7_port, SHIFT_5_6_port, SHIFT_5_5_port, 
      SHIFT_5_4_port, SHIFT_5_3_port, SHIFT_5_2_port, SHIFT_5_1_port, 
      SHIFT_5_0_port, SHIFT_4_39_port, SHIFT_4_38_port, SHIFT_4_37_port, 
      SHIFT_4_36_port, SHIFT_4_35_port, SHIFT_4_34_port, SHIFT_4_33_port, 
      SHIFT_4_32_port, SHIFT_4_31_port, SHIFT_4_30_port, SHIFT_4_29_port, 
      SHIFT_4_28_port, SHIFT_4_27_port, SHIFT_4_26_port, SHIFT_4_25_port, 
      SHIFT_4_24_port, SHIFT_4_23_port, SHIFT_4_22_port, SHIFT_4_21_port, 
      SHIFT_4_20_port, SHIFT_4_19_port, SHIFT_4_18_port, SHIFT_4_17_port, 
      SHIFT_4_16_port, SHIFT_4_15_port, SHIFT_4_14_port, SHIFT_4_13_port, 
      SHIFT_4_12_port, SHIFT_4_11_port, SHIFT_4_10_port, SHIFT_4_9_port, 
      SHIFT_4_8_port, SHIFT_4_7_port, SHIFT_4_6_port, SHIFT_4_5_port, 
      SHIFT_4_4_port, SHIFT_4_3_port, SHIFT_4_2_port, SHIFT_4_1_port, 
      SHIFT_4_0_port, SHIFT_3_37_port, SHIFT_3_36_port, SHIFT_3_35_port, 
      SHIFT_3_34_port, SHIFT_3_33_port, SHIFT_3_32_port, SHIFT_3_31_port, 
      SHIFT_3_30_port, SHIFT_3_29_port, SHIFT_3_28_port, SHIFT_3_27_port, 
      SHIFT_3_26_port, SHIFT_3_25_port, SHIFT_3_24_port, SHIFT_3_23_port, 
      SHIFT_3_22_port, SHIFT_3_21_port, SHIFT_3_20_port, SHIFT_3_19_port, 
      SHIFT_3_18_port, SHIFT_3_17_port, SHIFT_3_16_port, SHIFT_3_15_port, 
      SHIFT_3_14_port, SHIFT_3_13_port, SHIFT_3_12_port, SHIFT_3_11_port, 
      SHIFT_3_10_port, SHIFT_3_9_port, SHIFT_3_8_port, SHIFT_3_7_port, 
      SHIFT_3_6_port, SHIFT_3_5_port, SHIFT_3_4_port, SHIFT_3_3_port, 
      SHIFT_3_2_port, SHIFT_3_1_port, SHIFT_3_0_port, SHIFT_2_35_port, 
      SHIFT_2_34_port, SHIFT_2_33_port, SHIFT_2_32_port, SHIFT_2_31_port, 
      SHIFT_2_30_port, SHIFT_2_29_port, SHIFT_2_28_port, SHIFT_2_27_port, 
      SHIFT_2_26_port, SHIFT_2_25_port, SHIFT_2_24_port, SHIFT_2_23_port, 
      SHIFT_2_22_port, SHIFT_2_21_port, SHIFT_2_20_port, SHIFT_2_19_port, 
      SHIFT_2_18_port, SHIFT_2_17_port, SHIFT_2_16_port, SHIFT_2_15_port, 
      SHIFT_2_14_port, SHIFT_2_13_port, SHIFT_2_12_port, SHIFT_2_11_port, 
      SHIFT_2_10_port, SHIFT_2_9_port, SHIFT_2_8_port, SHIFT_2_7_port, 
      SHIFT_2_6_port, SHIFT_2_5_port, SHIFT_2_4_port, SHIFT_2_3_port, 
      SHIFT_2_2_port, SHIFT_2_1_port, SHIFT_2_0_port, SHIFT_1_33_port, 
      SHIFT_1_32_port, SHIFT_n_1_31_port, SHIFT_n_1_30_port, SHIFT_n_1_29_port,
      SHIFT_n_1_28_port, SHIFT_n_1_27_port, SHIFT_n_1_26_port, 
      SHIFT_n_1_25_port, SHIFT_n_1_24_port, SHIFT_n_1_23_port, 
      SHIFT_n_1_22_port, SHIFT_n_1_21_port, SHIFT_n_1_20_port, 
      SHIFT_n_1_19_port, SHIFT_n_1_18_port, SHIFT_n_1_17_port, 
      SHIFT_n_1_16_port, SHIFT_n_1_15_port, SHIFT_n_1_14_port, 
      SHIFT_n_1_13_port, SHIFT_n_1_12_port, SHIFT_n_1_11_port, 
      SHIFT_n_1_10_port, SHIFT_n_1_9_port, SHIFT_n_1_8_port, SHIFT_n_1_7_port, 
      SHIFT_n_1_6_port, SHIFT_n_1_5_port, SHIFT_n_1_4_port, SHIFT_n_1_3_port, 
      SHIFT_n_1_2_port, SHIFT_n_1_1_port, SHIFT_n_1_0_port, SHIFT_n_15_61_port,
      SHIFT_n_15_60_port, SHIFT_n_15_59_port, SHIFT_n_15_58_port, 
      SHIFT_n_15_57_port, SHIFT_n_15_56_port, SHIFT_n_15_55_port, 
      SHIFT_n_15_54_port, SHIFT_n_15_53_port, SHIFT_n_15_52_port, 
      SHIFT_n_15_51_port, SHIFT_n_15_50_port, SHIFT_n_15_49_port, 
      SHIFT_n_15_48_port, SHIFT_n_15_47_port, SHIFT_n_15_46_port, 
      SHIFT_n_15_45_port, SHIFT_n_15_44_port, SHIFT_n_15_43_port, 
      SHIFT_n_15_42_port, SHIFT_n_15_41_port, SHIFT_n_15_40_port, 
      SHIFT_n_15_39_port, SHIFT_n_15_38_port, SHIFT_n_15_37_port, 
      SHIFT_n_15_36_port, SHIFT_n_15_35_port, SHIFT_n_15_34_port, 
      SHIFT_n_15_33_port, SHIFT_n_15_32_port, SHIFT_n_15_31_port, 
      SHIFT_n_15_30_port, SHIFT_n_15_29_port, SHIFT_n_15_28_port, 
      SHIFT_n_15_27_port, SHIFT_n_15_26_port, SHIFT_n_15_25_port, 
      SHIFT_n_15_24_port, SHIFT_n_15_23_port, SHIFT_n_15_22_port, 
      SHIFT_n_15_21_port, SHIFT_n_15_20_port, SHIFT_n_15_19_port, 
      SHIFT_n_15_18_port, SHIFT_n_15_17_port, SHIFT_n_15_16_port, 
      SHIFT_n_15_15_port, SHIFT_n_15_14_port, SHIFT_n_15_13_port, 
      SHIFT_n_15_12_port, SHIFT_n_15_11_port, SHIFT_n_15_10_port, 
      SHIFT_n_15_9_port, SHIFT_n_15_8_port, SHIFT_n_15_7_port, 
      SHIFT_n_15_6_port, SHIFT_n_15_5_port, SHIFT_n_15_4_port, 
      SHIFT_n_15_3_port, SHIFT_n_15_2_port, SHIFT_n_15_1_port, 
      SHIFT_n_15_0_port, SHIFT_n_14_59_port, SHIFT_n_14_58_port, 
      SHIFT_n_14_57_port, SHIFT_n_14_56_port, SHIFT_n_14_55_port, 
      SHIFT_n_14_54_port, SHIFT_n_14_53_port, SHIFT_n_14_52_port, 
      SHIFT_n_14_51_port, SHIFT_n_14_50_port, SHIFT_n_14_49_port, 
      SHIFT_n_14_48_port, SHIFT_n_14_47_port, SHIFT_n_14_46_port, 
      SHIFT_n_14_45_port, SHIFT_n_14_44_port, SHIFT_n_14_43_port, 
      SHIFT_n_14_42_port, SHIFT_n_14_41_port, SHIFT_n_14_40_port, 
      SHIFT_n_14_39_port, SHIFT_n_14_38_port, SHIFT_n_14_37_port, 
      SHIFT_n_14_36_port, SHIFT_n_14_35_port, SHIFT_n_14_34_port, 
      SHIFT_n_14_33_port, SHIFT_n_14_32_port, SHIFT_n_14_31_port, 
      SHIFT_n_14_30_port, SHIFT_n_14_29_port, SHIFT_n_14_28_port, 
      SHIFT_n_14_27_port, SHIFT_n_14_26_port, SHIFT_n_14_25_port, 
      SHIFT_n_14_24_port, SHIFT_n_14_23_port, SHIFT_n_14_22_port, 
      SHIFT_n_14_21_port, SHIFT_n_14_20_port, SHIFT_n_14_19_port, 
      SHIFT_n_14_18_port, SHIFT_n_14_17_port, SHIFT_n_14_16_port, 
      SHIFT_n_14_15_port, SHIFT_n_14_14_port, SHIFT_n_14_13_port, 
      SHIFT_n_14_12_port, SHIFT_n_14_11_port, SHIFT_n_14_10_port, 
      SHIFT_n_14_9_port, SHIFT_n_14_8_port, SHIFT_n_14_7_port, 
      SHIFT_n_14_6_port, SHIFT_n_14_5_port, SHIFT_n_14_4_port, 
      SHIFT_n_14_3_port, SHIFT_n_14_2_port, SHIFT_n_14_1_port, 
      SHIFT_n_14_0_port, SHIFT_n_13_57_port, SHIFT_n_13_56_port, 
      SHIFT_n_13_55_port, SHIFT_n_13_54_port, SHIFT_n_13_53_port, 
      SHIFT_n_13_52_port, SHIFT_n_13_51_port, SHIFT_n_13_50_port, 
      SHIFT_n_13_49_port, SHIFT_n_13_48_port, SHIFT_n_13_47_port, 
      SHIFT_n_13_46_port, SHIFT_n_13_45_port, SHIFT_n_13_44_port, 
      SHIFT_n_13_43_port, SHIFT_n_13_42_port, SHIFT_n_13_41_port, 
      SHIFT_n_13_40_port, SHIFT_n_13_39_port, SHIFT_n_13_38_port, 
      SHIFT_n_13_37_port, SHIFT_n_13_36_port, SHIFT_n_13_35_port, 
      SHIFT_n_13_34_port, SHIFT_n_13_33_port, SHIFT_n_13_32_port, 
      SHIFT_n_13_31_port, SHIFT_n_13_30_port, SHIFT_n_13_29_port, 
      SHIFT_n_13_28_port, SHIFT_n_13_27_port, SHIFT_n_13_26_port, 
      SHIFT_n_13_25_port, SHIFT_n_13_24_port, SHIFT_n_13_23_port, 
      SHIFT_n_13_22_port, SHIFT_n_13_21_port, SHIFT_n_13_20_port, 
      SHIFT_n_13_19_port, SHIFT_n_13_18_port, SHIFT_n_13_17_port, 
      SHIFT_n_13_16_port, SHIFT_n_13_15_port, SHIFT_n_13_14_port, 
      SHIFT_n_13_13_port, SHIFT_n_13_12_port, SHIFT_n_13_11_port, 
      SHIFT_n_13_10_port, SHIFT_n_13_9_port, SHIFT_n_13_8_port, 
      SHIFT_n_13_7_port, SHIFT_n_13_6_port, SHIFT_n_13_5_port, 
      SHIFT_n_13_4_port, SHIFT_n_13_3_port, SHIFT_n_13_2_port, 
      SHIFT_n_13_1_port, SHIFT_n_13_0_port, SHIFT_n_12_55_port, 
      SHIFT_n_12_54_port, SHIFT_n_12_53_port, SHIFT_n_12_52_port, 
      SHIFT_n_12_51_port, SHIFT_n_12_50_port, SHIFT_n_12_49_port, 
      SHIFT_n_12_48_port, SHIFT_n_12_47_port, SHIFT_n_12_46_port, 
      SHIFT_n_12_45_port, SHIFT_n_12_44_port, SHIFT_n_12_43_port, 
      SHIFT_n_12_42_port, SHIFT_n_12_41_port, SHIFT_n_12_40_port, 
      SHIFT_n_12_39_port, SHIFT_n_12_38_port, SHIFT_n_12_37_port, 
      SHIFT_n_12_36_port, SHIFT_n_12_35_port, SHIFT_n_12_34_port, 
      SHIFT_n_12_33_port, SHIFT_n_12_32_port, SHIFT_n_12_31_port, 
      SHIFT_n_12_30_port, SHIFT_n_12_29_port, SHIFT_n_12_28_port, 
      SHIFT_n_12_27_port, SHIFT_n_12_26_port, SHIFT_n_12_25_port, 
      SHIFT_n_12_24_port, SHIFT_n_12_23_port, SHIFT_n_12_22_port, 
      SHIFT_n_12_21_port, SHIFT_n_12_20_port, SHIFT_n_12_19_port, 
      SHIFT_n_12_18_port, SHIFT_n_12_17_port, SHIFT_n_12_16_port, 
      SHIFT_n_12_15_port, SHIFT_n_12_14_port, SHIFT_n_12_13_port, 
      SHIFT_n_12_12_port, SHIFT_n_12_11_port, SHIFT_n_12_10_port, 
      SHIFT_n_12_9_port, SHIFT_n_12_8_port, SHIFT_n_12_7_port, 
      SHIFT_n_12_6_port, SHIFT_n_12_5_port, SHIFT_n_12_4_port, 
      SHIFT_n_12_3_port, SHIFT_n_12_2_port, SHIFT_n_12_1_port, 
      SHIFT_n_12_0_port, SHIFT_n_11_53_port, SHIFT_n_11_52_port, 
      SHIFT_n_11_51_port, SHIFT_n_11_50_port, SHIFT_n_11_49_port, 
      SHIFT_n_11_48_port, SHIFT_n_11_47_port, SHIFT_n_11_46_port, 
      SHIFT_n_11_45_port, SHIFT_n_11_44_port, SHIFT_n_11_43_port, 
      SHIFT_n_11_42_port, SHIFT_n_11_41_port, SHIFT_n_11_40_port, 
      SHIFT_n_11_39_port, SHIFT_n_11_38_port, SHIFT_n_11_37_port, 
      SHIFT_n_11_36_port, SHIFT_n_11_35_port, SHIFT_n_11_34_port, 
      SHIFT_n_11_33_port, SHIFT_n_11_32_port, SHIFT_n_11_31_port, 
      SHIFT_n_11_30_port, SHIFT_n_11_29_port, SHIFT_n_11_28_port, 
      SHIFT_n_11_27_port, SHIFT_n_11_26_port, SHIFT_n_11_25_port, 
      SHIFT_n_11_24_port, SHIFT_n_11_23_port, SHIFT_n_11_22_port, 
      SHIFT_n_11_21_port, SHIFT_n_11_20_port, SHIFT_n_11_19_port, 
      SHIFT_n_11_18_port, SHIFT_n_11_17_port, SHIFT_n_11_16_port, 
      SHIFT_n_11_15_port, SHIFT_n_11_14_port, SHIFT_n_11_13_port, 
      SHIFT_n_11_12_port, SHIFT_n_11_11_port, SHIFT_n_11_10_port, 
      SHIFT_n_11_9_port, SHIFT_n_11_8_port, SHIFT_n_11_7_port, 
      SHIFT_n_11_6_port, SHIFT_n_11_5_port, SHIFT_n_11_4_port, 
      SHIFT_n_11_3_port, SHIFT_n_11_2_port, SHIFT_n_11_1_port, 
      SHIFT_n_11_0_port, SHIFT_n_10_51_port, SHIFT_n_10_50_port, 
      SHIFT_n_10_49_port, SHIFT_n_10_48_port, SHIFT_n_10_47_port, 
      SHIFT_n_10_46_port, SHIFT_n_10_45_port, SHIFT_n_10_44_port, 
      SHIFT_n_10_43_port, SHIFT_n_10_42_port, SHIFT_n_10_41_port, 
      SHIFT_n_10_40_port, SHIFT_n_10_39_port, SHIFT_n_10_38_port, 
      SHIFT_n_10_37_port, SHIFT_n_10_36_port, SHIFT_n_10_35_port, 
      SHIFT_n_10_34_port, SHIFT_n_10_33_port, SHIFT_n_10_32_port, 
      SHIFT_n_10_31_port, SHIFT_n_10_30_port, SHIFT_n_10_29_port, 
      SHIFT_n_10_28_port, SHIFT_n_10_27_port, SHIFT_n_10_26_port, 
      SHIFT_n_10_25_port, SHIFT_n_10_24_port, SHIFT_n_10_23_port, 
      SHIFT_n_10_22_port, SHIFT_n_10_21_port, SHIFT_n_10_20_port, 
      SHIFT_n_10_19_port, SHIFT_n_10_18_port, SHIFT_n_10_17_port, 
      SHIFT_n_10_16_port, SHIFT_n_10_15_port, SHIFT_n_10_14_port, 
      SHIFT_n_10_13_port, SHIFT_n_10_12_port, SHIFT_n_10_11_port, 
      SHIFT_n_10_10_port, SHIFT_n_10_9_port, SHIFT_n_10_8_port, 
      SHIFT_n_10_7_port, SHIFT_n_10_6_port, SHIFT_n_10_5_port, 
      SHIFT_n_10_4_port, SHIFT_n_10_3_port, SHIFT_n_10_2_port, 
      SHIFT_n_10_1_port, SHIFT_n_10_0_port, SHIFT_n_9_49_port, 
      SHIFT_n_9_48_port, SHIFT_n_9_47_port, SHIFT_n_9_46_port, 
      SHIFT_n_9_45_port, SHIFT_n_9_44_port, SHIFT_n_9_43_port, 
      SHIFT_n_9_42_port, SHIFT_n_9_41_port, SHIFT_n_9_40_port, 
      SHIFT_n_9_39_port, SHIFT_n_9_38_port, SHIFT_n_9_37_port, 
      SHIFT_n_9_36_port, SHIFT_n_9_35_port, SHIFT_n_9_34_port, 
      SHIFT_n_9_33_port, SHIFT_n_9_32_port, SHIFT_n_9_31_port, 
      SHIFT_n_9_30_port, SHIFT_n_9_29_port, SHIFT_n_9_28_port, 
      SHIFT_n_9_27_port, SHIFT_n_9_26_port, SHIFT_n_9_25_port, 
      SHIFT_n_9_24_port, SHIFT_n_9_23_port, SHIFT_n_9_22_port, 
      SHIFT_n_9_21_port, SHIFT_n_9_20_port, SHIFT_n_9_19_port, 
      SHIFT_n_9_18_port, SHIFT_n_9_17_port, SHIFT_n_9_16_port, 
      SHIFT_n_9_15_port, SHIFT_n_9_14_port, SHIFT_n_9_13_port, 
      SHIFT_n_9_12_port, SHIFT_n_9_11_port, SHIFT_n_9_10_port, SHIFT_n_9_9_port
      , SHIFT_n_9_8_port, SHIFT_n_9_7_port, SHIFT_n_9_6_port, SHIFT_n_9_5_port,
      SHIFT_n_9_4_port, SHIFT_n_9_3_port, SHIFT_n_9_2_port, SHIFT_n_9_1_port, 
      SHIFT_n_9_0_port, SHIFT_n_8_47_port, SHIFT_n_8_46_port, SHIFT_n_8_45_port
      , SHIFT_n_8_44_port, SHIFT_n_8_43_port, SHIFT_n_8_42_port, 
      SHIFT_n_8_41_port, SHIFT_n_8_40_port, SHIFT_n_8_39_port, 
      SHIFT_n_8_38_port, SHIFT_n_8_37_port, SHIFT_n_8_36_port, 
      SHIFT_n_8_35_port, SHIFT_n_8_34_port, SHIFT_n_8_33_port, 
      SHIFT_n_8_32_port, SHIFT_n_8_31_port, SHIFT_n_8_30_port, 
      SHIFT_n_8_29_port, SHIFT_n_8_28_port, SHIFT_n_8_27_port, 
      SHIFT_n_8_26_port, SHIFT_n_8_25_port, SHIFT_n_8_24_port, 
      SHIFT_n_8_23_port, SHIFT_n_8_22_port, SHIFT_n_8_21_port, 
      SHIFT_n_8_20_port, SHIFT_n_8_19_port, SHIFT_n_8_18_port, 
      SHIFT_n_8_17_port, SHIFT_n_8_16_port, SHIFT_n_8_15_port, 
      SHIFT_n_8_14_port, SHIFT_n_8_13_port, SHIFT_n_8_12_port, 
      SHIFT_n_8_11_port, SHIFT_n_8_10_port, SHIFT_n_8_9_port, SHIFT_n_8_8_port,
      SHIFT_n_8_7_port, SHIFT_n_8_6_port, SHIFT_n_8_5_port, SHIFT_n_8_4_port, 
      SHIFT_n_8_3_port, SHIFT_n_8_2_port, SHIFT_n_8_1_port, SHIFT_n_8_0_port, 
      SHIFT_n_7_45_port, SHIFT_n_7_44_port, SHIFT_n_7_43_port, 
      SHIFT_n_7_42_port, SHIFT_n_7_41_port, SHIFT_n_7_40_port, 
      SHIFT_n_7_39_port, SHIFT_n_7_38_port, SHIFT_n_7_37_port, 
      SHIFT_n_7_36_port, SHIFT_n_7_35_port, SHIFT_n_7_34_port, 
      SHIFT_n_7_33_port, SHIFT_n_7_32_port, SHIFT_n_7_31_port, 
      SHIFT_n_7_30_port, SHIFT_n_7_29_port, SHIFT_n_7_28_port, 
      SHIFT_n_7_27_port, SHIFT_n_7_26_port, SHIFT_n_7_25_port, 
      SHIFT_n_7_24_port, SHIFT_n_7_23_port, SHIFT_n_7_22_port, 
      SHIFT_n_7_21_port, SHIFT_n_7_20_port, SHIFT_n_7_19_port, 
      SHIFT_n_7_18_port, SHIFT_n_7_17_port, SHIFT_n_7_16_port, 
      SHIFT_n_7_15_port, SHIFT_n_7_14_port, SHIFT_n_7_13_port, 
      SHIFT_n_7_12_port, SHIFT_n_7_11_port, SHIFT_n_7_10_port, SHIFT_n_7_9_port
      , SHIFT_n_7_8_port, SHIFT_n_7_7_port, SHIFT_n_7_6_port, SHIFT_n_7_5_port,
      SHIFT_n_7_4_port, SHIFT_n_7_3_port, SHIFT_n_7_2_port, SHIFT_n_7_1_port, 
      SHIFT_n_7_0_port, SHIFT_n_6_43_port, SHIFT_n_6_42_port, SHIFT_n_6_41_port
      , SHIFT_n_6_40_port, SHIFT_n_6_39_port, SHIFT_n_6_38_port, 
      SHIFT_n_6_37_port, SHIFT_n_6_36_port, SHIFT_n_6_35_port, 
      SHIFT_n_6_34_port, SHIFT_n_6_33_port, SHIFT_n_6_32_port, 
      SHIFT_n_6_31_port, SHIFT_n_6_30_port, SHIFT_n_6_29_port, 
      SHIFT_n_6_28_port, SHIFT_n_6_27_port, SHIFT_n_6_26_port, 
      SHIFT_n_6_25_port, SHIFT_n_6_24_port, SHIFT_n_6_23_port, 
      SHIFT_n_6_22_port, SHIFT_n_6_21_port, SHIFT_n_6_20_port, 
      SHIFT_n_6_19_port, SHIFT_n_6_18_port, SHIFT_n_6_17_port, 
      SHIFT_n_6_16_port, SHIFT_n_6_15_port, SHIFT_n_6_14_port, 
      SHIFT_n_6_13_port, SHIFT_n_6_12_port, SHIFT_n_6_11_port, 
      SHIFT_n_6_10_port, SHIFT_n_6_9_port, SHIFT_n_6_8_port, SHIFT_n_6_7_port, 
      SHIFT_n_6_6_port, SHIFT_n_6_5_port, SHIFT_n_6_4_port, SHIFT_n_6_3_port, 
      SHIFT_n_6_2_port, SHIFT_n_6_1_port, SHIFT_n_6_0_port, SHIFT_n_5_41_port, 
      SHIFT_n_5_40_port, SHIFT_n_5_39_port, SHIFT_n_5_38_port, 
      SHIFT_n_5_37_port, SHIFT_n_5_36_port, SHIFT_n_5_35_port, 
      SHIFT_n_5_34_port, SHIFT_n_5_33_port, SHIFT_n_5_32_port, 
      SHIFT_n_5_31_port, SHIFT_n_5_30_port, SHIFT_n_5_29_port, 
      SHIFT_n_5_28_port, SHIFT_n_5_27_port, SHIFT_n_5_26_port, 
      SHIFT_n_5_25_port, SHIFT_n_5_24_port, SHIFT_n_5_23_port, 
      SHIFT_n_5_22_port, SHIFT_n_5_21_port, SHIFT_n_5_20_port, 
      SHIFT_n_5_19_port, SHIFT_n_5_18_port, SHIFT_n_5_17_port, 
      SHIFT_n_5_16_port, SHIFT_n_5_15_port, SHIFT_n_5_14_port, 
      SHIFT_n_5_13_port, SHIFT_n_5_12_port, SHIFT_n_5_11_port, 
      SHIFT_n_5_10_port, SHIFT_n_5_9_port, SHIFT_n_5_8_port, SHIFT_n_5_7_port, 
      SHIFT_n_5_6_port, SHIFT_n_5_5_port, SHIFT_n_5_4_port, SHIFT_n_5_3_port, 
      SHIFT_n_5_2_port, SHIFT_n_5_1_port, SHIFT_n_5_0_port, SHIFT_n_4_39_port, 
      SHIFT_n_4_38_port, SHIFT_n_4_37_port, SHIFT_n_4_36_port, 
      SHIFT_n_4_35_port, SHIFT_n_4_34_port, SHIFT_n_4_33_port, 
      SHIFT_n_4_32_port, SHIFT_n_4_31_port, SHIFT_n_4_30_port, 
      SHIFT_n_4_29_port, SHIFT_n_4_28_port, SHIFT_n_4_27_port, 
      SHIFT_n_4_26_port, SHIFT_n_4_25_port, SHIFT_n_4_24_port, 
      SHIFT_n_4_23_port, SHIFT_n_4_22_port, SHIFT_n_4_21_port, 
      SHIFT_n_4_20_port, SHIFT_n_4_19_port, SHIFT_n_4_18_port, 
      SHIFT_n_4_17_port, SHIFT_n_4_16_port, SHIFT_n_4_15_port, 
      SHIFT_n_4_14_port, SHIFT_n_4_13_port, SHIFT_n_4_12_port, 
      SHIFT_n_4_11_port, SHIFT_n_4_10_port, SHIFT_n_4_9_port, SHIFT_n_4_8_port,
      SHIFT_n_4_7_port, SHIFT_n_4_6_port, SHIFT_n_4_5_port, SHIFT_n_4_4_port, 
      SHIFT_n_4_3_port, SHIFT_n_4_2_port, SHIFT_n_4_1_port, SHIFT_n_4_0_port, 
      SHIFT_n_3_37_port, SHIFT_n_3_36_port, SHIFT_n_3_35_port, 
      SHIFT_n_3_34_port, SHIFT_n_3_33_port, SHIFT_n_3_32_port, 
      SHIFT_n_3_31_port, SHIFT_n_3_30_port, SHIFT_n_3_29_port, 
      SHIFT_n_3_28_port, SHIFT_n_3_27_port, SHIFT_n_3_26_port, 
      SHIFT_n_3_25_port, SHIFT_n_3_24_port, SHIFT_n_3_23_port, 
      SHIFT_n_3_22_port, SHIFT_n_3_21_port, SHIFT_n_3_20_port, 
      SHIFT_n_3_19_port, SHIFT_n_3_18_port, SHIFT_n_3_17_port, 
      SHIFT_n_3_16_port, SHIFT_n_3_15_port, SHIFT_n_3_14_port, 
      SHIFT_n_3_13_port, SHIFT_n_3_12_port, SHIFT_n_3_11_port, 
      SHIFT_n_3_10_port, SHIFT_n_3_9_port, SHIFT_n_3_8_port, SHIFT_n_3_7_port, 
      SHIFT_n_3_6_port, SHIFT_n_3_5_port, SHIFT_n_3_4_port, SHIFT_n_3_3_port, 
      SHIFT_n_3_2_port, SHIFT_n_3_1_port, SHIFT_n_3_0_port, SHIFT_n_2_35_port, 
      SHIFT_n_2_34_port, SHIFT_n_2_33_port, SHIFT_n_2_32_port, 
      SHIFT_n_2_31_port, SHIFT_n_2_30_port, SHIFT_n_2_29_port, 
      SHIFT_n_2_28_port, SHIFT_n_2_27_port, SHIFT_n_2_26_port, 
      SHIFT_n_2_25_port, SHIFT_n_2_24_port, SHIFT_n_2_23_port, 
      SHIFT_n_2_22_port, SHIFT_n_2_21_port, SHIFT_n_2_20_port, 
      SHIFT_n_2_19_port, SHIFT_n_2_18_port, SHIFT_n_2_17_port, 
      SHIFT_n_2_16_port, SHIFT_n_2_15_port, SHIFT_n_2_14_port, 
      SHIFT_n_2_13_port, SHIFT_n_2_12_port, SHIFT_n_2_11_port, 
      SHIFT_n_2_10_port, SHIFT_n_2_9_port, SHIFT_n_2_8_port, SHIFT_n_2_7_port, 
      SHIFT_n_2_6_port, SHIFT_n_2_5_port, SHIFT_n_2_4_port, SHIFT_n_2_3_port, 
      SHIFT_n_2_2_port, SHIFT_n_2_1_port, SHIFT_n_2_0_port, SHIFT_n_1_33_port, 
      SHIFT_n_1_32_port, OTMP_8_15_port, OTMP_8_14_port, OTMP_8_13_port, 
      OTMP_8_12_port, OTMP_8_11_port, OTMP_8_10_port, OTMP_8_9_port, 
      OTMP_8_8_port, OTMP_8_7_port, OTMP_8_6_port, OTMP_8_5_port, OTMP_8_4_port
      , OTMP_8_3_port, OTMP_8_2_port, OTMP_8_1_port, OTMP_8_0_port, 
      OTMP_7_47_port, OTMP_7_46_port, OTMP_7_45_port, OTMP_7_44_port, 
      OTMP_7_43_port, OTMP_7_42_port, OTMP_7_41_port, OTMP_7_40_port, 
      OTMP_7_39_port, OTMP_7_38_port, OTMP_7_37_port, OTMP_7_36_port, 
      OTMP_7_35_port, OTMP_7_34_port, OTMP_7_33_port, OTMP_7_32_port, 
      OTMP_7_31_port, OTMP_7_30_port, OTMP_7_29_port, OTMP_7_28_port, 
      OTMP_7_27_port, OTMP_7_26_port, OTMP_7_25_port, OTMP_7_24_port, 
      OTMP_7_23_port, OTMP_7_22_port, OTMP_7_21_port, OTMP_7_20_port, 
      OTMP_7_19_port, OTMP_7_18_port, OTMP_7_17_port, OTMP_7_16_port, 
      OTMP_7_15_port, OTMP_7_14_port, OTMP_7_13_port, OTMP_7_12_port, 
      OTMP_7_11_port, OTMP_7_10_port, OTMP_7_9_port, OTMP_7_8_port, 
      OTMP_7_7_port, OTMP_7_6_port, OTMP_7_5_port, OTMP_7_4_port, OTMP_7_3_port
      , OTMP_7_2_port, OTMP_7_1_port, OTMP_7_0_port, OTMP_6_45_port, 
      OTMP_6_44_port, OTMP_6_43_port, OTMP_6_42_port, OTMP_6_41_port, 
      OTMP_6_40_port, OTMP_6_39_port, OTMP_6_38_port, OTMP_6_37_port, 
      OTMP_6_36_port, OTMP_6_35_port, OTMP_6_34_port, OTMP_6_33_port, 
      OTMP_6_32_port, OTMP_6_31_port, OTMP_6_30_port, OTMP_6_29_port, 
      OTMP_6_28_port, OTMP_6_27_port, OTMP_6_26_port, OTMP_6_25_port, 
      OTMP_6_24_port, OTMP_6_23_port, OTMP_6_22_port, OTMP_6_21_port, 
      OTMP_6_20_port, OTMP_6_19_port, OTMP_6_18_port, OTMP_6_17_port, 
      OTMP_6_16_port, OTMP_6_15_port, OTMP_6_14_port, OTMP_6_13_port, 
      OTMP_6_12_port, OTMP_6_11_port, OTMP_6_10_port, OTMP_6_9_port, 
      OTMP_6_8_port, OTMP_6_7_port, OTMP_6_6_port, OTMP_6_5_port, OTMP_6_4_port
      , OTMP_6_3_port, OTMP_6_2_port, OTMP_6_1_port, OTMP_6_0_port, 
      OTMP_5_43_port, OTMP_5_42_port, OTMP_5_41_port, OTMP_5_40_port, 
      OTMP_5_39_port, OTMP_5_38_port, OTMP_5_37_port, OTMP_5_36_port, 
      OTMP_5_35_port, OTMP_5_34_port, OTMP_5_33_port, OTMP_5_32_port, 
      OTMP_5_31_port, OTMP_5_30_port, OTMP_5_29_port, OTMP_5_28_port, 
      OTMP_5_27_port, OTMP_5_26_port, OTMP_5_25_port, OTMP_5_24_port, 
      OTMP_5_23_port, OTMP_5_22_port, OTMP_5_21_port, OTMP_5_20_port, 
      OTMP_5_19_port, OTMP_5_18_port, OTMP_5_17_port, OTMP_5_16_port, 
      OTMP_5_15_port, OTMP_5_14_port, OTMP_5_13_port, OTMP_5_12_port, 
      OTMP_5_11_port, OTMP_5_10_port, OTMP_5_9_port, OTMP_5_8_port, 
      OTMP_5_7_port, OTMP_5_6_port, OTMP_5_5_port, OTMP_5_4_port, OTMP_5_3_port
      , OTMP_5_2_port, OTMP_5_1_port, OTMP_5_0_port, OTMP_4_41_port, 
      OTMP_4_40_port, OTMP_4_39_port, OTMP_4_38_port, OTMP_4_37_port, 
      OTMP_4_36_port, OTMP_4_35_port, OTMP_4_34_port, OTMP_4_33_port, 
      OTMP_4_32_port, OTMP_4_31_port, OTMP_4_30_port, OTMP_4_29_port, 
      OTMP_4_28_port, OTMP_4_27_port, OTMP_4_26_port, OTMP_4_25_port, 
      OTMP_4_24_port, OTMP_4_23_port, OTMP_4_22_port, OTMP_4_21_port, 
      OTMP_4_20_port, OTMP_4_19_port, OTMP_4_18_port, OTMP_4_17_port, 
      OTMP_4_16_port, OTMP_4_15_port, OTMP_4_14_port, OTMP_4_13_port, 
      OTMP_4_12_port, OTMP_4_11_port, OTMP_4_10_port, OTMP_4_9_port, 
      OTMP_4_8_port, OTMP_4_7_port, OTMP_4_6_port, OTMP_4_5_port, OTMP_4_4_port
      , OTMP_4_3_port, OTMP_4_2_port, OTMP_4_1_port, OTMP_4_0_port, 
      OTMP_3_39_port, OTMP_3_38_port, OTMP_3_37_port, OTMP_3_36_port, 
      OTMP_3_35_port, OTMP_3_34_port, OTMP_3_33_port, OTMP_3_32_port, 
      OTMP_3_31_port, OTMP_3_30_port, OTMP_3_29_port, OTMP_3_28_port, 
      OTMP_3_27_port, OTMP_3_26_port, OTMP_3_25_port, OTMP_3_24_port, 
      OTMP_3_23_port, OTMP_3_22_port, OTMP_3_21_port, OTMP_3_20_port, 
      OTMP_3_19_port, OTMP_3_18_port, OTMP_3_17_port, OTMP_3_16_port, 
      OTMP_3_15_port, OTMP_3_14_port, OTMP_3_13_port, OTMP_3_12_port, 
      OTMP_3_11_port, OTMP_3_10_port, OTMP_3_9_port, OTMP_3_8_port, 
      OTMP_3_7_port, OTMP_3_6_port, OTMP_3_5_port, OTMP_3_4_port, OTMP_3_3_port
      , OTMP_3_2_port, OTMP_3_1_port, OTMP_3_0_port, OTMP_2_37_port, 
      OTMP_2_36_port, OTMP_2_35_port, OTMP_2_34_port, OTMP_2_33_port, 
      OTMP_2_32_port, OTMP_2_31_port, OTMP_2_30_port, OTMP_2_29_port, 
      OTMP_2_28_port, OTMP_2_27_port, OTMP_2_26_port, OTMP_2_25_port, 
      OTMP_2_24_port, OTMP_2_23_port, OTMP_2_22_port, OTMP_2_21_port, 
      OTMP_2_20_port, OTMP_2_19_port, OTMP_2_18_port, OTMP_2_17_port, 
      OTMP_2_16_port, OTMP_2_15_port, OTMP_2_14_port, OTMP_2_13_port, 
      OTMP_2_12_port, OTMP_2_11_port, OTMP_2_10_port, OTMP_2_9_port, 
      OTMP_2_8_port, OTMP_2_7_port, OTMP_2_6_port, OTMP_2_5_port, OTMP_2_4_port
      , OTMP_2_3_port, OTMP_2_2_port, OTMP_2_1_port, OTMP_2_0_port, 
      OTMP_1_35_port, OTMP_1_34_port, OTMP_1_33_port, OTMP_1_32_port, 
      OTMP_1_31_port, OTMP_1_30_port, OTMP_1_29_port, OTMP_1_28_port, 
      OTMP_1_27_port, OTMP_1_26_port, OTMP_1_25_port, OTMP_1_24_port, 
      OTMP_1_23_port, OTMP_1_22_port, OTMP_1_21_port, OTMP_1_20_port, 
      OTMP_1_19_port, OTMP_1_18_port, OTMP_1_17_port, OTMP_1_16_port, 
      OTMP_1_15_port, OTMP_1_14_port, OTMP_1_13_port, OTMP_1_12_port, 
      OTMP_1_11_port, OTMP_1_10_port, OTMP_1_9_port, OTMP_1_8_port, 
      OTMP_1_7_port, OTMP_1_6_port, OTMP_1_5_port, OTMP_1_4_port, OTMP_1_3_port
      , OTMP_1_2_port, OTMP_1_1_port, OTMP_1_0_port, OTMP_0_34_port, 
      OTMP_0_32_port, OTMP_0_31_port, OTMP_0_30_port, OTMP_0_29_port, 
      OTMP_0_28_port, OTMP_0_27_port, OTMP_0_26_port, OTMP_0_25_port, 
      OTMP_0_24_port, OTMP_0_23_port, OTMP_0_22_port, OTMP_0_21_port, 
      OTMP_0_20_port, OTMP_0_19_port, OTMP_0_18_port, OTMP_0_17_port, 
      OTMP_0_16_port, OTMP_0_15_port, OTMP_0_14_port, OTMP_0_13_port, 
      OTMP_0_12_port, OTMP_0_11_port, OTMP_0_10_port, OTMP_0_9_port, 
      OTMP_0_8_port, OTMP_0_7_port, OTMP_0_6_port, OTMP_0_5_port, OTMP_0_4_port
      , OTMP_0_3_port, OTMP_0_2_port, OTMP_0_1_port, OTMP_0_0_port, 
      OTMP_15_63_port, OTMP_15_62_port, OTMP_15_61_port, OTMP_15_60_port, 
      OTMP_15_59_port, OTMP_15_58_port, OTMP_15_57_port, OTMP_15_56_port, 
      OTMP_15_55_port, OTMP_15_54_port, OTMP_15_53_port, OTMP_15_52_port, 
      OTMP_15_51_port, OTMP_15_50_port, OTMP_15_49_port, OTMP_15_48_port, 
      OTMP_15_47_port, OTMP_15_46_port, OTMP_15_45_port, OTMP_15_44_port, 
      OTMP_15_43_port, OTMP_15_42_port, OTMP_15_41_port, OTMP_15_40_port, 
      OTMP_15_39_port, OTMP_15_38_port, OTMP_15_37_port, OTMP_15_36_port, 
      OTMP_15_35_port, OTMP_15_34_port, OTMP_15_33_port, OTMP_15_32_port, 
      OTMP_15_31_port, OTMP_15_30_port, OTMP_15_29_port, OTMP_15_28_port, 
      OTMP_15_27_port, OTMP_15_26_port, OTMP_15_25_port, OTMP_15_24_port, 
      OTMP_15_23_port, OTMP_15_22_port, OTMP_15_21_port, OTMP_15_20_port, 
      OTMP_15_19_port, OTMP_15_18_port, OTMP_15_17_port, OTMP_15_16_port, 
      OTMP_15_15_port, OTMP_15_14_port, OTMP_15_13_port, OTMP_15_12_port, 
      OTMP_15_11_port, OTMP_15_10_port, OTMP_15_9_port, OTMP_15_8_port, 
      OTMP_15_7_port, OTMP_15_6_port, OTMP_15_5_port, OTMP_15_4_port, 
      OTMP_15_3_port, OTMP_15_2_port, OTMP_15_1_port, OTMP_15_0_port, 
      OTMP_14_61_port, OTMP_14_60_port, OTMP_14_59_port, OTMP_14_58_port, 
      OTMP_14_57_port, OTMP_14_56_port, OTMP_14_55_port, OTMP_14_54_port, 
      OTMP_14_53_port, OTMP_14_52_port, OTMP_14_51_port, OTMP_14_50_port, 
      OTMP_14_49_port, OTMP_14_48_port, OTMP_14_47_port, OTMP_14_46_port, 
      OTMP_14_45_port, OTMP_14_44_port, OTMP_14_43_port, OTMP_14_42_port, 
      OTMP_14_41_port, OTMP_14_40_port, OTMP_14_39_port, OTMP_14_38_port, 
      OTMP_14_37_port, OTMP_14_36_port, OTMP_14_35_port, OTMP_14_34_port, 
      OTMP_14_33_port, OTMP_14_32_port, OTMP_14_31_port, OTMP_14_30_port, 
      OTMP_14_29_port, OTMP_14_28_port, OTMP_14_27_port, OTMP_14_26_port, 
      OTMP_14_25_port, OTMP_14_24_port, OTMP_14_23_port, OTMP_14_22_port, 
      OTMP_14_21_port, OTMP_14_20_port, OTMP_14_19_port, OTMP_14_18_port, 
      OTMP_14_17_port, OTMP_14_16_port, OTMP_14_15_port, OTMP_14_14_port, 
      OTMP_14_13_port, OTMP_14_12_port, OTMP_14_11_port, OTMP_14_10_port, 
      OTMP_14_9_port, OTMP_14_8_port, OTMP_14_7_port, OTMP_14_6_port, 
      OTMP_14_5_port, OTMP_14_4_port, OTMP_14_3_port, OTMP_14_2_port, 
      OTMP_14_1_port, OTMP_14_0_port, OTMP_13_59_port, OTMP_13_58_port, 
      OTMP_13_57_port, OTMP_13_56_port, OTMP_13_55_port, OTMP_13_54_port, 
      OTMP_13_53_port, OTMP_13_52_port, OTMP_13_51_port, OTMP_13_50_port, 
      OTMP_13_49_port, OTMP_13_48_port, OTMP_13_47_port, OTMP_13_46_port, 
      OTMP_13_45_port, OTMP_13_44_port, OTMP_13_43_port, OTMP_13_42_port, 
      OTMP_13_41_port, OTMP_13_40_port, OTMP_13_39_port, OTMP_13_38_port, 
      OTMP_13_37_port, OTMP_13_36_port, OTMP_13_35_port, OTMP_13_34_port, 
      OTMP_13_33_port, OTMP_13_32_port, OTMP_13_31_port, OTMP_13_30_port, 
      OTMP_13_29_port, OTMP_13_28_port, OTMP_13_27_port, OTMP_13_26_port, 
      OTMP_13_25_port, OTMP_13_24_port, OTMP_13_23_port, OTMP_13_22_port, 
      OTMP_13_21_port, OTMP_13_20_port, OTMP_13_19_port, OTMP_13_18_port, 
      OTMP_13_17_port, OTMP_13_16_port, OTMP_13_15_port, OTMP_13_14_port, 
      OTMP_13_13_port, OTMP_13_12_port, OTMP_13_11_port, OTMP_13_10_port, 
      OTMP_13_9_port, OTMP_13_8_port, OTMP_13_7_port, OTMP_13_6_port, 
      OTMP_13_5_port, OTMP_13_4_port, OTMP_13_3_port, OTMP_13_2_port, 
      OTMP_13_1_port, OTMP_13_0_port, OTMP_12_57_port, OTMP_12_56_port, 
      OTMP_12_55_port, OTMP_12_54_port, OTMP_12_53_port, OTMP_12_52_port, 
      OTMP_12_51_port, OTMP_12_50_port, OTMP_12_49_port, OTMP_12_48_port, 
      OTMP_12_47_port, OTMP_12_46_port, OTMP_12_45_port, OTMP_12_44_port, 
      OTMP_12_43_port, OTMP_12_42_port, OTMP_12_41_port, OTMP_12_40_port, 
      OTMP_12_39_port, OTMP_12_38_port, OTMP_12_37_port, OTMP_12_36_port, 
      OTMP_12_35_port, OTMP_12_34_port, OTMP_12_33_port, OTMP_12_32_port, 
      OTMP_12_31_port, OTMP_12_30_port, OTMP_12_29_port, OTMP_12_28_port, 
      OTMP_12_27_port, OTMP_12_26_port, OTMP_12_25_port, OTMP_12_24_port, 
      OTMP_12_23_port, OTMP_12_22_port, OTMP_12_21_port, OTMP_12_20_port, 
      OTMP_12_19_port, OTMP_12_18_port, OTMP_12_17_port, OTMP_12_16_port, 
      OTMP_12_15_port, OTMP_12_14_port, OTMP_12_13_port, OTMP_12_12_port, 
      OTMP_12_11_port, OTMP_12_10_port, OTMP_12_9_port, OTMP_12_8_port, 
      OTMP_12_7_port, OTMP_12_6_port, OTMP_12_5_port, OTMP_12_4_port, 
      OTMP_12_3_port, OTMP_12_2_port, OTMP_12_1_port, OTMP_12_0_port, 
      OTMP_11_55_port, OTMP_11_54_port, OTMP_11_53_port, OTMP_11_52_port, 
      OTMP_11_51_port, OTMP_11_50_port, OTMP_11_49_port, OTMP_11_48_port, 
      OTMP_11_47_port, OTMP_11_46_port, OTMP_11_45_port, OTMP_11_44_port, 
      OTMP_11_43_port, OTMP_11_42_port, OTMP_11_41_port, OTMP_11_40_port, 
      OTMP_11_39_port, OTMP_11_38_port, OTMP_11_37_port, OTMP_11_36_port, 
      OTMP_11_35_port, OTMP_11_34_port, OTMP_11_33_port, OTMP_11_32_port, 
      OTMP_11_31_port, OTMP_11_30_port, OTMP_11_29_port, OTMP_11_28_port, 
      OTMP_11_27_port, OTMP_11_26_port, OTMP_11_25_port, OTMP_11_24_port, 
      OTMP_11_23_port, OTMP_11_22_port, OTMP_11_21_port, OTMP_11_20_port, 
      OTMP_11_19_port, OTMP_11_18_port, OTMP_11_17_port, OTMP_11_16_port, 
      OTMP_11_15_port, OTMP_11_14_port, OTMP_11_13_port, OTMP_11_12_port, 
      OTMP_11_11_port, OTMP_11_10_port, OTMP_11_9_port, OTMP_11_8_port, 
      OTMP_11_7_port, OTMP_11_6_port, OTMP_11_5_port, OTMP_11_4_port, 
      OTMP_11_3_port, OTMP_11_2_port, OTMP_11_1_port, OTMP_11_0_port, 
      OTMP_10_53_port, OTMP_10_52_port, OTMP_10_51_port, OTMP_10_50_port, 
      OTMP_10_49_port, OTMP_10_48_port, OTMP_10_47_port, OTMP_10_46_port, 
      OTMP_10_45_port, OTMP_10_44_port, OTMP_10_43_port, OTMP_10_42_port, 
      OTMP_10_41_port, OTMP_10_40_port, OTMP_10_39_port, OTMP_10_38_port, 
      OTMP_10_37_port, OTMP_10_36_port, OTMP_10_35_port, OTMP_10_34_port, 
      OTMP_10_33_port, OTMP_10_32_port, OTMP_10_31_port, OTMP_10_30_port, 
      OTMP_10_29_port, OTMP_10_28_port, OTMP_10_27_port, OTMP_10_26_port, 
      OTMP_10_25_port, OTMP_10_24_port, OTMP_10_23_port, OTMP_10_22_port, 
      OTMP_10_21_port, OTMP_10_20_port, OTMP_10_19_port, OTMP_10_18_port, 
      OTMP_10_17_port, OTMP_10_16_port, OTMP_10_15_port, OTMP_10_14_port, 
      OTMP_10_13_port, OTMP_10_12_port, OTMP_10_11_port, OTMP_10_10_port, 
      OTMP_10_9_port, OTMP_10_8_port, OTMP_10_7_port, OTMP_10_6_port, 
      OTMP_10_5_port, OTMP_10_4_port, OTMP_10_3_port, OTMP_10_2_port, 
      OTMP_10_1_port, OTMP_10_0_port, OTMP_9_51_port, OTMP_9_50_port, 
      OTMP_9_49_port, OTMP_9_48_port, OTMP_9_47_port, OTMP_9_46_port, 
      OTMP_9_45_port, OTMP_9_44_port, OTMP_9_43_port, OTMP_9_42_port, 
      OTMP_9_41_port, OTMP_9_40_port, OTMP_9_39_port, OTMP_9_38_port, 
      OTMP_9_37_port, OTMP_9_36_port, OTMP_9_35_port, OTMP_9_34_port, 
      OTMP_9_33_port, OTMP_9_32_port, OTMP_9_31_port, OTMP_9_30_port, 
      OTMP_9_29_port, OTMP_9_28_port, OTMP_9_27_port, OTMP_9_26_port, 
      OTMP_9_25_port, OTMP_9_24_port, OTMP_9_23_port, OTMP_9_22_port, 
      OTMP_9_21_port, OTMP_9_20_port, OTMP_9_19_port, OTMP_9_18_port, 
      OTMP_9_17_port, OTMP_9_16_port, OTMP_9_15_port, OTMP_9_14_port, 
      OTMP_9_13_port, OTMP_9_12_port, OTMP_9_11_port, OTMP_9_10_port, 
      OTMP_9_9_port, OTMP_9_8_port, OTMP_9_7_port, OTMP_9_6_port, OTMP_9_5_port
      , OTMP_9_4_port, OTMP_9_3_port, OTMP_9_2_port, OTMP_9_1_port, 
      OTMP_9_0_port, OTMP_8_49_port, OTMP_8_48_port, OTMP_8_47_port, 
      OTMP_8_46_port, OTMP_8_45_port, OTMP_8_44_port, OTMP_8_43_port, 
      OTMP_8_42_port, OTMP_8_41_port, OTMP_8_40_port, OTMP_8_39_port, 
      OTMP_8_38_port, OTMP_8_37_port, OTMP_8_36_port, OTMP_8_35_port, 
      OTMP_8_34_port, OTMP_8_33_port, OTMP_8_32_port, OTMP_8_31_port, 
      OTMP_8_30_port, OTMP_8_29_port, OTMP_8_28_port, OTMP_8_27_port, 
      OTMP_8_26_port, OTMP_8_25_port, OTMP_8_24_port, OTMP_8_23_port, 
      OTMP_8_22_port, OTMP_8_21_port, OTMP_8_20_port, OTMP_8_19_port, 
      OTMP_8_18_port, OTMP_8_17_port, OTMP_8_16_port, PTMP_8_15_port, 
      PTMP_8_14_port, PTMP_8_13_port, PTMP_8_12_port, PTMP_8_11_port, 
      PTMP_8_10_port, PTMP_8_9_port, PTMP_8_8_port, PTMP_8_7_port, 
      PTMP_8_6_port, PTMP_8_5_port, PTMP_8_4_port, PTMP_8_3_port, PTMP_8_2_port
      , PTMP_8_1_port, PTMP_8_0_port, PTMP_7_49_port, PTMP_7_48_port, 
      PTMP_7_47_port, PTMP_7_46_port, PTMP_7_45_port, PTMP_7_44_port, 
      PTMP_7_43_port, PTMP_7_42_port, PTMP_7_41_port, PTMP_7_40_port, 
      PTMP_7_39_port, PTMP_7_38_port, PTMP_7_37_port, PTMP_7_36_port, 
      PTMP_7_35_port, PTMP_7_34_port, PTMP_7_33_port, PTMP_7_32_port, 
      PTMP_7_31_port, PTMP_7_30_port, PTMP_7_29_port, PTMP_7_28_port, 
      PTMP_7_27_port, PTMP_7_26_port, PTMP_7_25_port, PTMP_7_24_port, 
      PTMP_7_23_port, PTMP_7_22_port, PTMP_7_21_port, PTMP_7_20_port, 
      PTMP_7_19_port, PTMP_7_18_port, PTMP_7_17_port, PTMP_7_16_port, 
      PTMP_7_15_port, PTMP_7_14_port, PTMP_7_13_port, PTMP_7_12_port, 
      PTMP_7_11_port, PTMP_7_10_port, PTMP_7_9_port, PTMP_7_8_port, 
      PTMP_7_7_port, PTMP_7_6_port, PTMP_7_5_port, PTMP_7_4_port, PTMP_7_3_port
      , PTMP_7_2_port, PTMP_7_1_port, PTMP_7_0_port, PTMP_6_47_port, 
      PTMP_6_46_port, PTMP_6_45_port, PTMP_6_44_port, PTMP_6_43_port, 
      PTMP_6_42_port, PTMP_6_41_port, PTMP_6_40_port, PTMP_6_39_port, 
      PTMP_6_38_port, PTMP_6_37_port, PTMP_6_36_port, PTMP_6_35_port, 
      PTMP_6_34_port, PTMP_6_33_port, PTMP_6_32_port, PTMP_6_31_port, 
      PTMP_6_30_port, PTMP_6_29_port, PTMP_6_28_port, PTMP_6_27_port, 
      PTMP_6_26_port, PTMP_6_25_port, PTMP_6_24_port, PTMP_6_23_port, 
      PTMP_6_22_port, PTMP_6_21_port, PTMP_6_20_port, PTMP_6_19_port, 
      PTMP_6_18_port, PTMP_6_17_port, PTMP_6_16_port, PTMP_6_15_port, 
      PTMP_6_14_port, PTMP_6_13_port, PTMP_6_12_port, PTMP_6_11_port, 
      PTMP_6_10_port, PTMP_6_9_port, PTMP_6_8_port, PTMP_6_7_port, 
      PTMP_6_6_port, PTMP_6_5_port, PTMP_6_4_port, PTMP_6_3_port, PTMP_6_2_port
      , PTMP_6_1_port, PTMP_6_0_port, PTMP_5_45_port, PTMP_5_44_port, 
      PTMP_5_43_port, PTMP_5_42_port, PTMP_5_41_port, PTMP_5_40_port, 
      PTMP_5_39_port, PTMP_5_38_port, PTMP_5_37_port, PTMP_5_36_port, 
      PTMP_5_35_port, PTMP_5_34_port, PTMP_5_33_port, PTMP_5_32_port, 
      PTMP_5_31_port, PTMP_5_30_port, PTMP_5_29_port, PTMP_5_28_port, 
      PTMP_5_27_port, PTMP_5_26_port, PTMP_5_25_port, PTMP_5_24_port, 
      PTMP_5_23_port, PTMP_5_22_port, PTMP_5_21_port, PTMP_5_20_port, 
      PTMP_5_19_port, PTMP_5_18_port, PTMP_5_17_port, PTMP_5_16_port, 
      PTMP_5_15_port, PTMP_5_14_port, PTMP_5_13_port, PTMP_5_12_port, 
      PTMP_5_11_port, PTMP_5_10_port, PTMP_5_9_port, PTMP_5_8_port, 
      PTMP_5_7_port, PTMP_5_6_port, PTMP_5_5_port, PTMP_5_4_port, PTMP_5_3_port
      , PTMP_5_2_port, PTMP_5_1_port, PTMP_5_0_port, PTMP_4_43_port, 
      PTMP_4_42_port, PTMP_4_41_port, PTMP_4_40_port, PTMP_4_39_port, 
      PTMP_4_38_port, PTMP_4_37_port, PTMP_4_36_port, PTMP_4_35_port, 
      PTMP_4_34_port, PTMP_4_33_port, PTMP_4_32_port, PTMP_4_31_port, 
      PTMP_4_30_port, PTMP_4_29_port, PTMP_4_28_port, PTMP_4_27_port, 
      PTMP_4_26_port, PTMP_4_25_port, PTMP_4_24_port, PTMP_4_23_port, 
      PTMP_4_22_port, PTMP_4_21_port, PTMP_4_20_port, PTMP_4_19_port, 
      PTMP_4_18_port, PTMP_4_17_port, PTMP_4_16_port, PTMP_4_15_port, 
      PTMP_4_14_port, PTMP_4_13_port, PTMP_4_12_port, PTMP_4_11_port, 
      PTMP_4_10_port, PTMP_4_9_port, PTMP_4_8_port, PTMP_4_7_port, 
      PTMP_4_6_port, PTMP_4_5_port, PTMP_4_4_port, PTMP_4_3_port, PTMP_4_2_port
      , PTMP_4_1_port, PTMP_4_0_port, PTMP_3_41_port, PTMP_3_40_port, 
      PTMP_3_39_port, PTMP_3_38_port, PTMP_3_37_port, PTMP_3_36_port, 
      PTMP_3_35_port, PTMP_3_34_port, PTMP_3_33_port, PTMP_3_32_port, 
      PTMP_3_31_port, PTMP_3_30_port, PTMP_3_29_port, PTMP_3_28_port, 
      PTMP_3_27_port, PTMP_3_26_port, PTMP_3_25_port, PTMP_3_24_port, 
      PTMP_3_23_port, PTMP_3_22_port, PTMP_3_21_port, PTMP_3_20_port, 
      PTMP_3_19_port, PTMP_3_18_port, PTMP_3_17_port, PTMP_3_16_port, 
      PTMP_3_15_port, PTMP_3_14_port, PTMP_3_13_port, PTMP_3_12_port, 
      PTMP_3_11_port, PTMP_3_10_port, PTMP_3_9_port, PTMP_3_8_port, 
      PTMP_3_7_port, PTMP_3_6_port, PTMP_3_5_port, PTMP_3_4_port, PTMP_3_3_port
      , PTMP_3_2_port, PTMP_3_1_port, PTMP_3_0_port, PTMP_2_39_port, 
      PTMP_2_38_port, PTMP_2_37_port, PTMP_2_36_port, PTMP_2_35_port, 
      PTMP_2_34_port, PTMP_2_33_port, PTMP_2_32_port, PTMP_2_31_port, 
      PTMP_2_30_port, PTMP_2_29_port, PTMP_2_28_port, PTMP_2_27_port, 
      PTMP_2_26_port, PTMP_2_25_port, PTMP_2_24_port, PTMP_2_23_port, 
      PTMP_2_22_port, PTMP_2_21_port, PTMP_2_20_port, PTMP_2_19_port, 
      PTMP_2_18_port, PTMP_2_17_port, PTMP_2_16_port, PTMP_2_15_port, 
      PTMP_2_14_port, PTMP_2_13_port, PTMP_2_12_port, PTMP_2_11_port, 
      PTMP_2_10_port, PTMP_2_9_port, PTMP_2_8_port, PTMP_2_7_port, 
      PTMP_2_6_port, PTMP_2_5_port, PTMP_2_4_port, PTMP_2_3_port, PTMP_2_2_port
      , PTMP_2_1_port, PTMP_2_0_port, PTMP_1_37_port, PTMP_1_36_port, 
      PTMP_1_35_port, PTMP_1_34_port, PTMP_1_33_port, PTMP_1_32_port, 
      PTMP_1_31_port, PTMP_1_30_port, PTMP_1_29_port, PTMP_1_28_port, 
      PTMP_1_27_port, PTMP_1_26_port, PTMP_1_25_port, PTMP_1_24_port, 
      PTMP_1_23_port, PTMP_1_22_port, PTMP_1_21_port, PTMP_1_20_port, 
      PTMP_1_19_port, PTMP_1_18_port, PTMP_1_17_port, PTMP_1_16_port, 
      PTMP_1_15_port, PTMP_1_14_port, PTMP_1_13_port, PTMP_1_12_port, 
      PTMP_1_11_port, PTMP_1_10_port, PTMP_1_9_port, PTMP_1_8_port, 
      PTMP_1_7_port, PTMP_1_6_port, PTMP_1_5_port, PTMP_1_4_port, PTMP_1_3_port
      , PTMP_1_2_port, PTMP_1_1_port, PTMP_1_0_port, PTMP_0_36_port, 
      PTMP_0_34_port, PTMP_0_33_port, PTMP_0_32_port, PTMP_0_31_port, 
      PTMP_0_30_port, PTMP_0_29_port, PTMP_0_28_port, PTMP_0_27_port, 
      PTMP_0_26_port, PTMP_0_25_port, PTMP_0_24_port, PTMP_0_23_port, 
      PTMP_0_22_port, PTMP_0_21_port, PTMP_0_20_port, PTMP_0_19_port, 
      PTMP_0_18_port, PTMP_0_17_port, PTMP_0_16_port, PTMP_0_15_port, 
      PTMP_0_14_port, PTMP_0_13_port, PTMP_0_12_port, PTMP_0_11_port, 
      PTMP_0_10_port, PTMP_0_9_port, PTMP_0_8_port, PTMP_0_7_port, 
      PTMP_0_6_port, PTMP_0_5_port, PTMP_0_4_port, PTMP_0_3_port, PTMP_0_2_port
      , PTMP_0_1_port, PTMP_0_0_port, PTMP_13_61_port, PTMP_13_60_port, 
      PTMP_13_59_port, PTMP_13_58_port, PTMP_13_57_port, PTMP_13_56_port, 
      PTMP_13_55_port, PTMP_13_54_port, PTMP_13_53_port, PTMP_13_52_port, 
      PTMP_13_51_port, PTMP_13_50_port, PTMP_13_49_port, PTMP_13_48_port, 
      PTMP_13_47_port, PTMP_13_46_port, PTMP_13_45_port, PTMP_13_44_port, 
      PTMP_13_43_port, PTMP_13_42_port, PTMP_13_41_port, PTMP_13_40_port, 
      PTMP_13_39_port, PTMP_13_38_port, PTMP_13_37_port, PTMP_13_36_port, 
      PTMP_13_35_port, PTMP_13_34_port, PTMP_13_33_port, PTMP_13_32_port, 
      PTMP_13_31_port, PTMP_13_30_port, PTMP_13_29_port, PTMP_13_28_port, 
      PTMP_13_27_port, PTMP_13_26_port, PTMP_13_25_port, PTMP_13_24_port, 
      PTMP_13_23_port, PTMP_13_22_port, PTMP_13_21_port, PTMP_13_20_port, 
      PTMP_13_19_port, PTMP_13_18_port, PTMP_13_17_port, PTMP_13_16_port, 
      PTMP_13_15_port, PTMP_13_14_port, PTMP_13_13_port, PTMP_13_12_port, 
      PTMP_13_11_port, PTMP_13_10_port, PTMP_13_9_port, PTMP_13_8_port, 
      PTMP_13_7_port, PTMP_13_6_port, PTMP_13_5_port, PTMP_13_4_port, 
      PTMP_13_3_port, PTMP_13_2_port, PTMP_13_1_port, PTMP_13_0_port, 
      PTMP_12_59_port, PTMP_12_58_port, PTMP_12_57_port, PTMP_12_56_port, 
      PTMP_12_55_port, PTMP_12_54_port, PTMP_12_53_port, PTMP_12_52_port, 
      PTMP_12_51_port, PTMP_12_50_port, PTMP_12_49_port, PTMP_12_48_port, 
      PTMP_12_47_port, PTMP_12_46_port, PTMP_12_45_port, PTMP_12_44_port, 
      PTMP_12_43_port, PTMP_12_42_port, PTMP_12_41_port, PTMP_12_40_port, 
      PTMP_12_39_port, PTMP_12_38_port, PTMP_12_37_port, PTMP_12_36_port, 
      PTMP_12_35_port, PTMP_12_34_port, PTMP_12_33_port, PTMP_12_32_port, 
      PTMP_12_31_port, PTMP_12_30_port, PTMP_12_29_port, PTMP_12_28_port, 
      PTMP_12_27_port, PTMP_12_26_port, PTMP_12_25_port, PTMP_12_24_port, 
      PTMP_12_23_port, PTMP_12_22_port, PTMP_12_21_port, PTMP_12_20_port, 
      PTMP_12_19_port, PTMP_12_18_port, PTMP_12_17_port, PTMP_12_16_port, 
      PTMP_12_15_port, PTMP_12_14_port, PTMP_12_13_port, PTMP_12_12_port, 
      PTMP_12_11_port, PTMP_12_10_port, PTMP_12_9_port, PTMP_12_8_port, 
      PTMP_12_7_port, PTMP_12_6_port, PTMP_12_5_port, PTMP_12_4_port, 
      PTMP_12_3_port, PTMP_12_2_port, PTMP_12_1_port, PTMP_12_0_port, 
      PTMP_11_57_port, PTMP_11_56_port, PTMP_11_55_port, PTMP_11_54_port, 
      PTMP_11_53_port, PTMP_11_52_port, PTMP_11_51_port, PTMP_11_50_port, 
      PTMP_11_49_port, PTMP_11_48_port, PTMP_11_47_port, PTMP_11_46_port, 
      PTMP_11_45_port, PTMP_11_44_port, PTMP_11_43_port, PTMP_11_42_port, 
      PTMP_11_41_port, PTMP_11_40_port, PTMP_11_39_port, PTMP_11_38_port, 
      PTMP_11_37_port, PTMP_11_36_port, PTMP_11_35_port, PTMP_11_34_port, 
      PTMP_11_33_port, PTMP_11_32_port, PTMP_11_31_port, PTMP_11_30_port, 
      PTMP_11_29_port, PTMP_11_28_port, PTMP_11_27_port, PTMP_11_26_port, 
      PTMP_11_25_port, PTMP_11_24_port, PTMP_11_23_port, PTMP_11_22_port, 
      PTMP_11_21_port, PTMP_11_20_port, PTMP_11_19_port, PTMP_11_18_port, 
      PTMP_11_17_port, PTMP_11_16_port, PTMP_11_15_port, PTMP_11_14_port, 
      PTMP_11_13_port, PTMP_11_12_port, PTMP_11_11_port, PTMP_11_10_port, 
      PTMP_11_9_port, PTMP_11_8_port, PTMP_11_7_port, PTMP_11_6_port, 
      PTMP_11_5_port, PTMP_11_4_port, PTMP_11_3_port, PTMP_11_2_port, 
      PTMP_11_1_port, PTMP_11_0_port, PTMP_10_55_port, PTMP_10_54_port, 
      PTMP_10_53_port, PTMP_10_52_port, PTMP_10_51_port, PTMP_10_50_port, 
      PTMP_10_49_port, PTMP_10_48_port, PTMP_10_47_port, PTMP_10_46_port, 
      PTMP_10_45_port, PTMP_10_44_port, PTMP_10_43_port, PTMP_10_42_port, 
      PTMP_10_41_port, PTMP_10_40_port, PTMP_10_39_port, PTMP_10_38_port, 
      PTMP_10_37_port, PTMP_10_36_port, PTMP_10_35_port, PTMP_10_34_port, 
      PTMP_10_33_port, PTMP_10_32_port, PTMP_10_31_port, PTMP_10_30_port, 
      PTMP_10_29_port, PTMP_10_28_port, PTMP_10_27_port, PTMP_10_26_port, 
      PTMP_10_25_port, PTMP_10_24_port, PTMP_10_23_port, PTMP_10_22_port, 
      PTMP_10_21_port, PTMP_10_20_port, PTMP_10_19_port, PTMP_10_18_port, 
      PTMP_10_17_port, PTMP_10_16_port, PTMP_10_15_port, PTMP_10_14_port, 
      PTMP_10_13_port, PTMP_10_12_port, PTMP_10_11_port, PTMP_10_10_port, 
      PTMP_10_9_port, PTMP_10_8_port, PTMP_10_7_port, PTMP_10_6_port, 
      PTMP_10_5_port, PTMP_10_4_port, PTMP_10_3_port, PTMP_10_2_port, 
      PTMP_10_1_port, PTMP_10_0_port, PTMP_9_53_port, PTMP_9_52_port, 
      PTMP_9_51_port, PTMP_9_50_port, PTMP_9_49_port, PTMP_9_48_port, 
      PTMP_9_47_port, PTMP_9_46_port, PTMP_9_45_port, PTMP_9_44_port, 
      PTMP_9_43_port, PTMP_9_42_port, PTMP_9_41_port, PTMP_9_40_port, 
      PTMP_9_39_port, PTMP_9_38_port, PTMP_9_37_port, PTMP_9_36_port, 
      PTMP_9_35_port, PTMP_9_34_port, PTMP_9_33_port, PTMP_9_32_port, 
      PTMP_9_31_port, PTMP_9_30_port, PTMP_9_29_port, PTMP_9_28_port, 
      PTMP_9_27_port, PTMP_9_26_port, PTMP_9_25_port, PTMP_9_24_port, 
      PTMP_9_23_port, PTMP_9_22_port, PTMP_9_21_port, PTMP_9_20_port, 
      PTMP_9_19_port, PTMP_9_18_port, PTMP_9_17_port, PTMP_9_16_port, 
      PTMP_9_15_port, PTMP_9_14_port, PTMP_9_13_port, PTMP_9_12_port, 
      PTMP_9_11_port, PTMP_9_10_port, PTMP_9_9_port, PTMP_9_8_port, 
      PTMP_9_7_port, PTMP_9_6_port, PTMP_9_5_port, PTMP_9_4_port, PTMP_9_3_port
      , PTMP_9_2_port, PTMP_9_1_port, PTMP_9_0_port, PTMP_8_51_port, 
      PTMP_8_50_port, PTMP_8_49_port, PTMP_8_48_port, PTMP_8_47_port, 
      PTMP_8_46_port, PTMP_8_45_port, PTMP_8_44_port, PTMP_8_43_port, 
      PTMP_8_42_port, PTMP_8_41_port, PTMP_8_40_port, PTMP_8_39_port, 
      PTMP_8_38_port, PTMP_8_37_port, PTMP_8_36_port, PTMP_8_35_port, 
      PTMP_8_34_port, PTMP_8_33_port, PTMP_8_32_port, PTMP_8_31_port, 
      PTMP_8_30_port, PTMP_8_29_port, PTMP_8_28_port, PTMP_8_27_port, 
      PTMP_8_26_port, PTMP_8_25_port, PTMP_8_24_port, PTMP_8_23_port, 
      PTMP_8_22_port, PTMP_8_21_port, PTMP_8_20_port, PTMP_8_19_port, 
      PTMP_8_18_port, PTMP_8_17_port, PTMP_8_16_port, n4, n5, n6, n7, n8, n9, 
      n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n_1080, n_1081, n_1082,
      n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, 
      n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, 
      n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, 
      n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, 
      n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, 
      n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, 
      n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, 
      n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, 
      n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, 
      n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, 
      n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, 
      n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, 
      n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, 
      n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, 
      n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, 
      n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, 
      n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, 
      n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, 
      n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, 
      n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, 
      n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, 
      n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, 
      n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, 
      n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296 : std_logic;

begin
   
   X_Logic0_port <= '0';
   OTMP_15_0_port <= '0';
   SHIFT_n_15_0_port <= '0';
   SHIFT_n_15_1_port <= '0';
   SHIFT_15_0_port <= '0';
   SHIFT_15_1_port <= '0';
   OTMP_14_0_port <= '0';
   SHIFT_n_14_0_port <= '0';
   SHIFT_n_14_1_port <= '0';
   SHIFT_14_0_port <= '0';
   SHIFT_14_1_port <= '0';
   OTMP_13_0_port <= '0';
   SHIFT_n_13_0_port <= '0';
   SHIFT_n_13_1_port <= '0';
   SHIFT_13_0_port <= '0';
   SHIFT_13_1_port <= '0';
   OTMP_12_0_port <= '0';
   SHIFT_n_12_0_port <= '0';
   SHIFT_n_12_1_port <= '0';
   SHIFT_12_0_port <= '0';
   SHIFT_12_1_port <= '0';
   OTMP_11_0_port <= '0';
   SHIFT_n_11_0_port <= '0';
   SHIFT_n_11_1_port <= '0';
   SHIFT_11_0_port <= '0';
   SHIFT_11_1_port <= '0';
   OTMP_10_0_port <= '0';
   SHIFT_n_10_0_port <= '0';
   SHIFT_n_10_1_port <= '0';
   SHIFT_10_0_port <= '0';
   SHIFT_10_1_port <= '0';
   OTMP_9_0_port <= '0';
   SHIFT_n_9_0_port <= '0';
   SHIFT_n_9_1_port <= '0';
   SHIFT_9_0_port <= '0';
   SHIFT_9_1_port <= '0';
   OTMP_8_0_port <= '0';
   SHIFT_n_8_0_port <= '0';
   SHIFT_n_8_1_port <= '0';
   SHIFT_8_0_port <= '0';
   SHIFT_8_1_port <= '0';
   OTMP_7_0_port <= '0';
   SHIFT_n_7_0_port <= '0';
   SHIFT_n_7_1_port <= '0';
   SHIFT_7_0_port <= '0';
   SHIFT_7_1_port <= '0';
   OTMP_6_0_port <= '0';
   SHIFT_n_6_0_port <= '0';
   SHIFT_n_6_1_port <= '0';
   SHIFT_6_0_port <= '0';
   SHIFT_6_1_port <= '0';
   OTMP_5_0_port <= '0';
   SHIFT_n_5_0_port <= '0';
   SHIFT_n_5_1_port <= '0';
   SHIFT_5_0_port <= '0';
   SHIFT_5_1_port <= '0';
   OTMP_4_0_port <= '0';
   SHIFT_n_4_0_port <= '0';
   SHIFT_n_4_1_port <= '0';
   SHIFT_4_0_port <= '0';
   SHIFT_4_1_port <= '0';
   OTMP_3_0_port <= '0';
   SHIFT_n_3_0_port <= '0';
   SHIFT_n_3_1_port <= '0';
   SHIFT_3_0_port <= '0';
   SHIFT_3_1_port <= '0';
   OTMP_2_0_port <= '0';
   SHIFT_n_2_0_port <= '0';
   SHIFT_n_2_1_port <= '0';
   SHIFT_2_0_port <= '0';
   SHIFT_2_1_port <= '0';
   OTMP_1_0_port <= '0';
   SHIFT_n_1_0_port <= '0';
   SHIFT_1_0_port <= '0';
   n4 <= '0';
   n5 <= '0';
   ENC1 : BOOTHENC_NBIT34_i0 port map( A_s(33) => A(31), A_s(32) => A(31), 
                           A_s(31) => A(31), A_s(30) => A(30), A_s(29) => A(29)
                           , A_s(28) => A(28), A_s(27) => A(27), A_s(26) => 
                           A(26), A_s(25) => A(25), A_s(24) => A(24), A_s(23) 
                           => A(23), A_s(22) => A(22), A_s(21) => A(21), 
                           A_s(20) => A(20), A_s(19) => A(19), A_s(18) => A(18)
                           , A_s(17) => A(17), A_s(16) => A(16), A_s(15) => 
                           A(15), A_s(14) => A(14), A_s(13) => A(13), A_s(12) 
                           => A(12), A_s(11) => A(11), A_s(10) => A(10), A_s(9)
                           => A(9), A_s(8) => A(8), A_s(7) => A(7), A_s(6) => 
                           A(6), A_s(5) => A(5), A_s(4) => A(4), A_s(3) => A(3)
                           , A_s(2) => A(2), A_s(1) => n8, A_s(0) => A(0), 
                           A_ns(33) => A_n_65, A_ns(32) => A_n_65, A_ns(31) => 
                           A_n_65, A_ns(30) => A_n_30_port, A_ns(29) => 
                           A_n_29_port, A_ns(28) => A_n_28_port, A_ns(27) => 
                           A_n_27_port, A_ns(26) => A_n_26_port, A_ns(25) => 
                           A_n_25_port, A_ns(24) => A_n_24_port, A_ns(23) => 
                           A_n_23_port, A_ns(22) => A_n_22_port, A_ns(21) => 
                           A_n_21_port, A_ns(20) => A_n_20_port, A_ns(19) => 
                           A_n_19_port, A_ns(18) => A_n_18_port, A_ns(17) => 
                           A_n_17_port, A_ns(16) => A_n_16_port, A_ns(15) => 
                           A_n_15_port, A_ns(14) => A_n_14_port, A_ns(13) => 
                           A_n_13_port, A_ns(12) => A_n_12_port, A_ns(11) => 
                           A_n_11_port, A_ns(10) => A_n_10_port, A_ns(9) => 
                           A_n_9_port, A_ns(8) => A_n_8_port, A_ns(7) => 
                           A_n_7_port, A_ns(6) => A_n_6_port, A_ns(5) => 
                           A_n_5_port, A_ns(4) => A_n_4_port, A_ns(3) => 
                           A_n_3_port, A_ns(2) => A_n_2_port, A_ns(1) => 
                           A_n_1_port, A_ns(0) => A_n_0_port, B(33) => B(31), 
                           B(32) => B(31), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), O(33) => OTMP_0_34_port, O(32) 
                           => OTMP_0_32_port, O(31) => OTMP_0_31_port, O(30) =>
                           OTMP_0_30_port, O(29) => OTMP_0_29_port, O(28) => 
                           OTMP_0_28_port, O(27) => OTMP_0_27_port, O(26) => 
                           OTMP_0_26_port, O(25) => OTMP_0_25_port, O(24) => 
                           OTMP_0_24_port, O(23) => OTMP_0_23_port, O(22) => 
                           OTMP_0_22_port, O(21) => OTMP_0_21_port, O(20) => 
                           OTMP_0_20_port, O(19) => OTMP_0_19_port, O(18) => 
                           OTMP_0_18_port, O(17) => OTMP_0_17_port, O(16) => 
                           OTMP_0_16_port, O(15) => OTMP_0_15_port, O(14) => 
                           OTMP_0_14_port, O(13) => OTMP_0_13_port, O(12) => 
                           OTMP_0_12_port, O(11) => OTMP_0_11_port, O(10) => 
                           OTMP_0_10_port, O(9) => OTMP_0_9_port, O(8) => 
                           OTMP_0_8_port, O(7) => OTMP_0_7_port, O(6) => 
                           OTMP_0_6_port, O(5) => OTMP_0_5_port, O(4) => 
                           OTMP_0_4_port, O(3) => OTMP_0_3_port, O(2) => 
                           OTMP_0_2_port, O(1) => OTMP_0_1_port, O(0) => 
                           OTMP_0_0_port, A_so(33) => SHIFT_1_33_port, A_so(32)
                           => SHIFT_1_32_port, A_so(31) => SHIFT_1_31_port, 
                           A_so(30) => SHIFT_1_30_port, A_so(29) => 
                           SHIFT_1_29_port, A_so(28) => SHIFT_1_28_port, 
                           A_so(27) => SHIFT_1_27_port, A_so(26) => 
                           SHIFT_1_26_port, A_so(25) => SHIFT_1_25_port, 
                           A_so(24) => SHIFT_1_24_port, A_so(23) => 
                           SHIFT_1_23_port, A_so(22) => SHIFT_1_22_port, 
                           A_so(21) => SHIFT_1_21_port, A_so(20) => 
                           SHIFT_1_20_port, A_so(19) => SHIFT_1_19_port, 
                           A_so(18) => SHIFT_1_18_port, A_so(17) => 
                           SHIFT_1_17_port, A_so(16) => SHIFT_1_16_port, 
                           A_so(15) => SHIFT_1_15_port, A_so(14) => 
                           SHIFT_1_14_port, A_so(13) => SHIFT_1_13_port, 
                           A_so(12) => SHIFT_1_12_port, A_so(11) => 
                           SHIFT_1_11_port, A_so(10) => SHIFT_1_10_port, 
                           A_so(9) => SHIFT_1_9_port, A_so(8) => SHIFT_1_8_port
                           , A_so(7) => SHIFT_1_7_port, A_so(6) => 
                           SHIFT_1_6_port, A_so(5) => SHIFT_1_5_port, A_so(4) 
                           => SHIFT_1_4_port, A_so(3) => SHIFT_1_3_port, 
                           A_so(2) => SHIFT_1_2_port, A_so(1) => SHIFT_1_1_port
                           , A_so(0) => n_1080, A_nso(33) => SHIFT_n_1_33_port,
                           A_nso(32) => SHIFT_n_1_32_port, A_nso(31) => 
                           SHIFT_n_1_31_port, A_nso(30) => SHIFT_n_1_30_port, 
                           A_nso(29) => SHIFT_n_1_29_port, A_nso(28) => 
                           SHIFT_n_1_28_port, A_nso(27) => SHIFT_n_1_27_port, 
                           A_nso(26) => SHIFT_n_1_26_port, A_nso(25) => 
                           SHIFT_n_1_25_port, A_nso(24) => SHIFT_n_1_24_port, 
                           A_nso(23) => SHIFT_n_1_23_port, A_nso(22) => 
                           SHIFT_n_1_22_port, A_nso(21) => SHIFT_n_1_21_port, 
                           A_nso(20) => SHIFT_n_1_20_port, A_nso(19) => 
                           SHIFT_n_1_19_port, A_nso(18) => SHIFT_n_1_18_port, 
                           A_nso(17) => SHIFT_n_1_17_port, A_nso(16) => 
                           SHIFT_n_1_16_port, A_nso(15) => SHIFT_n_1_15_port, 
                           A_nso(14) => SHIFT_n_1_14_port, A_nso(13) => 
                           SHIFT_n_1_13_port, A_nso(12) => SHIFT_n_1_12_port, 
                           A_nso(11) => SHIFT_n_1_11_port, A_nso(10) => 
                           SHIFT_n_1_10_port, A_nso(9) => SHIFT_n_1_9_port, 
                           A_nso(8) => SHIFT_n_1_8_port, A_nso(7) => 
                           SHIFT_n_1_7_port, A_nso(6) => SHIFT_n_1_6_port, 
                           A_nso(5) => SHIFT_n_1_5_port, A_nso(4) => 
                           SHIFT_n_1_4_port, A_nso(3) => SHIFT_n_1_3_port, 
                           A_nso(2) => SHIFT_n_1_2_port, A_nso(1) => 
                           SHIFT_n_1_1_port, A_nso(0) => n_1081);
   ENC_1 : BOOTHENC_NBIT36_i2 port map( A_s(35) => SHIFT_1_33_port, A_s(34) => 
                           SHIFT_1_33_port, A_s(33) => SHIFT_1_33_port, A_s(32)
                           => SHIFT_1_32_port, A_s(31) => SHIFT_1_31_port, 
                           A_s(30) => SHIFT_1_30_port, A_s(29) => 
                           SHIFT_1_29_port, A_s(28) => SHIFT_1_28_port, A_s(27)
                           => SHIFT_1_27_port, A_s(26) => SHIFT_1_26_port, 
                           A_s(25) => SHIFT_1_25_port, A_s(24) => 
                           SHIFT_1_24_port, A_s(23) => SHIFT_1_23_port, A_s(22)
                           => SHIFT_1_22_port, A_s(21) => SHIFT_1_21_port, 
                           A_s(20) => SHIFT_1_20_port, A_s(19) => 
                           SHIFT_1_19_port, A_s(18) => SHIFT_1_18_port, A_s(17)
                           => SHIFT_1_17_port, A_s(16) => SHIFT_1_16_port, 
                           A_s(15) => SHIFT_1_15_port, A_s(14) => 
                           SHIFT_1_14_port, A_s(13) => SHIFT_1_13_port, A_s(12)
                           => SHIFT_1_12_port, A_s(11) => SHIFT_1_11_port, 
                           A_s(10) => SHIFT_1_10_port, A_s(9) => SHIFT_1_9_port
                           , A_s(8) => SHIFT_1_8_port, A_s(7) => SHIFT_1_7_port
                           , A_s(6) => SHIFT_1_6_port, A_s(5) => SHIFT_1_5_port
                           , A_s(4) => SHIFT_1_4_port, A_s(3) => SHIFT_1_3_port
                           , A_s(2) => SHIFT_1_2_port, A_s(1) => SHIFT_1_1_port
                           , A_s(0) => SHIFT_1_0_port, A_ns(35) => 
                           SHIFT_n_1_33_port, A_ns(34) => SHIFT_n_1_33_port, 
                           A_ns(33) => SHIFT_n_1_33_port, A_ns(32) => 
                           SHIFT_n_1_32_port, A_ns(31) => SHIFT_n_1_31_port, 
                           A_ns(30) => SHIFT_n_1_30_port, A_ns(29) => 
                           SHIFT_n_1_29_port, A_ns(28) => SHIFT_n_1_28_port, 
                           A_ns(27) => SHIFT_n_1_27_port, A_ns(26) => 
                           SHIFT_n_1_26_port, A_ns(25) => SHIFT_n_1_25_port, 
                           A_ns(24) => SHIFT_n_1_24_port, A_ns(23) => 
                           SHIFT_n_1_23_port, A_ns(22) => SHIFT_n_1_22_port, 
                           A_ns(21) => SHIFT_n_1_21_port, A_ns(20) => 
                           SHIFT_n_1_20_port, A_ns(19) => SHIFT_n_1_19_port, 
                           A_ns(18) => SHIFT_n_1_18_port, A_ns(17) => 
                           SHIFT_n_1_17_port, A_ns(16) => SHIFT_n_1_16_port, 
                           A_ns(15) => SHIFT_n_1_15_port, A_ns(14) => 
                           SHIFT_n_1_14_port, A_ns(13) => SHIFT_n_1_13_port, 
                           A_ns(12) => SHIFT_n_1_12_port, A_ns(11) => 
                           SHIFT_n_1_11_port, A_ns(10) => SHIFT_n_1_10_port, 
                           A_ns(9) => SHIFT_n_1_9_port, A_ns(8) => 
                           SHIFT_n_1_8_port, A_ns(7) => SHIFT_n_1_7_port, 
                           A_ns(6) => SHIFT_n_1_6_port, A_ns(5) => 
                           SHIFT_n_1_5_port, A_ns(4) => SHIFT_n_1_4_port, 
                           A_ns(3) => SHIFT_n_1_3_port, A_ns(2) => 
                           SHIFT_n_1_2_port, A_ns(1) => SHIFT_n_1_1_port, 
                           A_ns(0) => SHIFT_n_1_0_port, B(35) => B(31), B(34) 
                           => B(31), B(33) => B(31), B(32) => B(31), B(31) => 
                           B(31), B(30) => B(30), B(29) => B(29), B(28) => 
                           B(28), B(27) => B(27), B(26) => B(26), B(25) => 
                           B(25), B(24) => B(24), B(23) => B(23), B(22) => 
                           B(22), B(21) => B(21), B(20) => B(20), B(19) => 
                           B(19), B(18) => B(18), B(17) => B(17), B(16) => 
                           B(16), B(15) => B(15), B(14) => B(14), B(13) => 
                           B(13), B(12) => B(12), B(11) => B(11), B(10) => 
                           B(10), B(9) => B(9), B(8) => B(8), B(7) => B(7), 
                           B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3) => 
                           B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), 
                           O(35) => OTMP_1_35_port, O(34) => OTMP_1_34_port, 
                           O(33) => OTMP_1_33_port, O(32) => OTMP_1_32_port, 
                           O(31) => OTMP_1_31_port, O(30) => OTMP_1_30_port, 
                           O(29) => OTMP_1_29_port, O(28) => OTMP_1_28_port, 
                           O(27) => OTMP_1_27_port, O(26) => OTMP_1_26_port, 
                           O(25) => OTMP_1_25_port, O(24) => OTMP_1_24_port, 
                           O(23) => OTMP_1_23_port, O(22) => OTMP_1_22_port, 
                           O(21) => OTMP_1_21_port, O(20) => OTMP_1_20_port, 
                           O(19) => OTMP_1_19_port, O(18) => OTMP_1_18_port, 
                           O(17) => OTMP_1_17_port, O(16) => OTMP_1_16_port, 
                           O(15) => OTMP_1_15_port, O(14) => OTMP_1_14_port, 
                           O(13) => OTMP_1_13_port, O(12) => OTMP_1_12_port, 
                           O(11) => OTMP_1_11_port, O(10) => OTMP_1_10_port, 
                           O(9) => OTMP_1_9_port, O(8) => OTMP_1_8_port, O(7) 
                           => OTMP_1_7_port, O(6) => OTMP_1_6_port, O(5) => 
                           OTMP_1_5_port, O(4) => OTMP_1_4_port, O(3) => 
                           OTMP_1_3_port, O(2) => OTMP_1_2_port, O(1) => 
                           OTMP_1_1_port, O(0) => n_1082, A_so(35) => 
                           SHIFT_2_35_port, A_so(34) => SHIFT_2_34_port, 
                           A_so(33) => SHIFT_2_33_port, A_so(32) => 
                           SHIFT_2_32_port, A_so(31) => SHIFT_2_31_port, 
                           A_so(30) => SHIFT_2_30_port, A_so(29) => 
                           SHIFT_2_29_port, A_so(28) => SHIFT_2_28_port, 
                           A_so(27) => SHIFT_2_27_port, A_so(26) => 
                           SHIFT_2_26_port, A_so(25) => SHIFT_2_25_port, 
                           A_so(24) => SHIFT_2_24_port, A_so(23) => 
                           SHIFT_2_23_port, A_so(22) => SHIFT_2_22_port, 
                           A_so(21) => SHIFT_2_21_port, A_so(20) => 
                           SHIFT_2_20_port, A_so(19) => SHIFT_2_19_port, 
                           A_so(18) => SHIFT_2_18_port, A_so(17) => 
                           SHIFT_2_17_port, A_so(16) => SHIFT_2_16_port, 
                           A_so(15) => SHIFT_2_15_port, A_so(14) => 
                           SHIFT_2_14_port, A_so(13) => SHIFT_2_13_port, 
                           A_so(12) => SHIFT_2_12_port, A_so(11) => 
                           SHIFT_2_11_port, A_so(10) => SHIFT_2_10_port, 
                           A_so(9) => SHIFT_2_9_port, A_so(8) => SHIFT_2_8_port
                           , A_so(7) => SHIFT_2_7_port, A_so(6) => 
                           SHIFT_2_6_port, A_so(5) => SHIFT_2_5_port, A_so(4) 
                           => SHIFT_2_4_port, A_so(3) => SHIFT_2_3_port, 
                           A_so(2) => SHIFT_2_2_port, A_so(1) => n_1083, 
                           A_so(0) => n_1084, A_nso(35) => SHIFT_n_2_35_port, 
                           A_nso(34) => SHIFT_n_2_34_port, A_nso(33) => 
                           SHIFT_n_2_33_port, A_nso(32) => SHIFT_n_2_32_port, 
                           A_nso(31) => SHIFT_n_2_31_port, A_nso(30) => 
                           SHIFT_n_2_30_port, A_nso(29) => SHIFT_n_2_29_port, 
                           A_nso(28) => SHIFT_n_2_28_port, A_nso(27) => 
                           SHIFT_n_2_27_port, A_nso(26) => SHIFT_n_2_26_port, 
                           A_nso(25) => SHIFT_n_2_25_port, A_nso(24) => 
                           SHIFT_n_2_24_port, A_nso(23) => SHIFT_n_2_23_port, 
                           A_nso(22) => SHIFT_n_2_22_port, A_nso(21) => 
                           SHIFT_n_2_21_port, A_nso(20) => SHIFT_n_2_20_port, 
                           A_nso(19) => SHIFT_n_2_19_port, A_nso(18) => 
                           SHIFT_n_2_18_port, A_nso(17) => SHIFT_n_2_17_port, 
                           A_nso(16) => SHIFT_n_2_16_port, A_nso(15) => 
                           SHIFT_n_2_15_port, A_nso(14) => SHIFT_n_2_14_port, 
                           A_nso(13) => SHIFT_n_2_13_port, A_nso(12) => 
                           SHIFT_n_2_12_port, A_nso(11) => SHIFT_n_2_11_port, 
                           A_nso(10) => SHIFT_n_2_10_port, A_nso(9) => 
                           SHIFT_n_2_9_port, A_nso(8) => SHIFT_n_2_8_port, 
                           A_nso(7) => SHIFT_n_2_7_port, A_nso(6) => 
                           SHIFT_n_2_6_port, A_nso(5) => SHIFT_n_2_5_port, 
                           A_nso(4) => SHIFT_n_2_4_port, A_nso(3) => 
                           SHIFT_n_2_3_port, A_nso(2) => SHIFT_n_2_2_port, 
                           A_nso(1) => n_1085, A_nso(0) => n_1086);
   ENC_2 : BOOTHENC_NBIT38_i4 port map( A_s(37) => SHIFT_2_35_port, A_s(36) => 
                           SHIFT_2_35_port, A_s(35) => SHIFT_2_35_port, A_s(34)
                           => SHIFT_2_34_port, A_s(33) => SHIFT_2_33_port, 
                           A_s(32) => SHIFT_2_32_port, A_s(31) => 
                           SHIFT_2_31_port, A_s(30) => SHIFT_2_30_port, A_s(29)
                           => SHIFT_2_29_port, A_s(28) => SHIFT_2_28_port, 
                           A_s(27) => SHIFT_2_27_port, A_s(26) => 
                           SHIFT_2_26_port, A_s(25) => SHIFT_2_25_port, A_s(24)
                           => SHIFT_2_24_port, A_s(23) => SHIFT_2_23_port, 
                           A_s(22) => SHIFT_2_22_port, A_s(21) => 
                           SHIFT_2_21_port, A_s(20) => SHIFT_2_20_port, A_s(19)
                           => SHIFT_2_19_port, A_s(18) => SHIFT_2_18_port, 
                           A_s(17) => SHIFT_2_17_port, A_s(16) => 
                           SHIFT_2_16_port, A_s(15) => SHIFT_2_15_port, A_s(14)
                           => SHIFT_2_14_port, A_s(13) => SHIFT_2_13_port, 
                           A_s(12) => SHIFT_2_12_port, A_s(11) => 
                           SHIFT_2_11_port, A_s(10) => SHIFT_2_10_port, A_s(9) 
                           => SHIFT_2_9_port, A_s(8) => SHIFT_2_8_port, A_s(7) 
                           => SHIFT_2_7_port, A_s(6) => SHIFT_2_6_port, A_s(5) 
                           => SHIFT_2_5_port, A_s(4) => SHIFT_2_4_port, A_s(3) 
                           => SHIFT_2_3_port, A_s(2) => SHIFT_2_2_port, A_s(1) 
                           => SHIFT_2_1_port, A_s(0) => SHIFT_2_0_port, 
                           A_ns(37) => SHIFT_n_2_35_port, A_ns(36) => 
                           SHIFT_n_2_35_port, A_ns(35) => SHIFT_n_2_35_port, 
                           A_ns(34) => SHIFT_n_2_34_port, A_ns(33) => 
                           SHIFT_n_2_33_port, A_ns(32) => SHIFT_n_2_32_port, 
                           A_ns(31) => SHIFT_n_2_31_port, A_ns(30) => 
                           SHIFT_n_2_30_port, A_ns(29) => SHIFT_n_2_29_port, 
                           A_ns(28) => SHIFT_n_2_28_port, A_ns(27) => 
                           SHIFT_n_2_27_port, A_ns(26) => SHIFT_n_2_26_port, 
                           A_ns(25) => SHIFT_n_2_25_port, A_ns(24) => 
                           SHIFT_n_2_24_port, A_ns(23) => SHIFT_n_2_23_port, 
                           A_ns(22) => SHIFT_n_2_22_port, A_ns(21) => 
                           SHIFT_n_2_21_port, A_ns(20) => SHIFT_n_2_20_port, 
                           A_ns(19) => SHIFT_n_2_19_port, A_ns(18) => 
                           SHIFT_n_2_18_port, A_ns(17) => SHIFT_n_2_17_port, 
                           A_ns(16) => SHIFT_n_2_16_port, A_ns(15) => 
                           SHIFT_n_2_15_port, A_ns(14) => SHIFT_n_2_14_port, 
                           A_ns(13) => SHIFT_n_2_13_port, A_ns(12) => 
                           SHIFT_n_2_12_port, A_ns(11) => SHIFT_n_2_11_port, 
                           A_ns(10) => SHIFT_n_2_10_port, A_ns(9) => 
                           SHIFT_n_2_9_port, A_ns(8) => SHIFT_n_2_8_port, 
                           A_ns(7) => SHIFT_n_2_7_port, A_ns(6) => 
                           SHIFT_n_2_6_port, A_ns(5) => SHIFT_n_2_5_port, 
                           A_ns(4) => SHIFT_n_2_4_port, A_ns(3) => 
                           SHIFT_n_2_3_port, A_ns(2) => SHIFT_n_2_2_port, 
                           A_ns(1) => SHIFT_n_2_1_port, A_ns(0) => 
                           SHIFT_n_2_0_port, B(37) => B(31), B(36) => B(31), 
                           B(35) => B(31), B(34) => B(31), B(33) => B(31), 
                           B(32) => B(31), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), O(37) => OTMP_2_37_port, O(36) 
                           => OTMP_2_36_port, O(35) => OTMP_2_35_port, O(34) =>
                           OTMP_2_34_port, O(33) => OTMP_2_33_port, O(32) => 
                           OTMP_2_32_port, O(31) => OTMP_2_31_port, O(30) => 
                           OTMP_2_30_port, O(29) => OTMP_2_29_port, O(28) => 
                           OTMP_2_28_port, O(27) => OTMP_2_27_port, O(26) => 
                           OTMP_2_26_port, O(25) => OTMP_2_25_port, O(24) => 
                           OTMP_2_24_port, O(23) => OTMP_2_23_port, O(22) => 
                           OTMP_2_22_port, O(21) => OTMP_2_21_port, O(20) => 
                           OTMP_2_20_port, O(19) => OTMP_2_19_port, O(18) => 
                           OTMP_2_18_port, O(17) => OTMP_2_17_port, O(16) => 
                           OTMP_2_16_port, O(15) => OTMP_2_15_port, O(14) => 
                           OTMP_2_14_port, O(13) => OTMP_2_13_port, O(12) => 
                           OTMP_2_12_port, O(11) => OTMP_2_11_port, O(10) => 
                           OTMP_2_10_port, O(9) => OTMP_2_9_port, O(8) => 
                           OTMP_2_8_port, O(7) => OTMP_2_7_port, O(6) => 
                           OTMP_2_6_port, O(5) => OTMP_2_5_port, O(4) => 
                           OTMP_2_4_port, O(3) => OTMP_2_3_port, O(2) => 
                           OTMP_2_2_port, O(1) => OTMP_2_1_port, O(0) => n_1087
                           , A_so(37) => SHIFT_3_37_port, A_so(36) => 
                           SHIFT_3_36_port, A_so(35) => SHIFT_3_35_port, 
                           A_so(34) => SHIFT_3_34_port, A_so(33) => 
                           SHIFT_3_33_port, A_so(32) => SHIFT_3_32_port, 
                           A_so(31) => SHIFT_3_31_port, A_so(30) => 
                           SHIFT_3_30_port, A_so(29) => SHIFT_3_29_port, 
                           A_so(28) => SHIFT_3_28_port, A_so(27) => 
                           SHIFT_3_27_port, A_so(26) => SHIFT_3_26_port, 
                           A_so(25) => SHIFT_3_25_port, A_so(24) => 
                           SHIFT_3_24_port, A_so(23) => SHIFT_3_23_port, 
                           A_so(22) => SHIFT_3_22_port, A_so(21) => 
                           SHIFT_3_21_port, A_so(20) => SHIFT_3_20_port, 
                           A_so(19) => SHIFT_3_19_port, A_so(18) => 
                           SHIFT_3_18_port, A_so(17) => SHIFT_3_17_port, 
                           A_so(16) => SHIFT_3_16_port, A_so(15) => 
                           SHIFT_3_15_port, A_so(14) => SHIFT_3_14_port, 
                           A_so(13) => SHIFT_3_13_port, A_so(12) => 
                           SHIFT_3_12_port, A_so(11) => SHIFT_3_11_port, 
                           A_so(10) => SHIFT_3_10_port, A_so(9) => 
                           SHIFT_3_9_port, A_so(8) => SHIFT_3_8_port, A_so(7) 
                           => SHIFT_3_7_port, A_so(6) => SHIFT_3_6_port, 
                           A_so(5) => SHIFT_3_5_port, A_so(4) => SHIFT_3_4_port
                           , A_so(3) => SHIFT_3_3_port, A_so(2) => 
                           SHIFT_3_2_port, A_so(1) => n_1088, A_so(0) => n_1089
                           , A_nso(37) => SHIFT_n_3_37_port, A_nso(36) => 
                           SHIFT_n_3_36_port, A_nso(35) => SHIFT_n_3_35_port, 
                           A_nso(34) => SHIFT_n_3_34_port, A_nso(33) => 
                           SHIFT_n_3_33_port, A_nso(32) => SHIFT_n_3_32_port, 
                           A_nso(31) => SHIFT_n_3_31_port, A_nso(30) => 
                           SHIFT_n_3_30_port, A_nso(29) => SHIFT_n_3_29_port, 
                           A_nso(28) => SHIFT_n_3_28_port, A_nso(27) => 
                           SHIFT_n_3_27_port, A_nso(26) => SHIFT_n_3_26_port, 
                           A_nso(25) => SHIFT_n_3_25_port, A_nso(24) => 
                           SHIFT_n_3_24_port, A_nso(23) => SHIFT_n_3_23_port, 
                           A_nso(22) => SHIFT_n_3_22_port, A_nso(21) => 
                           SHIFT_n_3_21_port, A_nso(20) => SHIFT_n_3_20_port, 
                           A_nso(19) => SHIFT_n_3_19_port, A_nso(18) => 
                           SHIFT_n_3_18_port, A_nso(17) => SHIFT_n_3_17_port, 
                           A_nso(16) => SHIFT_n_3_16_port, A_nso(15) => 
                           SHIFT_n_3_15_port, A_nso(14) => SHIFT_n_3_14_port, 
                           A_nso(13) => SHIFT_n_3_13_port, A_nso(12) => 
                           SHIFT_n_3_12_port, A_nso(11) => SHIFT_n_3_11_port, 
                           A_nso(10) => SHIFT_n_3_10_port, A_nso(9) => 
                           SHIFT_n_3_9_port, A_nso(8) => SHIFT_n_3_8_port, 
                           A_nso(7) => SHIFT_n_3_7_port, A_nso(6) => 
                           SHIFT_n_3_6_port, A_nso(5) => SHIFT_n_3_5_port, 
                           A_nso(4) => SHIFT_n_3_4_port, A_nso(3) => 
                           SHIFT_n_3_3_port, A_nso(2) => SHIFT_n_3_2_port, 
                           A_nso(1) => n_1090, A_nso(0) => n_1091);
   ENC_3 : BOOTHENC_NBIT40_i6 port map( A_s(39) => n19, A_s(38) => n19, A_s(37)
                           => n19, A_s(36) => SHIFT_3_36_port, A_s(35) => 
                           SHIFT_3_35_port, A_s(34) => SHIFT_3_34_port, A_s(33)
                           => SHIFT_3_33_port, A_s(32) => SHIFT_3_32_port, 
                           A_s(31) => SHIFT_3_31_port, A_s(30) => 
                           SHIFT_3_30_port, A_s(29) => SHIFT_3_29_port, A_s(28)
                           => SHIFT_3_28_port, A_s(27) => SHIFT_3_27_port, 
                           A_s(26) => SHIFT_3_26_port, A_s(25) => 
                           SHIFT_3_25_port, A_s(24) => SHIFT_3_24_port, A_s(23)
                           => SHIFT_3_23_port, A_s(22) => SHIFT_3_22_port, 
                           A_s(21) => SHIFT_3_21_port, A_s(20) => 
                           SHIFT_3_20_port, A_s(19) => SHIFT_3_19_port, A_s(18)
                           => SHIFT_3_18_port, A_s(17) => SHIFT_3_17_port, 
                           A_s(16) => SHIFT_3_16_port, A_s(15) => 
                           SHIFT_3_15_port, A_s(14) => SHIFT_3_14_port, A_s(13)
                           => SHIFT_3_13_port, A_s(12) => SHIFT_3_12_port, 
                           A_s(11) => SHIFT_3_11_port, A_s(10) => 
                           SHIFT_3_10_port, A_s(9) => SHIFT_3_9_port, A_s(8) =>
                           SHIFT_3_8_port, A_s(7) => SHIFT_3_7_port, A_s(6) => 
                           SHIFT_3_6_port, A_s(5) => SHIFT_3_5_port, A_s(4) => 
                           SHIFT_3_4_port, A_s(3) => SHIFT_3_3_port, A_s(2) => 
                           SHIFT_3_2_port, A_s(1) => SHIFT_3_1_port, A_s(0) => 
                           SHIFT_3_0_port, A_ns(39) => SHIFT_n_3_37_port, 
                           A_ns(38) => SHIFT_n_3_37_port, A_ns(37) => 
                           SHIFT_n_3_37_port, A_ns(36) => SHIFT_n_3_36_port, 
                           A_ns(35) => SHIFT_n_3_35_port, A_ns(34) => 
                           SHIFT_n_3_34_port, A_ns(33) => SHIFT_n_3_33_port, 
                           A_ns(32) => SHIFT_n_3_32_port, A_ns(31) => 
                           SHIFT_n_3_31_port, A_ns(30) => SHIFT_n_3_30_port, 
                           A_ns(29) => SHIFT_n_3_29_port, A_ns(28) => 
                           SHIFT_n_3_28_port, A_ns(27) => SHIFT_n_3_27_port, 
                           A_ns(26) => SHIFT_n_3_26_port, A_ns(25) => 
                           SHIFT_n_3_25_port, A_ns(24) => SHIFT_n_3_24_port, 
                           A_ns(23) => SHIFT_n_3_23_port, A_ns(22) => 
                           SHIFT_n_3_22_port, A_ns(21) => SHIFT_n_3_21_port, 
                           A_ns(20) => SHIFT_n_3_20_port, A_ns(19) => 
                           SHIFT_n_3_19_port, A_ns(18) => SHIFT_n_3_18_port, 
                           A_ns(17) => SHIFT_n_3_17_port, A_ns(16) => 
                           SHIFT_n_3_16_port, A_ns(15) => SHIFT_n_3_15_port, 
                           A_ns(14) => SHIFT_n_3_14_port, A_ns(13) => 
                           SHIFT_n_3_13_port, A_ns(12) => SHIFT_n_3_12_port, 
                           A_ns(11) => SHIFT_n_3_11_port, A_ns(10) => 
                           SHIFT_n_3_10_port, A_ns(9) => SHIFT_n_3_9_port, 
                           A_ns(8) => SHIFT_n_3_8_port, A_ns(7) => 
                           SHIFT_n_3_7_port, A_ns(6) => SHIFT_n_3_6_port, 
                           A_ns(5) => SHIFT_n_3_5_port, A_ns(4) => 
                           SHIFT_n_3_4_port, A_ns(3) => SHIFT_n_3_3_port, 
                           A_ns(2) => SHIFT_n_3_2_port, A_ns(1) => 
                           SHIFT_n_3_1_port, A_ns(0) => SHIFT_n_3_0_port, B(39)
                           => B(31), B(38) => B(31), B(37) => B(31), B(36) => 
                           B(31), B(35) => B(31), B(34) => B(31), B(33) => 
                           B(31), B(32) => B(31), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), O(39) => OTMP_3_39_port, 
                           O(38) => OTMP_3_38_port, O(37) => OTMP_3_37_port, 
                           O(36) => OTMP_3_36_port, O(35) => OTMP_3_35_port, 
                           O(34) => OTMP_3_34_port, O(33) => OTMP_3_33_port, 
                           O(32) => OTMP_3_32_port, O(31) => OTMP_3_31_port, 
                           O(30) => OTMP_3_30_port, O(29) => OTMP_3_29_port, 
                           O(28) => OTMP_3_28_port, O(27) => OTMP_3_27_port, 
                           O(26) => OTMP_3_26_port, O(25) => OTMP_3_25_port, 
                           O(24) => OTMP_3_24_port, O(23) => OTMP_3_23_port, 
                           O(22) => OTMP_3_22_port, O(21) => OTMP_3_21_port, 
                           O(20) => OTMP_3_20_port, O(19) => OTMP_3_19_port, 
                           O(18) => OTMP_3_18_port, O(17) => OTMP_3_17_port, 
                           O(16) => OTMP_3_16_port, O(15) => OTMP_3_15_port, 
                           O(14) => OTMP_3_14_port, O(13) => OTMP_3_13_port, 
                           O(12) => OTMP_3_12_port, O(11) => OTMP_3_11_port, 
                           O(10) => OTMP_3_10_port, O(9) => OTMP_3_9_port, O(8)
                           => OTMP_3_8_port, O(7) => OTMP_3_7_port, O(6) => 
                           OTMP_3_6_port, O(5) => OTMP_3_5_port, O(4) => 
                           OTMP_3_4_port, O(3) => OTMP_3_3_port, O(2) => 
                           OTMP_3_2_port, O(1) => OTMP_3_1_port, O(0) => n_1092
                           , A_so(39) => SHIFT_4_39_port, A_so(38) => 
                           SHIFT_4_38_port, A_so(37) => SHIFT_4_37_port, 
                           A_so(36) => SHIFT_4_36_port, A_so(35) => 
                           SHIFT_4_35_port, A_so(34) => SHIFT_4_34_port, 
                           A_so(33) => SHIFT_4_33_port, A_so(32) => 
                           SHIFT_4_32_port, A_so(31) => SHIFT_4_31_port, 
                           A_so(30) => SHIFT_4_30_port, A_so(29) => 
                           SHIFT_4_29_port, A_so(28) => SHIFT_4_28_port, 
                           A_so(27) => SHIFT_4_27_port, A_so(26) => 
                           SHIFT_4_26_port, A_so(25) => SHIFT_4_25_port, 
                           A_so(24) => SHIFT_4_24_port, A_so(23) => 
                           SHIFT_4_23_port, A_so(22) => SHIFT_4_22_port, 
                           A_so(21) => SHIFT_4_21_port, A_so(20) => 
                           SHIFT_4_20_port, A_so(19) => SHIFT_4_19_port, 
                           A_so(18) => SHIFT_4_18_port, A_so(17) => 
                           SHIFT_4_17_port, A_so(16) => SHIFT_4_16_port, 
                           A_so(15) => SHIFT_4_15_port, A_so(14) => 
                           SHIFT_4_14_port, A_so(13) => SHIFT_4_13_port, 
                           A_so(12) => SHIFT_4_12_port, A_so(11) => 
                           SHIFT_4_11_port, A_so(10) => SHIFT_4_10_port, 
                           A_so(9) => SHIFT_4_9_port, A_so(8) => SHIFT_4_8_port
                           , A_so(7) => SHIFT_4_7_port, A_so(6) => 
                           SHIFT_4_6_port, A_so(5) => SHIFT_4_5_port, A_so(4) 
                           => SHIFT_4_4_port, A_so(3) => SHIFT_4_3_port, 
                           A_so(2) => SHIFT_4_2_port, A_so(1) => n_1093, 
                           A_so(0) => n_1094, A_nso(39) => SHIFT_n_4_39_port, 
                           A_nso(38) => SHIFT_n_4_38_port, A_nso(37) => 
                           SHIFT_n_4_37_port, A_nso(36) => SHIFT_n_4_36_port, 
                           A_nso(35) => SHIFT_n_4_35_port, A_nso(34) => 
                           SHIFT_n_4_34_port, A_nso(33) => SHIFT_n_4_33_port, 
                           A_nso(32) => SHIFT_n_4_32_port, A_nso(31) => 
                           SHIFT_n_4_31_port, A_nso(30) => SHIFT_n_4_30_port, 
                           A_nso(29) => SHIFT_n_4_29_port, A_nso(28) => 
                           SHIFT_n_4_28_port, A_nso(27) => SHIFT_n_4_27_port, 
                           A_nso(26) => SHIFT_n_4_26_port, A_nso(25) => 
                           SHIFT_n_4_25_port, A_nso(24) => SHIFT_n_4_24_port, 
                           A_nso(23) => SHIFT_n_4_23_port, A_nso(22) => 
                           SHIFT_n_4_22_port, A_nso(21) => SHIFT_n_4_21_port, 
                           A_nso(20) => SHIFT_n_4_20_port, A_nso(19) => 
                           SHIFT_n_4_19_port, A_nso(18) => SHIFT_n_4_18_port, 
                           A_nso(17) => SHIFT_n_4_17_port, A_nso(16) => 
                           SHIFT_n_4_16_port, A_nso(15) => SHIFT_n_4_15_port, 
                           A_nso(14) => SHIFT_n_4_14_port, A_nso(13) => 
                           SHIFT_n_4_13_port, A_nso(12) => SHIFT_n_4_12_port, 
                           A_nso(11) => SHIFT_n_4_11_port, A_nso(10) => 
                           SHIFT_n_4_10_port, A_nso(9) => SHIFT_n_4_9_port, 
                           A_nso(8) => SHIFT_n_4_8_port, A_nso(7) => 
                           SHIFT_n_4_7_port, A_nso(6) => SHIFT_n_4_6_port, 
                           A_nso(5) => SHIFT_n_4_5_port, A_nso(4) => 
                           SHIFT_n_4_4_port, A_nso(3) => SHIFT_n_4_3_port, 
                           A_nso(2) => SHIFT_n_4_2_port, A_nso(1) => n_1095, 
                           A_nso(0) => n_1096);
   ENC_4 : BOOTHENC_NBIT42_i8 port map( A_s(41) => SHIFT_4_39_port, A_s(40) => 
                           SHIFT_4_39_port, A_s(39) => SHIFT_4_39_port, A_s(38)
                           => SHIFT_4_38_port, A_s(37) => SHIFT_4_37_port, 
                           A_s(36) => SHIFT_4_36_port, A_s(35) => 
                           SHIFT_4_35_port, A_s(34) => SHIFT_4_34_port, A_s(33)
                           => SHIFT_4_33_port, A_s(32) => SHIFT_4_32_port, 
                           A_s(31) => SHIFT_4_31_port, A_s(30) => 
                           SHIFT_4_30_port, A_s(29) => SHIFT_4_29_port, A_s(28)
                           => SHIFT_4_28_port, A_s(27) => SHIFT_4_27_port, 
                           A_s(26) => SHIFT_4_26_port, A_s(25) => 
                           SHIFT_4_25_port, A_s(24) => SHIFT_4_24_port, A_s(23)
                           => SHIFT_4_23_port, A_s(22) => SHIFT_4_22_port, 
                           A_s(21) => SHIFT_4_21_port, A_s(20) => 
                           SHIFT_4_20_port, A_s(19) => SHIFT_4_19_port, A_s(18)
                           => SHIFT_4_18_port, A_s(17) => SHIFT_4_17_port, 
                           A_s(16) => SHIFT_4_16_port, A_s(15) => 
                           SHIFT_4_15_port, A_s(14) => SHIFT_4_14_port, A_s(13)
                           => SHIFT_4_13_port, A_s(12) => SHIFT_4_12_port, 
                           A_s(11) => SHIFT_4_11_port, A_s(10) => 
                           SHIFT_4_10_port, A_s(9) => SHIFT_4_9_port, A_s(8) =>
                           SHIFT_4_8_port, A_s(7) => SHIFT_4_7_port, A_s(6) => 
                           SHIFT_4_6_port, A_s(5) => SHIFT_4_5_port, A_s(4) => 
                           SHIFT_4_4_port, A_s(3) => SHIFT_4_3_port, A_s(2) => 
                           SHIFT_4_2_port, A_s(1) => SHIFT_4_1_port, A_s(0) => 
                           SHIFT_4_0_port, A_ns(41) => SHIFT_n_4_39_port, 
                           A_ns(40) => SHIFT_n_4_39_port, A_ns(39) => 
                           SHIFT_n_4_39_port, A_ns(38) => SHIFT_n_4_38_port, 
                           A_ns(37) => SHIFT_n_4_37_port, A_ns(36) => 
                           SHIFT_n_4_36_port, A_ns(35) => SHIFT_n_4_35_port, 
                           A_ns(34) => SHIFT_n_4_34_port, A_ns(33) => 
                           SHIFT_n_4_33_port, A_ns(32) => SHIFT_n_4_32_port, 
                           A_ns(31) => SHIFT_n_4_31_port, A_ns(30) => 
                           SHIFT_n_4_30_port, A_ns(29) => SHIFT_n_4_29_port, 
                           A_ns(28) => SHIFT_n_4_28_port, A_ns(27) => 
                           SHIFT_n_4_27_port, A_ns(26) => SHIFT_n_4_26_port, 
                           A_ns(25) => SHIFT_n_4_25_port, A_ns(24) => 
                           SHIFT_n_4_24_port, A_ns(23) => SHIFT_n_4_23_port, 
                           A_ns(22) => SHIFT_n_4_22_port, A_ns(21) => 
                           SHIFT_n_4_21_port, A_ns(20) => SHIFT_n_4_20_port, 
                           A_ns(19) => SHIFT_n_4_19_port, A_ns(18) => 
                           SHIFT_n_4_18_port, A_ns(17) => SHIFT_n_4_17_port, 
                           A_ns(16) => SHIFT_n_4_16_port, A_ns(15) => 
                           SHIFT_n_4_15_port, A_ns(14) => SHIFT_n_4_14_port, 
                           A_ns(13) => SHIFT_n_4_13_port, A_ns(12) => 
                           SHIFT_n_4_12_port, A_ns(11) => SHIFT_n_4_11_port, 
                           A_ns(10) => SHIFT_n_4_10_port, A_ns(9) => 
                           SHIFT_n_4_9_port, A_ns(8) => SHIFT_n_4_8_port, 
                           A_ns(7) => SHIFT_n_4_7_port, A_ns(6) => 
                           SHIFT_n_4_6_port, A_ns(5) => SHIFT_n_4_5_port, 
                           A_ns(4) => SHIFT_n_4_4_port, A_ns(3) => 
                           SHIFT_n_4_3_port, A_ns(2) => SHIFT_n_4_2_port, 
                           A_ns(1) => SHIFT_n_4_1_port, A_ns(0) => 
                           SHIFT_n_4_0_port, B(41) => B(31), B(40) => B(31), 
                           B(39) => B(31), B(38) => B(31), B(37) => B(31), 
                           B(36) => B(31), B(35) => B(31), B(34) => B(31), 
                           B(33) => B(31), B(32) => B(31), B(31) => B(31), 
                           B(30) => B(30), B(29) => B(29), B(28) => B(28), 
                           B(27) => B(27), B(26) => B(26), B(25) => B(25), 
                           B(24) => B(24), B(23) => B(23), B(22) => B(22), 
                           B(21) => B(21), B(20) => B(20), B(19) => B(19), 
                           B(18) => B(18), B(17) => B(17), B(16) => B(16), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => B(0), O(41) => 
                           OTMP_4_41_port, O(40) => OTMP_4_40_port, O(39) => 
                           OTMP_4_39_port, O(38) => OTMP_4_38_port, O(37) => 
                           OTMP_4_37_port, O(36) => OTMP_4_36_port, O(35) => 
                           OTMP_4_35_port, O(34) => OTMP_4_34_port, O(33) => 
                           OTMP_4_33_port, O(32) => OTMP_4_32_port, O(31) => 
                           OTMP_4_31_port, O(30) => OTMP_4_30_port, O(29) => 
                           OTMP_4_29_port, O(28) => OTMP_4_28_port, O(27) => 
                           OTMP_4_27_port, O(26) => OTMP_4_26_port, O(25) => 
                           OTMP_4_25_port, O(24) => OTMP_4_24_port, O(23) => 
                           OTMP_4_23_port, O(22) => OTMP_4_22_port, O(21) => 
                           OTMP_4_21_port, O(20) => OTMP_4_20_port, O(19) => 
                           OTMP_4_19_port, O(18) => OTMP_4_18_port, O(17) => 
                           OTMP_4_17_port, O(16) => OTMP_4_16_port, O(15) => 
                           OTMP_4_15_port, O(14) => OTMP_4_14_port, O(13) => 
                           OTMP_4_13_port, O(12) => OTMP_4_12_port, O(11) => 
                           OTMP_4_11_port, O(10) => OTMP_4_10_port, O(9) => 
                           OTMP_4_9_port, O(8) => OTMP_4_8_port, O(7) => 
                           OTMP_4_7_port, O(6) => OTMP_4_6_port, O(5) => 
                           OTMP_4_5_port, O(4) => OTMP_4_4_port, O(3) => 
                           OTMP_4_3_port, O(2) => OTMP_4_2_port, O(1) => 
                           OTMP_4_1_port, O(0) => n_1097, A_so(41) => 
                           SHIFT_5_41_port, A_so(40) => SHIFT_5_40_port, 
                           A_so(39) => SHIFT_5_39_port, A_so(38) => 
                           SHIFT_5_38_port, A_so(37) => SHIFT_5_37_port, 
                           A_so(36) => SHIFT_5_36_port, A_so(35) => 
                           SHIFT_5_35_port, A_so(34) => SHIFT_5_34_port, 
                           A_so(33) => SHIFT_5_33_port, A_so(32) => 
                           SHIFT_5_32_port, A_so(31) => SHIFT_5_31_port, 
                           A_so(30) => SHIFT_5_30_port, A_so(29) => 
                           SHIFT_5_29_port, A_so(28) => SHIFT_5_28_port, 
                           A_so(27) => SHIFT_5_27_port, A_so(26) => 
                           SHIFT_5_26_port, A_so(25) => SHIFT_5_25_port, 
                           A_so(24) => SHIFT_5_24_port, A_so(23) => 
                           SHIFT_5_23_port, A_so(22) => SHIFT_5_22_port, 
                           A_so(21) => SHIFT_5_21_port, A_so(20) => 
                           SHIFT_5_20_port, A_so(19) => SHIFT_5_19_port, 
                           A_so(18) => SHIFT_5_18_port, A_so(17) => 
                           SHIFT_5_17_port, A_so(16) => SHIFT_5_16_port, 
                           A_so(15) => SHIFT_5_15_port, A_so(14) => 
                           SHIFT_5_14_port, A_so(13) => SHIFT_5_13_port, 
                           A_so(12) => SHIFT_5_12_port, A_so(11) => 
                           SHIFT_5_11_port, A_so(10) => SHIFT_5_10_port, 
                           A_so(9) => SHIFT_5_9_port, A_so(8) => SHIFT_5_8_port
                           , A_so(7) => SHIFT_5_7_port, A_so(6) => 
                           SHIFT_5_6_port, A_so(5) => SHIFT_5_5_port, A_so(4) 
                           => SHIFT_5_4_port, A_so(3) => SHIFT_5_3_port, 
                           A_so(2) => SHIFT_5_2_port, A_so(1) => n_1098, 
                           A_so(0) => n_1099, A_nso(41) => SHIFT_n_5_41_port, 
                           A_nso(40) => SHIFT_n_5_40_port, A_nso(39) => 
                           SHIFT_n_5_39_port, A_nso(38) => SHIFT_n_5_38_port, 
                           A_nso(37) => SHIFT_n_5_37_port, A_nso(36) => 
                           SHIFT_n_5_36_port, A_nso(35) => SHIFT_n_5_35_port, 
                           A_nso(34) => SHIFT_n_5_34_port, A_nso(33) => 
                           SHIFT_n_5_33_port, A_nso(32) => SHIFT_n_5_32_port, 
                           A_nso(31) => SHIFT_n_5_31_port, A_nso(30) => 
                           SHIFT_n_5_30_port, A_nso(29) => SHIFT_n_5_29_port, 
                           A_nso(28) => SHIFT_n_5_28_port, A_nso(27) => 
                           SHIFT_n_5_27_port, A_nso(26) => SHIFT_n_5_26_port, 
                           A_nso(25) => SHIFT_n_5_25_port, A_nso(24) => 
                           SHIFT_n_5_24_port, A_nso(23) => SHIFT_n_5_23_port, 
                           A_nso(22) => SHIFT_n_5_22_port, A_nso(21) => 
                           SHIFT_n_5_21_port, A_nso(20) => SHIFT_n_5_20_port, 
                           A_nso(19) => SHIFT_n_5_19_port, A_nso(18) => 
                           SHIFT_n_5_18_port, A_nso(17) => SHIFT_n_5_17_port, 
                           A_nso(16) => SHIFT_n_5_16_port, A_nso(15) => 
                           SHIFT_n_5_15_port, A_nso(14) => SHIFT_n_5_14_port, 
                           A_nso(13) => SHIFT_n_5_13_port, A_nso(12) => 
                           SHIFT_n_5_12_port, A_nso(11) => SHIFT_n_5_11_port, 
                           A_nso(10) => SHIFT_n_5_10_port, A_nso(9) => 
                           SHIFT_n_5_9_port, A_nso(8) => SHIFT_n_5_8_port, 
                           A_nso(7) => SHIFT_n_5_7_port, A_nso(6) => 
                           SHIFT_n_5_6_port, A_nso(5) => SHIFT_n_5_5_port, 
                           A_nso(4) => SHIFT_n_5_4_port, A_nso(3) => 
                           SHIFT_n_5_3_port, A_nso(2) => SHIFT_n_5_2_port, 
                           A_nso(1) => n_1100, A_nso(0) => n_1101);
   ENC_5 : BOOTHENC_NBIT44_i10 port map( A_s(43) => SHIFT_5_41_port, A_s(42) =>
                           SHIFT_5_41_port, A_s(41) => SHIFT_5_41_port, A_s(40)
                           => SHIFT_5_40_port, A_s(39) => SHIFT_5_39_port, 
                           A_s(38) => SHIFT_5_38_port, A_s(37) => 
                           SHIFT_5_37_port, A_s(36) => SHIFT_5_36_port, A_s(35)
                           => SHIFT_5_35_port, A_s(34) => SHIFT_5_34_port, 
                           A_s(33) => SHIFT_5_33_port, A_s(32) => 
                           SHIFT_5_32_port, A_s(31) => SHIFT_5_31_port, A_s(30)
                           => SHIFT_5_30_port, A_s(29) => SHIFT_5_29_port, 
                           A_s(28) => SHIFT_5_28_port, A_s(27) => 
                           SHIFT_5_27_port, A_s(26) => SHIFT_5_26_port, A_s(25)
                           => SHIFT_5_25_port, A_s(24) => SHIFT_5_24_port, 
                           A_s(23) => SHIFT_5_23_port, A_s(22) => 
                           SHIFT_5_22_port, A_s(21) => SHIFT_5_21_port, A_s(20)
                           => SHIFT_5_20_port, A_s(19) => SHIFT_5_19_port, 
                           A_s(18) => SHIFT_5_18_port, A_s(17) => 
                           SHIFT_5_17_port, A_s(16) => SHIFT_5_16_port, A_s(15)
                           => SHIFT_5_15_port, A_s(14) => SHIFT_5_14_port, 
                           A_s(13) => SHIFT_5_13_port, A_s(12) => 
                           SHIFT_5_12_port, A_s(11) => SHIFT_5_11_port, A_s(10)
                           => SHIFT_5_10_port, A_s(9) => SHIFT_5_9_port, A_s(8)
                           => SHIFT_5_8_port, A_s(7) => SHIFT_5_7_port, A_s(6) 
                           => SHIFT_5_6_port, A_s(5) => SHIFT_5_5_port, A_s(4) 
                           => SHIFT_5_4_port, A_s(3) => SHIFT_5_3_port, A_s(2) 
                           => SHIFT_5_2_port, A_s(1) => SHIFT_5_1_port, A_s(0) 
                           => SHIFT_5_0_port, A_ns(43) => SHIFT_n_5_41_port, 
                           A_ns(42) => SHIFT_n_5_41_port, A_ns(41) => 
                           SHIFT_n_5_41_port, A_ns(40) => SHIFT_n_5_40_port, 
                           A_ns(39) => SHIFT_n_5_39_port, A_ns(38) => 
                           SHIFT_n_5_38_port, A_ns(37) => SHIFT_n_5_37_port, 
                           A_ns(36) => SHIFT_n_5_36_port, A_ns(35) => 
                           SHIFT_n_5_35_port, A_ns(34) => SHIFT_n_5_34_port, 
                           A_ns(33) => SHIFT_n_5_33_port, A_ns(32) => 
                           SHIFT_n_5_32_port, A_ns(31) => SHIFT_n_5_31_port, 
                           A_ns(30) => SHIFT_n_5_30_port, A_ns(29) => 
                           SHIFT_n_5_29_port, A_ns(28) => SHIFT_n_5_28_port, 
                           A_ns(27) => SHIFT_n_5_27_port, A_ns(26) => 
                           SHIFT_n_5_26_port, A_ns(25) => SHIFT_n_5_25_port, 
                           A_ns(24) => SHIFT_n_5_24_port, A_ns(23) => 
                           SHIFT_n_5_23_port, A_ns(22) => SHIFT_n_5_22_port, 
                           A_ns(21) => SHIFT_n_5_21_port, A_ns(20) => 
                           SHIFT_n_5_20_port, A_ns(19) => SHIFT_n_5_19_port, 
                           A_ns(18) => SHIFT_n_5_18_port, A_ns(17) => 
                           SHIFT_n_5_17_port, A_ns(16) => SHIFT_n_5_16_port, 
                           A_ns(15) => SHIFT_n_5_15_port, A_ns(14) => 
                           SHIFT_n_5_14_port, A_ns(13) => SHIFT_n_5_13_port, 
                           A_ns(12) => SHIFT_n_5_12_port, A_ns(11) => 
                           SHIFT_n_5_11_port, A_ns(10) => SHIFT_n_5_10_port, 
                           A_ns(9) => SHIFT_n_5_9_port, A_ns(8) => 
                           SHIFT_n_5_8_port, A_ns(7) => SHIFT_n_5_7_port, 
                           A_ns(6) => SHIFT_n_5_6_port, A_ns(5) => 
                           SHIFT_n_5_5_port, A_ns(4) => SHIFT_n_5_4_port, 
                           A_ns(3) => SHIFT_n_5_3_port, A_ns(2) => 
                           SHIFT_n_5_2_port, A_ns(1) => SHIFT_n_5_1_port, 
                           A_ns(0) => SHIFT_n_5_0_port, B(43) => B(31), B(42) 
                           => B(31), B(41) => B(31), B(40) => B(31), B(39) => 
                           B(31), B(38) => B(31), B(37) => B(31), B(36) => 
                           B(31), B(35) => B(31), B(34) => B(31), B(33) => 
                           B(31), B(32) => B(31), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), O(43) => OTMP_5_43_port, 
                           O(42) => OTMP_5_42_port, O(41) => OTMP_5_41_port, 
                           O(40) => OTMP_5_40_port, O(39) => OTMP_5_39_port, 
                           O(38) => OTMP_5_38_port, O(37) => OTMP_5_37_port, 
                           O(36) => OTMP_5_36_port, O(35) => OTMP_5_35_port, 
                           O(34) => OTMP_5_34_port, O(33) => OTMP_5_33_port, 
                           O(32) => OTMP_5_32_port, O(31) => OTMP_5_31_port, 
                           O(30) => OTMP_5_30_port, O(29) => OTMP_5_29_port, 
                           O(28) => OTMP_5_28_port, O(27) => OTMP_5_27_port, 
                           O(26) => OTMP_5_26_port, O(25) => OTMP_5_25_port, 
                           O(24) => OTMP_5_24_port, O(23) => OTMP_5_23_port, 
                           O(22) => OTMP_5_22_port, O(21) => OTMP_5_21_port, 
                           O(20) => OTMP_5_20_port, O(19) => OTMP_5_19_port, 
                           O(18) => OTMP_5_18_port, O(17) => OTMP_5_17_port, 
                           O(16) => OTMP_5_16_port, O(15) => OTMP_5_15_port, 
                           O(14) => OTMP_5_14_port, O(13) => OTMP_5_13_port, 
                           O(12) => OTMP_5_12_port, O(11) => OTMP_5_11_port, 
                           O(10) => OTMP_5_10_port, O(9) => OTMP_5_9_port, O(8)
                           => OTMP_5_8_port, O(7) => OTMP_5_7_port, O(6) => 
                           OTMP_5_6_port, O(5) => OTMP_5_5_port, O(4) => 
                           OTMP_5_4_port, O(3) => OTMP_5_3_port, O(2) => 
                           OTMP_5_2_port, O(1) => OTMP_5_1_port, O(0) => n_1102
                           , A_so(43) => SHIFT_6_43_port, A_so(42) => 
                           SHIFT_6_42_port, A_so(41) => SHIFT_6_41_port, 
                           A_so(40) => SHIFT_6_40_port, A_so(39) => 
                           SHIFT_6_39_port, A_so(38) => SHIFT_6_38_port, 
                           A_so(37) => SHIFT_6_37_port, A_so(36) => 
                           SHIFT_6_36_port, A_so(35) => SHIFT_6_35_port, 
                           A_so(34) => SHIFT_6_34_port, A_so(33) => 
                           SHIFT_6_33_port, A_so(32) => SHIFT_6_32_port, 
                           A_so(31) => SHIFT_6_31_port, A_so(30) => 
                           SHIFT_6_30_port, A_so(29) => SHIFT_6_29_port, 
                           A_so(28) => SHIFT_6_28_port, A_so(27) => 
                           SHIFT_6_27_port, A_so(26) => SHIFT_6_26_port, 
                           A_so(25) => SHIFT_6_25_port, A_so(24) => 
                           SHIFT_6_24_port, A_so(23) => SHIFT_6_23_port, 
                           A_so(22) => SHIFT_6_22_port, A_so(21) => 
                           SHIFT_6_21_port, A_so(20) => SHIFT_6_20_port, 
                           A_so(19) => SHIFT_6_19_port, A_so(18) => 
                           SHIFT_6_18_port, A_so(17) => SHIFT_6_17_port, 
                           A_so(16) => SHIFT_6_16_port, A_so(15) => 
                           SHIFT_6_15_port, A_so(14) => SHIFT_6_14_port, 
                           A_so(13) => SHIFT_6_13_port, A_so(12) => 
                           SHIFT_6_12_port, A_so(11) => SHIFT_6_11_port, 
                           A_so(10) => SHIFT_6_10_port, A_so(9) => 
                           SHIFT_6_9_port, A_so(8) => SHIFT_6_8_port, A_so(7) 
                           => SHIFT_6_7_port, A_so(6) => SHIFT_6_6_port, 
                           A_so(5) => SHIFT_6_5_port, A_so(4) => SHIFT_6_4_port
                           , A_so(3) => SHIFT_6_3_port, A_so(2) => 
                           SHIFT_6_2_port, A_so(1) => n_1103, A_so(0) => n_1104
                           , A_nso(43) => SHIFT_n_6_43_port, A_nso(42) => 
                           SHIFT_n_6_42_port, A_nso(41) => SHIFT_n_6_41_port, 
                           A_nso(40) => SHIFT_n_6_40_port, A_nso(39) => 
                           SHIFT_n_6_39_port, A_nso(38) => SHIFT_n_6_38_port, 
                           A_nso(37) => SHIFT_n_6_37_port, A_nso(36) => 
                           SHIFT_n_6_36_port, A_nso(35) => SHIFT_n_6_35_port, 
                           A_nso(34) => SHIFT_n_6_34_port, A_nso(33) => 
                           SHIFT_n_6_33_port, A_nso(32) => SHIFT_n_6_32_port, 
                           A_nso(31) => SHIFT_n_6_31_port, A_nso(30) => 
                           SHIFT_n_6_30_port, A_nso(29) => SHIFT_n_6_29_port, 
                           A_nso(28) => SHIFT_n_6_28_port, A_nso(27) => 
                           SHIFT_n_6_27_port, A_nso(26) => SHIFT_n_6_26_port, 
                           A_nso(25) => SHIFT_n_6_25_port, A_nso(24) => 
                           SHIFT_n_6_24_port, A_nso(23) => SHIFT_n_6_23_port, 
                           A_nso(22) => SHIFT_n_6_22_port, A_nso(21) => 
                           SHIFT_n_6_21_port, A_nso(20) => SHIFT_n_6_20_port, 
                           A_nso(19) => SHIFT_n_6_19_port, A_nso(18) => 
                           SHIFT_n_6_18_port, A_nso(17) => SHIFT_n_6_17_port, 
                           A_nso(16) => SHIFT_n_6_16_port, A_nso(15) => 
                           SHIFT_n_6_15_port, A_nso(14) => SHIFT_n_6_14_port, 
                           A_nso(13) => SHIFT_n_6_13_port, A_nso(12) => 
                           SHIFT_n_6_12_port, A_nso(11) => SHIFT_n_6_11_port, 
                           A_nso(10) => SHIFT_n_6_10_port, A_nso(9) => 
                           SHIFT_n_6_9_port, A_nso(8) => SHIFT_n_6_8_port, 
                           A_nso(7) => SHIFT_n_6_7_port, A_nso(6) => 
                           SHIFT_n_6_6_port, A_nso(5) => SHIFT_n_6_5_port, 
                           A_nso(4) => SHIFT_n_6_4_port, A_nso(3) => 
                           SHIFT_n_6_3_port, A_nso(2) => SHIFT_n_6_2_port, 
                           A_nso(1) => n_1105, A_nso(0) => n_1106);
   ENC_6 : BOOTHENC_NBIT46_i12 port map( A_s(45) => SHIFT_6_43_port, A_s(44) =>
                           SHIFT_6_43_port, A_s(43) => SHIFT_6_43_port, A_s(42)
                           => SHIFT_6_42_port, A_s(41) => SHIFT_6_41_port, 
                           A_s(40) => SHIFT_6_40_port, A_s(39) => 
                           SHIFT_6_39_port, A_s(38) => SHIFT_6_38_port, A_s(37)
                           => SHIFT_6_37_port, A_s(36) => SHIFT_6_36_port, 
                           A_s(35) => SHIFT_6_35_port, A_s(34) => 
                           SHIFT_6_34_port, A_s(33) => SHIFT_6_33_port, A_s(32)
                           => SHIFT_6_32_port, A_s(31) => SHIFT_6_31_port, 
                           A_s(30) => SHIFT_6_30_port, A_s(29) => 
                           SHIFT_6_29_port, A_s(28) => SHIFT_6_28_port, A_s(27)
                           => SHIFT_6_27_port, A_s(26) => SHIFT_6_26_port, 
                           A_s(25) => SHIFT_6_25_port, A_s(24) => 
                           SHIFT_6_24_port, A_s(23) => SHIFT_6_23_port, A_s(22)
                           => SHIFT_6_22_port, A_s(21) => SHIFT_6_21_port, 
                           A_s(20) => SHIFT_6_20_port, A_s(19) => 
                           SHIFT_6_19_port, A_s(18) => SHIFT_6_18_port, A_s(17)
                           => SHIFT_6_17_port, A_s(16) => SHIFT_6_16_port, 
                           A_s(15) => SHIFT_6_15_port, A_s(14) => 
                           SHIFT_6_14_port, A_s(13) => SHIFT_6_13_port, A_s(12)
                           => SHIFT_6_12_port, A_s(11) => SHIFT_6_11_port, 
                           A_s(10) => SHIFT_6_10_port, A_s(9) => SHIFT_6_9_port
                           , A_s(8) => SHIFT_6_8_port, A_s(7) => SHIFT_6_7_port
                           , A_s(6) => SHIFT_6_6_port, A_s(5) => SHIFT_6_5_port
                           , A_s(4) => SHIFT_6_4_port, A_s(3) => SHIFT_6_3_port
                           , A_s(2) => SHIFT_6_2_port, A_s(1) => SHIFT_6_1_port
                           , A_s(0) => SHIFT_6_0_port, A_ns(45) => 
                           SHIFT_n_6_43_port, A_ns(44) => SHIFT_n_6_43_port, 
                           A_ns(43) => SHIFT_n_6_43_port, A_ns(42) => 
                           SHIFT_n_6_42_port, A_ns(41) => SHIFT_n_6_41_port, 
                           A_ns(40) => SHIFT_n_6_40_port, A_ns(39) => 
                           SHIFT_n_6_39_port, A_ns(38) => SHIFT_n_6_38_port, 
                           A_ns(37) => SHIFT_n_6_37_port, A_ns(36) => 
                           SHIFT_n_6_36_port, A_ns(35) => SHIFT_n_6_35_port, 
                           A_ns(34) => SHIFT_n_6_34_port, A_ns(33) => 
                           SHIFT_n_6_33_port, A_ns(32) => SHIFT_n_6_32_port, 
                           A_ns(31) => SHIFT_n_6_31_port, A_ns(30) => 
                           SHIFT_n_6_30_port, A_ns(29) => SHIFT_n_6_29_port, 
                           A_ns(28) => SHIFT_n_6_28_port, A_ns(27) => 
                           SHIFT_n_6_27_port, A_ns(26) => SHIFT_n_6_26_port, 
                           A_ns(25) => SHIFT_n_6_25_port, A_ns(24) => 
                           SHIFT_n_6_24_port, A_ns(23) => SHIFT_n_6_23_port, 
                           A_ns(22) => SHIFT_n_6_22_port, A_ns(21) => 
                           SHIFT_n_6_21_port, A_ns(20) => SHIFT_n_6_20_port, 
                           A_ns(19) => SHIFT_n_6_19_port, A_ns(18) => 
                           SHIFT_n_6_18_port, A_ns(17) => SHIFT_n_6_17_port, 
                           A_ns(16) => SHIFT_n_6_16_port, A_ns(15) => 
                           SHIFT_n_6_15_port, A_ns(14) => SHIFT_n_6_14_port, 
                           A_ns(13) => SHIFT_n_6_13_port, A_ns(12) => 
                           SHIFT_n_6_12_port, A_ns(11) => SHIFT_n_6_11_port, 
                           A_ns(10) => SHIFT_n_6_10_port, A_ns(9) => 
                           SHIFT_n_6_9_port, A_ns(8) => SHIFT_n_6_8_port, 
                           A_ns(7) => SHIFT_n_6_7_port, A_ns(6) => 
                           SHIFT_n_6_6_port, A_ns(5) => SHIFT_n_6_5_port, 
                           A_ns(4) => SHIFT_n_6_4_port, A_ns(3) => 
                           SHIFT_n_6_3_port, A_ns(2) => SHIFT_n_6_2_port, 
                           A_ns(1) => SHIFT_n_6_1_port, A_ns(0) => 
                           SHIFT_n_6_0_port, B(45) => B(31), B(44) => B(31), 
                           B(43) => B(31), B(42) => B(31), B(41) => B(31), 
                           B(40) => B(31), B(39) => B(31), B(38) => B(31), 
                           B(37) => B(31), B(36) => B(31), B(35) => B(31), 
                           B(34) => B(31), B(33) => B(31), B(32) => B(31), 
                           B(31) => B(31), B(30) => B(30), B(29) => B(29), 
                           B(28) => B(28), B(27) => B(27), B(26) => B(26), 
                           B(25) => B(25), B(24) => B(24), B(23) => B(23), 
                           B(22) => B(22), B(21) => B(21), B(20) => B(20), 
                           B(19) => B(19), B(18) => B(18), B(17) => B(17), 
                           B(16) => B(16), B(15) => B(15), B(14) => B(14), 
                           B(13) => B(13), B(12) => B(12), B(11) => B(11), 
                           B(10) => B(10), B(9) => B(9), B(8) => B(8), B(7) => 
                           B(7), B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3)
                           => B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), 
                           O(45) => OTMP_6_45_port, O(44) => OTMP_6_44_port, 
                           O(43) => OTMP_6_43_port, O(42) => OTMP_6_42_port, 
                           O(41) => OTMP_6_41_port, O(40) => OTMP_6_40_port, 
                           O(39) => OTMP_6_39_port, O(38) => OTMP_6_38_port, 
                           O(37) => OTMP_6_37_port, O(36) => OTMP_6_36_port, 
                           O(35) => OTMP_6_35_port, O(34) => OTMP_6_34_port, 
                           O(33) => OTMP_6_33_port, O(32) => OTMP_6_32_port, 
                           O(31) => OTMP_6_31_port, O(30) => OTMP_6_30_port, 
                           O(29) => OTMP_6_29_port, O(28) => OTMP_6_28_port, 
                           O(27) => OTMP_6_27_port, O(26) => OTMP_6_26_port, 
                           O(25) => OTMP_6_25_port, O(24) => OTMP_6_24_port, 
                           O(23) => OTMP_6_23_port, O(22) => OTMP_6_22_port, 
                           O(21) => OTMP_6_21_port, O(20) => OTMP_6_20_port, 
                           O(19) => OTMP_6_19_port, O(18) => OTMP_6_18_port, 
                           O(17) => OTMP_6_17_port, O(16) => OTMP_6_16_port, 
                           O(15) => OTMP_6_15_port, O(14) => OTMP_6_14_port, 
                           O(13) => OTMP_6_13_port, O(12) => OTMP_6_12_port, 
                           O(11) => OTMP_6_11_port, O(10) => OTMP_6_10_port, 
                           O(9) => OTMP_6_9_port, O(8) => OTMP_6_8_port, O(7) 
                           => OTMP_6_7_port, O(6) => OTMP_6_6_port, O(5) => 
                           OTMP_6_5_port, O(4) => OTMP_6_4_port, O(3) => 
                           OTMP_6_3_port, O(2) => OTMP_6_2_port, O(1) => 
                           OTMP_6_1_port, O(0) => n_1107, A_so(45) => 
                           SHIFT_7_45_port, A_so(44) => SHIFT_7_44_port, 
                           A_so(43) => SHIFT_7_43_port, A_so(42) => 
                           SHIFT_7_42_port, A_so(41) => SHIFT_7_41_port, 
                           A_so(40) => SHIFT_7_40_port, A_so(39) => 
                           SHIFT_7_39_port, A_so(38) => SHIFT_7_38_port, 
                           A_so(37) => SHIFT_7_37_port, A_so(36) => 
                           SHIFT_7_36_port, A_so(35) => SHIFT_7_35_port, 
                           A_so(34) => SHIFT_7_34_port, A_so(33) => 
                           SHIFT_7_33_port, A_so(32) => SHIFT_7_32_port, 
                           A_so(31) => SHIFT_7_31_port, A_so(30) => 
                           SHIFT_7_30_port, A_so(29) => SHIFT_7_29_port, 
                           A_so(28) => SHIFT_7_28_port, A_so(27) => 
                           SHIFT_7_27_port, A_so(26) => SHIFT_7_26_port, 
                           A_so(25) => SHIFT_7_25_port, A_so(24) => 
                           SHIFT_7_24_port, A_so(23) => SHIFT_7_23_port, 
                           A_so(22) => SHIFT_7_22_port, A_so(21) => 
                           SHIFT_7_21_port, A_so(20) => SHIFT_7_20_port, 
                           A_so(19) => SHIFT_7_19_port, A_so(18) => 
                           SHIFT_7_18_port, A_so(17) => SHIFT_7_17_port, 
                           A_so(16) => SHIFT_7_16_port, A_so(15) => 
                           SHIFT_7_15_port, A_so(14) => SHIFT_7_14_port, 
                           A_so(13) => SHIFT_7_13_port, A_so(12) => 
                           SHIFT_7_12_port, A_so(11) => SHIFT_7_11_port, 
                           A_so(10) => SHIFT_7_10_port, A_so(9) => 
                           SHIFT_7_9_port, A_so(8) => SHIFT_7_8_port, A_so(7) 
                           => SHIFT_7_7_port, A_so(6) => SHIFT_7_6_port, 
                           A_so(5) => SHIFT_7_5_port, A_so(4) => SHIFT_7_4_port
                           , A_so(3) => SHIFT_7_3_port, A_so(2) => 
                           SHIFT_7_2_port, A_so(1) => n_1108, A_so(0) => n_1109
                           , A_nso(45) => SHIFT_n_7_45_port, A_nso(44) => 
                           SHIFT_n_7_44_port, A_nso(43) => SHIFT_n_7_43_port, 
                           A_nso(42) => SHIFT_n_7_42_port, A_nso(41) => 
                           SHIFT_n_7_41_port, A_nso(40) => SHIFT_n_7_40_port, 
                           A_nso(39) => SHIFT_n_7_39_port, A_nso(38) => 
                           SHIFT_n_7_38_port, A_nso(37) => SHIFT_n_7_37_port, 
                           A_nso(36) => SHIFT_n_7_36_port, A_nso(35) => 
                           SHIFT_n_7_35_port, A_nso(34) => SHIFT_n_7_34_port, 
                           A_nso(33) => SHIFT_n_7_33_port, A_nso(32) => 
                           SHIFT_n_7_32_port, A_nso(31) => SHIFT_n_7_31_port, 
                           A_nso(30) => SHIFT_n_7_30_port, A_nso(29) => 
                           SHIFT_n_7_29_port, A_nso(28) => SHIFT_n_7_28_port, 
                           A_nso(27) => SHIFT_n_7_27_port, A_nso(26) => 
                           SHIFT_n_7_26_port, A_nso(25) => SHIFT_n_7_25_port, 
                           A_nso(24) => SHIFT_n_7_24_port, A_nso(23) => 
                           SHIFT_n_7_23_port, A_nso(22) => SHIFT_n_7_22_port, 
                           A_nso(21) => SHIFT_n_7_21_port, A_nso(20) => 
                           SHIFT_n_7_20_port, A_nso(19) => SHIFT_n_7_19_port, 
                           A_nso(18) => SHIFT_n_7_18_port, A_nso(17) => 
                           SHIFT_n_7_17_port, A_nso(16) => SHIFT_n_7_16_port, 
                           A_nso(15) => SHIFT_n_7_15_port, A_nso(14) => 
                           SHIFT_n_7_14_port, A_nso(13) => SHIFT_n_7_13_port, 
                           A_nso(12) => SHIFT_n_7_12_port, A_nso(11) => 
                           SHIFT_n_7_11_port, A_nso(10) => SHIFT_n_7_10_port, 
                           A_nso(9) => SHIFT_n_7_9_port, A_nso(8) => 
                           SHIFT_n_7_8_port, A_nso(7) => SHIFT_n_7_7_port, 
                           A_nso(6) => SHIFT_n_7_6_port, A_nso(5) => 
                           SHIFT_n_7_5_port, A_nso(4) => SHIFT_n_7_4_port, 
                           A_nso(3) => SHIFT_n_7_3_port, A_nso(2) => 
                           SHIFT_n_7_2_port, A_nso(1) => n_1110, A_nso(0) => 
                           n_1111);
   ENC_7 : BOOTHENC_NBIT48_i14 port map( A_s(47) => SHIFT_7_45_port, A_s(46) =>
                           SHIFT_7_45_port, A_s(45) => SHIFT_7_45_port, A_s(44)
                           => SHIFT_7_44_port, A_s(43) => SHIFT_7_43_port, 
                           A_s(42) => SHIFT_7_42_port, A_s(41) => 
                           SHIFT_7_41_port, A_s(40) => SHIFT_7_40_port, A_s(39)
                           => SHIFT_7_39_port, A_s(38) => SHIFT_7_38_port, 
                           A_s(37) => SHIFT_7_37_port, A_s(36) => 
                           SHIFT_7_36_port, A_s(35) => SHIFT_7_35_port, A_s(34)
                           => SHIFT_7_34_port, A_s(33) => SHIFT_7_33_port, 
                           A_s(32) => SHIFT_7_32_port, A_s(31) => 
                           SHIFT_7_31_port, A_s(30) => SHIFT_7_30_port, A_s(29)
                           => SHIFT_7_29_port, A_s(28) => SHIFT_7_28_port, 
                           A_s(27) => SHIFT_7_27_port, A_s(26) => 
                           SHIFT_7_26_port, A_s(25) => SHIFT_7_25_port, A_s(24)
                           => SHIFT_7_24_port, A_s(23) => SHIFT_7_23_port, 
                           A_s(22) => SHIFT_7_22_port, A_s(21) => 
                           SHIFT_7_21_port, A_s(20) => SHIFT_7_20_port, A_s(19)
                           => SHIFT_7_19_port, A_s(18) => SHIFT_7_18_port, 
                           A_s(17) => SHIFT_7_17_port, A_s(16) => 
                           SHIFT_7_16_port, A_s(15) => SHIFT_7_15_port, A_s(14)
                           => SHIFT_7_14_port, A_s(13) => SHIFT_7_13_port, 
                           A_s(12) => SHIFT_7_12_port, A_s(11) => 
                           SHIFT_7_11_port, A_s(10) => SHIFT_7_10_port, A_s(9) 
                           => SHIFT_7_9_port, A_s(8) => SHIFT_7_8_port, A_s(7) 
                           => SHIFT_7_7_port, A_s(6) => SHIFT_7_6_port, A_s(5) 
                           => SHIFT_7_5_port, A_s(4) => SHIFT_7_4_port, A_s(3) 
                           => SHIFT_7_3_port, A_s(2) => SHIFT_7_2_port, A_s(1) 
                           => SHIFT_7_1_port, A_s(0) => SHIFT_7_0_port, 
                           A_ns(47) => SHIFT_n_7_45_port, A_ns(46) => 
                           SHIFT_n_7_45_port, A_ns(45) => SHIFT_n_7_45_port, 
                           A_ns(44) => SHIFT_n_7_44_port, A_ns(43) => 
                           SHIFT_n_7_43_port, A_ns(42) => SHIFT_n_7_42_port, 
                           A_ns(41) => SHIFT_n_7_41_port, A_ns(40) => 
                           SHIFT_n_7_40_port, A_ns(39) => SHIFT_n_7_39_port, 
                           A_ns(38) => SHIFT_n_7_38_port, A_ns(37) => 
                           SHIFT_n_7_37_port, A_ns(36) => SHIFT_n_7_36_port, 
                           A_ns(35) => SHIFT_n_7_35_port, A_ns(34) => 
                           SHIFT_n_7_34_port, A_ns(33) => SHIFT_n_7_33_port, 
                           A_ns(32) => SHIFT_n_7_32_port, A_ns(31) => 
                           SHIFT_n_7_31_port, A_ns(30) => SHIFT_n_7_30_port, 
                           A_ns(29) => SHIFT_n_7_29_port, A_ns(28) => 
                           SHIFT_n_7_28_port, A_ns(27) => SHIFT_n_7_27_port, 
                           A_ns(26) => SHIFT_n_7_26_port, A_ns(25) => 
                           SHIFT_n_7_25_port, A_ns(24) => SHIFT_n_7_24_port, 
                           A_ns(23) => SHIFT_n_7_23_port, A_ns(22) => 
                           SHIFT_n_7_22_port, A_ns(21) => SHIFT_n_7_21_port, 
                           A_ns(20) => SHIFT_n_7_20_port, A_ns(19) => 
                           SHIFT_n_7_19_port, A_ns(18) => SHIFT_n_7_18_port, 
                           A_ns(17) => SHIFT_n_7_17_port, A_ns(16) => 
                           SHIFT_n_7_16_port, A_ns(15) => SHIFT_n_7_15_port, 
                           A_ns(14) => SHIFT_n_7_14_port, A_ns(13) => 
                           SHIFT_n_7_13_port, A_ns(12) => SHIFT_n_7_12_port, 
                           A_ns(11) => SHIFT_n_7_11_port, A_ns(10) => 
                           SHIFT_n_7_10_port, A_ns(9) => SHIFT_n_7_9_port, 
                           A_ns(8) => SHIFT_n_7_8_port, A_ns(7) => 
                           SHIFT_n_7_7_port, A_ns(6) => SHIFT_n_7_6_port, 
                           A_ns(5) => SHIFT_n_7_5_port, A_ns(4) => 
                           SHIFT_n_7_4_port, A_ns(3) => SHIFT_n_7_3_port, 
                           A_ns(2) => SHIFT_n_7_2_port, A_ns(1) => 
                           SHIFT_n_7_1_port, A_ns(0) => SHIFT_n_7_0_port, B(47)
                           => B(31), B(46) => B(31), B(45) => B(31), B(44) => 
                           B(31), B(43) => B(31), B(42) => B(31), B(41) => 
                           B(31), B(40) => B(31), B(39) => B(31), B(38) => 
                           B(31), B(37) => B(31), B(36) => B(31), B(35) => 
                           B(31), B(34) => B(31), B(33) => B(31), B(32) => 
                           B(31), B(31) => B(31), B(30) => B(30), B(29) => 
                           B(29), B(28) => B(28), B(27) => B(27), B(26) => 
                           B(26), B(25) => B(25), B(24) => B(24), B(23) => 
                           B(23), B(22) => B(22), B(21) => B(21), B(20) => 
                           B(20), B(19) => B(19), B(18) => B(18), B(17) => 
                           B(17), B(16) => B(16), B(15) => B(15), B(14) => 
                           B(14), B(13) => B(13), B(12) => B(12), B(11) => 
                           B(11), B(10) => B(10), B(9) => B(9), B(8) => B(8), 
                           B(7) => B(7), B(6) => B(6), B(5) => B(5), B(4) => 
                           B(4), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), O(47) => OTMP_7_47_port, O(46) => 
                           OTMP_7_46_port, O(45) => OTMP_7_45_port, O(44) => 
                           OTMP_7_44_port, O(43) => OTMP_7_43_port, O(42) => 
                           OTMP_7_42_port, O(41) => OTMP_7_41_port, O(40) => 
                           OTMP_7_40_port, O(39) => OTMP_7_39_port, O(38) => 
                           OTMP_7_38_port, O(37) => OTMP_7_37_port, O(36) => 
                           OTMP_7_36_port, O(35) => OTMP_7_35_port, O(34) => 
                           OTMP_7_34_port, O(33) => OTMP_7_33_port, O(32) => 
                           OTMP_7_32_port, O(31) => OTMP_7_31_port, O(30) => 
                           OTMP_7_30_port, O(29) => OTMP_7_29_port, O(28) => 
                           OTMP_7_28_port, O(27) => OTMP_7_27_port, O(26) => 
                           OTMP_7_26_port, O(25) => OTMP_7_25_port, O(24) => 
                           OTMP_7_24_port, O(23) => OTMP_7_23_port, O(22) => 
                           OTMP_7_22_port, O(21) => OTMP_7_21_port, O(20) => 
                           OTMP_7_20_port, O(19) => OTMP_7_19_port, O(18) => 
                           OTMP_7_18_port, O(17) => OTMP_7_17_port, O(16) => 
                           OTMP_7_16_port, O(15) => OTMP_7_15_port, O(14) => 
                           OTMP_7_14_port, O(13) => OTMP_7_13_port, O(12) => 
                           OTMP_7_12_port, O(11) => OTMP_7_11_port, O(10) => 
                           OTMP_7_10_port, O(9) => OTMP_7_9_port, O(8) => 
                           OTMP_7_8_port, O(7) => OTMP_7_7_port, O(6) => 
                           OTMP_7_6_port, O(5) => OTMP_7_5_port, O(4) => 
                           OTMP_7_4_port, O(3) => OTMP_7_3_port, O(2) => 
                           OTMP_7_2_port, O(1) => OTMP_7_1_port, O(0) => n_1112
                           , A_so(47) => SHIFT_8_47_port, A_so(46) => 
                           SHIFT_8_46_port, A_so(45) => SHIFT_8_45_port, 
                           A_so(44) => SHIFT_8_44_port, A_so(43) => 
                           SHIFT_8_43_port, A_so(42) => SHIFT_8_42_port, 
                           A_so(41) => SHIFT_8_41_port, A_so(40) => 
                           SHIFT_8_40_port, A_so(39) => SHIFT_8_39_port, 
                           A_so(38) => SHIFT_8_38_port, A_so(37) => 
                           SHIFT_8_37_port, A_so(36) => SHIFT_8_36_port, 
                           A_so(35) => SHIFT_8_35_port, A_so(34) => 
                           SHIFT_8_34_port, A_so(33) => SHIFT_8_33_port, 
                           A_so(32) => SHIFT_8_32_port, A_so(31) => 
                           SHIFT_8_31_port, A_so(30) => SHIFT_8_30_port, 
                           A_so(29) => SHIFT_8_29_port, A_so(28) => 
                           SHIFT_8_28_port, A_so(27) => SHIFT_8_27_port, 
                           A_so(26) => SHIFT_8_26_port, A_so(25) => 
                           SHIFT_8_25_port, A_so(24) => SHIFT_8_24_port, 
                           A_so(23) => SHIFT_8_23_port, A_so(22) => 
                           SHIFT_8_22_port, A_so(21) => SHIFT_8_21_port, 
                           A_so(20) => SHIFT_8_20_port, A_so(19) => 
                           SHIFT_8_19_port, A_so(18) => SHIFT_8_18_port, 
                           A_so(17) => SHIFT_8_17_port, A_so(16) => 
                           SHIFT_8_16_port, A_so(15) => SHIFT_8_15_port, 
                           A_so(14) => SHIFT_8_14_port, A_so(13) => 
                           SHIFT_8_13_port, A_so(12) => SHIFT_8_12_port, 
                           A_so(11) => SHIFT_8_11_port, A_so(10) => 
                           SHIFT_8_10_port, A_so(9) => SHIFT_8_9_port, A_so(8) 
                           => SHIFT_8_8_port, A_so(7) => SHIFT_8_7_port, 
                           A_so(6) => SHIFT_8_6_port, A_so(5) => SHIFT_8_5_port
                           , A_so(4) => SHIFT_8_4_port, A_so(3) => 
                           SHIFT_8_3_port, A_so(2) => SHIFT_8_2_port, A_so(1) 
                           => n_1113, A_so(0) => n_1114, A_nso(47) => 
                           SHIFT_n_8_47_port, A_nso(46) => SHIFT_n_8_46_port, 
                           A_nso(45) => SHIFT_n_8_45_port, A_nso(44) => 
                           SHIFT_n_8_44_port, A_nso(43) => SHIFT_n_8_43_port, 
                           A_nso(42) => SHIFT_n_8_42_port, A_nso(41) => 
                           SHIFT_n_8_41_port, A_nso(40) => SHIFT_n_8_40_port, 
                           A_nso(39) => SHIFT_n_8_39_port, A_nso(38) => 
                           SHIFT_n_8_38_port, A_nso(37) => SHIFT_n_8_37_port, 
                           A_nso(36) => SHIFT_n_8_36_port, A_nso(35) => 
                           SHIFT_n_8_35_port, A_nso(34) => SHIFT_n_8_34_port, 
                           A_nso(33) => SHIFT_n_8_33_port, A_nso(32) => 
                           SHIFT_n_8_32_port, A_nso(31) => SHIFT_n_8_31_port, 
                           A_nso(30) => SHIFT_n_8_30_port, A_nso(29) => 
                           SHIFT_n_8_29_port, A_nso(28) => SHIFT_n_8_28_port, 
                           A_nso(27) => SHIFT_n_8_27_port, A_nso(26) => 
                           SHIFT_n_8_26_port, A_nso(25) => SHIFT_n_8_25_port, 
                           A_nso(24) => SHIFT_n_8_24_port, A_nso(23) => 
                           SHIFT_n_8_23_port, A_nso(22) => SHIFT_n_8_22_port, 
                           A_nso(21) => SHIFT_n_8_21_port, A_nso(20) => 
                           SHIFT_n_8_20_port, A_nso(19) => SHIFT_n_8_19_port, 
                           A_nso(18) => SHIFT_n_8_18_port, A_nso(17) => 
                           SHIFT_n_8_17_port, A_nso(16) => SHIFT_n_8_16_port, 
                           A_nso(15) => SHIFT_n_8_15_port, A_nso(14) => 
                           SHIFT_n_8_14_port, A_nso(13) => SHIFT_n_8_13_port, 
                           A_nso(12) => SHIFT_n_8_12_port, A_nso(11) => 
                           SHIFT_n_8_11_port, A_nso(10) => SHIFT_n_8_10_port, 
                           A_nso(9) => SHIFT_n_8_9_port, A_nso(8) => 
                           SHIFT_n_8_8_port, A_nso(7) => SHIFT_n_8_7_port, 
                           A_nso(6) => SHIFT_n_8_6_port, A_nso(5) => 
                           SHIFT_n_8_5_port, A_nso(4) => SHIFT_n_8_4_port, 
                           A_nso(3) => SHIFT_n_8_3_port, A_nso(2) => 
                           SHIFT_n_8_2_port, A_nso(1) => n_1115, A_nso(0) => 
                           n_1116);
   ENC_8 : BOOTHENC_NBIT50_i16 port map( A_s(49) => SHIFT_8_47_port, A_s(48) =>
                           SHIFT_8_47_port, A_s(47) => SHIFT_8_47_port, A_s(46)
                           => SHIFT_8_46_port, A_s(45) => SHIFT_8_45_port, 
                           A_s(44) => SHIFT_8_44_port, A_s(43) => 
                           SHIFT_8_43_port, A_s(42) => SHIFT_8_42_port, A_s(41)
                           => SHIFT_8_41_port, A_s(40) => SHIFT_8_40_port, 
                           A_s(39) => SHIFT_8_39_port, A_s(38) => 
                           SHIFT_8_38_port, A_s(37) => SHIFT_8_37_port, A_s(36)
                           => SHIFT_8_36_port, A_s(35) => SHIFT_8_35_port, 
                           A_s(34) => SHIFT_8_34_port, A_s(33) => 
                           SHIFT_8_33_port, A_s(32) => SHIFT_8_32_port, A_s(31)
                           => SHIFT_8_31_port, A_s(30) => SHIFT_8_30_port, 
                           A_s(29) => SHIFT_8_29_port, A_s(28) => 
                           SHIFT_8_28_port, A_s(27) => SHIFT_8_27_port, A_s(26)
                           => SHIFT_8_26_port, A_s(25) => SHIFT_8_25_port, 
                           A_s(24) => SHIFT_8_24_port, A_s(23) => 
                           SHIFT_8_23_port, A_s(22) => SHIFT_8_22_port, A_s(21)
                           => SHIFT_8_21_port, A_s(20) => SHIFT_8_20_port, 
                           A_s(19) => SHIFT_8_19_port, A_s(18) => 
                           SHIFT_8_18_port, A_s(17) => SHIFT_8_17_port, A_s(16)
                           => SHIFT_8_16_port, A_s(15) => SHIFT_8_15_port, 
                           A_s(14) => SHIFT_8_14_port, A_s(13) => 
                           SHIFT_8_13_port, A_s(12) => SHIFT_8_12_port, A_s(11)
                           => SHIFT_8_11_port, A_s(10) => SHIFT_8_10_port, 
                           A_s(9) => SHIFT_8_9_port, A_s(8) => SHIFT_8_8_port, 
                           A_s(7) => SHIFT_8_7_port, A_s(6) => SHIFT_8_6_port, 
                           A_s(5) => SHIFT_8_5_port, A_s(4) => SHIFT_8_4_port, 
                           A_s(3) => SHIFT_8_3_port, A_s(2) => SHIFT_8_2_port, 
                           A_s(1) => SHIFT_8_1_port, A_s(0) => SHIFT_8_0_port, 
                           A_ns(49) => SHIFT_n_8_47_port, A_ns(48) => 
                           SHIFT_n_8_47_port, A_ns(47) => SHIFT_n_8_47_port, 
                           A_ns(46) => SHIFT_n_8_46_port, A_ns(45) => 
                           SHIFT_n_8_45_port, A_ns(44) => SHIFT_n_8_44_port, 
                           A_ns(43) => SHIFT_n_8_43_port, A_ns(42) => 
                           SHIFT_n_8_42_port, A_ns(41) => SHIFT_n_8_41_port, 
                           A_ns(40) => SHIFT_n_8_40_port, A_ns(39) => 
                           SHIFT_n_8_39_port, A_ns(38) => SHIFT_n_8_38_port, 
                           A_ns(37) => SHIFT_n_8_37_port, A_ns(36) => 
                           SHIFT_n_8_36_port, A_ns(35) => SHIFT_n_8_35_port, 
                           A_ns(34) => SHIFT_n_8_34_port, A_ns(33) => 
                           SHIFT_n_8_33_port, A_ns(32) => SHIFT_n_8_32_port, 
                           A_ns(31) => SHIFT_n_8_31_port, A_ns(30) => 
                           SHIFT_n_8_30_port, A_ns(29) => SHIFT_n_8_29_port, 
                           A_ns(28) => SHIFT_n_8_28_port, A_ns(27) => 
                           SHIFT_n_8_27_port, A_ns(26) => SHIFT_n_8_26_port, 
                           A_ns(25) => SHIFT_n_8_25_port, A_ns(24) => 
                           SHIFT_n_8_24_port, A_ns(23) => SHIFT_n_8_23_port, 
                           A_ns(22) => SHIFT_n_8_22_port, A_ns(21) => 
                           SHIFT_n_8_21_port, A_ns(20) => SHIFT_n_8_20_port, 
                           A_ns(19) => SHIFT_n_8_19_port, A_ns(18) => 
                           SHIFT_n_8_18_port, A_ns(17) => SHIFT_n_8_17_port, 
                           A_ns(16) => SHIFT_n_8_16_port, A_ns(15) => 
                           SHIFT_n_8_15_port, A_ns(14) => SHIFT_n_8_14_port, 
                           A_ns(13) => SHIFT_n_8_13_port, A_ns(12) => 
                           SHIFT_n_8_12_port, A_ns(11) => SHIFT_n_8_11_port, 
                           A_ns(10) => SHIFT_n_8_10_port, A_ns(9) => 
                           SHIFT_n_8_9_port, A_ns(8) => SHIFT_n_8_8_port, 
                           A_ns(7) => SHIFT_n_8_7_port, A_ns(6) => 
                           SHIFT_n_8_6_port, A_ns(5) => SHIFT_n_8_5_port, 
                           A_ns(4) => SHIFT_n_8_4_port, A_ns(3) => 
                           SHIFT_n_8_3_port, A_ns(2) => SHIFT_n_8_2_port, 
                           A_ns(1) => SHIFT_n_8_1_port, A_ns(0) => 
                           SHIFT_n_8_0_port, B(49) => B(31), B(48) => B(31), 
                           B(47) => B(31), B(46) => B(31), B(45) => B(31), 
                           B(44) => B(31), B(43) => B(31), B(42) => B(31), 
                           B(41) => B(31), B(40) => B(31), B(39) => B(31), 
                           B(38) => B(31), B(37) => B(31), B(36) => B(31), 
                           B(35) => B(31), B(34) => B(31), B(33) => B(31), 
                           B(32) => B(31), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), O(49) => OTMP_8_49_port, O(48) 
                           => OTMP_8_48_port, O(47) => OTMP_8_47_port, O(46) =>
                           OTMP_8_46_port, O(45) => OTMP_8_45_port, O(44) => 
                           OTMP_8_44_port, O(43) => OTMP_8_43_port, O(42) => 
                           OTMP_8_42_port, O(41) => OTMP_8_41_port, O(40) => 
                           OTMP_8_40_port, O(39) => OTMP_8_39_port, O(38) => 
                           OTMP_8_38_port, O(37) => OTMP_8_37_port, O(36) => 
                           OTMP_8_36_port, O(35) => OTMP_8_35_port, O(34) => 
                           OTMP_8_34_port, O(33) => OTMP_8_33_port, O(32) => 
                           OTMP_8_32_port, O(31) => OTMP_8_31_port, O(30) => 
                           OTMP_8_30_port, O(29) => OTMP_8_29_port, O(28) => 
                           OTMP_8_28_port, O(27) => OTMP_8_27_port, O(26) => 
                           OTMP_8_26_port, O(25) => OTMP_8_25_port, O(24) => 
                           OTMP_8_24_port, O(23) => OTMP_8_23_port, O(22) => 
                           OTMP_8_22_port, O(21) => OTMP_8_21_port, O(20) => 
                           OTMP_8_20_port, O(19) => OTMP_8_19_port, O(18) => 
                           OTMP_8_18_port, O(17) => OTMP_8_17_port, O(16) => 
                           OTMP_8_16_port, O(15) => OTMP_8_15_port, O(14) => 
                           OTMP_8_14_port, O(13) => OTMP_8_13_port, O(12) => 
                           OTMP_8_12_port, O(11) => OTMP_8_11_port, O(10) => 
                           OTMP_8_10_port, O(9) => OTMP_8_9_port, O(8) => 
                           OTMP_8_8_port, O(7) => OTMP_8_7_port, O(6) => 
                           OTMP_8_6_port, O(5) => OTMP_8_5_port, O(4) => 
                           OTMP_8_4_port, O(3) => OTMP_8_3_port, O(2) => 
                           OTMP_8_2_port, O(1) => OTMP_8_1_port, O(0) => n_1117
                           , A_so(49) => SHIFT_9_49_port, A_so(48) => 
                           SHIFT_9_48_port, A_so(47) => SHIFT_9_47_port, 
                           A_so(46) => SHIFT_9_46_port, A_so(45) => 
                           SHIFT_9_45_port, A_so(44) => SHIFT_9_44_port, 
                           A_so(43) => SHIFT_9_43_port, A_so(42) => 
                           SHIFT_9_42_port, A_so(41) => SHIFT_9_41_port, 
                           A_so(40) => SHIFT_9_40_port, A_so(39) => 
                           SHIFT_9_39_port, A_so(38) => SHIFT_9_38_port, 
                           A_so(37) => SHIFT_9_37_port, A_so(36) => 
                           SHIFT_9_36_port, A_so(35) => SHIFT_9_35_port, 
                           A_so(34) => SHIFT_9_34_port, A_so(33) => 
                           SHIFT_9_33_port, A_so(32) => SHIFT_9_32_port, 
                           A_so(31) => SHIFT_9_31_port, A_so(30) => 
                           SHIFT_9_30_port, A_so(29) => SHIFT_9_29_port, 
                           A_so(28) => SHIFT_9_28_port, A_so(27) => 
                           SHIFT_9_27_port, A_so(26) => SHIFT_9_26_port, 
                           A_so(25) => SHIFT_9_25_port, A_so(24) => 
                           SHIFT_9_24_port, A_so(23) => SHIFT_9_23_port, 
                           A_so(22) => SHIFT_9_22_port, A_so(21) => 
                           SHIFT_9_21_port, A_so(20) => SHIFT_9_20_port, 
                           A_so(19) => SHIFT_9_19_port, A_so(18) => 
                           SHIFT_9_18_port, A_so(17) => SHIFT_9_17_port, 
                           A_so(16) => SHIFT_9_16_port, A_so(15) => 
                           SHIFT_9_15_port, A_so(14) => SHIFT_9_14_port, 
                           A_so(13) => SHIFT_9_13_port, A_so(12) => 
                           SHIFT_9_12_port, A_so(11) => SHIFT_9_11_port, 
                           A_so(10) => SHIFT_9_10_port, A_so(9) => 
                           SHIFT_9_9_port, A_so(8) => SHIFT_9_8_port, A_so(7) 
                           => SHIFT_9_7_port, A_so(6) => SHIFT_9_6_port, 
                           A_so(5) => SHIFT_9_5_port, A_so(4) => SHIFT_9_4_port
                           , A_so(3) => SHIFT_9_3_port, A_so(2) => 
                           SHIFT_9_2_port, A_so(1) => n_1118, A_so(0) => n_1119
                           , A_nso(49) => SHIFT_n_9_49_port, A_nso(48) => 
                           SHIFT_n_9_48_port, A_nso(47) => SHIFT_n_9_47_port, 
                           A_nso(46) => SHIFT_n_9_46_port, A_nso(45) => 
                           SHIFT_n_9_45_port, A_nso(44) => SHIFT_n_9_44_port, 
                           A_nso(43) => SHIFT_n_9_43_port, A_nso(42) => 
                           SHIFT_n_9_42_port, A_nso(41) => SHIFT_n_9_41_port, 
                           A_nso(40) => SHIFT_n_9_40_port, A_nso(39) => 
                           SHIFT_n_9_39_port, A_nso(38) => SHIFT_n_9_38_port, 
                           A_nso(37) => SHIFT_n_9_37_port, A_nso(36) => 
                           SHIFT_n_9_36_port, A_nso(35) => SHIFT_n_9_35_port, 
                           A_nso(34) => SHIFT_n_9_34_port, A_nso(33) => 
                           SHIFT_n_9_33_port, A_nso(32) => SHIFT_n_9_32_port, 
                           A_nso(31) => SHIFT_n_9_31_port, A_nso(30) => 
                           SHIFT_n_9_30_port, A_nso(29) => SHIFT_n_9_29_port, 
                           A_nso(28) => SHIFT_n_9_28_port, A_nso(27) => 
                           SHIFT_n_9_27_port, A_nso(26) => SHIFT_n_9_26_port, 
                           A_nso(25) => SHIFT_n_9_25_port, A_nso(24) => 
                           SHIFT_n_9_24_port, A_nso(23) => SHIFT_n_9_23_port, 
                           A_nso(22) => SHIFT_n_9_22_port, A_nso(21) => 
                           SHIFT_n_9_21_port, A_nso(20) => SHIFT_n_9_20_port, 
                           A_nso(19) => SHIFT_n_9_19_port, A_nso(18) => 
                           SHIFT_n_9_18_port, A_nso(17) => SHIFT_n_9_17_port, 
                           A_nso(16) => SHIFT_n_9_16_port, A_nso(15) => 
                           SHIFT_n_9_15_port, A_nso(14) => SHIFT_n_9_14_port, 
                           A_nso(13) => SHIFT_n_9_13_port, A_nso(12) => 
                           SHIFT_n_9_12_port, A_nso(11) => SHIFT_n_9_11_port, 
                           A_nso(10) => SHIFT_n_9_10_port, A_nso(9) => 
                           SHIFT_n_9_9_port, A_nso(8) => SHIFT_n_9_8_port, 
                           A_nso(7) => SHIFT_n_9_7_port, A_nso(6) => 
                           SHIFT_n_9_6_port, A_nso(5) => SHIFT_n_9_5_port, 
                           A_nso(4) => SHIFT_n_9_4_port, A_nso(3) => 
                           SHIFT_n_9_3_port, A_nso(2) => SHIFT_n_9_2_port, 
                           A_nso(1) => n_1120, A_nso(0) => n_1121);
   ENC_9 : BOOTHENC_NBIT52_i18 port map( A_s(51) => SHIFT_9_49_port, A_s(50) =>
                           SHIFT_9_49_port, A_s(49) => SHIFT_9_49_port, A_s(48)
                           => SHIFT_9_48_port, A_s(47) => SHIFT_9_47_port, 
                           A_s(46) => SHIFT_9_46_port, A_s(45) => 
                           SHIFT_9_45_port, A_s(44) => SHIFT_9_44_port, A_s(43)
                           => SHIFT_9_43_port, A_s(42) => SHIFT_9_42_port, 
                           A_s(41) => SHIFT_9_41_port, A_s(40) => 
                           SHIFT_9_40_port, A_s(39) => SHIFT_9_39_port, A_s(38)
                           => SHIFT_9_38_port, A_s(37) => SHIFT_9_37_port, 
                           A_s(36) => SHIFT_9_36_port, A_s(35) => 
                           SHIFT_9_35_port, A_s(34) => SHIFT_9_34_port, A_s(33)
                           => SHIFT_9_33_port, A_s(32) => SHIFT_9_32_port, 
                           A_s(31) => SHIFT_9_31_port, A_s(30) => 
                           SHIFT_9_30_port, A_s(29) => SHIFT_9_29_port, A_s(28)
                           => SHIFT_9_28_port, A_s(27) => SHIFT_9_27_port, 
                           A_s(26) => SHIFT_9_26_port, A_s(25) => 
                           SHIFT_9_25_port, A_s(24) => SHIFT_9_24_port, A_s(23)
                           => SHIFT_9_23_port, A_s(22) => SHIFT_9_22_port, 
                           A_s(21) => SHIFT_9_21_port, A_s(20) => 
                           SHIFT_9_20_port, A_s(19) => SHIFT_9_19_port, A_s(18)
                           => SHIFT_9_18_port, A_s(17) => SHIFT_9_17_port, 
                           A_s(16) => SHIFT_9_16_port, A_s(15) => 
                           SHIFT_9_15_port, A_s(14) => SHIFT_9_14_port, A_s(13)
                           => SHIFT_9_13_port, A_s(12) => SHIFT_9_12_port, 
                           A_s(11) => SHIFT_9_11_port, A_s(10) => 
                           SHIFT_9_10_port, A_s(9) => SHIFT_9_9_port, A_s(8) =>
                           SHIFT_9_8_port, A_s(7) => SHIFT_9_7_port, A_s(6) => 
                           SHIFT_9_6_port, A_s(5) => SHIFT_9_5_port, A_s(4) => 
                           SHIFT_9_4_port, A_s(3) => SHIFT_9_3_port, A_s(2) => 
                           SHIFT_9_2_port, A_s(1) => SHIFT_9_1_port, A_s(0) => 
                           SHIFT_9_0_port, A_ns(51) => SHIFT_n_9_49_port, 
                           A_ns(50) => SHIFT_n_9_49_port, A_ns(49) => 
                           SHIFT_n_9_49_port, A_ns(48) => SHIFT_n_9_48_port, 
                           A_ns(47) => SHIFT_n_9_47_port, A_ns(46) => 
                           SHIFT_n_9_46_port, A_ns(45) => SHIFT_n_9_45_port, 
                           A_ns(44) => SHIFT_n_9_44_port, A_ns(43) => 
                           SHIFT_n_9_43_port, A_ns(42) => SHIFT_n_9_42_port, 
                           A_ns(41) => SHIFT_n_9_41_port, A_ns(40) => 
                           SHIFT_n_9_40_port, A_ns(39) => SHIFT_n_9_39_port, 
                           A_ns(38) => SHIFT_n_9_38_port, A_ns(37) => 
                           SHIFT_n_9_37_port, A_ns(36) => SHIFT_n_9_36_port, 
                           A_ns(35) => SHIFT_n_9_35_port, A_ns(34) => 
                           SHIFT_n_9_34_port, A_ns(33) => SHIFT_n_9_33_port, 
                           A_ns(32) => SHIFT_n_9_32_port, A_ns(31) => 
                           SHIFT_n_9_31_port, A_ns(30) => SHIFT_n_9_30_port, 
                           A_ns(29) => SHIFT_n_9_29_port, A_ns(28) => 
                           SHIFT_n_9_28_port, A_ns(27) => SHIFT_n_9_27_port, 
                           A_ns(26) => SHIFT_n_9_26_port, A_ns(25) => 
                           SHIFT_n_9_25_port, A_ns(24) => SHIFT_n_9_24_port, 
                           A_ns(23) => SHIFT_n_9_23_port, A_ns(22) => 
                           SHIFT_n_9_22_port, A_ns(21) => SHIFT_n_9_21_port, 
                           A_ns(20) => SHIFT_n_9_20_port, A_ns(19) => 
                           SHIFT_n_9_19_port, A_ns(18) => SHIFT_n_9_18_port, 
                           A_ns(17) => SHIFT_n_9_17_port, A_ns(16) => 
                           SHIFT_n_9_16_port, A_ns(15) => SHIFT_n_9_15_port, 
                           A_ns(14) => SHIFT_n_9_14_port, A_ns(13) => 
                           SHIFT_n_9_13_port, A_ns(12) => SHIFT_n_9_12_port, 
                           A_ns(11) => SHIFT_n_9_11_port, A_ns(10) => 
                           SHIFT_n_9_10_port, A_ns(9) => SHIFT_n_9_9_port, 
                           A_ns(8) => SHIFT_n_9_8_port, A_ns(7) => 
                           SHIFT_n_9_7_port, A_ns(6) => SHIFT_n_9_6_port, 
                           A_ns(5) => SHIFT_n_9_5_port, A_ns(4) => 
                           SHIFT_n_9_4_port, A_ns(3) => SHIFT_n_9_3_port, 
                           A_ns(2) => SHIFT_n_9_2_port, A_ns(1) => 
                           SHIFT_n_9_1_port, A_ns(0) => SHIFT_n_9_0_port, B(51)
                           => B(31), B(50) => B(31), B(49) => B(31), B(48) => 
                           B(31), B(47) => B(31), B(46) => B(31), B(45) => 
                           B(31), B(44) => B(31), B(43) => B(31), B(42) => 
                           B(31), B(41) => B(31), B(40) => B(31), B(39) => 
                           B(31), B(38) => B(31), B(37) => B(31), B(36) => 
                           B(31), B(35) => B(31), B(34) => B(31), B(33) => 
                           B(31), B(32) => B(31), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), O(51) => OTMP_9_51_port, 
                           O(50) => OTMP_9_50_port, O(49) => OTMP_9_49_port, 
                           O(48) => OTMP_9_48_port, O(47) => OTMP_9_47_port, 
                           O(46) => OTMP_9_46_port, O(45) => OTMP_9_45_port, 
                           O(44) => OTMP_9_44_port, O(43) => OTMP_9_43_port, 
                           O(42) => OTMP_9_42_port, O(41) => OTMP_9_41_port, 
                           O(40) => OTMP_9_40_port, O(39) => OTMP_9_39_port, 
                           O(38) => OTMP_9_38_port, O(37) => OTMP_9_37_port, 
                           O(36) => OTMP_9_36_port, O(35) => OTMP_9_35_port, 
                           O(34) => OTMP_9_34_port, O(33) => OTMP_9_33_port, 
                           O(32) => OTMP_9_32_port, O(31) => OTMP_9_31_port, 
                           O(30) => OTMP_9_30_port, O(29) => OTMP_9_29_port, 
                           O(28) => OTMP_9_28_port, O(27) => OTMP_9_27_port, 
                           O(26) => OTMP_9_26_port, O(25) => OTMP_9_25_port, 
                           O(24) => OTMP_9_24_port, O(23) => OTMP_9_23_port, 
                           O(22) => OTMP_9_22_port, O(21) => OTMP_9_21_port, 
                           O(20) => OTMP_9_20_port, O(19) => OTMP_9_19_port, 
                           O(18) => OTMP_9_18_port, O(17) => OTMP_9_17_port, 
                           O(16) => OTMP_9_16_port, O(15) => OTMP_9_15_port, 
                           O(14) => OTMP_9_14_port, O(13) => OTMP_9_13_port, 
                           O(12) => OTMP_9_12_port, O(11) => OTMP_9_11_port, 
                           O(10) => OTMP_9_10_port, O(9) => OTMP_9_9_port, O(8)
                           => OTMP_9_8_port, O(7) => OTMP_9_7_port, O(6) => 
                           OTMP_9_6_port, O(5) => OTMP_9_5_port, O(4) => 
                           OTMP_9_4_port, O(3) => OTMP_9_3_port, O(2) => 
                           OTMP_9_2_port, O(1) => OTMP_9_1_port, O(0) => n_1122
                           , A_so(51) => SHIFT_10_51_port, A_so(50) => 
                           SHIFT_10_50_port, A_so(49) => SHIFT_10_49_port, 
                           A_so(48) => SHIFT_10_48_port, A_so(47) => 
                           SHIFT_10_47_port, A_so(46) => SHIFT_10_46_port, 
                           A_so(45) => SHIFT_10_45_port, A_so(44) => 
                           SHIFT_10_44_port, A_so(43) => SHIFT_10_43_port, 
                           A_so(42) => SHIFT_10_42_port, A_so(41) => 
                           SHIFT_10_41_port, A_so(40) => SHIFT_10_40_port, 
                           A_so(39) => SHIFT_10_39_port, A_so(38) => 
                           SHIFT_10_38_port, A_so(37) => SHIFT_10_37_port, 
                           A_so(36) => SHIFT_10_36_port, A_so(35) => 
                           SHIFT_10_35_port, A_so(34) => SHIFT_10_34_port, 
                           A_so(33) => SHIFT_10_33_port, A_so(32) => 
                           SHIFT_10_32_port, A_so(31) => SHIFT_10_31_port, 
                           A_so(30) => SHIFT_10_30_port, A_so(29) => 
                           SHIFT_10_29_port, A_so(28) => SHIFT_10_28_port, 
                           A_so(27) => SHIFT_10_27_port, A_so(26) => 
                           SHIFT_10_26_port, A_so(25) => SHIFT_10_25_port, 
                           A_so(24) => SHIFT_10_24_port, A_so(23) => 
                           SHIFT_10_23_port, A_so(22) => SHIFT_10_22_port, 
                           A_so(21) => SHIFT_10_21_port, A_so(20) => 
                           SHIFT_10_20_port, A_so(19) => SHIFT_10_19_port, 
                           A_so(18) => SHIFT_10_18_port, A_so(17) => 
                           SHIFT_10_17_port, A_so(16) => SHIFT_10_16_port, 
                           A_so(15) => SHIFT_10_15_port, A_so(14) => 
                           SHIFT_10_14_port, A_so(13) => SHIFT_10_13_port, 
                           A_so(12) => SHIFT_10_12_port, A_so(11) => 
                           SHIFT_10_11_port, A_so(10) => SHIFT_10_10_port, 
                           A_so(9) => SHIFT_10_9_port, A_so(8) => 
                           SHIFT_10_8_port, A_so(7) => SHIFT_10_7_port, A_so(6)
                           => SHIFT_10_6_port, A_so(5) => SHIFT_10_5_port, 
                           A_so(4) => SHIFT_10_4_port, A_so(3) => 
                           SHIFT_10_3_port, A_so(2) => SHIFT_10_2_port, A_so(1)
                           => n_1123, A_so(0) => n_1124, A_nso(51) => 
                           SHIFT_n_10_51_port, A_nso(50) => SHIFT_n_10_50_port,
                           A_nso(49) => SHIFT_n_10_49_port, A_nso(48) => 
                           SHIFT_n_10_48_port, A_nso(47) => SHIFT_n_10_47_port,
                           A_nso(46) => SHIFT_n_10_46_port, A_nso(45) => 
                           SHIFT_n_10_45_port, A_nso(44) => SHIFT_n_10_44_port,
                           A_nso(43) => SHIFT_n_10_43_port, A_nso(42) => 
                           SHIFT_n_10_42_port, A_nso(41) => SHIFT_n_10_41_port,
                           A_nso(40) => SHIFT_n_10_40_port, A_nso(39) => 
                           SHIFT_n_10_39_port, A_nso(38) => SHIFT_n_10_38_port,
                           A_nso(37) => SHIFT_n_10_37_port, A_nso(36) => 
                           SHIFT_n_10_36_port, A_nso(35) => SHIFT_n_10_35_port,
                           A_nso(34) => SHIFT_n_10_34_port, A_nso(33) => 
                           SHIFT_n_10_33_port, A_nso(32) => SHIFT_n_10_32_port,
                           A_nso(31) => SHIFT_n_10_31_port, A_nso(30) => 
                           SHIFT_n_10_30_port, A_nso(29) => SHIFT_n_10_29_port,
                           A_nso(28) => SHIFT_n_10_28_port, A_nso(27) => 
                           SHIFT_n_10_27_port, A_nso(26) => SHIFT_n_10_26_port,
                           A_nso(25) => SHIFT_n_10_25_port, A_nso(24) => 
                           SHIFT_n_10_24_port, A_nso(23) => SHIFT_n_10_23_port,
                           A_nso(22) => SHIFT_n_10_22_port, A_nso(21) => 
                           SHIFT_n_10_21_port, A_nso(20) => SHIFT_n_10_20_port,
                           A_nso(19) => SHIFT_n_10_19_port, A_nso(18) => 
                           SHIFT_n_10_18_port, A_nso(17) => SHIFT_n_10_17_port,
                           A_nso(16) => SHIFT_n_10_16_port, A_nso(15) => 
                           SHIFT_n_10_15_port, A_nso(14) => SHIFT_n_10_14_port,
                           A_nso(13) => SHIFT_n_10_13_port, A_nso(12) => 
                           SHIFT_n_10_12_port, A_nso(11) => SHIFT_n_10_11_port,
                           A_nso(10) => SHIFT_n_10_10_port, A_nso(9) => 
                           SHIFT_n_10_9_port, A_nso(8) => SHIFT_n_10_8_port, 
                           A_nso(7) => SHIFT_n_10_7_port, A_nso(6) => 
                           SHIFT_n_10_6_port, A_nso(5) => SHIFT_n_10_5_port, 
                           A_nso(4) => SHIFT_n_10_4_port, A_nso(3) => 
                           SHIFT_n_10_3_port, A_nso(2) => SHIFT_n_10_2_port, 
                           A_nso(1) => n_1125, A_nso(0) => n_1126);
   ENC_10 : BOOTHENC_NBIT54_i20 port map( A_s(53) => SHIFT_10_51_port, A_s(52) 
                           => SHIFT_10_51_port, A_s(51) => SHIFT_10_51_port, 
                           A_s(50) => SHIFT_10_50_port, A_s(49) => 
                           SHIFT_10_49_port, A_s(48) => SHIFT_10_48_port, 
                           A_s(47) => SHIFT_10_47_port, A_s(46) => 
                           SHIFT_10_46_port, A_s(45) => SHIFT_10_45_port, 
                           A_s(44) => SHIFT_10_44_port, A_s(43) => 
                           SHIFT_10_43_port, A_s(42) => SHIFT_10_42_port, 
                           A_s(41) => SHIFT_10_41_port, A_s(40) => 
                           SHIFT_10_40_port, A_s(39) => SHIFT_10_39_port, 
                           A_s(38) => SHIFT_10_38_port, A_s(37) => 
                           SHIFT_10_37_port, A_s(36) => SHIFT_10_36_port, 
                           A_s(35) => SHIFT_10_35_port, A_s(34) => 
                           SHIFT_10_34_port, A_s(33) => SHIFT_10_33_port, 
                           A_s(32) => SHIFT_10_32_port, A_s(31) => 
                           SHIFT_10_31_port, A_s(30) => SHIFT_10_30_port, 
                           A_s(29) => SHIFT_10_29_port, A_s(28) => 
                           SHIFT_10_28_port, A_s(27) => SHIFT_10_27_port, 
                           A_s(26) => SHIFT_10_26_port, A_s(25) => 
                           SHIFT_10_25_port, A_s(24) => SHIFT_10_24_port, 
                           A_s(23) => SHIFT_10_23_port, A_s(22) => 
                           SHIFT_10_22_port, A_s(21) => SHIFT_10_21_port, 
                           A_s(20) => SHIFT_10_20_port, A_s(19) => 
                           SHIFT_10_19_port, A_s(18) => SHIFT_10_18_port, 
                           A_s(17) => SHIFT_10_17_port, A_s(16) => 
                           SHIFT_10_16_port, A_s(15) => SHIFT_10_15_port, 
                           A_s(14) => SHIFT_10_14_port, A_s(13) => 
                           SHIFT_10_13_port, A_s(12) => SHIFT_10_12_port, 
                           A_s(11) => SHIFT_10_11_port, A_s(10) => 
                           SHIFT_10_10_port, A_s(9) => SHIFT_10_9_port, A_s(8) 
                           => SHIFT_10_8_port, A_s(7) => SHIFT_10_7_port, 
                           A_s(6) => SHIFT_10_6_port, A_s(5) => SHIFT_10_5_port
                           , A_s(4) => SHIFT_10_4_port, A_s(3) => 
                           SHIFT_10_3_port, A_s(2) => SHIFT_10_2_port, A_s(1) 
                           => SHIFT_10_1_port, A_s(0) => SHIFT_10_0_port, 
                           A_ns(53) => SHIFT_n_10_51_port, A_ns(52) => 
                           SHIFT_n_10_51_port, A_ns(51) => SHIFT_n_10_51_port, 
                           A_ns(50) => SHIFT_n_10_50_port, A_ns(49) => 
                           SHIFT_n_10_49_port, A_ns(48) => SHIFT_n_10_48_port, 
                           A_ns(47) => SHIFT_n_10_47_port, A_ns(46) => 
                           SHIFT_n_10_46_port, A_ns(45) => SHIFT_n_10_45_port, 
                           A_ns(44) => SHIFT_n_10_44_port, A_ns(43) => 
                           SHIFT_n_10_43_port, A_ns(42) => SHIFT_n_10_42_port, 
                           A_ns(41) => SHIFT_n_10_41_port, A_ns(40) => 
                           SHIFT_n_10_40_port, A_ns(39) => SHIFT_n_10_39_port, 
                           A_ns(38) => SHIFT_n_10_38_port, A_ns(37) => 
                           SHIFT_n_10_37_port, A_ns(36) => SHIFT_n_10_36_port, 
                           A_ns(35) => SHIFT_n_10_35_port, A_ns(34) => 
                           SHIFT_n_10_34_port, A_ns(33) => SHIFT_n_10_33_port, 
                           A_ns(32) => SHIFT_n_10_32_port, A_ns(31) => 
                           SHIFT_n_10_31_port, A_ns(30) => SHIFT_n_10_30_port, 
                           A_ns(29) => SHIFT_n_10_29_port, A_ns(28) => 
                           SHIFT_n_10_28_port, A_ns(27) => SHIFT_n_10_27_port, 
                           A_ns(26) => SHIFT_n_10_26_port, A_ns(25) => 
                           SHIFT_n_10_25_port, A_ns(24) => SHIFT_n_10_24_port, 
                           A_ns(23) => SHIFT_n_10_23_port, A_ns(22) => 
                           SHIFT_n_10_22_port, A_ns(21) => SHIFT_n_10_21_port, 
                           A_ns(20) => SHIFT_n_10_20_port, A_ns(19) => 
                           SHIFT_n_10_19_port, A_ns(18) => SHIFT_n_10_18_port, 
                           A_ns(17) => SHIFT_n_10_17_port, A_ns(16) => 
                           SHIFT_n_10_16_port, A_ns(15) => SHIFT_n_10_15_port, 
                           A_ns(14) => SHIFT_n_10_14_port, A_ns(13) => 
                           SHIFT_n_10_13_port, A_ns(12) => SHIFT_n_10_12_port, 
                           A_ns(11) => SHIFT_n_10_11_port, A_ns(10) => 
                           SHIFT_n_10_10_port, A_ns(9) => SHIFT_n_10_9_port, 
                           A_ns(8) => SHIFT_n_10_8_port, A_ns(7) => 
                           SHIFT_n_10_7_port, A_ns(6) => SHIFT_n_10_6_port, 
                           A_ns(5) => SHIFT_n_10_5_port, A_ns(4) => 
                           SHIFT_n_10_4_port, A_ns(3) => SHIFT_n_10_3_port, 
                           A_ns(2) => SHIFT_n_10_2_port, A_ns(1) => 
                           SHIFT_n_10_1_port, A_ns(0) => SHIFT_n_10_0_port, 
                           B(53) => B(31), B(52) => B(31), B(51) => B(31), 
                           B(50) => B(31), B(49) => B(31), B(48) => B(31), 
                           B(47) => B(31), B(46) => B(31), B(45) => B(31), 
                           B(44) => B(31), B(43) => B(31), B(42) => B(31), 
                           B(41) => B(31), B(40) => B(31), B(39) => B(31), 
                           B(38) => B(31), B(37) => B(31), B(36) => B(31), 
                           B(35) => B(31), B(34) => B(31), B(33) => B(31), 
                           B(32) => B(31), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), O(53) => OTMP_10_53_port, O(52) 
                           => OTMP_10_52_port, O(51) => OTMP_10_51_port, O(50) 
                           => OTMP_10_50_port, O(49) => OTMP_10_49_port, O(48) 
                           => OTMP_10_48_port, O(47) => OTMP_10_47_port, O(46) 
                           => OTMP_10_46_port, O(45) => OTMP_10_45_port, O(44) 
                           => OTMP_10_44_port, O(43) => OTMP_10_43_port, O(42) 
                           => OTMP_10_42_port, O(41) => OTMP_10_41_port, O(40) 
                           => OTMP_10_40_port, O(39) => OTMP_10_39_port, O(38) 
                           => OTMP_10_38_port, O(37) => OTMP_10_37_port, O(36) 
                           => OTMP_10_36_port, O(35) => OTMP_10_35_port, O(34) 
                           => OTMP_10_34_port, O(33) => OTMP_10_33_port, O(32) 
                           => OTMP_10_32_port, O(31) => OTMP_10_31_port, O(30) 
                           => OTMP_10_30_port, O(29) => OTMP_10_29_port, O(28) 
                           => OTMP_10_28_port, O(27) => OTMP_10_27_port, O(26) 
                           => OTMP_10_26_port, O(25) => OTMP_10_25_port, O(24) 
                           => OTMP_10_24_port, O(23) => OTMP_10_23_port, O(22) 
                           => OTMP_10_22_port, O(21) => OTMP_10_21_port, O(20) 
                           => OTMP_10_20_port, O(19) => OTMP_10_19_port, O(18) 
                           => OTMP_10_18_port, O(17) => OTMP_10_17_port, O(16) 
                           => OTMP_10_16_port, O(15) => OTMP_10_15_port, O(14) 
                           => OTMP_10_14_port, O(13) => OTMP_10_13_port, O(12) 
                           => OTMP_10_12_port, O(11) => OTMP_10_11_port, O(10) 
                           => OTMP_10_10_port, O(9) => OTMP_10_9_port, O(8) => 
                           OTMP_10_8_port, O(7) => OTMP_10_7_port, O(6) => 
                           OTMP_10_6_port, O(5) => OTMP_10_5_port, O(4) => 
                           OTMP_10_4_port, O(3) => OTMP_10_3_port, O(2) => 
                           OTMP_10_2_port, O(1) => OTMP_10_1_port, O(0) => 
                           n_1127, A_so(53) => SHIFT_11_53_port, A_so(52) => 
                           SHIFT_11_52_port, A_so(51) => SHIFT_11_51_port, 
                           A_so(50) => SHIFT_11_50_port, A_so(49) => 
                           SHIFT_11_49_port, A_so(48) => SHIFT_11_48_port, 
                           A_so(47) => SHIFT_11_47_port, A_so(46) => 
                           SHIFT_11_46_port, A_so(45) => SHIFT_11_45_port, 
                           A_so(44) => SHIFT_11_44_port, A_so(43) => 
                           SHIFT_11_43_port, A_so(42) => SHIFT_11_42_port, 
                           A_so(41) => SHIFT_11_41_port, A_so(40) => 
                           SHIFT_11_40_port, A_so(39) => SHIFT_11_39_port, 
                           A_so(38) => SHIFT_11_38_port, A_so(37) => 
                           SHIFT_11_37_port, A_so(36) => SHIFT_11_36_port, 
                           A_so(35) => SHIFT_11_35_port, A_so(34) => 
                           SHIFT_11_34_port, A_so(33) => SHIFT_11_33_port, 
                           A_so(32) => SHIFT_11_32_port, A_so(31) => 
                           SHIFT_11_31_port, A_so(30) => SHIFT_11_30_port, 
                           A_so(29) => SHIFT_11_29_port, A_so(28) => 
                           SHIFT_11_28_port, A_so(27) => SHIFT_11_27_port, 
                           A_so(26) => SHIFT_11_26_port, A_so(25) => 
                           SHIFT_11_25_port, A_so(24) => SHIFT_11_24_port, 
                           A_so(23) => SHIFT_11_23_port, A_so(22) => 
                           SHIFT_11_22_port, A_so(21) => SHIFT_11_21_port, 
                           A_so(20) => SHIFT_11_20_port, A_so(19) => 
                           SHIFT_11_19_port, A_so(18) => SHIFT_11_18_port, 
                           A_so(17) => SHIFT_11_17_port, A_so(16) => 
                           SHIFT_11_16_port, A_so(15) => SHIFT_11_15_port, 
                           A_so(14) => SHIFT_11_14_port, A_so(13) => 
                           SHIFT_11_13_port, A_so(12) => SHIFT_11_12_port, 
                           A_so(11) => SHIFT_11_11_port, A_so(10) => 
                           SHIFT_11_10_port, A_so(9) => SHIFT_11_9_port, 
                           A_so(8) => SHIFT_11_8_port, A_so(7) => 
                           SHIFT_11_7_port, A_so(6) => SHIFT_11_6_port, A_so(5)
                           => SHIFT_11_5_port, A_so(4) => SHIFT_11_4_port, 
                           A_so(3) => SHIFT_11_3_port, A_so(2) => 
                           SHIFT_11_2_port, A_so(1) => n_1128, A_so(0) => 
                           n_1129, A_nso(53) => SHIFT_n_11_53_port, A_nso(52) 
                           => SHIFT_n_11_52_port, A_nso(51) => 
                           SHIFT_n_11_51_port, A_nso(50) => SHIFT_n_11_50_port,
                           A_nso(49) => SHIFT_n_11_49_port, A_nso(48) => 
                           SHIFT_n_11_48_port, A_nso(47) => SHIFT_n_11_47_port,
                           A_nso(46) => SHIFT_n_11_46_port, A_nso(45) => 
                           SHIFT_n_11_45_port, A_nso(44) => SHIFT_n_11_44_port,
                           A_nso(43) => SHIFT_n_11_43_port, A_nso(42) => 
                           SHIFT_n_11_42_port, A_nso(41) => SHIFT_n_11_41_port,
                           A_nso(40) => SHIFT_n_11_40_port, A_nso(39) => 
                           SHIFT_n_11_39_port, A_nso(38) => SHIFT_n_11_38_port,
                           A_nso(37) => SHIFT_n_11_37_port, A_nso(36) => 
                           SHIFT_n_11_36_port, A_nso(35) => SHIFT_n_11_35_port,
                           A_nso(34) => SHIFT_n_11_34_port, A_nso(33) => 
                           SHIFT_n_11_33_port, A_nso(32) => SHIFT_n_11_32_port,
                           A_nso(31) => SHIFT_n_11_31_port, A_nso(30) => 
                           SHIFT_n_11_30_port, A_nso(29) => SHIFT_n_11_29_port,
                           A_nso(28) => SHIFT_n_11_28_port, A_nso(27) => 
                           SHIFT_n_11_27_port, A_nso(26) => SHIFT_n_11_26_port,
                           A_nso(25) => SHIFT_n_11_25_port, A_nso(24) => 
                           SHIFT_n_11_24_port, A_nso(23) => SHIFT_n_11_23_port,
                           A_nso(22) => SHIFT_n_11_22_port, A_nso(21) => 
                           SHIFT_n_11_21_port, A_nso(20) => SHIFT_n_11_20_port,
                           A_nso(19) => SHIFT_n_11_19_port, A_nso(18) => 
                           SHIFT_n_11_18_port, A_nso(17) => SHIFT_n_11_17_port,
                           A_nso(16) => SHIFT_n_11_16_port, A_nso(15) => 
                           SHIFT_n_11_15_port, A_nso(14) => SHIFT_n_11_14_port,
                           A_nso(13) => SHIFT_n_11_13_port, A_nso(12) => 
                           SHIFT_n_11_12_port, A_nso(11) => SHIFT_n_11_11_port,
                           A_nso(10) => SHIFT_n_11_10_port, A_nso(9) => 
                           SHIFT_n_11_9_port, A_nso(8) => SHIFT_n_11_8_port, 
                           A_nso(7) => SHIFT_n_11_7_port, A_nso(6) => 
                           SHIFT_n_11_6_port, A_nso(5) => SHIFT_n_11_5_port, 
                           A_nso(4) => SHIFT_n_11_4_port, A_nso(3) => 
                           SHIFT_n_11_3_port, A_nso(2) => SHIFT_n_11_2_port, 
                           A_nso(1) => n_1130, A_nso(0) => n_1131);
   ENC_11 : BOOTHENC_NBIT56_i22 port map( A_s(55) => SHIFT_11_53_port, A_s(54) 
                           => SHIFT_11_53_port, A_s(53) => SHIFT_11_53_port, 
                           A_s(52) => SHIFT_11_52_port, A_s(51) => 
                           SHIFT_11_51_port, A_s(50) => SHIFT_11_50_port, 
                           A_s(49) => SHIFT_11_49_port, A_s(48) => 
                           SHIFT_11_48_port, A_s(47) => SHIFT_11_47_port, 
                           A_s(46) => SHIFT_11_46_port, A_s(45) => 
                           SHIFT_11_45_port, A_s(44) => SHIFT_11_44_port, 
                           A_s(43) => SHIFT_11_43_port, A_s(42) => 
                           SHIFT_11_42_port, A_s(41) => SHIFT_11_41_port, 
                           A_s(40) => SHIFT_11_40_port, A_s(39) => 
                           SHIFT_11_39_port, A_s(38) => SHIFT_11_38_port, 
                           A_s(37) => SHIFT_11_37_port, A_s(36) => 
                           SHIFT_11_36_port, A_s(35) => SHIFT_11_35_port, 
                           A_s(34) => SHIFT_11_34_port, A_s(33) => 
                           SHIFT_11_33_port, A_s(32) => SHIFT_11_32_port, 
                           A_s(31) => SHIFT_11_31_port, A_s(30) => 
                           SHIFT_11_30_port, A_s(29) => SHIFT_11_29_port, 
                           A_s(28) => SHIFT_11_28_port, A_s(27) => 
                           SHIFT_11_27_port, A_s(26) => SHIFT_11_26_port, 
                           A_s(25) => SHIFT_11_25_port, A_s(24) => 
                           SHIFT_11_24_port, A_s(23) => SHIFT_11_23_port, 
                           A_s(22) => SHIFT_11_22_port, A_s(21) => 
                           SHIFT_11_21_port, A_s(20) => SHIFT_11_20_port, 
                           A_s(19) => SHIFT_11_19_port, A_s(18) => 
                           SHIFT_11_18_port, A_s(17) => SHIFT_11_17_port, 
                           A_s(16) => SHIFT_11_16_port, A_s(15) => 
                           SHIFT_11_15_port, A_s(14) => SHIFT_11_14_port, 
                           A_s(13) => SHIFT_11_13_port, A_s(12) => 
                           SHIFT_11_12_port, A_s(11) => SHIFT_11_11_port, 
                           A_s(10) => SHIFT_11_10_port, A_s(9) => 
                           SHIFT_11_9_port, A_s(8) => SHIFT_11_8_port, A_s(7) 
                           => SHIFT_11_7_port, A_s(6) => SHIFT_11_6_port, 
                           A_s(5) => SHIFT_11_5_port, A_s(4) => SHIFT_11_4_port
                           , A_s(3) => SHIFT_11_3_port, A_s(2) => 
                           SHIFT_11_2_port, A_s(1) => SHIFT_11_1_port, A_s(0) 
                           => SHIFT_11_0_port, A_ns(55) => SHIFT_n_11_53_port, 
                           A_ns(54) => SHIFT_n_11_53_port, A_ns(53) => 
                           SHIFT_n_11_53_port, A_ns(52) => SHIFT_n_11_52_port, 
                           A_ns(51) => SHIFT_n_11_51_port, A_ns(50) => 
                           SHIFT_n_11_50_port, A_ns(49) => SHIFT_n_11_49_port, 
                           A_ns(48) => SHIFT_n_11_48_port, A_ns(47) => 
                           SHIFT_n_11_47_port, A_ns(46) => SHIFT_n_11_46_port, 
                           A_ns(45) => SHIFT_n_11_45_port, A_ns(44) => 
                           SHIFT_n_11_44_port, A_ns(43) => SHIFT_n_11_43_port, 
                           A_ns(42) => SHIFT_n_11_42_port, A_ns(41) => 
                           SHIFT_n_11_41_port, A_ns(40) => SHIFT_n_11_40_port, 
                           A_ns(39) => SHIFT_n_11_39_port, A_ns(38) => 
                           SHIFT_n_11_38_port, A_ns(37) => SHIFT_n_11_37_port, 
                           A_ns(36) => SHIFT_n_11_36_port, A_ns(35) => 
                           SHIFT_n_11_35_port, A_ns(34) => SHIFT_n_11_34_port, 
                           A_ns(33) => SHIFT_n_11_33_port, A_ns(32) => 
                           SHIFT_n_11_32_port, A_ns(31) => SHIFT_n_11_31_port, 
                           A_ns(30) => SHIFT_n_11_30_port, A_ns(29) => 
                           SHIFT_n_11_29_port, A_ns(28) => SHIFT_n_11_28_port, 
                           A_ns(27) => SHIFT_n_11_27_port, A_ns(26) => 
                           SHIFT_n_11_26_port, A_ns(25) => SHIFT_n_11_25_port, 
                           A_ns(24) => SHIFT_n_11_24_port, A_ns(23) => 
                           SHIFT_n_11_23_port, A_ns(22) => SHIFT_n_11_22_port, 
                           A_ns(21) => SHIFT_n_11_21_port, A_ns(20) => 
                           SHIFT_n_11_20_port, A_ns(19) => SHIFT_n_11_19_port, 
                           A_ns(18) => SHIFT_n_11_18_port, A_ns(17) => 
                           SHIFT_n_11_17_port, A_ns(16) => SHIFT_n_11_16_port, 
                           A_ns(15) => SHIFT_n_11_15_port, A_ns(14) => 
                           SHIFT_n_11_14_port, A_ns(13) => SHIFT_n_11_13_port, 
                           A_ns(12) => SHIFT_n_11_12_port, A_ns(11) => 
                           SHIFT_n_11_11_port, A_ns(10) => SHIFT_n_11_10_port, 
                           A_ns(9) => SHIFT_n_11_9_port, A_ns(8) => 
                           SHIFT_n_11_8_port, A_ns(7) => SHIFT_n_11_7_port, 
                           A_ns(6) => SHIFT_n_11_6_port, A_ns(5) => 
                           SHIFT_n_11_5_port, A_ns(4) => SHIFT_n_11_4_port, 
                           A_ns(3) => SHIFT_n_11_3_port, A_ns(2) => 
                           SHIFT_n_11_2_port, A_ns(1) => SHIFT_n_11_1_port, 
                           A_ns(0) => SHIFT_n_11_0_port, B(55) => B(31), B(54) 
                           => B(31), B(53) => B(31), B(52) => B(31), B(51) => 
                           B(31), B(50) => B(31), B(49) => B(31), B(48) => 
                           B(31), B(47) => B(31), B(46) => B(31), B(45) => 
                           B(31), B(44) => B(31), B(43) => B(31), B(42) => 
                           B(31), B(41) => B(31), B(40) => B(31), B(39) => 
                           B(31), B(38) => B(31), B(37) => B(31), B(36) => 
                           B(31), B(35) => B(31), B(34) => B(31), B(33) => 
                           B(31), B(32) => B(31), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), O(55) => OTMP_11_55_port, 
                           O(54) => OTMP_11_54_port, O(53) => OTMP_11_53_port, 
                           O(52) => OTMP_11_52_port, O(51) => OTMP_11_51_port, 
                           O(50) => OTMP_11_50_port, O(49) => OTMP_11_49_port, 
                           O(48) => OTMP_11_48_port, O(47) => OTMP_11_47_port, 
                           O(46) => OTMP_11_46_port, O(45) => OTMP_11_45_port, 
                           O(44) => OTMP_11_44_port, O(43) => OTMP_11_43_port, 
                           O(42) => OTMP_11_42_port, O(41) => OTMP_11_41_port, 
                           O(40) => OTMP_11_40_port, O(39) => OTMP_11_39_port, 
                           O(38) => OTMP_11_38_port, O(37) => OTMP_11_37_port, 
                           O(36) => OTMP_11_36_port, O(35) => OTMP_11_35_port, 
                           O(34) => OTMP_11_34_port, O(33) => OTMP_11_33_port, 
                           O(32) => OTMP_11_32_port, O(31) => OTMP_11_31_port, 
                           O(30) => OTMP_11_30_port, O(29) => OTMP_11_29_port, 
                           O(28) => OTMP_11_28_port, O(27) => OTMP_11_27_port, 
                           O(26) => OTMP_11_26_port, O(25) => OTMP_11_25_port, 
                           O(24) => OTMP_11_24_port, O(23) => OTMP_11_23_port, 
                           O(22) => OTMP_11_22_port, O(21) => OTMP_11_21_port, 
                           O(20) => OTMP_11_20_port, O(19) => OTMP_11_19_port, 
                           O(18) => OTMP_11_18_port, O(17) => OTMP_11_17_port, 
                           O(16) => OTMP_11_16_port, O(15) => OTMP_11_15_port, 
                           O(14) => OTMP_11_14_port, O(13) => OTMP_11_13_port, 
                           O(12) => OTMP_11_12_port, O(11) => OTMP_11_11_port, 
                           O(10) => OTMP_11_10_port, O(9) => OTMP_11_9_port, 
                           O(8) => OTMP_11_8_port, O(7) => OTMP_11_7_port, O(6)
                           => OTMP_11_6_port, O(5) => OTMP_11_5_port, O(4) => 
                           OTMP_11_4_port, O(3) => OTMP_11_3_port, O(2) => 
                           OTMP_11_2_port, O(1) => OTMP_11_1_port, O(0) => 
                           n_1132, A_so(55) => SHIFT_12_55_port, A_so(54) => 
                           SHIFT_12_54_port, A_so(53) => SHIFT_12_53_port, 
                           A_so(52) => SHIFT_12_52_port, A_so(51) => 
                           SHIFT_12_51_port, A_so(50) => SHIFT_12_50_port, 
                           A_so(49) => SHIFT_12_49_port, A_so(48) => 
                           SHIFT_12_48_port, A_so(47) => SHIFT_12_47_port, 
                           A_so(46) => SHIFT_12_46_port, A_so(45) => 
                           SHIFT_12_45_port, A_so(44) => SHIFT_12_44_port, 
                           A_so(43) => SHIFT_12_43_port, A_so(42) => 
                           SHIFT_12_42_port, A_so(41) => SHIFT_12_41_port, 
                           A_so(40) => SHIFT_12_40_port, A_so(39) => 
                           SHIFT_12_39_port, A_so(38) => SHIFT_12_38_port, 
                           A_so(37) => SHIFT_12_37_port, A_so(36) => 
                           SHIFT_12_36_port, A_so(35) => SHIFT_12_35_port, 
                           A_so(34) => SHIFT_12_34_port, A_so(33) => 
                           SHIFT_12_33_port, A_so(32) => SHIFT_12_32_port, 
                           A_so(31) => SHIFT_12_31_port, A_so(30) => 
                           SHIFT_12_30_port, A_so(29) => SHIFT_12_29_port, 
                           A_so(28) => SHIFT_12_28_port, A_so(27) => 
                           SHIFT_12_27_port, A_so(26) => SHIFT_12_26_port, 
                           A_so(25) => SHIFT_12_25_port, A_so(24) => 
                           SHIFT_12_24_port, A_so(23) => SHIFT_12_23_port, 
                           A_so(22) => SHIFT_12_22_port, A_so(21) => 
                           SHIFT_12_21_port, A_so(20) => SHIFT_12_20_port, 
                           A_so(19) => SHIFT_12_19_port, A_so(18) => 
                           SHIFT_12_18_port, A_so(17) => SHIFT_12_17_port, 
                           A_so(16) => SHIFT_12_16_port, A_so(15) => 
                           SHIFT_12_15_port, A_so(14) => SHIFT_12_14_port, 
                           A_so(13) => SHIFT_12_13_port, A_so(12) => 
                           SHIFT_12_12_port, A_so(11) => SHIFT_12_11_port, 
                           A_so(10) => SHIFT_12_10_port, A_so(9) => 
                           SHIFT_12_9_port, A_so(8) => SHIFT_12_8_port, A_so(7)
                           => SHIFT_12_7_port, A_so(6) => SHIFT_12_6_port, 
                           A_so(5) => SHIFT_12_5_port, A_so(4) => 
                           SHIFT_12_4_port, A_so(3) => SHIFT_12_3_port, A_so(2)
                           => SHIFT_12_2_port, A_so(1) => n_1133, A_so(0) => 
                           n_1134, A_nso(55) => SHIFT_n_12_55_port, A_nso(54) 
                           => SHIFT_n_12_54_port, A_nso(53) => 
                           SHIFT_n_12_53_port, A_nso(52) => SHIFT_n_12_52_port,
                           A_nso(51) => SHIFT_n_12_51_port, A_nso(50) => 
                           SHIFT_n_12_50_port, A_nso(49) => SHIFT_n_12_49_port,
                           A_nso(48) => SHIFT_n_12_48_port, A_nso(47) => 
                           SHIFT_n_12_47_port, A_nso(46) => SHIFT_n_12_46_port,
                           A_nso(45) => SHIFT_n_12_45_port, A_nso(44) => 
                           SHIFT_n_12_44_port, A_nso(43) => SHIFT_n_12_43_port,
                           A_nso(42) => SHIFT_n_12_42_port, A_nso(41) => 
                           SHIFT_n_12_41_port, A_nso(40) => SHIFT_n_12_40_port,
                           A_nso(39) => SHIFT_n_12_39_port, A_nso(38) => 
                           SHIFT_n_12_38_port, A_nso(37) => SHIFT_n_12_37_port,
                           A_nso(36) => SHIFT_n_12_36_port, A_nso(35) => 
                           SHIFT_n_12_35_port, A_nso(34) => SHIFT_n_12_34_port,
                           A_nso(33) => SHIFT_n_12_33_port, A_nso(32) => 
                           SHIFT_n_12_32_port, A_nso(31) => SHIFT_n_12_31_port,
                           A_nso(30) => SHIFT_n_12_30_port, A_nso(29) => 
                           SHIFT_n_12_29_port, A_nso(28) => SHIFT_n_12_28_port,
                           A_nso(27) => SHIFT_n_12_27_port, A_nso(26) => 
                           SHIFT_n_12_26_port, A_nso(25) => SHIFT_n_12_25_port,
                           A_nso(24) => SHIFT_n_12_24_port, A_nso(23) => 
                           SHIFT_n_12_23_port, A_nso(22) => SHIFT_n_12_22_port,
                           A_nso(21) => SHIFT_n_12_21_port, A_nso(20) => 
                           SHIFT_n_12_20_port, A_nso(19) => SHIFT_n_12_19_port,
                           A_nso(18) => SHIFT_n_12_18_port, A_nso(17) => 
                           SHIFT_n_12_17_port, A_nso(16) => SHIFT_n_12_16_port,
                           A_nso(15) => SHIFT_n_12_15_port, A_nso(14) => 
                           SHIFT_n_12_14_port, A_nso(13) => SHIFT_n_12_13_port,
                           A_nso(12) => SHIFT_n_12_12_port, A_nso(11) => 
                           SHIFT_n_12_11_port, A_nso(10) => SHIFT_n_12_10_port,
                           A_nso(9) => SHIFT_n_12_9_port, A_nso(8) => 
                           SHIFT_n_12_8_port, A_nso(7) => SHIFT_n_12_7_port, 
                           A_nso(6) => SHIFT_n_12_6_port, A_nso(5) => 
                           SHIFT_n_12_5_port, A_nso(4) => SHIFT_n_12_4_port, 
                           A_nso(3) => SHIFT_n_12_3_port, A_nso(2) => 
                           SHIFT_n_12_2_port, A_nso(1) => n_1135, A_nso(0) => 
                           n_1136);
   ENC_12 : BOOTHENC_NBIT58_i24 port map( A_s(57) => SHIFT_12_55_port, A_s(56) 
                           => SHIFT_12_55_port, A_s(55) => SHIFT_12_55_port, 
                           A_s(54) => SHIFT_12_54_port, A_s(53) => 
                           SHIFT_12_53_port, A_s(52) => SHIFT_12_52_port, 
                           A_s(51) => SHIFT_12_51_port, A_s(50) => 
                           SHIFT_12_50_port, A_s(49) => SHIFT_12_49_port, 
                           A_s(48) => SHIFT_12_48_port, A_s(47) => 
                           SHIFT_12_47_port, A_s(46) => SHIFT_12_46_port, 
                           A_s(45) => SHIFT_12_45_port, A_s(44) => 
                           SHIFT_12_44_port, A_s(43) => SHIFT_12_43_port, 
                           A_s(42) => SHIFT_12_42_port, A_s(41) => 
                           SHIFT_12_41_port, A_s(40) => SHIFT_12_40_port, 
                           A_s(39) => SHIFT_12_39_port, A_s(38) => 
                           SHIFT_12_38_port, A_s(37) => SHIFT_12_37_port, 
                           A_s(36) => SHIFT_12_36_port, A_s(35) => 
                           SHIFT_12_35_port, A_s(34) => SHIFT_12_34_port, 
                           A_s(33) => SHIFT_12_33_port, A_s(32) => 
                           SHIFT_12_32_port, A_s(31) => SHIFT_12_31_port, 
                           A_s(30) => SHIFT_12_30_port, A_s(29) => 
                           SHIFT_12_29_port, A_s(28) => SHIFT_12_28_port, 
                           A_s(27) => SHIFT_12_27_port, A_s(26) => 
                           SHIFT_12_26_port, A_s(25) => SHIFT_12_25_port, 
                           A_s(24) => SHIFT_12_24_port, A_s(23) => 
                           SHIFT_12_23_port, A_s(22) => SHIFT_12_22_port, 
                           A_s(21) => SHIFT_12_21_port, A_s(20) => 
                           SHIFT_12_20_port, A_s(19) => SHIFT_12_19_port, 
                           A_s(18) => SHIFT_12_18_port, A_s(17) => 
                           SHIFT_12_17_port, A_s(16) => SHIFT_12_16_port, 
                           A_s(15) => SHIFT_12_15_port, A_s(14) => 
                           SHIFT_12_14_port, A_s(13) => SHIFT_12_13_port, 
                           A_s(12) => SHIFT_12_12_port, A_s(11) => 
                           SHIFT_12_11_port, A_s(10) => SHIFT_12_10_port, 
                           A_s(9) => SHIFT_12_9_port, A_s(8) => SHIFT_12_8_port
                           , A_s(7) => SHIFT_12_7_port, A_s(6) => 
                           SHIFT_12_6_port, A_s(5) => SHIFT_12_5_port, A_s(4) 
                           => SHIFT_12_4_port, A_s(3) => SHIFT_12_3_port, 
                           A_s(2) => SHIFT_12_2_port, A_s(1) => SHIFT_12_1_port
                           , A_s(0) => SHIFT_12_0_port, A_ns(57) => 
                           SHIFT_n_12_55_port, A_ns(56) => SHIFT_n_12_55_port, 
                           A_ns(55) => SHIFT_n_12_55_port, A_ns(54) => 
                           SHIFT_n_12_54_port, A_ns(53) => SHIFT_n_12_53_port, 
                           A_ns(52) => SHIFT_n_12_52_port, A_ns(51) => 
                           SHIFT_n_12_51_port, A_ns(50) => SHIFT_n_12_50_port, 
                           A_ns(49) => SHIFT_n_12_49_port, A_ns(48) => 
                           SHIFT_n_12_48_port, A_ns(47) => SHIFT_n_12_47_port, 
                           A_ns(46) => SHIFT_n_12_46_port, A_ns(45) => 
                           SHIFT_n_12_45_port, A_ns(44) => SHIFT_n_12_44_port, 
                           A_ns(43) => SHIFT_n_12_43_port, A_ns(42) => 
                           SHIFT_n_12_42_port, A_ns(41) => SHIFT_n_12_41_port, 
                           A_ns(40) => SHIFT_n_12_40_port, A_ns(39) => 
                           SHIFT_n_12_39_port, A_ns(38) => SHIFT_n_12_38_port, 
                           A_ns(37) => SHIFT_n_12_37_port, A_ns(36) => 
                           SHIFT_n_12_36_port, A_ns(35) => SHIFT_n_12_35_port, 
                           A_ns(34) => SHIFT_n_12_34_port, A_ns(33) => 
                           SHIFT_n_12_33_port, A_ns(32) => SHIFT_n_12_32_port, 
                           A_ns(31) => SHIFT_n_12_31_port, A_ns(30) => 
                           SHIFT_n_12_30_port, A_ns(29) => SHIFT_n_12_29_port, 
                           A_ns(28) => SHIFT_n_12_28_port, A_ns(27) => 
                           SHIFT_n_12_27_port, A_ns(26) => SHIFT_n_12_26_port, 
                           A_ns(25) => SHIFT_n_12_25_port, A_ns(24) => 
                           SHIFT_n_12_24_port, A_ns(23) => SHIFT_n_12_23_port, 
                           A_ns(22) => SHIFT_n_12_22_port, A_ns(21) => 
                           SHIFT_n_12_21_port, A_ns(20) => SHIFT_n_12_20_port, 
                           A_ns(19) => SHIFT_n_12_19_port, A_ns(18) => 
                           SHIFT_n_12_18_port, A_ns(17) => SHIFT_n_12_17_port, 
                           A_ns(16) => SHIFT_n_12_16_port, A_ns(15) => 
                           SHIFT_n_12_15_port, A_ns(14) => SHIFT_n_12_14_port, 
                           A_ns(13) => SHIFT_n_12_13_port, A_ns(12) => 
                           SHIFT_n_12_12_port, A_ns(11) => SHIFT_n_12_11_port, 
                           A_ns(10) => SHIFT_n_12_10_port, A_ns(9) => 
                           SHIFT_n_12_9_port, A_ns(8) => SHIFT_n_12_8_port, 
                           A_ns(7) => SHIFT_n_12_7_port, A_ns(6) => 
                           SHIFT_n_12_6_port, A_ns(5) => SHIFT_n_12_5_port, 
                           A_ns(4) => SHIFT_n_12_4_port, A_ns(3) => 
                           SHIFT_n_12_3_port, A_ns(2) => SHIFT_n_12_2_port, 
                           A_ns(1) => SHIFT_n_12_1_port, A_ns(0) => 
                           SHIFT_n_12_0_port, B(57) => B(31), B(56) => B(31), 
                           B(55) => B(31), B(54) => B(31), B(53) => B(31), 
                           B(52) => B(31), B(51) => B(31), B(50) => B(31), 
                           B(49) => B(31), B(48) => B(31), B(47) => B(31), 
                           B(46) => B(31), B(45) => B(31), B(44) => B(31), 
                           B(43) => B(31), B(42) => B(31), B(41) => B(31), 
                           B(40) => B(31), B(39) => B(31), B(38) => B(31), 
                           B(37) => B(31), B(36) => B(31), B(35) => B(31), 
                           B(34) => B(31), B(33) => B(31), B(32) => B(31), 
                           B(31) => B(31), B(30) => B(30), B(29) => B(29), 
                           B(28) => B(28), B(27) => B(27), B(26) => B(26), 
                           B(25) => B(25), B(24) => B(24), B(23) => B(23), 
                           B(22) => B(22), B(21) => B(21), B(20) => B(20), 
                           B(19) => B(19), B(18) => B(18), B(17) => B(17), 
                           B(16) => B(16), B(15) => B(15), B(14) => B(14), 
                           B(13) => B(13), B(12) => B(12), B(11) => B(11), 
                           B(10) => B(10), B(9) => B(9), B(8) => B(8), B(7) => 
                           B(7), B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3)
                           => B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), 
                           O(57) => OTMP_12_57_port, O(56) => OTMP_12_56_port, 
                           O(55) => OTMP_12_55_port, O(54) => OTMP_12_54_port, 
                           O(53) => OTMP_12_53_port, O(52) => OTMP_12_52_port, 
                           O(51) => OTMP_12_51_port, O(50) => OTMP_12_50_port, 
                           O(49) => OTMP_12_49_port, O(48) => OTMP_12_48_port, 
                           O(47) => OTMP_12_47_port, O(46) => OTMP_12_46_port, 
                           O(45) => OTMP_12_45_port, O(44) => OTMP_12_44_port, 
                           O(43) => OTMP_12_43_port, O(42) => OTMP_12_42_port, 
                           O(41) => OTMP_12_41_port, O(40) => OTMP_12_40_port, 
                           O(39) => OTMP_12_39_port, O(38) => OTMP_12_38_port, 
                           O(37) => OTMP_12_37_port, O(36) => OTMP_12_36_port, 
                           O(35) => OTMP_12_35_port, O(34) => OTMP_12_34_port, 
                           O(33) => OTMP_12_33_port, O(32) => OTMP_12_32_port, 
                           O(31) => OTMP_12_31_port, O(30) => OTMP_12_30_port, 
                           O(29) => OTMP_12_29_port, O(28) => OTMP_12_28_port, 
                           O(27) => OTMP_12_27_port, O(26) => OTMP_12_26_port, 
                           O(25) => OTMP_12_25_port, O(24) => OTMP_12_24_port, 
                           O(23) => OTMP_12_23_port, O(22) => OTMP_12_22_port, 
                           O(21) => OTMP_12_21_port, O(20) => OTMP_12_20_port, 
                           O(19) => OTMP_12_19_port, O(18) => OTMP_12_18_port, 
                           O(17) => OTMP_12_17_port, O(16) => OTMP_12_16_port, 
                           O(15) => OTMP_12_15_port, O(14) => OTMP_12_14_port, 
                           O(13) => OTMP_12_13_port, O(12) => OTMP_12_12_port, 
                           O(11) => OTMP_12_11_port, O(10) => OTMP_12_10_port, 
                           O(9) => OTMP_12_9_port, O(8) => OTMP_12_8_port, O(7)
                           => OTMP_12_7_port, O(6) => OTMP_12_6_port, O(5) => 
                           OTMP_12_5_port, O(4) => OTMP_12_4_port, O(3) => 
                           OTMP_12_3_port, O(2) => OTMP_12_2_port, O(1) => 
                           OTMP_12_1_port, O(0) => n_1137, A_so(57) => 
                           SHIFT_13_57_port, A_so(56) => SHIFT_13_56_port, 
                           A_so(55) => SHIFT_13_55_port, A_so(54) => 
                           SHIFT_13_54_port, A_so(53) => SHIFT_13_53_port, 
                           A_so(52) => SHIFT_13_52_port, A_so(51) => 
                           SHIFT_13_51_port, A_so(50) => SHIFT_13_50_port, 
                           A_so(49) => SHIFT_13_49_port, A_so(48) => 
                           SHIFT_13_48_port, A_so(47) => SHIFT_13_47_port, 
                           A_so(46) => SHIFT_13_46_port, A_so(45) => 
                           SHIFT_13_45_port, A_so(44) => SHIFT_13_44_port, 
                           A_so(43) => SHIFT_13_43_port, A_so(42) => 
                           SHIFT_13_42_port, A_so(41) => SHIFT_13_41_port, 
                           A_so(40) => SHIFT_13_40_port, A_so(39) => 
                           SHIFT_13_39_port, A_so(38) => SHIFT_13_38_port, 
                           A_so(37) => SHIFT_13_37_port, A_so(36) => 
                           SHIFT_13_36_port, A_so(35) => SHIFT_13_35_port, 
                           A_so(34) => SHIFT_13_34_port, A_so(33) => 
                           SHIFT_13_33_port, A_so(32) => SHIFT_13_32_port, 
                           A_so(31) => SHIFT_13_31_port, A_so(30) => 
                           SHIFT_13_30_port, A_so(29) => SHIFT_13_29_port, 
                           A_so(28) => SHIFT_13_28_port, A_so(27) => 
                           SHIFT_13_27_port, A_so(26) => SHIFT_13_26_port, 
                           A_so(25) => SHIFT_13_25_port, A_so(24) => 
                           SHIFT_13_24_port, A_so(23) => SHIFT_13_23_port, 
                           A_so(22) => SHIFT_13_22_port, A_so(21) => 
                           SHIFT_13_21_port, A_so(20) => SHIFT_13_20_port, 
                           A_so(19) => SHIFT_13_19_port, A_so(18) => 
                           SHIFT_13_18_port, A_so(17) => SHIFT_13_17_port, 
                           A_so(16) => SHIFT_13_16_port, A_so(15) => 
                           SHIFT_13_15_port, A_so(14) => SHIFT_13_14_port, 
                           A_so(13) => SHIFT_13_13_port, A_so(12) => 
                           SHIFT_13_12_port, A_so(11) => SHIFT_13_11_port, 
                           A_so(10) => SHIFT_13_10_port, A_so(9) => 
                           SHIFT_13_9_port, A_so(8) => SHIFT_13_8_port, A_so(7)
                           => SHIFT_13_7_port, A_so(6) => SHIFT_13_6_port, 
                           A_so(5) => SHIFT_13_5_port, A_so(4) => 
                           SHIFT_13_4_port, A_so(3) => SHIFT_13_3_port, A_so(2)
                           => SHIFT_13_2_port, A_so(1) => n_1138, A_so(0) => 
                           n_1139, A_nso(57) => SHIFT_n_13_57_port, A_nso(56) 
                           => SHIFT_n_13_56_port, A_nso(55) => 
                           SHIFT_n_13_55_port, A_nso(54) => SHIFT_n_13_54_port,
                           A_nso(53) => SHIFT_n_13_53_port, A_nso(52) => 
                           SHIFT_n_13_52_port, A_nso(51) => SHIFT_n_13_51_port,
                           A_nso(50) => SHIFT_n_13_50_port, A_nso(49) => 
                           SHIFT_n_13_49_port, A_nso(48) => SHIFT_n_13_48_port,
                           A_nso(47) => SHIFT_n_13_47_port, A_nso(46) => 
                           SHIFT_n_13_46_port, A_nso(45) => SHIFT_n_13_45_port,
                           A_nso(44) => SHIFT_n_13_44_port, A_nso(43) => 
                           SHIFT_n_13_43_port, A_nso(42) => SHIFT_n_13_42_port,
                           A_nso(41) => SHIFT_n_13_41_port, A_nso(40) => 
                           SHIFT_n_13_40_port, A_nso(39) => SHIFT_n_13_39_port,
                           A_nso(38) => SHIFT_n_13_38_port, A_nso(37) => 
                           SHIFT_n_13_37_port, A_nso(36) => SHIFT_n_13_36_port,
                           A_nso(35) => SHIFT_n_13_35_port, A_nso(34) => 
                           SHIFT_n_13_34_port, A_nso(33) => SHIFT_n_13_33_port,
                           A_nso(32) => SHIFT_n_13_32_port, A_nso(31) => 
                           SHIFT_n_13_31_port, A_nso(30) => SHIFT_n_13_30_port,
                           A_nso(29) => SHIFT_n_13_29_port, A_nso(28) => 
                           SHIFT_n_13_28_port, A_nso(27) => SHIFT_n_13_27_port,
                           A_nso(26) => SHIFT_n_13_26_port, A_nso(25) => 
                           SHIFT_n_13_25_port, A_nso(24) => SHIFT_n_13_24_port,
                           A_nso(23) => SHIFT_n_13_23_port, A_nso(22) => 
                           SHIFT_n_13_22_port, A_nso(21) => SHIFT_n_13_21_port,
                           A_nso(20) => SHIFT_n_13_20_port, A_nso(19) => 
                           SHIFT_n_13_19_port, A_nso(18) => SHIFT_n_13_18_port,
                           A_nso(17) => SHIFT_n_13_17_port, A_nso(16) => 
                           SHIFT_n_13_16_port, A_nso(15) => SHIFT_n_13_15_port,
                           A_nso(14) => SHIFT_n_13_14_port, A_nso(13) => 
                           SHIFT_n_13_13_port, A_nso(12) => SHIFT_n_13_12_port,
                           A_nso(11) => SHIFT_n_13_11_port, A_nso(10) => 
                           SHIFT_n_13_10_port, A_nso(9) => SHIFT_n_13_9_port, 
                           A_nso(8) => SHIFT_n_13_8_port, A_nso(7) => 
                           SHIFT_n_13_7_port, A_nso(6) => SHIFT_n_13_6_port, 
                           A_nso(5) => SHIFT_n_13_5_port, A_nso(4) => 
                           SHIFT_n_13_4_port, A_nso(3) => SHIFT_n_13_3_port, 
                           A_nso(2) => SHIFT_n_13_2_port, A_nso(1) => n_1140, 
                           A_nso(0) => n_1141);
   ENC_13 : BOOTHENC_NBIT60_i26 port map( A_s(59) => SHIFT_13_57_port, A_s(58) 
                           => SHIFT_13_57_port, A_s(57) => SHIFT_13_57_port, 
                           A_s(56) => SHIFT_13_56_port, A_s(55) => 
                           SHIFT_13_55_port, A_s(54) => SHIFT_13_54_port, 
                           A_s(53) => SHIFT_13_53_port, A_s(52) => 
                           SHIFT_13_52_port, A_s(51) => SHIFT_13_51_port, 
                           A_s(50) => SHIFT_13_50_port, A_s(49) => 
                           SHIFT_13_49_port, A_s(48) => SHIFT_13_48_port, 
                           A_s(47) => SHIFT_13_47_port, A_s(46) => 
                           SHIFT_13_46_port, A_s(45) => SHIFT_13_45_port, 
                           A_s(44) => SHIFT_13_44_port, A_s(43) => 
                           SHIFT_13_43_port, A_s(42) => SHIFT_13_42_port, 
                           A_s(41) => SHIFT_13_41_port, A_s(40) => 
                           SHIFT_13_40_port, A_s(39) => SHIFT_13_39_port, 
                           A_s(38) => SHIFT_13_38_port, A_s(37) => 
                           SHIFT_13_37_port, A_s(36) => SHIFT_13_36_port, 
                           A_s(35) => SHIFT_13_35_port, A_s(34) => 
                           SHIFT_13_34_port, A_s(33) => SHIFT_13_33_port, 
                           A_s(32) => SHIFT_13_32_port, A_s(31) => 
                           SHIFT_13_31_port, A_s(30) => SHIFT_13_30_port, 
                           A_s(29) => SHIFT_13_29_port, A_s(28) => 
                           SHIFT_13_28_port, A_s(27) => SHIFT_13_27_port, 
                           A_s(26) => SHIFT_13_26_port, A_s(25) => 
                           SHIFT_13_25_port, A_s(24) => SHIFT_13_24_port, 
                           A_s(23) => SHIFT_13_23_port, A_s(22) => 
                           SHIFT_13_22_port, A_s(21) => SHIFT_13_21_port, 
                           A_s(20) => SHIFT_13_20_port, A_s(19) => 
                           SHIFT_13_19_port, A_s(18) => SHIFT_13_18_port, 
                           A_s(17) => SHIFT_13_17_port, A_s(16) => 
                           SHIFT_13_16_port, A_s(15) => SHIFT_13_15_port, 
                           A_s(14) => SHIFT_13_14_port, A_s(13) => 
                           SHIFT_13_13_port, A_s(12) => SHIFT_13_12_port, 
                           A_s(11) => SHIFT_13_11_port, A_s(10) => 
                           SHIFT_13_10_port, A_s(9) => SHIFT_13_9_port, A_s(8) 
                           => SHIFT_13_8_port, A_s(7) => SHIFT_13_7_port, 
                           A_s(6) => SHIFT_13_6_port, A_s(5) => SHIFT_13_5_port
                           , A_s(4) => SHIFT_13_4_port, A_s(3) => 
                           SHIFT_13_3_port, A_s(2) => SHIFT_13_2_port, A_s(1) 
                           => SHIFT_13_1_port, A_s(0) => SHIFT_13_0_port, 
                           A_ns(59) => SHIFT_n_13_57_port, A_ns(58) => 
                           SHIFT_n_13_57_port, A_ns(57) => SHIFT_n_13_57_port, 
                           A_ns(56) => SHIFT_n_13_56_port, A_ns(55) => 
                           SHIFT_n_13_55_port, A_ns(54) => SHIFT_n_13_54_port, 
                           A_ns(53) => SHIFT_n_13_53_port, A_ns(52) => 
                           SHIFT_n_13_52_port, A_ns(51) => SHIFT_n_13_51_port, 
                           A_ns(50) => SHIFT_n_13_50_port, A_ns(49) => 
                           SHIFT_n_13_49_port, A_ns(48) => SHIFT_n_13_48_port, 
                           A_ns(47) => SHIFT_n_13_47_port, A_ns(46) => 
                           SHIFT_n_13_46_port, A_ns(45) => SHIFT_n_13_45_port, 
                           A_ns(44) => SHIFT_n_13_44_port, A_ns(43) => 
                           SHIFT_n_13_43_port, A_ns(42) => SHIFT_n_13_42_port, 
                           A_ns(41) => SHIFT_n_13_41_port, A_ns(40) => 
                           SHIFT_n_13_40_port, A_ns(39) => SHIFT_n_13_39_port, 
                           A_ns(38) => SHIFT_n_13_38_port, A_ns(37) => 
                           SHIFT_n_13_37_port, A_ns(36) => SHIFT_n_13_36_port, 
                           A_ns(35) => SHIFT_n_13_35_port, A_ns(34) => 
                           SHIFT_n_13_34_port, A_ns(33) => SHIFT_n_13_33_port, 
                           A_ns(32) => SHIFT_n_13_32_port, A_ns(31) => 
                           SHIFT_n_13_31_port, A_ns(30) => SHIFT_n_13_30_port, 
                           A_ns(29) => SHIFT_n_13_29_port, A_ns(28) => 
                           SHIFT_n_13_28_port, A_ns(27) => SHIFT_n_13_27_port, 
                           A_ns(26) => SHIFT_n_13_26_port, A_ns(25) => 
                           SHIFT_n_13_25_port, A_ns(24) => SHIFT_n_13_24_port, 
                           A_ns(23) => SHIFT_n_13_23_port, A_ns(22) => 
                           SHIFT_n_13_22_port, A_ns(21) => SHIFT_n_13_21_port, 
                           A_ns(20) => SHIFT_n_13_20_port, A_ns(19) => 
                           SHIFT_n_13_19_port, A_ns(18) => SHIFT_n_13_18_port, 
                           A_ns(17) => SHIFT_n_13_17_port, A_ns(16) => 
                           SHIFT_n_13_16_port, A_ns(15) => SHIFT_n_13_15_port, 
                           A_ns(14) => SHIFT_n_13_14_port, A_ns(13) => 
                           SHIFT_n_13_13_port, A_ns(12) => SHIFT_n_13_12_port, 
                           A_ns(11) => SHIFT_n_13_11_port, A_ns(10) => 
                           SHIFT_n_13_10_port, A_ns(9) => SHIFT_n_13_9_port, 
                           A_ns(8) => SHIFT_n_13_8_port, A_ns(7) => 
                           SHIFT_n_13_7_port, A_ns(6) => SHIFT_n_13_6_port, 
                           A_ns(5) => SHIFT_n_13_5_port, A_ns(4) => 
                           SHIFT_n_13_4_port, A_ns(3) => SHIFT_n_13_3_port, 
                           A_ns(2) => SHIFT_n_13_2_port, A_ns(1) => 
                           SHIFT_n_13_1_port, A_ns(0) => SHIFT_n_13_0_port, 
                           B(59) => B(31), B(58) => B(31), B(57) => B(31), 
                           B(56) => B(31), B(55) => B(31), B(54) => B(31), 
                           B(53) => B(31), B(52) => B(31), B(51) => B(31), 
                           B(50) => B(31), B(49) => B(31), B(48) => B(31), 
                           B(47) => B(31), B(46) => B(31), B(45) => B(31), 
                           B(44) => B(31), B(43) => B(31), B(42) => B(31), 
                           B(41) => B(31), B(40) => B(31), B(39) => B(31), 
                           B(38) => B(31), B(37) => B(31), B(36) => B(31), 
                           B(35) => B(31), B(34) => B(31), B(33) => B(31), 
                           B(32) => B(31), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), O(59) => OTMP_13_59_port, O(58) 
                           => OTMP_13_58_port, O(57) => OTMP_13_57_port, O(56) 
                           => OTMP_13_56_port, O(55) => OTMP_13_55_port, O(54) 
                           => OTMP_13_54_port, O(53) => OTMP_13_53_port, O(52) 
                           => OTMP_13_52_port, O(51) => OTMP_13_51_port, O(50) 
                           => OTMP_13_50_port, O(49) => OTMP_13_49_port, O(48) 
                           => OTMP_13_48_port, O(47) => OTMP_13_47_port, O(46) 
                           => OTMP_13_46_port, O(45) => OTMP_13_45_port, O(44) 
                           => OTMP_13_44_port, O(43) => OTMP_13_43_port, O(42) 
                           => OTMP_13_42_port, O(41) => OTMP_13_41_port, O(40) 
                           => OTMP_13_40_port, O(39) => OTMP_13_39_port, O(38) 
                           => OTMP_13_38_port, O(37) => OTMP_13_37_port, O(36) 
                           => OTMP_13_36_port, O(35) => OTMP_13_35_port, O(34) 
                           => OTMP_13_34_port, O(33) => OTMP_13_33_port, O(32) 
                           => OTMP_13_32_port, O(31) => OTMP_13_31_port, O(30) 
                           => OTMP_13_30_port, O(29) => OTMP_13_29_port, O(28) 
                           => OTMP_13_28_port, O(27) => OTMP_13_27_port, O(26) 
                           => OTMP_13_26_port, O(25) => OTMP_13_25_port, O(24) 
                           => OTMP_13_24_port, O(23) => OTMP_13_23_port, O(22) 
                           => OTMP_13_22_port, O(21) => OTMP_13_21_port, O(20) 
                           => OTMP_13_20_port, O(19) => OTMP_13_19_port, O(18) 
                           => OTMP_13_18_port, O(17) => OTMP_13_17_port, O(16) 
                           => OTMP_13_16_port, O(15) => OTMP_13_15_port, O(14) 
                           => OTMP_13_14_port, O(13) => OTMP_13_13_port, O(12) 
                           => OTMP_13_12_port, O(11) => OTMP_13_11_port, O(10) 
                           => OTMP_13_10_port, O(9) => OTMP_13_9_port, O(8) => 
                           OTMP_13_8_port, O(7) => OTMP_13_7_port, O(6) => 
                           OTMP_13_6_port, O(5) => OTMP_13_5_port, O(4) => 
                           OTMP_13_4_port, O(3) => OTMP_13_3_port, O(2) => 
                           OTMP_13_2_port, O(1) => OTMP_13_1_port, O(0) => 
                           n_1142, A_so(59) => SHIFT_14_59_port, A_so(58) => 
                           SHIFT_14_58_port, A_so(57) => SHIFT_14_57_port, 
                           A_so(56) => SHIFT_14_56_port, A_so(55) => 
                           SHIFT_14_55_port, A_so(54) => SHIFT_14_54_port, 
                           A_so(53) => SHIFT_14_53_port, A_so(52) => 
                           SHIFT_14_52_port, A_so(51) => SHIFT_14_51_port, 
                           A_so(50) => SHIFT_14_50_port, A_so(49) => 
                           SHIFT_14_49_port, A_so(48) => SHIFT_14_48_port, 
                           A_so(47) => SHIFT_14_47_port, A_so(46) => 
                           SHIFT_14_46_port, A_so(45) => SHIFT_14_45_port, 
                           A_so(44) => SHIFT_14_44_port, A_so(43) => 
                           SHIFT_14_43_port, A_so(42) => SHIFT_14_42_port, 
                           A_so(41) => SHIFT_14_41_port, A_so(40) => 
                           SHIFT_14_40_port, A_so(39) => SHIFT_14_39_port, 
                           A_so(38) => SHIFT_14_38_port, A_so(37) => 
                           SHIFT_14_37_port, A_so(36) => SHIFT_14_36_port, 
                           A_so(35) => SHIFT_14_35_port, A_so(34) => 
                           SHIFT_14_34_port, A_so(33) => SHIFT_14_33_port, 
                           A_so(32) => SHIFT_14_32_port, A_so(31) => 
                           SHIFT_14_31_port, A_so(30) => SHIFT_14_30_port, 
                           A_so(29) => SHIFT_14_29_port, A_so(28) => 
                           SHIFT_14_28_port, A_so(27) => SHIFT_14_27_port, 
                           A_so(26) => SHIFT_14_26_port, A_so(25) => 
                           SHIFT_14_25_port, A_so(24) => SHIFT_14_24_port, 
                           A_so(23) => SHIFT_14_23_port, A_so(22) => 
                           SHIFT_14_22_port, A_so(21) => SHIFT_14_21_port, 
                           A_so(20) => SHIFT_14_20_port, A_so(19) => 
                           SHIFT_14_19_port, A_so(18) => SHIFT_14_18_port, 
                           A_so(17) => SHIFT_14_17_port, A_so(16) => 
                           SHIFT_14_16_port, A_so(15) => SHIFT_14_15_port, 
                           A_so(14) => SHIFT_14_14_port, A_so(13) => 
                           SHIFT_14_13_port, A_so(12) => SHIFT_14_12_port, 
                           A_so(11) => SHIFT_14_11_port, A_so(10) => 
                           SHIFT_14_10_port, A_so(9) => SHIFT_14_9_port, 
                           A_so(8) => SHIFT_14_8_port, A_so(7) => 
                           SHIFT_14_7_port, A_so(6) => SHIFT_14_6_port, A_so(5)
                           => SHIFT_14_5_port, A_so(4) => SHIFT_14_4_port, 
                           A_so(3) => SHIFT_14_3_port, A_so(2) => 
                           SHIFT_14_2_port, A_so(1) => n_1143, A_so(0) => 
                           n_1144, A_nso(59) => SHIFT_n_14_59_port, A_nso(58) 
                           => SHIFT_n_14_58_port, A_nso(57) => 
                           SHIFT_n_14_57_port, A_nso(56) => SHIFT_n_14_56_port,
                           A_nso(55) => SHIFT_n_14_55_port, A_nso(54) => 
                           SHIFT_n_14_54_port, A_nso(53) => SHIFT_n_14_53_port,
                           A_nso(52) => SHIFT_n_14_52_port, A_nso(51) => 
                           SHIFT_n_14_51_port, A_nso(50) => SHIFT_n_14_50_port,
                           A_nso(49) => SHIFT_n_14_49_port, A_nso(48) => 
                           SHIFT_n_14_48_port, A_nso(47) => SHIFT_n_14_47_port,
                           A_nso(46) => SHIFT_n_14_46_port, A_nso(45) => 
                           SHIFT_n_14_45_port, A_nso(44) => SHIFT_n_14_44_port,
                           A_nso(43) => SHIFT_n_14_43_port, A_nso(42) => 
                           SHIFT_n_14_42_port, A_nso(41) => SHIFT_n_14_41_port,
                           A_nso(40) => SHIFT_n_14_40_port, A_nso(39) => 
                           SHIFT_n_14_39_port, A_nso(38) => SHIFT_n_14_38_port,
                           A_nso(37) => SHIFT_n_14_37_port, A_nso(36) => 
                           SHIFT_n_14_36_port, A_nso(35) => SHIFT_n_14_35_port,
                           A_nso(34) => SHIFT_n_14_34_port, A_nso(33) => 
                           SHIFT_n_14_33_port, A_nso(32) => SHIFT_n_14_32_port,
                           A_nso(31) => SHIFT_n_14_31_port, A_nso(30) => 
                           SHIFT_n_14_30_port, A_nso(29) => SHIFT_n_14_29_port,
                           A_nso(28) => SHIFT_n_14_28_port, A_nso(27) => 
                           SHIFT_n_14_27_port, A_nso(26) => SHIFT_n_14_26_port,
                           A_nso(25) => SHIFT_n_14_25_port, A_nso(24) => 
                           SHIFT_n_14_24_port, A_nso(23) => SHIFT_n_14_23_port,
                           A_nso(22) => SHIFT_n_14_22_port, A_nso(21) => 
                           SHIFT_n_14_21_port, A_nso(20) => SHIFT_n_14_20_port,
                           A_nso(19) => SHIFT_n_14_19_port, A_nso(18) => 
                           SHIFT_n_14_18_port, A_nso(17) => SHIFT_n_14_17_port,
                           A_nso(16) => SHIFT_n_14_16_port, A_nso(15) => 
                           SHIFT_n_14_15_port, A_nso(14) => SHIFT_n_14_14_port,
                           A_nso(13) => SHIFT_n_14_13_port, A_nso(12) => 
                           SHIFT_n_14_12_port, A_nso(11) => SHIFT_n_14_11_port,
                           A_nso(10) => SHIFT_n_14_10_port, A_nso(9) => 
                           SHIFT_n_14_9_port, A_nso(8) => SHIFT_n_14_8_port, 
                           A_nso(7) => SHIFT_n_14_7_port, A_nso(6) => 
                           SHIFT_n_14_6_port, A_nso(5) => SHIFT_n_14_5_port, 
                           A_nso(4) => SHIFT_n_14_4_port, A_nso(3) => 
                           SHIFT_n_14_3_port, A_nso(2) => SHIFT_n_14_2_port, 
                           A_nso(1) => n_1145, A_nso(0) => n_1146);
   ENC_14 : BOOTHENC_NBIT62_i28 port map( A_s(61) => SHIFT_14_59_port, A_s(60) 
                           => SHIFT_14_59_port, A_s(59) => SHIFT_14_59_port, 
                           A_s(58) => SHIFT_14_58_port, A_s(57) => 
                           SHIFT_14_57_port, A_s(56) => SHIFT_14_56_port, 
                           A_s(55) => SHIFT_14_55_port, A_s(54) => 
                           SHIFT_14_54_port, A_s(53) => SHIFT_14_53_port, 
                           A_s(52) => SHIFT_14_52_port, A_s(51) => 
                           SHIFT_14_51_port, A_s(50) => SHIFT_14_50_port, 
                           A_s(49) => SHIFT_14_49_port, A_s(48) => 
                           SHIFT_14_48_port, A_s(47) => SHIFT_14_47_port, 
                           A_s(46) => SHIFT_14_46_port, A_s(45) => 
                           SHIFT_14_45_port, A_s(44) => SHIFT_14_44_port, 
                           A_s(43) => SHIFT_14_43_port, A_s(42) => 
                           SHIFT_14_42_port, A_s(41) => SHIFT_14_41_port, 
                           A_s(40) => SHIFT_14_40_port, A_s(39) => 
                           SHIFT_14_39_port, A_s(38) => SHIFT_14_38_port, 
                           A_s(37) => SHIFT_14_37_port, A_s(36) => 
                           SHIFT_14_36_port, A_s(35) => SHIFT_14_35_port, 
                           A_s(34) => SHIFT_14_34_port, A_s(33) => 
                           SHIFT_14_33_port, A_s(32) => SHIFT_14_32_port, 
                           A_s(31) => SHIFT_14_31_port, A_s(30) => 
                           SHIFT_14_30_port, A_s(29) => SHIFT_14_29_port, 
                           A_s(28) => SHIFT_14_28_port, A_s(27) => 
                           SHIFT_14_27_port, A_s(26) => SHIFT_14_26_port, 
                           A_s(25) => SHIFT_14_25_port, A_s(24) => 
                           SHIFT_14_24_port, A_s(23) => SHIFT_14_23_port, 
                           A_s(22) => SHIFT_14_22_port, A_s(21) => 
                           SHIFT_14_21_port, A_s(20) => SHIFT_14_20_port, 
                           A_s(19) => SHIFT_14_19_port, A_s(18) => 
                           SHIFT_14_18_port, A_s(17) => SHIFT_14_17_port, 
                           A_s(16) => SHIFT_14_16_port, A_s(15) => 
                           SHIFT_14_15_port, A_s(14) => SHIFT_14_14_port, 
                           A_s(13) => SHIFT_14_13_port, A_s(12) => 
                           SHIFT_14_12_port, A_s(11) => SHIFT_14_11_port, 
                           A_s(10) => SHIFT_14_10_port, A_s(9) => 
                           SHIFT_14_9_port, A_s(8) => SHIFT_14_8_port, A_s(7) 
                           => SHIFT_14_7_port, A_s(6) => SHIFT_14_6_port, 
                           A_s(5) => SHIFT_14_5_port, A_s(4) => SHIFT_14_4_port
                           , A_s(3) => SHIFT_14_3_port, A_s(2) => 
                           SHIFT_14_2_port, A_s(1) => SHIFT_14_1_port, A_s(0) 
                           => SHIFT_14_0_port, A_ns(61) => SHIFT_n_14_59_port, 
                           A_ns(60) => SHIFT_n_14_59_port, A_ns(59) => 
                           SHIFT_n_14_59_port, A_ns(58) => SHIFT_n_14_58_port, 
                           A_ns(57) => SHIFT_n_14_57_port, A_ns(56) => 
                           SHIFT_n_14_56_port, A_ns(55) => SHIFT_n_14_55_port, 
                           A_ns(54) => SHIFT_n_14_54_port, A_ns(53) => 
                           SHIFT_n_14_53_port, A_ns(52) => SHIFT_n_14_52_port, 
                           A_ns(51) => SHIFT_n_14_51_port, A_ns(50) => 
                           SHIFT_n_14_50_port, A_ns(49) => SHIFT_n_14_49_port, 
                           A_ns(48) => SHIFT_n_14_48_port, A_ns(47) => 
                           SHIFT_n_14_47_port, A_ns(46) => SHIFT_n_14_46_port, 
                           A_ns(45) => SHIFT_n_14_45_port, A_ns(44) => 
                           SHIFT_n_14_44_port, A_ns(43) => SHIFT_n_14_43_port, 
                           A_ns(42) => SHIFT_n_14_42_port, A_ns(41) => 
                           SHIFT_n_14_41_port, A_ns(40) => SHIFT_n_14_40_port, 
                           A_ns(39) => SHIFT_n_14_39_port, A_ns(38) => 
                           SHIFT_n_14_38_port, A_ns(37) => SHIFT_n_14_37_port, 
                           A_ns(36) => SHIFT_n_14_36_port, A_ns(35) => 
                           SHIFT_n_14_35_port, A_ns(34) => SHIFT_n_14_34_port, 
                           A_ns(33) => SHIFT_n_14_33_port, A_ns(32) => 
                           SHIFT_n_14_32_port, A_ns(31) => SHIFT_n_14_31_port, 
                           A_ns(30) => SHIFT_n_14_30_port, A_ns(29) => 
                           SHIFT_n_14_29_port, A_ns(28) => SHIFT_n_14_28_port, 
                           A_ns(27) => SHIFT_n_14_27_port, A_ns(26) => 
                           SHIFT_n_14_26_port, A_ns(25) => SHIFT_n_14_25_port, 
                           A_ns(24) => SHIFT_n_14_24_port, A_ns(23) => 
                           SHIFT_n_14_23_port, A_ns(22) => SHIFT_n_14_22_port, 
                           A_ns(21) => SHIFT_n_14_21_port, A_ns(20) => 
                           SHIFT_n_14_20_port, A_ns(19) => SHIFT_n_14_19_port, 
                           A_ns(18) => SHIFT_n_14_18_port, A_ns(17) => 
                           SHIFT_n_14_17_port, A_ns(16) => SHIFT_n_14_16_port, 
                           A_ns(15) => SHIFT_n_14_15_port, A_ns(14) => 
                           SHIFT_n_14_14_port, A_ns(13) => SHIFT_n_14_13_port, 
                           A_ns(12) => SHIFT_n_14_12_port, A_ns(11) => 
                           SHIFT_n_14_11_port, A_ns(10) => SHIFT_n_14_10_port, 
                           A_ns(9) => SHIFT_n_14_9_port, A_ns(8) => 
                           SHIFT_n_14_8_port, A_ns(7) => SHIFT_n_14_7_port, 
                           A_ns(6) => SHIFT_n_14_6_port, A_ns(5) => 
                           SHIFT_n_14_5_port, A_ns(4) => SHIFT_n_14_4_port, 
                           A_ns(3) => SHIFT_n_14_3_port, A_ns(2) => 
                           SHIFT_n_14_2_port, A_ns(1) => SHIFT_n_14_1_port, 
                           A_ns(0) => SHIFT_n_14_0_port, B(61) => B(31), B(60) 
                           => B(31), B(59) => B(31), B(58) => B(31), B(57) => 
                           B(31), B(56) => B(31), B(55) => B(31), B(54) => 
                           B(31), B(53) => B(31), B(52) => B(31), B(51) => 
                           B(31), B(50) => B(31), B(49) => B(31), B(48) => 
                           B(31), B(47) => B(31), B(46) => B(31), B(45) => 
                           B(31), B(44) => B(31), B(43) => B(31), B(42) => 
                           B(31), B(41) => B(31), B(40) => B(31), B(39) => 
                           B(31), B(38) => B(31), B(37) => B(31), B(36) => 
                           B(31), B(35) => B(31), B(34) => B(31), B(33) => 
                           B(31), B(32) => B(31), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), O(61) => OTMP_14_61_port, 
                           O(60) => OTMP_14_60_port, O(59) => OTMP_14_59_port, 
                           O(58) => OTMP_14_58_port, O(57) => OTMP_14_57_port, 
                           O(56) => OTMP_14_56_port, O(55) => OTMP_14_55_port, 
                           O(54) => OTMP_14_54_port, O(53) => OTMP_14_53_port, 
                           O(52) => OTMP_14_52_port, O(51) => OTMP_14_51_port, 
                           O(50) => OTMP_14_50_port, O(49) => OTMP_14_49_port, 
                           O(48) => OTMP_14_48_port, O(47) => OTMP_14_47_port, 
                           O(46) => OTMP_14_46_port, O(45) => OTMP_14_45_port, 
                           O(44) => OTMP_14_44_port, O(43) => OTMP_14_43_port, 
                           O(42) => OTMP_14_42_port, O(41) => OTMP_14_41_port, 
                           O(40) => OTMP_14_40_port, O(39) => OTMP_14_39_port, 
                           O(38) => OTMP_14_38_port, O(37) => OTMP_14_37_port, 
                           O(36) => OTMP_14_36_port, O(35) => OTMP_14_35_port, 
                           O(34) => OTMP_14_34_port, O(33) => OTMP_14_33_port, 
                           O(32) => OTMP_14_32_port, O(31) => OTMP_14_31_port, 
                           O(30) => OTMP_14_30_port, O(29) => OTMP_14_29_port, 
                           O(28) => OTMP_14_28_port, O(27) => OTMP_14_27_port, 
                           O(26) => OTMP_14_26_port, O(25) => OTMP_14_25_port, 
                           O(24) => OTMP_14_24_port, O(23) => OTMP_14_23_port, 
                           O(22) => OTMP_14_22_port, O(21) => OTMP_14_21_port, 
                           O(20) => OTMP_14_20_port, O(19) => OTMP_14_19_port, 
                           O(18) => OTMP_14_18_port, O(17) => OTMP_14_17_port, 
                           O(16) => OTMP_14_16_port, O(15) => OTMP_14_15_port, 
                           O(14) => OTMP_14_14_port, O(13) => OTMP_14_13_port, 
                           O(12) => OTMP_14_12_port, O(11) => OTMP_14_11_port, 
                           O(10) => OTMP_14_10_port, O(9) => OTMP_14_9_port, 
                           O(8) => OTMP_14_8_port, O(7) => OTMP_14_7_port, O(6)
                           => OTMP_14_6_port, O(5) => OTMP_14_5_port, O(4) => 
                           OTMP_14_4_port, O(3) => OTMP_14_3_port, O(2) => 
                           OTMP_14_2_port, O(1) => OTMP_14_1_port, O(0) => 
                           n_1147, A_so(61) => SHIFT_15_61_port, A_so(60) => 
                           SHIFT_15_60_port, A_so(59) => SHIFT_15_59_port, 
                           A_so(58) => SHIFT_15_58_port, A_so(57) => 
                           SHIFT_15_57_port, A_so(56) => SHIFT_15_56_port, 
                           A_so(55) => SHIFT_15_55_port, A_so(54) => 
                           SHIFT_15_54_port, A_so(53) => SHIFT_15_53_port, 
                           A_so(52) => SHIFT_15_52_port, A_so(51) => 
                           SHIFT_15_51_port, A_so(50) => SHIFT_15_50_port, 
                           A_so(49) => SHIFT_15_49_port, A_so(48) => 
                           SHIFT_15_48_port, A_so(47) => SHIFT_15_47_port, 
                           A_so(46) => SHIFT_15_46_port, A_so(45) => 
                           SHIFT_15_45_port, A_so(44) => SHIFT_15_44_port, 
                           A_so(43) => SHIFT_15_43_port, A_so(42) => 
                           SHIFT_15_42_port, A_so(41) => SHIFT_15_41_port, 
                           A_so(40) => SHIFT_15_40_port, A_so(39) => 
                           SHIFT_15_39_port, A_so(38) => SHIFT_15_38_port, 
                           A_so(37) => SHIFT_15_37_port, A_so(36) => 
                           SHIFT_15_36_port, A_so(35) => SHIFT_15_35_port, 
                           A_so(34) => SHIFT_15_34_port, A_so(33) => 
                           SHIFT_15_33_port, A_so(32) => SHIFT_15_32_port, 
                           A_so(31) => SHIFT_15_31_port, A_so(30) => 
                           SHIFT_15_30_port, A_so(29) => SHIFT_15_29_port, 
                           A_so(28) => SHIFT_15_28_port, A_so(27) => 
                           SHIFT_15_27_port, A_so(26) => SHIFT_15_26_port, 
                           A_so(25) => SHIFT_15_25_port, A_so(24) => 
                           SHIFT_15_24_port, A_so(23) => SHIFT_15_23_port, 
                           A_so(22) => SHIFT_15_22_port, A_so(21) => 
                           SHIFT_15_21_port, A_so(20) => SHIFT_15_20_port, 
                           A_so(19) => SHIFT_15_19_port, A_so(18) => 
                           SHIFT_15_18_port, A_so(17) => SHIFT_15_17_port, 
                           A_so(16) => SHIFT_15_16_port, A_so(15) => 
                           SHIFT_15_15_port, A_so(14) => SHIFT_15_14_port, 
                           A_so(13) => SHIFT_15_13_port, A_so(12) => 
                           SHIFT_15_12_port, A_so(11) => SHIFT_15_11_port, 
                           A_so(10) => SHIFT_15_10_port, A_so(9) => 
                           SHIFT_15_9_port, A_so(8) => SHIFT_15_8_port, A_so(7)
                           => SHIFT_15_7_port, A_so(6) => SHIFT_15_6_port, 
                           A_so(5) => SHIFT_15_5_port, A_so(4) => 
                           SHIFT_15_4_port, A_so(3) => SHIFT_15_3_port, A_so(2)
                           => SHIFT_15_2_port, A_so(1) => n_1148, A_so(0) => 
                           n_1149, A_nso(61) => SHIFT_n_15_61_port, A_nso(60) 
                           => SHIFT_n_15_60_port, A_nso(59) => 
                           SHIFT_n_15_59_port, A_nso(58) => SHIFT_n_15_58_port,
                           A_nso(57) => SHIFT_n_15_57_port, A_nso(56) => 
                           SHIFT_n_15_56_port, A_nso(55) => SHIFT_n_15_55_port,
                           A_nso(54) => SHIFT_n_15_54_port, A_nso(53) => 
                           SHIFT_n_15_53_port, A_nso(52) => SHIFT_n_15_52_port,
                           A_nso(51) => SHIFT_n_15_51_port, A_nso(50) => 
                           SHIFT_n_15_50_port, A_nso(49) => SHIFT_n_15_49_port,
                           A_nso(48) => SHIFT_n_15_48_port, A_nso(47) => 
                           SHIFT_n_15_47_port, A_nso(46) => SHIFT_n_15_46_port,
                           A_nso(45) => SHIFT_n_15_45_port, A_nso(44) => 
                           SHIFT_n_15_44_port, A_nso(43) => SHIFT_n_15_43_port,
                           A_nso(42) => SHIFT_n_15_42_port, A_nso(41) => 
                           SHIFT_n_15_41_port, A_nso(40) => SHIFT_n_15_40_port,
                           A_nso(39) => SHIFT_n_15_39_port, A_nso(38) => 
                           SHIFT_n_15_38_port, A_nso(37) => SHIFT_n_15_37_port,
                           A_nso(36) => SHIFT_n_15_36_port, A_nso(35) => 
                           SHIFT_n_15_35_port, A_nso(34) => SHIFT_n_15_34_port,
                           A_nso(33) => SHIFT_n_15_33_port, A_nso(32) => 
                           SHIFT_n_15_32_port, A_nso(31) => SHIFT_n_15_31_port,
                           A_nso(30) => SHIFT_n_15_30_port, A_nso(29) => 
                           SHIFT_n_15_29_port, A_nso(28) => SHIFT_n_15_28_port,
                           A_nso(27) => SHIFT_n_15_27_port, A_nso(26) => 
                           SHIFT_n_15_26_port, A_nso(25) => SHIFT_n_15_25_port,
                           A_nso(24) => SHIFT_n_15_24_port, A_nso(23) => 
                           SHIFT_n_15_23_port, A_nso(22) => SHIFT_n_15_22_port,
                           A_nso(21) => SHIFT_n_15_21_port, A_nso(20) => 
                           SHIFT_n_15_20_port, A_nso(19) => SHIFT_n_15_19_port,
                           A_nso(18) => SHIFT_n_15_18_port, A_nso(17) => 
                           SHIFT_n_15_17_port, A_nso(16) => SHIFT_n_15_16_port,
                           A_nso(15) => SHIFT_n_15_15_port, A_nso(14) => 
                           SHIFT_n_15_14_port, A_nso(13) => SHIFT_n_15_13_port,
                           A_nso(12) => SHIFT_n_15_12_port, A_nso(11) => 
                           SHIFT_n_15_11_port, A_nso(10) => SHIFT_n_15_10_port,
                           A_nso(9) => SHIFT_n_15_9_port, A_nso(8) => 
                           SHIFT_n_15_8_port, A_nso(7) => SHIFT_n_15_7_port, 
                           A_nso(6) => SHIFT_n_15_6_port, A_nso(5) => 
                           SHIFT_n_15_5_port, A_nso(4) => SHIFT_n_15_4_port, 
                           A_nso(3) => SHIFT_n_15_3_port, A_nso(2) => 
                           SHIFT_n_15_2_port, A_nso(1) => n_1150, A_nso(0) => 
                           n_1151);
   ENC_15 : BOOTHENC_NBIT64_i30 port map( A_s(63) => SHIFT_15_61_port, A_s(62) 
                           => SHIFT_15_61_port, A_s(61) => SHIFT_15_61_port, 
                           A_s(60) => SHIFT_15_60_port, A_s(59) => 
                           SHIFT_15_59_port, A_s(58) => SHIFT_15_58_port, 
                           A_s(57) => SHIFT_15_57_port, A_s(56) => 
                           SHIFT_15_56_port, A_s(55) => SHIFT_15_55_port, 
                           A_s(54) => SHIFT_15_54_port, A_s(53) => 
                           SHIFT_15_53_port, A_s(52) => SHIFT_15_52_port, 
                           A_s(51) => SHIFT_15_51_port, A_s(50) => 
                           SHIFT_15_50_port, A_s(49) => SHIFT_15_49_port, 
                           A_s(48) => SHIFT_15_48_port, A_s(47) => 
                           SHIFT_15_47_port, A_s(46) => SHIFT_15_46_port, 
                           A_s(45) => SHIFT_15_45_port, A_s(44) => 
                           SHIFT_15_44_port, A_s(43) => SHIFT_15_43_port, 
                           A_s(42) => SHIFT_15_42_port, A_s(41) => 
                           SHIFT_15_41_port, A_s(40) => SHIFT_15_40_port, 
                           A_s(39) => SHIFT_15_39_port, A_s(38) => 
                           SHIFT_15_38_port, A_s(37) => SHIFT_15_37_port, 
                           A_s(36) => SHIFT_15_36_port, A_s(35) => 
                           SHIFT_15_35_port, A_s(34) => SHIFT_15_34_port, 
                           A_s(33) => SHIFT_15_33_port, A_s(32) => 
                           SHIFT_15_32_port, A_s(31) => SHIFT_15_31_port, 
                           A_s(30) => SHIFT_15_30_port, A_s(29) => 
                           SHIFT_15_29_port, A_s(28) => SHIFT_15_28_port, 
                           A_s(27) => SHIFT_15_27_port, A_s(26) => 
                           SHIFT_15_26_port, A_s(25) => SHIFT_15_25_port, 
                           A_s(24) => SHIFT_15_24_port, A_s(23) => 
                           SHIFT_15_23_port, A_s(22) => SHIFT_15_22_port, 
                           A_s(21) => SHIFT_15_21_port, A_s(20) => 
                           SHIFT_15_20_port, A_s(19) => SHIFT_15_19_port, 
                           A_s(18) => SHIFT_15_18_port, A_s(17) => 
                           SHIFT_15_17_port, A_s(16) => SHIFT_15_16_port, 
                           A_s(15) => SHIFT_15_15_port, A_s(14) => 
                           SHIFT_15_14_port, A_s(13) => SHIFT_15_13_port, 
                           A_s(12) => SHIFT_15_12_port, A_s(11) => 
                           SHIFT_15_11_port, A_s(10) => SHIFT_15_10_port, 
                           A_s(9) => SHIFT_15_9_port, A_s(8) => SHIFT_15_8_port
                           , A_s(7) => SHIFT_15_7_port, A_s(6) => 
                           SHIFT_15_6_port, A_s(5) => SHIFT_15_5_port, A_s(4) 
                           => SHIFT_15_4_port, A_s(3) => SHIFT_15_3_port, 
                           A_s(2) => SHIFT_15_2_port, A_s(1) => SHIFT_15_1_port
                           , A_s(0) => SHIFT_15_0_port, A_ns(63) => 
                           SHIFT_n_15_61_port, A_ns(62) => SHIFT_n_15_61_port, 
                           A_ns(61) => SHIFT_n_15_61_port, A_ns(60) => 
                           SHIFT_n_15_60_port, A_ns(59) => SHIFT_n_15_59_port, 
                           A_ns(58) => SHIFT_n_15_58_port, A_ns(57) => 
                           SHIFT_n_15_57_port, A_ns(56) => SHIFT_n_15_56_port, 
                           A_ns(55) => SHIFT_n_15_55_port, A_ns(54) => 
                           SHIFT_n_15_54_port, A_ns(53) => SHIFT_n_15_53_port, 
                           A_ns(52) => SHIFT_n_15_52_port, A_ns(51) => 
                           SHIFT_n_15_51_port, A_ns(50) => SHIFT_n_15_50_port, 
                           A_ns(49) => SHIFT_n_15_49_port, A_ns(48) => 
                           SHIFT_n_15_48_port, A_ns(47) => SHIFT_n_15_47_port, 
                           A_ns(46) => SHIFT_n_15_46_port, A_ns(45) => 
                           SHIFT_n_15_45_port, A_ns(44) => SHIFT_n_15_44_port, 
                           A_ns(43) => SHIFT_n_15_43_port, A_ns(42) => 
                           SHIFT_n_15_42_port, A_ns(41) => SHIFT_n_15_41_port, 
                           A_ns(40) => SHIFT_n_15_40_port, A_ns(39) => 
                           SHIFT_n_15_39_port, A_ns(38) => SHIFT_n_15_38_port, 
                           A_ns(37) => SHIFT_n_15_37_port, A_ns(36) => 
                           SHIFT_n_15_36_port, A_ns(35) => SHIFT_n_15_35_port, 
                           A_ns(34) => SHIFT_n_15_34_port, A_ns(33) => 
                           SHIFT_n_15_33_port, A_ns(32) => SHIFT_n_15_32_port, 
                           A_ns(31) => SHIFT_n_15_31_port, A_ns(30) => 
                           SHIFT_n_15_30_port, A_ns(29) => SHIFT_n_15_29_port, 
                           A_ns(28) => SHIFT_n_15_28_port, A_ns(27) => 
                           SHIFT_n_15_27_port, A_ns(26) => SHIFT_n_15_26_port, 
                           A_ns(25) => SHIFT_n_15_25_port, A_ns(24) => 
                           SHIFT_n_15_24_port, A_ns(23) => SHIFT_n_15_23_port, 
                           A_ns(22) => SHIFT_n_15_22_port, A_ns(21) => 
                           SHIFT_n_15_21_port, A_ns(20) => SHIFT_n_15_20_port, 
                           A_ns(19) => SHIFT_n_15_19_port, A_ns(18) => 
                           SHIFT_n_15_18_port, A_ns(17) => SHIFT_n_15_17_port, 
                           A_ns(16) => SHIFT_n_15_16_port, A_ns(15) => 
                           SHIFT_n_15_15_port, A_ns(14) => SHIFT_n_15_14_port, 
                           A_ns(13) => SHIFT_n_15_13_port, A_ns(12) => 
                           SHIFT_n_15_12_port, A_ns(11) => SHIFT_n_15_11_port, 
                           A_ns(10) => SHIFT_n_15_10_port, A_ns(9) => 
                           SHIFT_n_15_9_port, A_ns(8) => SHIFT_n_15_8_port, 
                           A_ns(7) => SHIFT_n_15_7_port, A_ns(6) => 
                           SHIFT_n_15_6_port, A_ns(5) => SHIFT_n_15_5_port, 
                           A_ns(4) => SHIFT_n_15_4_port, A_ns(3) => 
                           SHIFT_n_15_3_port, A_ns(2) => SHIFT_n_15_2_port, 
                           A_ns(1) => SHIFT_n_15_1_port, A_ns(0) => 
                           SHIFT_n_15_0_port, B(63) => B(31), B(62) => B(31), 
                           B(61) => B(31), B(60) => B(31), B(59) => B(31), 
                           B(58) => B(31), B(57) => B(31), B(56) => B(31), 
                           B(55) => B(31), B(54) => B(31), B(53) => B(31), 
                           B(52) => B(31), B(51) => B(31), B(50) => B(31), 
                           B(49) => B(31), B(48) => B(31), B(47) => B(31), 
                           B(46) => B(31), B(45) => B(31), B(44) => B(31), 
                           B(43) => B(31), B(42) => B(31), B(41) => B(31), 
                           B(40) => B(31), B(39) => B(31), B(38) => B(31), 
                           B(37) => B(31), B(36) => B(31), B(35) => B(31), 
                           B(34) => B(31), B(33) => B(31), B(32) => B(31), 
                           B(31) => B(31), B(30) => B(30), B(29) => B(29), 
                           B(28) => B(28), B(27) => B(27), B(26) => B(26), 
                           B(25) => B(25), B(24) => B(24), B(23) => B(23), 
                           B(22) => B(22), B(21) => B(21), B(20) => B(20), 
                           B(19) => B(19), B(18) => B(18), B(17) => B(17), 
                           B(16) => B(16), B(15) => B(15), B(14) => B(14), 
                           B(13) => B(13), B(12) => B(12), B(11) => B(11), 
                           B(10) => B(10), B(9) => B(9), B(8) => B(8), B(7) => 
                           B(7), B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3)
                           => B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), 
                           O(63) => OTMP_15_63_port, O(62) => OTMP_15_62_port, 
                           O(61) => OTMP_15_61_port, O(60) => OTMP_15_60_port, 
                           O(59) => OTMP_15_59_port, O(58) => OTMP_15_58_port, 
                           O(57) => OTMP_15_57_port, O(56) => OTMP_15_56_port, 
                           O(55) => OTMP_15_55_port, O(54) => OTMP_15_54_port, 
                           O(53) => OTMP_15_53_port, O(52) => OTMP_15_52_port, 
                           O(51) => OTMP_15_51_port, O(50) => OTMP_15_50_port, 
                           O(49) => OTMP_15_49_port, O(48) => OTMP_15_48_port, 
                           O(47) => OTMP_15_47_port, O(46) => OTMP_15_46_port, 
                           O(45) => OTMP_15_45_port, O(44) => OTMP_15_44_port, 
                           O(43) => OTMP_15_43_port, O(42) => OTMP_15_42_port, 
                           O(41) => OTMP_15_41_port, O(40) => OTMP_15_40_port, 
                           O(39) => OTMP_15_39_port, O(38) => OTMP_15_38_port, 
                           O(37) => OTMP_15_37_port, O(36) => OTMP_15_36_port, 
                           O(35) => OTMP_15_35_port, O(34) => OTMP_15_34_port, 
                           O(33) => OTMP_15_33_port, O(32) => OTMP_15_32_port, 
                           O(31) => OTMP_15_31_port, O(30) => OTMP_15_30_port, 
                           O(29) => OTMP_15_29_port, O(28) => OTMP_15_28_port, 
                           O(27) => OTMP_15_27_port, O(26) => OTMP_15_26_port, 
                           O(25) => OTMP_15_25_port, O(24) => OTMP_15_24_port, 
                           O(23) => OTMP_15_23_port, O(22) => OTMP_15_22_port, 
                           O(21) => OTMP_15_21_port, O(20) => OTMP_15_20_port, 
                           O(19) => OTMP_15_19_port, O(18) => OTMP_15_18_port, 
                           O(17) => OTMP_15_17_port, O(16) => OTMP_15_16_port, 
                           O(15) => OTMP_15_15_port, O(14) => OTMP_15_14_port, 
                           O(13) => OTMP_15_13_port, O(12) => OTMP_15_12_port, 
                           O(11) => OTMP_15_11_port, O(10) => OTMP_15_10_port, 
                           O(9) => OTMP_15_9_port, O(8) => OTMP_15_8_port, O(7)
                           => OTMP_15_7_port, O(6) => OTMP_15_6_port, O(5) => 
                           OTMP_15_5_port, O(4) => OTMP_15_4_port, O(3) => 
                           OTMP_15_3_port, O(2) => OTMP_15_2_port, O(1) => 
                           OTMP_15_1_port, O(0) => n_1152, A_so(63) => n_1153, 
                           A_so(62) => n_1154, A_so(61) => n_1155, A_so(60) => 
                           n_1156, A_so(59) => n_1157, A_so(58) => n_1158, 
                           A_so(57) => n_1159, A_so(56) => n_1160, A_so(55) => 
                           n_1161, A_so(54) => n_1162, A_so(53) => n_1163, 
                           A_so(52) => n_1164, A_so(51) => n_1165, A_so(50) => 
                           n_1166, A_so(49) => n_1167, A_so(48) => n_1168, 
                           A_so(47) => n_1169, A_so(46) => n_1170, A_so(45) => 
                           n_1171, A_so(44) => n_1172, A_so(43) => n_1173, 
                           A_so(42) => n_1174, A_so(41) => n_1175, A_so(40) => 
                           n_1176, A_so(39) => n_1177, A_so(38) => n_1178, 
                           A_so(37) => n_1179, A_so(36) => n_1180, A_so(35) => 
                           n_1181, A_so(34) => n_1182, A_so(33) => n_1183, 
                           A_so(32) => n_1184, A_so(31) => n_1185, A_so(30) => 
                           n_1186, A_so(29) => n_1187, A_so(28) => n_1188, 
                           A_so(27) => n_1189, A_so(26) => n_1190, A_so(25) => 
                           n_1191, A_so(24) => n_1192, A_so(23) => n_1193, 
                           A_so(22) => n_1194, A_so(21) => n_1195, A_so(20) => 
                           n_1196, A_so(19) => n_1197, A_so(18) => n_1198, 
                           A_so(17) => n_1199, A_so(16) => n_1200, A_so(15) => 
                           n_1201, A_so(14) => n_1202, A_so(13) => n_1203, 
                           A_so(12) => n_1204, A_so(11) => n_1205, A_so(10) => 
                           n_1206, A_so(9) => n_1207, A_so(8) => n_1208, 
                           A_so(7) => n_1209, A_so(6) => n_1210, A_so(5) => 
                           n_1211, A_so(4) => n_1212, A_so(3) => n_1213, 
                           A_so(2) => n_1214, A_so(1) => n_1215, A_so(0) => 
                           n_1216, A_nso(63) => n_1217, A_nso(62) => n_1218, 
                           A_nso(61) => n_1219, A_nso(60) => n_1220, A_nso(59) 
                           => n_1221, A_nso(58) => n_1222, A_nso(57) => n_1223,
                           A_nso(56) => n_1224, A_nso(55) => n_1225, A_nso(54) 
                           => n_1226, A_nso(53) => n_1227, A_nso(52) => n_1228,
                           A_nso(51) => n_1229, A_nso(50) => n_1230, A_nso(49) 
                           => n_1231, A_nso(48) => n_1232, A_nso(47) => n_1233,
                           A_nso(46) => n_1234, A_nso(45) => n_1235, A_nso(44) 
                           => n_1236, A_nso(43) => n_1237, A_nso(42) => n_1238,
                           A_nso(41) => n_1239, A_nso(40) => n_1240, A_nso(39) 
                           => n_1241, A_nso(38) => n_1242, A_nso(37) => n_1243,
                           A_nso(36) => n_1244, A_nso(35) => n_1245, A_nso(34) 
                           => n_1246, A_nso(33) => n_1247, A_nso(32) => n_1248,
                           A_nso(31) => n_1249, A_nso(30) => n_1250, A_nso(29) 
                           => n_1251, A_nso(28) => n_1252, A_nso(27) => n_1253,
                           A_nso(26) => n_1254, A_nso(25) => n_1255, A_nso(24) 
                           => n_1256, A_nso(23) => n_1257, A_nso(22) => n_1258,
                           A_nso(21) => n_1259, A_nso(20) => n_1260, A_nso(19) 
                           => n_1261, A_nso(18) => n_1262, A_nso(17) => n_1263,
                           A_nso(16) => n_1264, A_nso(15) => n_1265, A_nso(14) 
                           => n_1266, A_nso(13) => n_1267, A_nso(12) => n_1268,
                           A_nso(11) => n_1269, A_nso(10) => n_1270, A_nso(9) 
                           => n_1271, A_nso(8) => n_1272, A_nso(7) => n_1273, 
                           A_nso(6) => n_1274, A_nso(5) => n_1275, A_nso(4) => 
                           n_1276, A_nso(3) => n_1277, A_nso(2) => n_1278, 
                           A_nso(1) => n_1279, A_nso(0) => n_1280);
   ADDER1 : RCA_NBIT36 port map( A(35) => OTMP_0_34_port, A(34) => 
                           OTMP_0_34_port, A(33) => OTMP_0_34_port, A(32) => 
                           OTMP_0_32_port, A(31) => OTMP_0_31_port, A(30) => 
                           OTMP_0_30_port, A(29) => OTMP_0_29_port, A(28) => 
                           OTMP_0_28_port, A(27) => OTMP_0_27_port, A(26) => 
                           OTMP_0_26_port, A(25) => OTMP_0_25_port, A(24) => 
                           OTMP_0_24_port, A(23) => OTMP_0_23_port, A(22) => 
                           OTMP_0_22_port, A(21) => OTMP_0_21_port, A(20) => 
                           OTMP_0_20_port, A(19) => OTMP_0_19_port, A(18) => 
                           OTMP_0_18_port, A(17) => OTMP_0_17_port, A(16) => 
                           OTMP_0_16_port, A(15) => OTMP_0_15_port, A(14) => 
                           OTMP_0_14_port, A(13) => OTMP_0_13_port, A(12) => 
                           OTMP_0_12_port, A(11) => OTMP_0_11_port, A(10) => 
                           OTMP_0_10_port, A(9) => OTMP_0_9_port, A(8) => 
                           OTMP_0_8_port, A(7) => OTMP_0_7_port, A(6) => 
                           OTMP_0_6_port, A(5) => OTMP_0_5_port, A(4) => 
                           OTMP_0_4_port, A(3) => OTMP_0_3_port, A(2) => 
                           OTMP_0_2_port, A(1) => OTMP_0_1_port, A(0) => 
                           OTMP_0_0_port, B(35) => OTMP_1_35_port, B(34) => 
                           OTMP_1_34_port, B(33) => OTMP_1_33_port, B(32) => 
                           OTMP_1_32_port, B(31) => OTMP_1_31_port, B(30) => 
                           OTMP_1_30_port, B(29) => OTMP_1_29_port, B(28) => 
                           OTMP_1_28_port, B(27) => OTMP_1_27_port, B(26) => 
                           OTMP_1_26_port, B(25) => OTMP_1_25_port, B(24) => 
                           OTMP_1_24_port, B(23) => OTMP_1_23_port, B(22) => 
                           OTMP_1_22_port, B(21) => OTMP_1_21_port, B(20) => 
                           OTMP_1_20_port, B(19) => OTMP_1_19_port, B(18) => 
                           OTMP_1_18_port, B(17) => OTMP_1_17_port, B(16) => 
                           OTMP_1_16_port, B(15) => OTMP_1_15_port, B(14) => 
                           OTMP_1_14_port, B(13) => OTMP_1_13_port, B(12) => 
                           OTMP_1_12_port, B(11) => OTMP_1_11_port, B(10) => 
                           OTMP_1_10_port, B(9) => OTMP_1_9_port, B(8) => 
                           OTMP_1_8_port, B(7) => OTMP_1_7_port, B(6) => 
                           OTMP_1_6_port, B(5) => OTMP_1_5_port, B(4) => 
                           OTMP_1_4_port, B(3) => OTMP_1_3_port, B(2) => 
                           OTMP_1_2_port, B(1) => OTMP_1_1_port, B(0) => 
                           OTMP_1_0_port, Ci => X_Logic0_port, S(35) => 
                           PTMP_0_36_port, S(34) => PTMP_0_34_port, S(33) => 
                           PTMP_0_33_port, S(32) => PTMP_0_32_port, S(31) => 
                           PTMP_0_31_port, S(30) => PTMP_0_30_port, S(29) => 
                           PTMP_0_29_port, S(28) => PTMP_0_28_port, S(27) => 
                           PTMP_0_27_port, S(26) => PTMP_0_26_port, S(25) => 
                           PTMP_0_25_port, S(24) => PTMP_0_24_port, S(23) => 
                           PTMP_0_23_port, S(22) => PTMP_0_22_port, S(21) => 
                           PTMP_0_21_port, S(20) => PTMP_0_20_port, S(19) => 
                           PTMP_0_19_port, S(18) => PTMP_0_18_port, S(17) => 
                           PTMP_0_17_port, S(16) => PTMP_0_16_port, S(15) => 
                           PTMP_0_15_port, S(14) => PTMP_0_14_port, S(13) => 
                           PTMP_0_13_port, S(12) => PTMP_0_12_port, S(11) => 
                           PTMP_0_11_port, S(10) => PTMP_0_10_port, S(9) => 
                           PTMP_0_9_port, S(8) => PTMP_0_8_port, S(7) => 
                           PTMP_0_7_port, S(6) => PTMP_0_6_port, S(5) => 
                           PTMP_0_5_port, S(4) => PTMP_0_4_port, S(3) => 
                           PTMP_0_3_port, S(2) => PTMP_0_2_port, S(1) => 
                           PTMP_0_1_port, S(0) => PTMP_0_0_port, Co => n_1281);
   ADDER_2 : RCA_NBIT38 port map( A(37) => PTMP_0_36_port, A(36) => 
                           PTMP_0_36_port, A(35) => PTMP_0_36_port, A(34) => 
                           PTMP_0_34_port, A(33) => PTMP_0_33_port, A(32) => 
                           PTMP_0_32_port, A(31) => PTMP_0_31_port, A(30) => 
                           PTMP_0_30_port, A(29) => PTMP_0_29_port, A(28) => 
                           PTMP_0_28_port, A(27) => PTMP_0_27_port, A(26) => 
                           PTMP_0_26_port, A(25) => PTMP_0_25_port, A(24) => 
                           PTMP_0_24_port, A(23) => PTMP_0_23_port, A(22) => 
                           PTMP_0_22_port, A(21) => PTMP_0_21_port, A(20) => 
                           PTMP_0_20_port, A(19) => PTMP_0_19_port, A(18) => 
                           PTMP_0_18_port, A(17) => PTMP_0_17_port, A(16) => 
                           PTMP_0_16_port, A(15) => PTMP_0_15_port, A(14) => 
                           PTMP_0_14_port, A(13) => PTMP_0_13_port, A(12) => 
                           PTMP_0_12_port, A(11) => PTMP_0_11_port, A(10) => 
                           PTMP_0_10_port, A(9) => PTMP_0_9_port, A(8) => 
                           PTMP_0_8_port, A(7) => PTMP_0_7_port, A(6) => 
                           PTMP_0_6_port, A(5) => PTMP_0_5_port, A(4) => 
                           PTMP_0_4_port, A(3) => PTMP_0_3_port, A(2) => 
                           PTMP_0_2_port, A(1) => PTMP_0_1_port, A(0) => 
                           PTMP_0_0_port, B(37) => OTMP_2_37_port, B(36) => 
                           OTMP_2_36_port, B(35) => OTMP_2_35_port, B(34) => 
                           OTMP_2_34_port, B(33) => OTMP_2_33_port, B(32) => 
                           OTMP_2_32_port, B(31) => OTMP_2_31_port, B(30) => 
                           OTMP_2_30_port, B(29) => OTMP_2_29_port, B(28) => 
                           OTMP_2_28_port, B(27) => OTMP_2_27_port, B(26) => 
                           OTMP_2_26_port, B(25) => OTMP_2_25_port, B(24) => 
                           OTMP_2_24_port, B(23) => OTMP_2_23_port, B(22) => 
                           OTMP_2_22_port, B(21) => OTMP_2_21_port, B(20) => 
                           OTMP_2_20_port, B(19) => OTMP_2_19_port, B(18) => 
                           OTMP_2_18_port, B(17) => OTMP_2_17_port, B(16) => 
                           OTMP_2_16_port, B(15) => OTMP_2_15_port, B(14) => 
                           OTMP_2_14_port, B(13) => OTMP_2_13_port, B(12) => 
                           OTMP_2_12_port, B(11) => OTMP_2_11_port, B(10) => 
                           OTMP_2_10_port, B(9) => OTMP_2_9_port, B(8) => 
                           OTMP_2_8_port, B(7) => OTMP_2_7_port, B(6) => 
                           OTMP_2_6_port, B(5) => OTMP_2_5_port, B(4) => 
                           OTMP_2_4_port, B(3) => OTMP_2_3_port, B(2) => 
                           OTMP_2_2_port, B(1) => OTMP_2_1_port, B(0) => 
                           OTMP_2_0_port, Ci => X_Logic0_port, S(37) => 
                           PTMP_1_37_port, S(36) => PTMP_1_36_port, S(35) => 
                           PTMP_1_35_port, S(34) => PTMP_1_34_port, S(33) => 
                           PTMP_1_33_port, S(32) => PTMP_1_32_port, S(31) => 
                           PTMP_1_31_port, S(30) => PTMP_1_30_port, S(29) => 
                           PTMP_1_29_port, S(28) => PTMP_1_28_port, S(27) => 
                           PTMP_1_27_port, S(26) => PTMP_1_26_port, S(25) => 
                           PTMP_1_25_port, S(24) => PTMP_1_24_port, S(23) => 
                           PTMP_1_23_port, S(22) => PTMP_1_22_port, S(21) => 
                           PTMP_1_21_port, S(20) => PTMP_1_20_port, S(19) => 
                           PTMP_1_19_port, S(18) => PTMP_1_18_port, S(17) => 
                           PTMP_1_17_port, S(16) => PTMP_1_16_port, S(15) => 
                           PTMP_1_15_port, S(14) => PTMP_1_14_port, S(13) => 
                           PTMP_1_13_port, S(12) => PTMP_1_12_port, S(11) => 
                           PTMP_1_11_port, S(10) => PTMP_1_10_port, S(9) => 
                           PTMP_1_9_port, S(8) => PTMP_1_8_port, S(7) => 
                           PTMP_1_7_port, S(6) => PTMP_1_6_port, S(5) => 
                           PTMP_1_5_port, S(4) => PTMP_1_4_port, S(3) => 
                           PTMP_1_3_port, S(2) => PTMP_1_2_port, S(1) => 
                           PTMP_1_1_port, S(0) => PTMP_1_0_port, Co => n_1282);
   ADDER_3 : RCA_NBIT40 port map( A(39) => PTMP_1_37_port, A(38) => 
                           PTMP_1_37_port, A(37) => PTMP_1_37_port, A(36) => 
                           PTMP_1_36_port, A(35) => PTMP_1_35_port, A(34) => 
                           PTMP_1_34_port, A(33) => PTMP_1_33_port, A(32) => 
                           PTMP_1_32_port, A(31) => PTMP_1_31_port, A(30) => 
                           PTMP_1_30_port, A(29) => PTMP_1_29_port, A(28) => 
                           PTMP_1_28_port, A(27) => PTMP_1_27_port, A(26) => 
                           PTMP_1_26_port, A(25) => PTMP_1_25_port, A(24) => 
                           PTMP_1_24_port, A(23) => PTMP_1_23_port, A(22) => 
                           PTMP_1_22_port, A(21) => PTMP_1_21_port, A(20) => 
                           PTMP_1_20_port, A(19) => PTMP_1_19_port, A(18) => 
                           PTMP_1_18_port, A(17) => PTMP_1_17_port, A(16) => 
                           PTMP_1_16_port, A(15) => PTMP_1_15_port, A(14) => 
                           PTMP_1_14_port, A(13) => PTMP_1_13_port, A(12) => 
                           PTMP_1_12_port, A(11) => PTMP_1_11_port, A(10) => 
                           PTMP_1_10_port, A(9) => PTMP_1_9_port, A(8) => 
                           PTMP_1_8_port, A(7) => PTMP_1_7_port, A(6) => 
                           PTMP_1_6_port, A(5) => PTMP_1_5_port, A(4) => 
                           PTMP_1_4_port, A(3) => PTMP_1_3_port, A(2) => 
                           PTMP_1_2_port, A(1) => PTMP_1_1_port, A(0) => 
                           PTMP_1_0_port, B(39) => OTMP_3_39_port, B(38) => 
                           OTMP_3_38_port, B(37) => OTMP_3_37_port, B(36) => 
                           OTMP_3_36_port, B(35) => OTMP_3_35_port, B(34) => 
                           OTMP_3_34_port, B(33) => OTMP_3_33_port, B(32) => 
                           OTMP_3_32_port, B(31) => OTMP_3_31_port, B(30) => 
                           OTMP_3_30_port, B(29) => OTMP_3_29_port, B(28) => 
                           OTMP_3_28_port, B(27) => OTMP_3_27_port, B(26) => 
                           OTMP_3_26_port, B(25) => OTMP_3_25_port, B(24) => 
                           OTMP_3_24_port, B(23) => OTMP_3_23_port, B(22) => 
                           OTMP_3_22_port, B(21) => OTMP_3_21_port, B(20) => 
                           OTMP_3_20_port, B(19) => OTMP_3_19_port, B(18) => 
                           OTMP_3_18_port, B(17) => OTMP_3_17_port, B(16) => 
                           OTMP_3_16_port, B(15) => OTMP_3_15_port, B(14) => 
                           OTMP_3_14_port, B(13) => OTMP_3_13_port, B(12) => 
                           OTMP_3_12_port, B(11) => OTMP_3_11_port, B(10) => 
                           OTMP_3_10_port, B(9) => OTMP_3_9_port, B(8) => 
                           OTMP_3_8_port, B(7) => OTMP_3_7_port, B(6) => 
                           OTMP_3_6_port, B(5) => OTMP_3_5_port, B(4) => 
                           OTMP_3_4_port, B(3) => OTMP_3_3_port, B(2) => 
                           OTMP_3_2_port, B(1) => OTMP_3_1_port, B(0) => 
                           OTMP_3_0_port, Ci => X_Logic0_port, S(39) => 
                           PTMP_2_39_port, S(38) => PTMP_2_38_port, S(37) => 
                           PTMP_2_37_port, S(36) => PTMP_2_36_port, S(35) => 
                           PTMP_2_35_port, S(34) => PTMP_2_34_port, S(33) => 
                           PTMP_2_33_port, S(32) => PTMP_2_32_port, S(31) => 
                           PTMP_2_31_port, S(30) => PTMP_2_30_port, S(29) => 
                           PTMP_2_29_port, S(28) => PTMP_2_28_port, S(27) => 
                           PTMP_2_27_port, S(26) => PTMP_2_26_port, S(25) => 
                           PTMP_2_25_port, S(24) => PTMP_2_24_port, S(23) => 
                           PTMP_2_23_port, S(22) => PTMP_2_22_port, S(21) => 
                           PTMP_2_21_port, S(20) => PTMP_2_20_port, S(19) => 
                           PTMP_2_19_port, S(18) => PTMP_2_18_port, S(17) => 
                           PTMP_2_17_port, S(16) => PTMP_2_16_port, S(15) => 
                           PTMP_2_15_port, S(14) => PTMP_2_14_port, S(13) => 
                           PTMP_2_13_port, S(12) => PTMP_2_12_port, S(11) => 
                           PTMP_2_11_port, S(10) => PTMP_2_10_port, S(9) => 
                           PTMP_2_9_port, S(8) => PTMP_2_8_port, S(7) => 
                           PTMP_2_7_port, S(6) => PTMP_2_6_port, S(5) => 
                           PTMP_2_5_port, S(4) => PTMP_2_4_port, S(3) => 
                           PTMP_2_3_port, S(2) => PTMP_2_2_port, S(1) => 
                           PTMP_2_1_port, S(0) => PTMP_2_0_port, Co => n_1283);
   ADDER_4 : RCA_NBIT42 port map( A(41) => n13, A(40) => n13, A(39) => 
                           PTMP_2_39_port, A(38) => PTMP_2_38_port, A(37) => 
                           PTMP_2_37_port, A(36) => PTMP_2_36_port, A(35) => 
                           PTMP_2_35_port, A(34) => PTMP_2_34_port, A(33) => 
                           PTMP_2_33_port, A(32) => PTMP_2_32_port, A(31) => 
                           PTMP_2_31_port, A(30) => PTMP_2_30_port, A(29) => 
                           PTMP_2_29_port, A(28) => PTMP_2_28_port, A(27) => 
                           PTMP_2_27_port, A(26) => PTMP_2_26_port, A(25) => 
                           PTMP_2_25_port, A(24) => PTMP_2_24_port, A(23) => 
                           PTMP_2_23_port, A(22) => PTMP_2_22_port, A(21) => 
                           PTMP_2_21_port, A(20) => PTMP_2_20_port, A(19) => 
                           PTMP_2_19_port, A(18) => PTMP_2_18_port, A(17) => 
                           PTMP_2_17_port, A(16) => PTMP_2_16_port, A(15) => 
                           PTMP_2_15_port, A(14) => PTMP_2_14_port, A(13) => 
                           PTMP_2_13_port, A(12) => PTMP_2_12_port, A(11) => 
                           PTMP_2_11_port, A(10) => PTMP_2_10_port, A(9) => 
                           PTMP_2_9_port, A(8) => PTMP_2_8_port, A(7) => 
                           PTMP_2_7_port, A(6) => PTMP_2_6_port, A(5) => 
                           PTMP_2_5_port, A(4) => PTMP_2_4_port, A(3) => 
                           PTMP_2_3_port, A(2) => PTMP_2_2_port, A(1) => 
                           PTMP_2_1_port, A(0) => PTMP_2_0_port, B(41) => 
                           OTMP_4_41_port, B(40) => OTMP_4_40_port, B(39) => 
                           OTMP_4_39_port, B(38) => OTMP_4_38_port, B(37) => 
                           OTMP_4_37_port, B(36) => OTMP_4_36_port, B(35) => 
                           OTMP_4_35_port, B(34) => OTMP_4_34_port, B(33) => 
                           OTMP_4_33_port, B(32) => OTMP_4_32_port, B(31) => 
                           OTMP_4_31_port, B(30) => OTMP_4_30_port, B(29) => 
                           OTMP_4_29_port, B(28) => OTMP_4_28_port, B(27) => 
                           OTMP_4_27_port, B(26) => OTMP_4_26_port, B(25) => 
                           OTMP_4_25_port, B(24) => OTMP_4_24_port, B(23) => 
                           OTMP_4_23_port, B(22) => OTMP_4_22_port, B(21) => 
                           OTMP_4_21_port, B(20) => OTMP_4_20_port, B(19) => 
                           OTMP_4_19_port, B(18) => OTMP_4_18_port, B(17) => 
                           OTMP_4_17_port, B(16) => OTMP_4_16_port, B(15) => 
                           OTMP_4_15_port, B(14) => OTMP_4_14_port, B(13) => 
                           OTMP_4_13_port, B(12) => OTMP_4_12_port, B(11) => 
                           OTMP_4_11_port, B(10) => OTMP_4_10_port, B(9) => 
                           OTMP_4_9_port, B(8) => OTMP_4_8_port, B(7) => 
                           OTMP_4_7_port, B(6) => OTMP_4_6_port, B(5) => 
                           OTMP_4_5_port, B(4) => OTMP_4_4_port, B(3) => 
                           OTMP_4_3_port, B(2) => OTMP_4_2_port, B(1) => 
                           OTMP_4_1_port, B(0) => OTMP_4_0_port, Ci => 
                           X_Logic0_port, S(41) => PTMP_3_41_port, S(40) => 
                           PTMP_3_40_port, S(39) => PTMP_3_39_port, S(38) => 
                           PTMP_3_38_port, S(37) => PTMP_3_37_port, S(36) => 
                           PTMP_3_36_port, S(35) => PTMP_3_35_port, S(34) => 
                           PTMP_3_34_port, S(33) => PTMP_3_33_port, S(32) => 
                           PTMP_3_32_port, S(31) => PTMP_3_31_port, S(30) => 
                           PTMP_3_30_port, S(29) => PTMP_3_29_port, S(28) => 
                           PTMP_3_28_port, S(27) => PTMP_3_27_port, S(26) => 
                           PTMP_3_26_port, S(25) => PTMP_3_25_port, S(24) => 
                           PTMP_3_24_port, S(23) => PTMP_3_23_port, S(22) => 
                           PTMP_3_22_port, S(21) => PTMP_3_21_port, S(20) => 
                           PTMP_3_20_port, S(19) => PTMP_3_19_port, S(18) => 
                           PTMP_3_18_port, S(17) => PTMP_3_17_port, S(16) => 
                           PTMP_3_16_port, S(15) => PTMP_3_15_port, S(14) => 
                           PTMP_3_14_port, S(13) => PTMP_3_13_port, S(12) => 
                           PTMP_3_12_port, S(11) => PTMP_3_11_port, S(10) => 
                           PTMP_3_10_port, S(9) => PTMP_3_9_port, S(8) => 
                           PTMP_3_8_port, S(7) => PTMP_3_7_port, S(6) => 
                           PTMP_3_6_port, S(5) => PTMP_3_5_port, S(4) => 
                           PTMP_3_4_port, S(3) => PTMP_3_3_port, S(2) => 
                           PTMP_3_2_port, S(1) => PTMP_3_1_port, S(0) => 
                           PTMP_3_0_port, Co => n_1284);
   ADDER_5 : RCA_NBIT44 port map( A(43) => n7, A(42) => n7, A(41) => 
                           PTMP_3_41_port, A(40) => PTMP_3_40_port, A(39) => 
                           PTMP_3_39_port, A(38) => PTMP_3_38_port, A(37) => 
                           PTMP_3_37_port, A(36) => PTMP_3_36_port, A(35) => 
                           PTMP_3_35_port, A(34) => PTMP_3_34_port, A(33) => 
                           PTMP_3_33_port, A(32) => PTMP_3_32_port, A(31) => 
                           PTMP_3_31_port, A(30) => PTMP_3_30_port, A(29) => 
                           PTMP_3_29_port, A(28) => PTMP_3_28_port, A(27) => 
                           PTMP_3_27_port, A(26) => PTMP_3_26_port, A(25) => 
                           PTMP_3_25_port, A(24) => PTMP_3_24_port, A(23) => 
                           PTMP_3_23_port, A(22) => PTMP_3_22_port, A(21) => 
                           PTMP_3_21_port, A(20) => PTMP_3_20_port, A(19) => 
                           PTMP_3_19_port, A(18) => PTMP_3_18_port, A(17) => 
                           PTMP_3_17_port, A(16) => PTMP_3_16_port, A(15) => 
                           PTMP_3_15_port, A(14) => PTMP_3_14_port, A(13) => 
                           PTMP_3_13_port, A(12) => PTMP_3_12_port, A(11) => 
                           PTMP_3_11_port, A(10) => PTMP_3_10_port, A(9) => 
                           PTMP_3_9_port, A(8) => PTMP_3_8_port, A(7) => 
                           PTMP_3_7_port, A(6) => PTMP_3_6_port, A(5) => 
                           PTMP_3_5_port, A(4) => PTMP_3_4_port, A(3) => 
                           PTMP_3_3_port, A(2) => PTMP_3_2_port, A(1) => 
                           PTMP_3_1_port, A(0) => PTMP_3_0_port, B(43) => 
                           OTMP_5_43_port, B(42) => OTMP_5_42_port, B(41) => 
                           OTMP_5_41_port, B(40) => OTMP_5_40_port, B(39) => 
                           OTMP_5_39_port, B(38) => OTMP_5_38_port, B(37) => 
                           OTMP_5_37_port, B(36) => OTMP_5_36_port, B(35) => 
                           OTMP_5_35_port, B(34) => OTMP_5_34_port, B(33) => 
                           OTMP_5_33_port, B(32) => OTMP_5_32_port, B(31) => 
                           OTMP_5_31_port, B(30) => OTMP_5_30_port, B(29) => 
                           OTMP_5_29_port, B(28) => OTMP_5_28_port, B(27) => 
                           OTMP_5_27_port, B(26) => OTMP_5_26_port, B(25) => 
                           OTMP_5_25_port, B(24) => OTMP_5_24_port, B(23) => 
                           OTMP_5_23_port, B(22) => OTMP_5_22_port, B(21) => 
                           OTMP_5_21_port, B(20) => OTMP_5_20_port, B(19) => 
                           OTMP_5_19_port, B(18) => OTMP_5_18_port, B(17) => 
                           OTMP_5_17_port, B(16) => OTMP_5_16_port, B(15) => 
                           OTMP_5_15_port, B(14) => OTMP_5_14_port, B(13) => 
                           OTMP_5_13_port, B(12) => OTMP_5_12_port, B(11) => 
                           OTMP_5_11_port, B(10) => OTMP_5_10_port, B(9) => 
                           OTMP_5_9_port, B(8) => OTMP_5_8_port, B(7) => 
                           OTMP_5_7_port, B(6) => OTMP_5_6_port, B(5) => 
                           OTMP_5_5_port, B(4) => OTMP_5_4_port, B(3) => 
                           OTMP_5_3_port, B(2) => OTMP_5_2_port, B(1) => 
                           OTMP_5_1_port, B(0) => OTMP_5_0_port, Ci => 
                           X_Logic0_port, S(43) => PTMP_4_43_port, S(42) => 
                           PTMP_4_42_port, S(41) => PTMP_4_41_port, S(40) => 
                           PTMP_4_40_port, S(39) => PTMP_4_39_port, S(38) => 
                           PTMP_4_38_port, S(37) => PTMP_4_37_port, S(36) => 
                           PTMP_4_36_port, S(35) => PTMP_4_35_port, S(34) => 
                           PTMP_4_34_port, S(33) => PTMP_4_33_port, S(32) => 
                           PTMP_4_32_port, S(31) => PTMP_4_31_port, S(30) => 
                           PTMP_4_30_port, S(29) => PTMP_4_29_port, S(28) => 
                           PTMP_4_28_port, S(27) => PTMP_4_27_port, S(26) => 
                           PTMP_4_26_port, S(25) => PTMP_4_25_port, S(24) => 
                           PTMP_4_24_port, S(23) => PTMP_4_23_port, S(22) => 
                           PTMP_4_22_port, S(21) => PTMP_4_21_port, S(20) => 
                           PTMP_4_20_port, S(19) => PTMP_4_19_port, S(18) => 
                           PTMP_4_18_port, S(17) => PTMP_4_17_port, S(16) => 
                           PTMP_4_16_port, S(15) => PTMP_4_15_port, S(14) => 
                           PTMP_4_14_port, S(13) => PTMP_4_13_port, S(12) => 
                           PTMP_4_12_port, S(11) => PTMP_4_11_port, S(10) => 
                           PTMP_4_10_port, S(9) => PTMP_4_9_port, S(8) => 
                           PTMP_4_8_port, S(7) => PTMP_4_7_port, S(6) => 
                           PTMP_4_6_port, S(5) => PTMP_4_5_port, S(4) => 
                           PTMP_4_4_port, S(3) => PTMP_4_3_port, S(2) => 
                           PTMP_4_2_port, S(1) => PTMP_4_1_port, S(0) => 
                           PTMP_4_0_port, Co => n_1285);
   ADDER_6 : RCA_NBIT46 port map( A(45) => n12, A(44) => n12, A(43) => 
                           PTMP_4_43_port, A(42) => PTMP_4_42_port, A(41) => 
                           PTMP_4_41_port, A(40) => PTMP_4_40_port, A(39) => 
                           PTMP_4_39_port, A(38) => PTMP_4_38_port, A(37) => 
                           PTMP_4_37_port, A(36) => PTMP_4_36_port, A(35) => 
                           PTMP_4_35_port, A(34) => PTMP_4_34_port, A(33) => 
                           PTMP_4_33_port, A(32) => PTMP_4_32_port, A(31) => 
                           PTMP_4_31_port, A(30) => PTMP_4_30_port, A(29) => 
                           PTMP_4_29_port, A(28) => PTMP_4_28_port, A(27) => 
                           PTMP_4_27_port, A(26) => PTMP_4_26_port, A(25) => 
                           PTMP_4_25_port, A(24) => PTMP_4_24_port, A(23) => 
                           PTMP_4_23_port, A(22) => PTMP_4_22_port, A(21) => 
                           PTMP_4_21_port, A(20) => PTMP_4_20_port, A(19) => 
                           PTMP_4_19_port, A(18) => PTMP_4_18_port, A(17) => 
                           PTMP_4_17_port, A(16) => PTMP_4_16_port, A(15) => 
                           PTMP_4_15_port, A(14) => PTMP_4_14_port, A(13) => 
                           PTMP_4_13_port, A(12) => PTMP_4_12_port, A(11) => 
                           PTMP_4_11_port, A(10) => PTMP_4_10_port, A(9) => 
                           PTMP_4_9_port, A(8) => PTMP_4_8_port, A(7) => 
                           PTMP_4_7_port, A(6) => PTMP_4_6_port, A(5) => 
                           PTMP_4_5_port, A(4) => PTMP_4_4_port, A(3) => 
                           PTMP_4_3_port, A(2) => PTMP_4_2_port, A(1) => 
                           PTMP_4_1_port, A(0) => PTMP_4_0_port, B(45) => 
                           OTMP_6_45_port, B(44) => OTMP_6_44_port, B(43) => 
                           OTMP_6_43_port, B(42) => OTMP_6_42_port, B(41) => 
                           OTMP_6_41_port, B(40) => OTMP_6_40_port, B(39) => 
                           OTMP_6_39_port, B(38) => OTMP_6_38_port, B(37) => 
                           OTMP_6_37_port, B(36) => OTMP_6_36_port, B(35) => 
                           OTMP_6_35_port, B(34) => OTMP_6_34_port, B(33) => 
                           OTMP_6_33_port, B(32) => OTMP_6_32_port, B(31) => 
                           OTMP_6_31_port, B(30) => OTMP_6_30_port, B(29) => 
                           OTMP_6_29_port, B(28) => OTMP_6_28_port, B(27) => 
                           OTMP_6_27_port, B(26) => OTMP_6_26_port, B(25) => 
                           OTMP_6_25_port, B(24) => OTMP_6_24_port, B(23) => 
                           OTMP_6_23_port, B(22) => OTMP_6_22_port, B(21) => 
                           OTMP_6_21_port, B(20) => OTMP_6_20_port, B(19) => 
                           OTMP_6_19_port, B(18) => OTMP_6_18_port, B(17) => 
                           OTMP_6_17_port, B(16) => OTMP_6_16_port, B(15) => 
                           OTMP_6_15_port, B(14) => OTMP_6_14_port, B(13) => 
                           OTMP_6_13_port, B(12) => OTMP_6_12_port, B(11) => 
                           OTMP_6_11_port, B(10) => OTMP_6_10_port, B(9) => 
                           OTMP_6_9_port, B(8) => OTMP_6_8_port, B(7) => 
                           OTMP_6_7_port, B(6) => OTMP_6_6_port, B(5) => 
                           OTMP_6_5_port, B(4) => OTMP_6_4_port, B(3) => 
                           OTMP_6_3_port, B(2) => OTMP_6_2_port, B(1) => 
                           OTMP_6_1_port, B(0) => OTMP_6_0_port, Ci => 
                           X_Logic0_port, S(45) => PTMP_5_45_port, S(44) => 
                           PTMP_5_44_port, S(43) => PTMP_5_43_port, S(42) => 
                           PTMP_5_42_port, S(41) => PTMP_5_41_port, S(40) => 
                           PTMP_5_40_port, S(39) => PTMP_5_39_port, S(38) => 
                           PTMP_5_38_port, S(37) => PTMP_5_37_port, S(36) => 
                           PTMP_5_36_port, S(35) => PTMP_5_35_port, S(34) => 
                           PTMP_5_34_port, S(33) => PTMP_5_33_port, S(32) => 
                           PTMP_5_32_port, S(31) => PTMP_5_31_port, S(30) => 
                           PTMP_5_30_port, S(29) => PTMP_5_29_port, S(28) => 
                           PTMP_5_28_port, S(27) => PTMP_5_27_port, S(26) => 
                           PTMP_5_26_port, S(25) => PTMP_5_25_port, S(24) => 
                           PTMP_5_24_port, S(23) => PTMP_5_23_port, S(22) => 
                           PTMP_5_22_port, S(21) => PTMP_5_21_port, S(20) => 
                           PTMP_5_20_port, S(19) => PTMP_5_19_port, S(18) => 
                           PTMP_5_18_port, S(17) => PTMP_5_17_port, S(16) => 
                           PTMP_5_16_port, S(15) => PTMP_5_15_port, S(14) => 
                           PTMP_5_14_port, S(13) => PTMP_5_13_port, S(12) => 
                           PTMP_5_12_port, S(11) => PTMP_5_11_port, S(10) => 
                           PTMP_5_10_port, S(9) => PTMP_5_9_port, S(8) => 
                           PTMP_5_8_port, S(7) => PTMP_5_7_port, S(6) => 
                           PTMP_5_6_port, S(5) => PTMP_5_5_port, S(4) => 
                           PTMP_5_4_port, S(3) => PTMP_5_3_port, S(2) => 
                           PTMP_5_2_port, S(1) => PTMP_5_1_port, S(0) => 
                           PTMP_5_0_port, Co => n_1286);
   ADDER_7 : RCA_NBIT48 port map( A(47) => n14, A(46) => n14, A(45) => 
                           PTMP_5_45_port, A(44) => PTMP_5_44_port, A(43) => 
                           PTMP_5_43_port, A(42) => PTMP_5_42_port, A(41) => 
                           PTMP_5_41_port, A(40) => PTMP_5_40_port, A(39) => 
                           PTMP_5_39_port, A(38) => PTMP_5_38_port, A(37) => 
                           PTMP_5_37_port, A(36) => PTMP_5_36_port, A(35) => 
                           PTMP_5_35_port, A(34) => PTMP_5_34_port, A(33) => 
                           PTMP_5_33_port, A(32) => PTMP_5_32_port, A(31) => 
                           PTMP_5_31_port, A(30) => PTMP_5_30_port, A(29) => 
                           PTMP_5_29_port, A(28) => PTMP_5_28_port, A(27) => 
                           PTMP_5_27_port, A(26) => PTMP_5_26_port, A(25) => 
                           PTMP_5_25_port, A(24) => PTMP_5_24_port, A(23) => 
                           PTMP_5_23_port, A(22) => PTMP_5_22_port, A(21) => 
                           PTMP_5_21_port, A(20) => PTMP_5_20_port, A(19) => 
                           PTMP_5_19_port, A(18) => PTMP_5_18_port, A(17) => 
                           PTMP_5_17_port, A(16) => PTMP_5_16_port, A(15) => 
                           PTMP_5_15_port, A(14) => PTMP_5_14_port, A(13) => 
                           PTMP_5_13_port, A(12) => PTMP_5_12_port, A(11) => 
                           PTMP_5_11_port, A(10) => PTMP_5_10_port, A(9) => 
                           PTMP_5_9_port, A(8) => PTMP_5_8_port, A(7) => 
                           PTMP_5_7_port, A(6) => PTMP_5_6_port, A(5) => 
                           PTMP_5_5_port, A(4) => PTMP_5_4_port, A(3) => 
                           PTMP_5_3_port, A(2) => PTMP_5_2_port, A(1) => 
                           PTMP_5_1_port, A(0) => PTMP_5_0_port, B(47) => 
                           OTMP_7_47_port, B(46) => OTMP_7_46_port, B(45) => 
                           OTMP_7_45_port, B(44) => OTMP_7_44_port, B(43) => 
                           OTMP_7_43_port, B(42) => OTMP_7_42_port, B(41) => 
                           OTMP_7_41_port, B(40) => OTMP_7_40_port, B(39) => 
                           OTMP_7_39_port, B(38) => OTMP_7_38_port, B(37) => 
                           OTMP_7_37_port, B(36) => OTMP_7_36_port, B(35) => 
                           OTMP_7_35_port, B(34) => OTMP_7_34_port, B(33) => 
                           OTMP_7_33_port, B(32) => OTMP_7_32_port, B(31) => 
                           OTMP_7_31_port, B(30) => OTMP_7_30_port, B(29) => 
                           OTMP_7_29_port, B(28) => OTMP_7_28_port, B(27) => 
                           OTMP_7_27_port, B(26) => OTMP_7_26_port, B(25) => 
                           OTMP_7_25_port, B(24) => OTMP_7_24_port, B(23) => 
                           OTMP_7_23_port, B(22) => OTMP_7_22_port, B(21) => 
                           OTMP_7_21_port, B(20) => OTMP_7_20_port, B(19) => 
                           OTMP_7_19_port, B(18) => OTMP_7_18_port, B(17) => 
                           OTMP_7_17_port, B(16) => OTMP_7_16_port, B(15) => 
                           OTMP_7_15_port, B(14) => OTMP_7_14_port, B(13) => 
                           OTMP_7_13_port, B(12) => OTMP_7_12_port, B(11) => 
                           OTMP_7_11_port, B(10) => OTMP_7_10_port, B(9) => 
                           OTMP_7_9_port, B(8) => OTMP_7_8_port, B(7) => 
                           OTMP_7_7_port, B(6) => OTMP_7_6_port, B(5) => 
                           OTMP_7_5_port, B(4) => OTMP_7_4_port, B(3) => 
                           OTMP_7_3_port, B(2) => OTMP_7_2_port, B(1) => 
                           OTMP_7_1_port, B(0) => OTMP_7_0_port, Ci => 
                           X_Logic0_port, S(47) => PTMP_6_47_port, S(46) => 
                           PTMP_6_46_port, S(45) => PTMP_6_45_port, S(44) => 
                           PTMP_6_44_port, S(43) => PTMP_6_43_port, S(42) => 
                           PTMP_6_42_port, S(41) => PTMP_6_41_port, S(40) => 
                           PTMP_6_40_port, S(39) => PTMP_6_39_port, S(38) => 
                           PTMP_6_38_port, S(37) => PTMP_6_37_port, S(36) => 
                           PTMP_6_36_port, S(35) => PTMP_6_35_port, S(34) => 
                           PTMP_6_34_port, S(33) => PTMP_6_33_port, S(32) => 
                           PTMP_6_32_port, S(31) => PTMP_6_31_port, S(30) => 
                           PTMP_6_30_port, S(29) => PTMP_6_29_port, S(28) => 
                           PTMP_6_28_port, S(27) => PTMP_6_27_port, S(26) => 
                           PTMP_6_26_port, S(25) => PTMP_6_25_port, S(24) => 
                           PTMP_6_24_port, S(23) => PTMP_6_23_port, S(22) => 
                           PTMP_6_22_port, S(21) => PTMP_6_21_port, S(20) => 
                           PTMP_6_20_port, S(19) => PTMP_6_19_port, S(18) => 
                           PTMP_6_18_port, S(17) => PTMP_6_17_port, S(16) => 
                           PTMP_6_16_port, S(15) => PTMP_6_15_port, S(14) => 
                           PTMP_6_14_port, S(13) => PTMP_6_13_port, S(12) => 
                           PTMP_6_12_port, S(11) => PTMP_6_11_port, S(10) => 
                           PTMP_6_10_port, S(9) => PTMP_6_9_port, S(8) => 
                           PTMP_6_8_port, S(7) => PTMP_6_7_port, S(6) => 
                           PTMP_6_6_port, S(5) => PTMP_6_5_port, S(4) => 
                           PTMP_6_4_port, S(3) => PTMP_6_3_port, S(2) => 
                           PTMP_6_2_port, S(1) => PTMP_6_1_port, S(0) => 
                           PTMP_6_0_port, Co => n_1287);
   ADDER_8 : RCA_NBIT50 port map( A(49) => n17, A(48) => n17, A(47) => 
                           PTMP_6_47_port, A(46) => PTMP_6_46_port, A(45) => 
                           PTMP_6_45_port, A(44) => PTMP_6_44_port, A(43) => 
                           PTMP_6_43_port, A(42) => PTMP_6_42_port, A(41) => 
                           PTMP_6_41_port, A(40) => PTMP_6_40_port, A(39) => 
                           PTMP_6_39_port, A(38) => PTMP_6_38_port, A(37) => 
                           PTMP_6_37_port, A(36) => PTMP_6_36_port, A(35) => 
                           PTMP_6_35_port, A(34) => PTMP_6_34_port, A(33) => 
                           PTMP_6_33_port, A(32) => PTMP_6_32_port, A(31) => 
                           PTMP_6_31_port, A(30) => PTMP_6_30_port, A(29) => 
                           PTMP_6_29_port, A(28) => PTMP_6_28_port, A(27) => 
                           PTMP_6_27_port, A(26) => PTMP_6_26_port, A(25) => 
                           PTMP_6_25_port, A(24) => PTMP_6_24_port, A(23) => 
                           PTMP_6_23_port, A(22) => PTMP_6_22_port, A(21) => 
                           PTMP_6_21_port, A(20) => PTMP_6_20_port, A(19) => 
                           PTMP_6_19_port, A(18) => PTMP_6_18_port, A(17) => 
                           PTMP_6_17_port, A(16) => PTMP_6_16_port, A(15) => 
                           PTMP_6_15_port, A(14) => PTMP_6_14_port, A(13) => 
                           PTMP_6_13_port, A(12) => PTMP_6_12_port, A(11) => 
                           PTMP_6_11_port, A(10) => PTMP_6_10_port, A(9) => 
                           PTMP_6_9_port, A(8) => PTMP_6_8_port, A(7) => 
                           PTMP_6_7_port, A(6) => PTMP_6_6_port, A(5) => 
                           PTMP_6_5_port, A(4) => PTMP_6_4_port, A(3) => 
                           PTMP_6_3_port, A(2) => PTMP_6_2_port, A(1) => 
                           PTMP_6_1_port, A(0) => PTMP_6_0_port, B(49) => 
                           OTMP_8_49_port, B(48) => OTMP_8_48_port, B(47) => 
                           OTMP_8_47_port, B(46) => OTMP_8_46_port, B(45) => 
                           OTMP_8_45_port, B(44) => OTMP_8_44_port, B(43) => 
                           OTMP_8_43_port, B(42) => OTMP_8_42_port, B(41) => 
                           OTMP_8_41_port, B(40) => OTMP_8_40_port, B(39) => 
                           OTMP_8_39_port, B(38) => OTMP_8_38_port, B(37) => 
                           OTMP_8_37_port, B(36) => OTMP_8_36_port, B(35) => 
                           OTMP_8_35_port, B(34) => OTMP_8_34_port, B(33) => 
                           OTMP_8_33_port, B(32) => OTMP_8_32_port, B(31) => 
                           OTMP_8_31_port, B(30) => OTMP_8_30_port, B(29) => 
                           OTMP_8_29_port, B(28) => OTMP_8_28_port, B(27) => 
                           OTMP_8_27_port, B(26) => OTMP_8_26_port, B(25) => 
                           OTMP_8_25_port, B(24) => OTMP_8_24_port, B(23) => 
                           OTMP_8_23_port, B(22) => OTMP_8_22_port, B(21) => 
                           OTMP_8_21_port, B(20) => OTMP_8_20_port, B(19) => 
                           OTMP_8_19_port, B(18) => OTMP_8_18_port, B(17) => 
                           OTMP_8_17_port, B(16) => OTMP_8_16_port, B(15) => 
                           OTMP_8_15_port, B(14) => OTMP_8_14_port, B(13) => 
                           OTMP_8_13_port, B(12) => OTMP_8_12_port, B(11) => 
                           OTMP_8_11_port, B(10) => OTMP_8_10_port, B(9) => 
                           OTMP_8_9_port, B(8) => OTMP_8_8_port, B(7) => 
                           OTMP_8_7_port, B(6) => OTMP_8_6_port, B(5) => 
                           OTMP_8_5_port, B(4) => OTMP_8_4_port, B(3) => 
                           OTMP_8_3_port, B(2) => OTMP_8_2_port, B(1) => 
                           OTMP_8_1_port, B(0) => OTMP_8_0_port, Ci => 
                           X_Logic0_port, S(49) => PTMP_7_49_port, S(48) => 
                           PTMP_7_48_port, S(47) => PTMP_7_47_port, S(46) => 
                           PTMP_7_46_port, S(45) => PTMP_7_45_port, S(44) => 
                           PTMP_7_44_port, S(43) => PTMP_7_43_port, S(42) => 
                           PTMP_7_42_port, S(41) => PTMP_7_41_port, S(40) => 
                           PTMP_7_40_port, S(39) => PTMP_7_39_port, S(38) => 
                           PTMP_7_38_port, S(37) => PTMP_7_37_port, S(36) => 
                           PTMP_7_36_port, S(35) => PTMP_7_35_port, S(34) => 
                           PTMP_7_34_port, S(33) => PTMP_7_33_port, S(32) => 
                           PTMP_7_32_port, S(31) => PTMP_7_31_port, S(30) => 
                           PTMP_7_30_port, S(29) => PTMP_7_29_port, S(28) => 
                           PTMP_7_28_port, S(27) => PTMP_7_27_port, S(26) => 
                           PTMP_7_26_port, S(25) => PTMP_7_25_port, S(24) => 
                           PTMP_7_24_port, S(23) => PTMP_7_23_port, S(22) => 
                           PTMP_7_22_port, S(21) => PTMP_7_21_port, S(20) => 
                           PTMP_7_20_port, S(19) => PTMP_7_19_port, S(18) => 
                           PTMP_7_18_port, S(17) => PTMP_7_17_port, S(16) => 
                           PTMP_7_16_port, S(15) => PTMP_7_15_port, S(14) => 
                           PTMP_7_14_port, S(13) => PTMP_7_13_port, S(12) => 
                           PTMP_7_12_port, S(11) => PTMP_7_11_port, S(10) => 
                           PTMP_7_10_port, S(9) => PTMP_7_9_port, S(8) => 
                           PTMP_7_8_port, S(7) => PTMP_7_7_port, S(6) => 
                           PTMP_7_6_port, S(5) => PTMP_7_5_port, S(4) => 
                           PTMP_7_4_port, S(3) => PTMP_7_3_port, S(2) => 
                           PTMP_7_2_port, S(1) => PTMP_7_1_port, S(0) => 
                           PTMP_7_0_port, Co => n_1288);
   ADDER_9 : RCA_NBIT52 port map( A(51) => n16, A(50) => n16, A(49) => 
                           PTMP_7_49_port, A(48) => PTMP_7_48_port, A(47) => 
                           PTMP_7_47_port, A(46) => PTMP_7_46_port, A(45) => 
                           PTMP_7_45_port, A(44) => PTMP_7_44_port, A(43) => 
                           PTMP_7_43_port, A(42) => PTMP_7_42_port, A(41) => 
                           PTMP_7_41_port, A(40) => PTMP_7_40_port, A(39) => 
                           PTMP_7_39_port, A(38) => PTMP_7_38_port, A(37) => 
                           PTMP_7_37_port, A(36) => PTMP_7_36_port, A(35) => 
                           PTMP_7_35_port, A(34) => PTMP_7_34_port, A(33) => 
                           PTMP_7_33_port, A(32) => PTMP_7_32_port, A(31) => 
                           PTMP_7_31_port, A(30) => PTMP_7_30_port, A(29) => 
                           PTMP_7_29_port, A(28) => PTMP_7_28_port, A(27) => 
                           PTMP_7_27_port, A(26) => PTMP_7_26_port, A(25) => 
                           PTMP_7_25_port, A(24) => PTMP_7_24_port, A(23) => 
                           PTMP_7_23_port, A(22) => PTMP_7_22_port, A(21) => 
                           PTMP_7_21_port, A(20) => PTMP_7_20_port, A(19) => 
                           PTMP_7_19_port, A(18) => PTMP_7_18_port, A(17) => 
                           PTMP_7_17_port, A(16) => PTMP_7_16_port, A(15) => 
                           PTMP_7_15_port, A(14) => PTMP_7_14_port, A(13) => 
                           PTMP_7_13_port, A(12) => PTMP_7_12_port, A(11) => 
                           PTMP_7_11_port, A(10) => PTMP_7_10_port, A(9) => 
                           PTMP_7_9_port, A(8) => PTMP_7_8_port, A(7) => 
                           PTMP_7_7_port, A(6) => PTMP_7_6_port, A(5) => 
                           PTMP_7_5_port, A(4) => PTMP_7_4_port, A(3) => 
                           PTMP_7_3_port, A(2) => PTMP_7_2_port, A(1) => 
                           PTMP_7_1_port, A(0) => PTMP_7_0_port, B(51) => 
                           OTMP_9_51_port, B(50) => OTMP_9_50_port, B(49) => 
                           OTMP_9_49_port, B(48) => OTMP_9_48_port, B(47) => 
                           OTMP_9_47_port, B(46) => OTMP_9_46_port, B(45) => 
                           OTMP_9_45_port, B(44) => OTMP_9_44_port, B(43) => 
                           OTMP_9_43_port, B(42) => OTMP_9_42_port, B(41) => 
                           OTMP_9_41_port, B(40) => OTMP_9_40_port, B(39) => 
                           OTMP_9_39_port, B(38) => OTMP_9_38_port, B(37) => 
                           OTMP_9_37_port, B(36) => OTMP_9_36_port, B(35) => 
                           OTMP_9_35_port, B(34) => OTMP_9_34_port, B(33) => 
                           OTMP_9_33_port, B(32) => OTMP_9_32_port, B(31) => 
                           OTMP_9_31_port, B(30) => OTMP_9_30_port, B(29) => 
                           OTMP_9_29_port, B(28) => OTMP_9_28_port, B(27) => 
                           OTMP_9_27_port, B(26) => OTMP_9_26_port, B(25) => 
                           OTMP_9_25_port, B(24) => OTMP_9_24_port, B(23) => 
                           OTMP_9_23_port, B(22) => OTMP_9_22_port, B(21) => 
                           OTMP_9_21_port, B(20) => OTMP_9_20_port, B(19) => 
                           OTMP_9_19_port, B(18) => OTMP_9_18_port, B(17) => 
                           OTMP_9_17_port, B(16) => OTMP_9_16_port, B(15) => 
                           OTMP_9_15_port, B(14) => OTMP_9_14_port, B(13) => 
                           OTMP_9_13_port, B(12) => OTMP_9_12_port, B(11) => 
                           OTMP_9_11_port, B(10) => OTMP_9_10_port, B(9) => 
                           OTMP_9_9_port, B(8) => OTMP_9_8_port, B(7) => 
                           OTMP_9_7_port, B(6) => OTMP_9_6_port, B(5) => 
                           OTMP_9_5_port, B(4) => OTMP_9_4_port, B(3) => 
                           OTMP_9_3_port, B(2) => OTMP_9_2_port, B(1) => 
                           OTMP_9_1_port, B(0) => OTMP_9_0_port, Ci => 
                           X_Logic0_port, S(51) => PTMP_8_51_port, S(50) => 
                           PTMP_8_50_port, S(49) => PTMP_8_49_port, S(48) => 
                           PTMP_8_48_port, S(47) => PTMP_8_47_port, S(46) => 
                           PTMP_8_46_port, S(45) => PTMP_8_45_port, S(44) => 
                           PTMP_8_44_port, S(43) => PTMP_8_43_port, S(42) => 
                           PTMP_8_42_port, S(41) => PTMP_8_41_port, S(40) => 
                           PTMP_8_40_port, S(39) => PTMP_8_39_port, S(38) => 
                           PTMP_8_38_port, S(37) => PTMP_8_37_port, S(36) => 
                           PTMP_8_36_port, S(35) => PTMP_8_35_port, S(34) => 
                           PTMP_8_34_port, S(33) => PTMP_8_33_port, S(32) => 
                           PTMP_8_32_port, S(31) => PTMP_8_31_port, S(30) => 
                           PTMP_8_30_port, S(29) => PTMP_8_29_port, S(28) => 
                           PTMP_8_28_port, S(27) => PTMP_8_27_port, S(26) => 
                           PTMP_8_26_port, S(25) => PTMP_8_25_port, S(24) => 
                           PTMP_8_24_port, S(23) => PTMP_8_23_port, S(22) => 
                           PTMP_8_22_port, S(21) => PTMP_8_21_port, S(20) => 
                           PTMP_8_20_port, S(19) => PTMP_8_19_port, S(18) => 
                           PTMP_8_18_port, S(17) => PTMP_8_17_port, S(16) => 
                           PTMP_8_16_port, S(15) => PTMP_8_15_port, S(14) => 
                           PTMP_8_14_port, S(13) => PTMP_8_13_port, S(12) => 
                           PTMP_8_12_port, S(11) => PTMP_8_11_port, S(10) => 
                           PTMP_8_10_port, S(9) => PTMP_8_9_port, S(8) => 
                           PTMP_8_8_port, S(7) => PTMP_8_7_port, S(6) => 
                           PTMP_8_6_port, S(5) => PTMP_8_5_port, S(4) => 
                           PTMP_8_4_port, S(3) => PTMP_8_3_port, S(2) => 
                           PTMP_8_2_port, S(1) => PTMP_8_1_port, S(0) => 
                           PTMP_8_0_port, Co => n_1289);
   ADDER_10 : RCA_NBIT54 port map( A(53) => n11, A(52) => n6, A(51) => 
                           PTMP_8_51_port, A(50) => PTMP_8_50_port, A(49) => 
                           PTMP_8_49_port, A(48) => PTMP_8_48_port, A(47) => 
                           PTMP_8_47_port, A(46) => PTMP_8_46_port, A(45) => 
                           PTMP_8_45_port, A(44) => PTMP_8_44_port, A(43) => 
                           PTMP_8_43_port, A(42) => PTMP_8_42_port, A(41) => 
                           PTMP_8_41_port, A(40) => PTMP_8_40_port, A(39) => 
                           PTMP_8_39_port, A(38) => PTMP_8_38_port, A(37) => 
                           PTMP_8_37_port, A(36) => PTMP_8_36_port, A(35) => 
                           PTMP_8_35_port, A(34) => PTMP_8_34_port, A(33) => 
                           PTMP_8_33_port, A(32) => PTMP_8_32_port, A(31) => 
                           PTMP_8_31_port, A(30) => PTMP_8_30_port, A(29) => 
                           PTMP_8_29_port, A(28) => PTMP_8_28_port, A(27) => 
                           PTMP_8_27_port, A(26) => PTMP_8_26_port, A(25) => 
                           PTMP_8_25_port, A(24) => PTMP_8_24_port, A(23) => 
                           PTMP_8_23_port, A(22) => PTMP_8_22_port, A(21) => 
                           PTMP_8_21_port, A(20) => PTMP_8_20_port, A(19) => 
                           PTMP_8_19_port, A(18) => PTMP_8_18_port, A(17) => 
                           PTMP_8_17_port, A(16) => PTMP_8_16_port, A(15) => 
                           PTMP_8_15_port, A(14) => PTMP_8_14_port, A(13) => 
                           PTMP_8_13_port, A(12) => PTMP_8_12_port, A(11) => 
                           PTMP_8_11_port, A(10) => PTMP_8_10_port, A(9) => 
                           PTMP_8_9_port, A(8) => PTMP_8_8_port, A(7) => 
                           PTMP_8_7_port, A(6) => PTMP_8_6_port, A(5) => 
                           PTMP_8_5_port, A(4) => PTMP_8_4_port, A(3) => 
                           PTMP_8_3_port, A(2) => PTMP_8_2_port, A(1) => 
                           PTMP_8_1_port, A(0) => PTMP_8_0_port, B(53) => 
                           OTMP_10_53_port, B(52) => OTMP_10_52_port, B(51) => 
                           OTMP_10_51_port, B(50) => OTMP_10_50_port, B(49) => 
                           OTMP_10_49_port, B(48) => OTMP_10_48_port, B(47) => 
                           OTMP_10_47_port, B(46) => OTMP_10_46_port, B(45) => 
                           OTMP_10_45_port, B(44) => OTMP_10_44_port, B(43) => 
                           OTMP_10_43_port, B(42) => OTMP_10_42_port, B(41) => 
                           OTMP_10_41_port, B(40) => OTMP_10_40_port, B(39) => 
                           OTMP_10_39_port, B(38) => OTMP_10_38_port, B(37) => 
                           OTMP_10_37_port, B(36) => OTMP_10_36_port, B(35) => 
                           OTMP_10_35_port, B(34) => OTMP_10_34_port, B(33) => 
                           OTMP_10_33_port, B(32) => OTMP_10_32_port, B(31) => 
                           OTMP_10_31_port, B(30) => OTMP_10_30_port, B(29) => 
                           OTMP_10_29_port, B(28) => OTMP_10_28_port, B(27) => 
                           OTMP_10_27_port, B(26) => OTMP_10_26_port, B(25) => 
                           OTMP_10_25_port, B(24) => OTMP_10_24_port, B(23) => 
                           OTMP_10_23_port, B(22) => OTMP_10_22_port, B(21) => 
                           OTMP_10_21_port, B(20) => OTMP_10_20_port, B(19) => 
                           OTMP_10_19_port, B(18) => OTMP_10_18_port, B(17) => 
                           OTMP_10_17_port, B(16) => OTMP_10_16_port, B(15) => 
                           OTMP_10_15_port, B(14) => OTMP_10_14_port, B(13) => 
                           OTMP_10_13_port, B(12) => OTMP_10_12_port, B(11) => 
                           OTMP_10_11_port, B(10) => OTMP_10_10_port, B(9) => 
                           OTMP_10_9_port, B(8) => OTMP_10_8_port, B(7) => 
                           OTMP_10_7_port, B(6) => OTMP_10_6_port, B(5) => 
                           OTMP_10_5_port, B(4) => OTMP_10_4_port, B(3) => 
                           OTMP_10_3_port, B(2) => OTMP_10_2_port, B(1) => 
                           OTMP_10_1_port, B(0) => OTMP_10_0_port, Ci => 
                           X_Logic0_port, S(53) => PTMP_9_53_port, S(52) => 
                           PTMP_9_52_port, S(51) => PTMP_9_51_port, S(50) => 
                           PTMP_9_50_port, S(49) => PTMP_9_49_port, S(48) => 
                           PTMP_9_48_port, S(47) => PTMP_9_47_port, S(46) => 
                           PTMP_9_46_port, S(45) => PTMP_9_45_port, S(44) => 
                           PTMP_9_44_port, S(43) => PTMP_9_43_port, S(42) => 
                           PTMP_9_42_port, S(41) => PTMP_9_41_port, S(40) => 
                           PTMP_9_40_port, S(39) => PTMP_9_39_port, S(38) => 
                           PTMP_9_38_port, S(37) => PTMP_9_37_port, S(36) => 
                           PTMP_9_36_port, S(35) => PTMP_9_35_port, S(34) => 
                           PTMP_9_34_port, S(33) => PTMP_9_33_port, S(32) => 
                           PTMP_9_32_port, S(31) => PTMP_9_31_port, S(30) => 
                           PTMP_9_30_port, S(29) => PTMP_9_29_port, S(28) => 
                           PTMP_9_28_port, S(27) => PTMP_9_27_port, S(26) => 
                           PTMP_9_26_port, S(25) => PTMP_9_25_port, S(24) => 
                           PTMP_9_24_port, S(23) => PTMP_9_23_port, S(22) => 
                           PTMP_9_22_port, S(21) => PTMP_9_21_port, S(20) => 
                           PTMP_9_20_port, S(19) => PTMP_9_19_port, S(18) => 
                           PTMP_9_18_port, S(17) => PTMP_9_17_port, S(16) => 
                           PTMP_9_16_port, S(15) => PTMP_9_15_port, S(14) => 
                           PTMP_9_14_port, S(13) => PTMP_9_13_port, S(12) => 
                           PTMP_9_12_port, S(11) => PTMP_9_11_port, S(10) => 
                           PTMP_9_10_port, S(9) => PTMP_9_9_port, S(8) => 
                           PTMP_9_8_port, S(7) => PTMP_9_7_port, S(6) => 
                           PTMP_9_6_port, S(5) => PTMP_9_5_port, S(4) => 
                           PTMP_9_4_port, S(3) => PTMP_9_3_port, S(2) => 
                           PTMP_9_2_port, S(1) => PTMP_9_1_port, S(0) => 
                           PTMP_9_0_port, Co => n_1290);
   ADDER_11 : RCA_NBIT56 port map( A(55) => PTMP_9_53_port, A(54) => n10, A(53)
                           => PTMP_9_53_port, A(52) => PTMP_9_52_port, A(51) =>
                           PTMP_9_51_port, A(50) => PTMP_9_50_port, A(49) => 
                           PTMP_9_49_port, A(48) => PTMP_9_48_port, A(47) => 
                           PTMP_9_47_port, A(46) => PTMP_9_46_port, A(45) => 
                           PTMP_9_45_port, A(44) => PTMP_9_44_port, A(43) => 
                           PTMP_9_43_port, A(42) => PTMP_9_42_port, A(41) => 
                           PTMP_9_41_port, A(40) => PTMP_9_40_port, A(39) => 
                           PTMP_9_39_port, A(38) => PTMP_9_38_port, A(37) => 
                           PTMP_9_37_port, A(36) => PTMP_9_36_port, A(35) => 
                           PTMP_9_35_port, A(34) => PTMP_9_34_port, A(33) => 
                           PTMP_9_33_port, A(32) => PTMP_9_32_port, A(31) => 
                           PTMP_9_31_port, A(30) => PTMP_9_30_port, A(29) => 
                           PTMP_9_29_port, A(28) => PTMP_9_28_port, A(27) => 
                           PTMP_9_27_port, A(26) => PTMP_9_26_port, A(25) => 
                           PTMP_9_25_port, A(24) => PTMP_9_24_port, A(23) => 
                           PTMP_9_23_port, A(22) => PTMP_9_22_port, A(21) => 
                           PTMP_9_21_port, A(20) => PTMP_9_20_port, A(19) => 
                           PTMP_9_19_port, A(18) => PTMP_9_18_port, A(17) => 
                           PTMP_9_17_port, A(16) => PTMP_9_16_port, A(15) => 
                           PTMP_9_15_port, A(14) => PTMP_9_14_port, A(13) => 
                           PTMP_9_13_port, A(12) => PTMP_9_12_port, A(11) => 
                           PTMP_9_11_port, A(10) => PTMP_9_10_port, A(9) => 
                           PTMP_9_9_port, A(8) => PTMP_9_8_port, A(7) => 
                           PTMP_9_7_port, A(6) => PTMP_9_6_port, A(5) => 
                           PTMP_9_5_port, A(4) => PTMP_9_4_port, A(3) => 
                           PTMP_9_3_port, A(2) => PTMP_9_2_port, A(1) => 
                           PTMP_9_1_port, A(0) => PTMP_9_0_port, B(55) => 
                           OTMP_11_55_port, B(54) => OTMP_11_54_port, B(53) => 
                           OTMP_11_53_port, B(52) => OTMP_11_52_port, B(51) => 
                           OTMP_11_51_port, B(50) => OTMP_11_50_port, B(49) => 
                           OTMP_11_49_port, B(48) => OTMP_11_48_port, B(47) => 
                           OTMP_11_47_port, B(46) => OTMP_11_46_port, B(45) => 
                           OTMP_11_45_port, B(44) => OTMP_11_44_port, B(43) => 
                           OTMP_11_43_port, B(42) => OTMP_11_42_port, B(41) => 
                           OTMP_11_41_port, B(40) => OTMP_11_40_port, B(39) => 
                           OTMP_11_39_port, B(38) => OTMP_11_38_port, B(37) => 
                           OTMP_11_37_port, B(36) => OTMP_11_36_port, B(35) => 
                           OTMP_11_35_port, B(34) => OTMP_11_34_port, B(33) => 
                           OTMP_11_33_port, B(32) => OTMP_11_32_port, B(31) => 
                           OTMP_11_31_port, B(30) => OTMP_11_30_port, B(29) => 
                           OTMP_11_29_port, B(28) => OTMP_11_28_port, B(27) => 
                           OTMP_11_27_port, B(26) => OTMP_11_26_port, B(25) => 
                           OTMP_11_25_port, B(24) => OTMP_11_24_port, B(23) => 
                           OTMP_11_23_port, B(22) => OTMP_11_22_port, B(21) => 
                           OTMP_11_21_port, B(20) => OTMP_11_20_port, B(19) => 
                           OTMP_11_19_port, B(18) => OTMP_11_18_port, B(17) => 
                           OTMP_11_17_port, B(16) => OTMP_11_16_port, B(15) => 
                           OTMP_11_15_port, B(14) => OTMP_11_14_port, B(13) => 
                           OTMP_11_13_port, B(12) => OTMP_11_12_port, B(11) => 
                           OTMP_11_11_port, B(10) => OTMP_11_10_port, B(9) => 
                           OTMP_11_9_port, B(8) => OTMP_11_8_port, B(7) => 
                           OTMP_11_7_port, B(6) => OTMP_11_6_port, B(5) => 
                           OTMP_11_5_port, B(4) => OTMP_11_4_port, B(3) => 
                           OTMP_11_3_port, B(2) => OTMP_11_2_port, B(1) => 
                           OTMP_11_1_port, B(0) => OTMP_11_0_port, Ci => 
                           X_Logic0_port, S(55) => PTMP_10_55_port, S(54) => 
                           PTMP_10_54_port, S(53) => PTMP_10_53_port, S(52) => 
                           PTMP_10_52_port, S(51) => PTMP_10_51_port, S(50) => 
                           PTMP_10_50_port, S(49) => PTMP_10_49_port, S(48) => 
                           PTMP_10_48_port, S(47) => PTMP_10_47_port, S(46) => 
                           PTMP_10_46_port, S(45) => PTMP_10_45_port, S(44) => 
                           PTMP_10_44_port, S(43) => PTMP_10_43_port, S(42) => 
                           PTMP_10_42_port, S(41) => PTMP_10_41_port, S(40) => 
                           PTMP_10_40_port, S(39) => PTMP_10_39_port, S(38) => 
                           PTMP_10_38_port, S(37) => PTMP_10_37_port, S(36) => 
                           PTMP_10_36_port, S(35) => PTMP_10_35_port, S(34) => 
                           PTMP_10_34_port, S(33) => PTMP_10_33_port, S(32) => 
                           PTMP_10_32_port, S(31) => PTMP_10_31_port, S(30) => 
                           PTMP_10_30_port, S(29) => PTMP_10_29_port, S(28) => 
                           PTMP_10_28_port, S(27) => PTMP_10_27_port, S(26) => 
                           PTMP_10_26_port, S(25) => PTMP_10_25_port, S(24) => 
                           PTMP_10_24_port, S(23) => PTMP_10_23_port, S(22) => 
                           PTMP_10_22_port, S(21) => PTMP_10_21_port, S(20) => 
                           PTMP_10_20_port, S(19) => PTMP_10_19_port, S(18) => 
                           PTMP_10_18_port, S(17) => PTMP_10_17_port, S(16) => 
                           PTMP_10_16_port, S(15) => PTMP_10_15_port, S(14) => 
                           PTMP_10_14_port, S(13) => PTMP_10_13_port, S(12) => 
                           PTMP_10_12_port, S(11) => PTMP_10_11_port, S(10) => 
                           PTMP_10_10_port, S(9) => PTMP_10_9_port, S(8) => 
                           PTMP_10_8_port, S(7) => PTMP_10_7_port, S(6) => 
                           PTMP_10_6_port, S(5) => PTMP_10_5_port, S(4) => 
                           PTMP_10_4_port, S(3) => PTMP_10_3_port, S(2) => 
                           PTMP_10_2_port, S(1) => PTMP_10_1_port, S(0) => 
                           PTMP_10_0_port, Co => n_1291);
   ADDER_12 : RCA_NBIT58 port map( A(57) => n15, A(56) => n15, A(55) => 
                           PTMP_10_55_port, A(54) => PTMP_10_54_port, A(53) => 
                           PTMP_10_53_port, A(52) => PTMP_10_52_port, A(51) => 
                           PTMP_10_51_port, A(50) => PTMP_10_50_port, A(49) => 
                           PTMP_10_49_port, A(48) => PTMP_10_48_port, A(47) => 
                           PTMP_10_47_port, A(46) => PTMP_10_46_port, A(45) => 
                           PTMP_10_45_port, A(44) => PTMP_10_44_port, A(43) => 
                           PTMP_10_43_port, A(42) => PTMP_10_42_port, A(41) => 
                           PTMP_10_41_port, A(40) => PTMP_10_40_port, A(39) => 
                           PTMP_10_39_port, A(38) => PTMP_10_38_port, A(37) => 
                           PTMP_10_37_port, A(36) => PTMP_10_36_port, A(35) => 
                           PTMP_10_35_port, A(34) => PTMP_10_34_port, A(33) => 
                           PTMP_10_33_port, A(32) => PTMP_10_32_port, A(31) => 
                           PTMP_10_31_port, A(30) => PTMP_10_30_port, A(29) => 
                           PTMP_10_29_port, A(28) => PTMP_10_28_port, A(27) => 
                           PTMP_10_27_port, A(26) => PTMP_10_26_port, A(25) => 
                           PTMP_10_25_port, A(24) => PTMP_10_24_port, A(23) => 
                           PTMP_10_23_port, A(22) => PTMP_10_22_port, A(21) => 
                           PTMP_10_21_port, A(20) => PTMP_10_20_port, A(19) => 
                           PTMP_10_19_port, A(18) => PTMP_10_18_port, A(17) => 
                           PTMP_10_17_port, A(16) => PTMP_10_16_port, A(15) => 
                           PTMP_10_15_port, A(14) => PTMP_10_14_port, A(13) => 
                           PTMP_10_13_port, A(12) => PTMP_10_12_port, A(11) => 
                           PTMP_10_11_port, A(10) => PTMP_10_10_port, A(9) => 
                           PTMP_10_9_port, A(8) => PTMP_10_8_port, A(7) => 
                           PTMP_10_7_port, A(6) => PTMP_10_6_port, A(5) => 
                           PTMP_10_5_port, A(4) => PTMP_10_4_port, A(3) => 
                           PTMP_10_3_port, A(2) => PTMP_10_2_port, A(1) => 
                           PTMP_10_1_port, A(0) => PTMP_10_0_port, B(57) => 
                           OTMP_12_57_port, B(56) => OTMP_12_56_port, B(55) => 
                           OTMP_12_55_port, B(54) => OTMP_12_54_port, B(53) => 
                           OTMP_12_53_port, B(52) => OTMP_12_52_port, B(51) => 
                           OTMP_12_51_port, B(50) => OTMP_12_50_port, B(49) => 
                           OTMP_12_49_port, B(48) => OTMP_12_48_port, B(47) => 
                           OTMP_12_47_port, B(46) => OTMP_12_46_port, B(45) => 
                           OTMP_12_45_port, B(44) => OTMP_12_44_port, B(43) => 
                           OTMP_12_43_port, B(42) => OTMP_12_42_port, B(41) => 
                           OTMP_12_41_port, B(40) => OTMP_12_40_port, B(39) => 
                           OTMP_12_39_port, B(38) => OTMP_12_38_port, B(37) => 
                           OTMP_12_37_port, B(36) => OTMP_12_36_port, B(35) => 
                           OTMP_12_35_port, B(34) => OTMP_12_34_port, B(33) => 
                           OTMP_12_33_port, B(32) => OTMP_12_32_port, B(31) => 
                           OTMP_12_31_port, B(30) => OTMP_12_30_port, B(29) => 
                           OTMP_12_29_port, B(28) => OTMP_12_28_port, B(27) => 
                           OTMP_12_27_port, B(26) => OTMP_12_26_port, B(25) => 
                           OTMP_12_25_port, B(24) => OTMP_12_24_port, B(23) => 
                           OTMP_12_23_port, B(22) => OTMP_12_22_port, B(21) => 
                           OTMP_12_21_port, B(20) => OTMP_12_20_port, B(19) => 
                           OTMP_12_19_port, B(18) => OTMP_12_18_port, B(17) => 
                           OTMP_12_17_port, B(16) => OTMP_12_16_port, B(15) => 
                           OTMP_12_15_port, B(14) => OTMP_12_14_port, B(13) => 
                           OTMP_12_13_port, B(12) => OTMP_12_12_port, B(11) => 
                           OTMP_12_11_port, B(10) => OTMP_12_10_port, B(9) => 
                           OTMP_12_9_port, B(8) => OTMP_12_8_port, B(7) => 
                           OTMP_12_7_port, B(6) => OTMP_12_6_port, B(5) => 
                           OTMP_12_5_port, B(4) => OTMP_12_4_port, B(3) => 
                           OTMP_12_3_port, B(2) => OTMP_12_2_port, B(1) => 
                           OTMP_12_1_port, B(0) => OTMP_12_0_port, Ci => 
                           X_Logic0_port, S(57) => PTMP_11_57_port, S(56) => 
                           PTMP_11_56_port, S(55) => PTMP_11_55_port, S(54) => 
                           PTMP_11_54_port, S(53) => PTMP_11_53_port, S(52) => 
                           PTMP_11_52_port, S(51) => PTMP_11_51_port, S(50) => 
                           PTMP_11_50_port, S(49) => PTMP_11_49_port, S(48) => 
                           PTMP_11_48_port, S(47) => PTMP_11_47_port, S(46) => 
                           PTMP_11_46_port, S(45) => PTMP_11_45_port, S(44) => 
                           PTMP_11_44_port, S(43) => PTMP_11_43_port, S(42) => 
                           PTMP_11_42_port, S(41) => PTMP_11_41_port, S(40) => 
                           PTMP_11_40_port, S(39) => PTMP_11_39_port, S(38) => 
                           PTMP_11_38_port, S(37) => PTMP_11_37_port, S(36) => 
                           PTMP_11_36_port, S(35) => PTMP_11_35_port, S(34) => 
                           PTMP_11_34_port, S(33) => PTMP_11_33_port, S(32) => 
                           PTMP_11_32_port, S(31) => PTMP_11_31_port, S(30) => 
                           PTMP_11_30_port, S(29) => PTMP_11_29_port, S(28) => 
                           PTMP_11_28_port, S(27) => PTMP_11_27_port, S(26) => 
                           PTMP_11_26_port, S(25) => PTMP_11_25_port, S(24) => 
                           PTMP_11_24_port, S(23) => PTMP_11_23_port, S(22) => 
                           PTMP_11_22_port, S(21) => PTMP_11_21_port, S(20) => 
                           PTMP_11_20_port, S(19) => PTMP_11_19_port, S(18) => 
                           PTMP_11_18_port, S(17) => PTMP_11_17_port, S(16) => 
                           PTMP_11_16_port, S(15) => PTMP_11_15_port, S(14) => 
                           PTMP_11_14_port, S(13) => PTMP_11_13_port, S(12) => 
                           PTMP_11_12_port, S(11) => PTMP_11_11_port, S(10) => 
                           PTMP_11_10_port, S(9) => PTMP_11_9_port, S(8) => 
                           PTMP_11_8_port, S(7) => PTMP_11_7_port, S(6) => 
                           PTMP_11_6_port, S(5) => PTMP_11_5_port, S(4) => 
                           PTMP_11_4_port, S(3) => PTMP_11_3_port, S(2) => 
                           PTMP_11_2_port, S(1) => PTMP_11_1_port, S(0) => 
                           PTMP_11_0_port, Co => n_1292);
   ADDER_13 : RCA_NBIT60 port map( A(59) => n18, A(58) => n18, A(57) => 
                           PTMP_11_57_port, A(56) => PTMP_11_56_port, A(55) => 
                           PTMP_11_55_port, A(54) => PTMP_11_54_port, A(53) => 
                           PTMP_11_53_port, A(52) => PTMP_11_52_port, A(51) => 
                           PTMP_11_51_port, A(50) => PTMP_11_50_port, A(49) => 
                           PTMP_11_49_port, A(48) => PTMP_11_48_port, A(47) => 
                           PTMP_11_47_port, A(46) => PTMP_11_46_port, A(45) => 
                           PTMP_11_45_port, A(44) => PTMP_11_44_port, A(43) => 
                           PTMP_11_43_port, A(42) => PTMP_11_42_port, A(41) => 
                           PTMP_11_41_port, A(40) => PTMP_11_40_port, A(39) => 
                           PTMP_11_39_port, A(38) => PTMP_11_38_port, A(37) => 
                           PTMP_11_37_port, A(36) => PTMP_11_36_port, A(35) => 
                           PTMP_11_35_port, A(34) => PTMP_11_34_port, A(33) => 
                           PTMP_11_33_port, A(32) => PTMP_11_32_port, A(31) => 
                           PTMP_11_31_port, A(30) => PTMP_11_30_port, A(29) => 
                           PTMP_11_29_port, A(28) => PTMP_11_28_port, A(27) => 
                           PTMP_11_27_port, A(26) => PTMP_11_26_port, A(25) => 
                           PTMP_11_25_port, A(24) => PTMP_11_24_port, A(23) => 
                           PTMP_11_23_port, A(22) => PTMP_11_22_port, A(21) => 
                           PTMP_11_21_port, A(20) => PTMP_11_20_port, A(19) => 
                           PTMP_11_19_port, A(18) => PTMP_11_18_port, A(17) => 
                           PTMP_11_17_port, A(16) => PTMP_11_16_port, A(15) => 
                           PTMP_11_15_port, A(14) => PTMP_11_14_port, A(13) => 
                           PTMP_11_13_port, A(12) => PTMP_11_12_port, A(11) => 
                           PTMP_11_11_port, A(10) => PTMP_11_10_port, A(9) => 
                           PTMP_11_9_port, A(8) => PTMP_11_8_port, A(7) => 
                           PTMP_11_7_port, A(6) => PTMP_11_6_port, A(5) => 
                           PTMP_11_5_port, A(4) => PTMP_11_4_port, A(3) => 
                           PTMP_11_3_port, A(2) => PTMP_11_2_port, A(1) => 
                           PTMP_11_1_port, A(0) => PTMP_11_0_port, B(59) => 
                           OTMP_13_59_port, B(58) => OTMP_13_58_port, B(57) => 
                           OTMP_13_57_port, B(56) => OTMP_13_56_port, B(55) => 
                           OTMP_13_55_port, B(54) => OTMP_13_54_port, B(53) => 
                           OTMP_13_53_port, B(52) => OTMP_13_52_port, B(51) => 
                           OTMP_13_51_port, B(50) => OTMP_13_50_port, B(49) => 
                           OTMP_13_49_port, B(48) => OTMP_13_48_port, B(47) => 
                           OTMP_13_47_port, B(46) => OTMP_13_46_port, B(45) => 
                           OTMP_13_45_port, B(44) => OTMP_13_44_port, B(43) => 
                           OTMP_13_43_port, B(42) => OTMP_13_42_port, B(41) => 
                           OTMP_13_41_port, B(40) => OTMP_13_40_port, B(39) => 
                           OTMP_13_39_port, B(38) => OTMP_13_38_port, B(37) => 
                           OTMP_13_37_port, B(36) => OTMP_13_36_port, B(35) => 
                           OTMP_13_35_port, B(34) => OTMP_13_34_port, B(33) => 
                           OTMP_13_33_port, B(32) => OTMP_13_32_port, B(31) => 
                           OTMP_13_31_port, B(30) => OTMP_13_30_port, B(29) => 
                           OTMP_13_29_port, B(28) => OTMP_13_28_port, B(27) => 
                           OTMP_13_27_port, B(26) => OTMP_13_26_port, B(25) => 
                           OTMP_13_25_port, B(24) => OTMP_13_24_port, B(23) => 
                           OTMP_13_23_port, B(22) => OTMP_13_22_port, B(21) => 
                           OTMP_13_21_port, B(20) => OTMP_13_20_port, B(19) => 
                           OTMP_13_19_port, B(18) => OTMP_13_18_port, B(17) => 
                           OTMP_13_17_port, B(16) => OTMP_13_16_port, B(15) => 
                           OTMP_13_15_port, B(14) => OTMP_13_14_port, B(13) => 
                           OTMP_13_13_port, B(12) => OTMP_13_12_port, B(11) => 
                           OTMP_13_11_port, B(10) => OTMP_13_10_port, B(9) => 
                           OTMP_13_9_port, B(8) => OTMP_13_8_port, B(7) => 
                           OTMP_13_7_port, B(6) => OTMP_13_6_port, B(5) => 
                           OTMP_13_5_port, B(4) => OTMP_13_4_port, B(3) => 
                           OTMP_13_3_port, B(2) => OTMP_13_2_port, B(1) => 
                           OTMP_13_1_port, B(0) => OTMP_13_0_port, Ci => 
                           X_Logic0_port, S(59) => PTMP_12_59_port, S(58) => 
                           PTMP_12_58_port, S(57) => PTMP_12_57_port, S(56) => 
                           PTMP_12_56_port, S(55) => PTMP_12_55_port, S(54) => 
                           PTMP_12_54_port, S(53) => PTMP_12_53_port, S(52) => 
                           PTMP_12_52_port, S(51) => PTMP_12_51_port, S(50) => 
                           PTMP_12_50_port, S(49) => PTMP_12_49_port, S(48) => 
                           PTMP_12_48_port, S(47) => PTMP_12_47_port, S(46) => 
                           PTMP_12_46_port, S(45) => PTMP_12_45_port, S(44) => 
                           PTMP_12_44_port, S(43) => PTMP_12_43_port, S(42) => 
                           PTMP_12_42_port, S(41) => PTMP_12_41_port, S(40) => 
                           PTMP_12_40_port, S(39) => PTMP_12_39_port, S(38) => 
                           PTMP_12_38_port, S(37) => PTMP_12_37_port, S(36) => 
                           PTMP_12_36_port, S(35) => PTMP_12_35_port, S(34) => 
                           PTMP_12_34_port, S(33) => PTMP_12_33_port, S(32) => 
                           PTMP_12_32_port, S(31) => PTMP_12_31_port, S(30) => 
                           PTMP_12_30_port, S(29) => PTMP_12_29_port, S(28) => 
                           PTMP_12_28_port, S(27) => PTMP_12_27_port, S(26) => 
                           PTMP_12_26_port, S(25) => PTMP_12_25_port, S(24) => 
                           PTMP_12_24_port, S(23) => PTMP_12_23_port, S(22) => 
                           PTMP_12_22_port, S(21) => PTMP_12_21_port, S(20) => 
                           PTMP_12_20_port, S(19) => PTMP_12_19_port, S(18) => 
                           PTMP_12_18_port, S(17) => PTMP_12_17_port, S(16) => 
                           PTMP_12_16_port, S(15) => PTMP_12_15_port, S(14) => 
                           PTMP_12_14_port, S(13) => PTMP_12_13_port, S(12) => 
                           PTMP_12_12_port, S(11) => PTMP_12_11_port, S(10) => 
                           PTMP_12_10_port, S(9) => PTMP_12_9_port, S(8) => 
                           PTMP_12_8_port, S(7) => PTMP_12_7_port, S(6) => 
                           PTMP_12_6_port, S(5) => PTMP_12_5_port, S(4) => 
                           PTMP_12_4_port, S(3) => PTMP_12_3_port, S(2) => 
                           PTMP_12_2_port, S(1) => PTMP_12_1_port, S(0) => 
                           PTMP_12_0_port, Co => n_1293);
   ADDER_14 : RCA_NBIT62 port map( A(61) => PTMP_12_59_port, A(60) => 
                           PTMP_12_59_port, A(59) => PTMP_12_59_port, A(58) => 
                           PTMP_12_58_port, A(57) => PTMP_12_57_port, A(56) => 
                           PTMP_12_56_port, A(55) => PTMP_12_55_port, A(54) => 
                           PTMP_12_54_port, A(53) => PTMP_12_53_port, A(52) => 
                           PTMP_12_52_port, A(51) => PTMP_12_51_port, A(50) => 
                           PTMP_12_50_port, A(49) => PTMP_12_49_port, A(48) => 
                           PTMP_12_48_port, A(47) => PTMP_12_47_port, A(46) => 
                           PTMP_12_46_port, A(45) => PTMP_12_45_port, A(44) => 
                           PTMP_12_44_port, A(43) => PTMP_12_43_port, A(42) => 
                           PTMP_12_42_port, A(41) => PTMP_12_41_port, A(40) => 
                           PTMP_12_40_port, A(39) => PTMP_12_39_port, A(38) => 
                           PTMP_12_38_port, A(37) => PTMP_12_37_port, A(36) => 
                           PTMP_12_36_port, A(35) => PTMP_12_35_port, A(34) => 
                           PTMP_12_34_port, A(33) => PTMP_12_33_port, A(32) => 
                           PTMP_12_32_port, A(31) => PTMP_12_31_port, A(30) => 
                           PTMP_12_30_port, A(29) => PTMP_12_29_port, A(28) => 
                           PTMP_12_28_port, A(27) => PTMP_12_27_port, A(26) => 
                           PTMP_12_26_port, A(25) => PTMP_12_25_port, A(24) => 
                           PTMP_12_24_port, A(23) => PTMP_12_23_port, A(22) => 
                           PTMP_12_22_port, A(21) => PTMP_12_21_port, A(20) => 
                           PTMP_12_20_port, A(19) => PTMP_12_19_port, A(18) => 
                           PTMP_12_18_port, A(17) => PTMP_12_17_port, A(16) => 
                           PTMP_12_16_port, A(15) => PTMP_12_15_port, A(14) => 
                           PTMP_12_14_port, A(13) => PTMP_12_13_port, A(12) => 
                           PTMP_12_12_port, A(11) => PTMP_12_11_port, A(10) => 
                           PTMP_12_10_port, A(9) => PTMP_12_9_port, A(8) => 
                           PTMP_12_8_port, A(7) => PTMP_12_7_port, A(6) => 
                           PTMP_12_6_port, A(5) => PTMP_12_5_port, A(4) => 
                           PTMP_12_4_port, A(3) => PTMP_12_3_port, A(2) => 
                           PTMP_12_2_port, A(1) => PTMP_12_1_port, A(0) => 
                           PTMP_12_0_port, B(61) => OTMP_14_61_port, B(60) => 
                           OTMP_14_60_port, B(59) => OTMP_14_59_port, B(58) => 
                           OTMP_14_58_port, B(57) => OTMP_14_57_port, B(56) => 
                           OTMP_14_56_port, B(55) => OTMP_14_55_port, B(54) => 
                           OTMP_14_54_port, B(53) => OTMP_14_53_port, B(52) => 
                           OTMP_14_52_port, B(51) => OTMP_14_51_port, B(50) => 
                           OTMP_14_50_port, B(49) => OTMP_14_49_port, B(48) => 
                           OTMP_14_48_port, B(47) => OTMP_14_47_port, B(46) => 
                           OTMP_14_46_port, B(45) => OTMP_14_45_port, B(44) => 
                           OTMP_14_44_port, B(43) => OTMP_14_43_port, B(42) => 
                           OTMP_14_42_port, B(41) => OTMP_14_41_port, B(40) => 
                           OTMP_14_40_port, B(39) => OTMP_14_39_port, B(38) => 
                           OTMP_14_38_port, B(37) => OTMP_14_37_port, B(36) => 
                           OTMP_14_36_port, B(35) => OTMP_14_35_port, B(34) => 
                           OTMP_14_34_port, B(33) => OTMP_14_33_port, B(32) => 
                           OTMP_14_32_port, B(31) => OTMP_14_31_port, B(30) => 
                           OTMP_14_30_port, B(29) => OTMP_14_29_port, B(28) => 
                           OTMP_14_28_port, B(27) => OTMP_14_27_port, B(26) => 
                           OTMP_14_26_port, B(25) => OTMP_14_25_port, B(24) => 
                           OTMP_14_24_port, B(23) => OTMP_14_23_port, B(22) => 
                           OTMP_14_22_port, B(21) => OTMP_14_21_port, B(20) => 
                           OTMP_14_20_port, B(19) => OTMP_14_19_port, B(18) => 
                           OTMP_14_18_port, B(17) => OTMP_14_17_port, B(16) => 
                           OTMP_14_16_port, B(15) => OTMP_14_15_port, B(14) => 
                           OTMP_14_14_port, B(13) => OTMP_14_13_port, B(12) => 
                           OTMP_14_12_port, B(11) => OTMP_14_11_port, B(10) => 
                           OTMP_14_10_port, B(9) => OTMP_14_9_port, B(8) => 
                           OTMP_14_8_port, B(7) => OTMP_14_7_port, B(6) => 
                           OTMP_14_6_port, B(5) => OTMP_14_5_port, B(4) => 
                           OTMP_14_4_port, B(3) => OTMP_14_3_port, B(2) => 
                           OTMP_14_2_port, B(1) => OTMP_14_1_port, B(0) => 
                           OTMP_14_0_port, Ci => X_Logic0_port, S(61) => 
                           PTMP_13_61_port, S(60) => PTMP_13_60_port, S(59) => 
                           PTMP_13_59_port, S(58) => PTMP_13_58_port, S(57) => 
                           PTMP_13_57_port, S(56) => PTMP_13_56_port, S(55) => 
                           PTMP_13_55_port, S(54) => PTMP_13_54_port, S(53) => 
                           PTMP_13_53_port, S(52) => PTMP_13_52_port, S(51) => 
                           PTMP_13_51_port, S(50) => PTMP_13_50_port, S(49) => 
                           PTMP_13_49_port, S(48) => PTMP_13_48_port, S(47) => 
                           PTMP_13_47_port, S(46) => PTMP_13_46_port, S(45) => 
                           PTMP_13_45_port, S(44) => PTMP_13_44_port, S(43) => 
                           PTMP_13_43_port, S(42) => PTMP_13_42_port, S(41) => 
                           PTMP_13_41_port, S(40) => PTMP_13_40_port, S(39) => 
                           PTMP_13_39_port, S(38) => PTMP_13_38_port, S(37) => 
                           PTMP_13_37_port, S(36) => PTMP_13_36_port, S(35) => 
                           PTMP_13_35_port, S(34) => PTMP_13_34_port, S(33) => 
                           PTMP_13_33_port, S(32) => PTMP_13_32_port, S(31) => 
                           PTMP_13_31_port, S(30) => PTMP_13_30_port, S(29) => 
                           PTMP_13_29_port, S(28) => PTMP_13_28_port, S(27) => 
                           PTMP_13_27_port, S(26) => PTMP_13_26_port, S(25) => 
                           PTMP_13_25_port, S(24) => PTMP_13_24_port, S(23) => 
                           PTMP_13_23_port, S(22) => PTMP_13_22_port, S(21) => 
                           PTMP_13_21_port, S(20) => PTMP_13_20_port, S(19) => 
                           PTMP_13_19_port, S(18) => PTMP_13_18_port, S(17) => 
                           PTMP_13_17_port, S(16) => PTMP_13_16_port, S(15) => 
                           PTMP_13_15_port, S(14) => PTMP_13_14_port, S(13) => 
                           PTMP_13_13_port, S(12) => PTMP_13_12_port, S(11) => 
                           PTMP_13_11_port, S(10) => PTMP_13_10_port, S(9) => 
                           PTMP_13_9_port, S(8) => PTMP_13_8_port, S(7) => 
                           PTMP_13_7_port, S(6) => PTMP_13_6_port, S(5) => 
                           PTMP_13_5_port, S(4) => PTMP_13_4_port, S(3) => 
                           PTMP_13_3_port, S(2) => PTMP_13_2_port, S(1) => 
                           PTMP_13_1_port, S(0) => PTMP_13_0_port, Co => n_1294
                           );
   ADDER_15 : RCA_NBIT64 port map( A(63) => n9, A(62) => n9, A(61) => 
                           PTMP_13_61_port, A(60) => PTMP_13_60_port, A(59) => 
                           PTMP_13_59_port, A(58) => PTMP_13_58_port, A(57) => 
                           PTMP_13_57_port, A(56) => PTMP_13_56_port, A(55) => 
                           PTMP_13_55_port, A(54) => PTMP_13_54_port, A(53) => 
                           PTMP_13_53_port, A(52) => PTMP_13_52_port, A(51) => 
                           PTMP_13_51_port, A(50) => PTMP_13_50_port, A(49) => 
                           PTMP_13_49_port, A(48) => PTMP_13_48_port, A(47) => 
                           PTMP_13_47_port, A(46) => PTMP_13_46_port, A(45) => 
                           PTMP_13_45_port, A(44) => PTMP_13_44_port, A(43) => 
                           PTMP_13_43_port, A(42) => PTMP_13_42_port, A(41) => 
                           PTMP_13_41_port, A(40) => PTMP_13_40_port, A(39) => 
                           PTMP_13_39_port, A(38) => PTMP_13_38_port, A(37) => 
                           PTMP_13_37_port, A(36) => PTMP_13_36_port, A(35) => 
                           PTMP_13_35_port, A(34) => PTMP_13_34_port, A(33) => 
                           PTMP_13_33_port, A(32) => PTMP_13_32_port, A(31) => 
                           PTMP_13_31_port, A(30) => PTMP_13_30_port, A(29) => 
                           PTMP_13_29_port, A(28) => PTMP_13_28_port, A(27) => 
                           PTMP_13_27_port, A(26) => PTMP_13_26_port, A(25) => 
                           PTMP_13_25_port, A(24) => PTMP_13_24_port, A(23) => 
                           PTMP_13_23_port, A(22) => PTMP_13_22_port, A(21) => 
                           PTMP_13_21_port, A(20) => PTMP_13_20_port, A(19) => 
                           PTMP_13_19_port, A(18) => PTMP_13_18_port, A(17) => 
                           PTMP_13_17_port, A(16) => PTMP_13_16_port, A(15) => 
                           PTMP_13_15_port, A(14) => PTMP_13_14_port, A(13) => 
                           PTMP_13_13_port, A(12) => PTMP_13_12_port, A(11) => 
                           PTMP_13_11_port, A(10) => PTMP_13_10_port, A(9) => 
                           PTMP_13_9_port, A(8) => PTMP_13_8_port, A(7) => 
                           PTMP_13_7_port, A(6) => PTMP_13_6_port, A(5) => 
                           PTMP_13_5_port, A(4) => PTMP_13_4_port, A(3) => 
                           PTMP_13_3_port, A(2) => PTMP_13_2_port, A(1) => 
                           PTMP_13_1_port, A(0) => PTMP_13_0_port, B(63) => 
                           OTMP_15_63_port, B(62) => OTMP_15_62_port, B(61) => 
                           OTMP_15_61_port, B(60) => OTMP_15_60_port, B(59) => 
                           OTMP_15_59_port, B(58) => OTMP_15_58_port, B(57) => 
                           OTMP_15_57_port, B(56) => OTMP_15_56_port, B(55) => 
                           OTMP_15_55_port, B(54) => OTMP_15_54_port, B(53) => 
                           OTMP_15_53_port, B(52) => OTMP_15_52_port, B(51) => 
                           OTMP_15_51_port, B(50) => OTMP_15_50_port, B(49) => 
                           OTMP_15_49_port, B(48) => OTMP_15_48_port, B(47) => 
                           OTMP_15_47_port, B(46) => OTMP_15_46_port, B(45) => 
                           OTMP_15_45_port, B(44) => OTMP_15_44_port, B(43) => 
                           OTMP_15_43_port, B(42) => OTMP_15_42_port, B(41) => 
                           OTMP_15_41_port, B(40) => OTMP_15_40_port, B(39) => 
                           OTMP_15_39_port, B(38) => OTMP_15_38_port, B(37) => 
                           OTMP_15_37_port, B(36) => OTMP_15_36_port, B(35) => 
                           OTMP_15_35_port, B(34) => OTMP_15_34_port, B(33) => 
                           OTMP_15_33_port, B(32) => OTMP_15_32_port, B(31) => 
                           OTMP_15_31_port, B(30) => OTMP_15_30_port, B(29) => 
                           OTMP_15_29_port, B(28) => OTMP_15_28_port, B(27) => 
                           OTMP_15_27_port, B(26) => OTMP_15_26_port, B(25) => 
                           OTMP_15_25_port, B(24) => OTMP_15_24_port, B(23) => 
                           OTMP_15_23_port, B(22) => OTMP_15_22_port, B(21) => 
                           OTMP_15_21_port, B(20) => OTMP_15_20_port, B(19) => 
                           OTMP_15_19_port, B(18) => OTMP_15_18_port, B(17) => 
                           OTMP_15_17_port, B(16) => OTMP_15_16_port, B(15) => 
                           OTMP_15_15_port, B(14) => OTMP_15_14_port, B(13) => 
                           OTMP_15_13_port, B(12) => OTMP_15_12_port, B(11) => 
                           OTMP_15_11_port, B(10) => OTMP_15_10_port, B(9) => 
                           OTMP_15_9_port, B(8) => OTMP_15_8_port, B(7) => 
                           OTMP_15_7_port, B(6) => OTMP_15_6_port, B(5) => 
                           OTMP_15_5_port, B(4) => OTMP_15_4_port, B(3) => 
                           OTMP_15_3_port, B(2) => OTMP_15_2_port, B(1) => 
                           OTMP_15_1_port, B(0) => OTMP_15_0_port, Ci => 
                           X_Logic0_port, S(63) => S(63), S(62) => S(62), S(61)
                           => S(61), S(60) => S(60), S(59) => S(59), S(58) => 
                           S(58), S(57) => S(57), S(56) => S(56), S(55) => 
                           S(55), S(54) => S(54), S(53) => S(53), S(52) => 
                           S(52), S(51) => S(51), S(50) => S(50), S(49) => 
                           S(49), S(48) => S(48), S(47) => S(47), S(46) => 
                           S(46), S(45) => S(45), S(44) => S(44), S(43) => 
                           S(43), S(42) => S(42), S(41) => S(41), S(40) => 
                           S(40), S(39) => S(39), S(38) => S(38), S(37) => 
                           S(37), S(36) => S(36), S(35) => S(35), S(34) => 
                           S(34), S(33) => S(33), S(32) => S(32), S(31) => 
                           S(31), S(30) => S(30), S(29) => S(29), S(28) => 
                           S(28), S(27) => S(27), S(26) => S(26), S(25) => 
                           S(25), S(24) => S(24), S(23) => S(23), S(22) => 
                           S(22), S(21) => S(21), S(20) => S(20), S(19) => 
                           S(19), S(18) => S(18), S(17) => S(17), S(16) => 
                           S(16), S(15) => S(15), S(14) => S(14), S(13) => 
                           S(13), S(12) => S(12), S(11) => S(11), S(10) => 
                           S(10), S(9) => S(9), S(8) => S(8), S(7) => S(7), 
                           S(6) => S(6), S(5) => S(5), S(4) => S(4), S(3) => 
                           S(3), S(2) => S(2), S(1) => S(1), S(0) => S(0), Co 
                           => n_1295);
   sub_101 : BOOTHMUL_NBIT32_DW01_sub_0 port map( A(31) => n4, A(30) => n4, 
                           A(29) => n4, A(28) => n4, A(27) => n4, A(26) => n4, 
                           A(25) => n4, A(24) => n4, A(23) => n4, A(22) => n4, 
                           A(21) => n4, A(20) => n4, A(19) => n4, A(18) => n4, 
                           A(17) => n4, A(16) => n4, A(15) => n4, A(14) => n4, 
                           A(13) => n4, A(12) => n4, A(11) => n4, A(10) => n4, 
                           A(9) => n4, A(8) => n4, A(7) => n4, A(6) => n4, A(5)
                           => n4, A(4) => n4, A(3) => n4, A(2) => n4, A(1) => 
                           n4, A(0) => n4, B(31) => A(31), B(30) => A(30), 
                           B(29) => A(29), B(28) => A(28), B(27) => A(27), 
                           B(26) => A(26), B(25) => A(25), B(24) => A(24), 
                           B(23) => A(23), B(22) => A(22), B(21) => A(21), 
                           B(20) => A(20), B(19) => A(19), B(18) => A(18), 
                           B(17) => A(17), B(16) => A(16), B(15) => A(15), 
                           B(14) => A(14), B(13) => A(13), B(12) => A(12), 
                           B(11) => A(11), B(10) => A(10), B(9) => A(9), B(8) 
                           => A(8), B(7) => A(7), B(6) => A(6), B(5) => A(5), 
                           B(4) => A(4), B(3) => A(3), B(2) => A(2), B(1) => 
                           A(1), B(0) => A(0), CI => n5, DIFF(31) => A_n_65, 
                           DIFF(30) => A_n_30_port, DIFF(29) => A_n_29_port, 
                           DIFF(28) => A_n_28_port, DIFF(27) => A_n_27_port, 
                           DIFF(26) => A_n_26_port, DIFF(25) => A_n_25_port, 
                           DIFF(24) => A_n_24_port, DIFF(23) => A_n_23_port, 
                           DIFF(22) => A_n_22_port, DIFF(21) => A_n_21_port, 
                           DIFF(20) => A_n_20_port, DIFF(19) => A_n_19_port, 
                           DIFF(18) => A_n_18_port, DIFF(17) => A_n_17_port, 
                           DIFF(16) => A_n_16_port, DIFF(15) => A_n_15_port, 
                           DIFF(14) => A_n_14_port, DIFF(13) => A_n_13_port, 
                           DIFF(12) => A_n_12_port, DIFF(11) => A_n_11_port, 
                           DIFF(10) => A_n_10_port, DIFF(9) => A_n_9_port, 
                           DIFF(8) => A_n_8_port, DIFF(7) => A_n_7_port, 
                           DIFF(6) => A_n_6_port, DIFF(5) => A_n_5_port, 
                           DIFF(4) => A_n_4_port, DIFF(3) => A_n_3_port, 
                           DIFF(2) => A_n_2_port, DIFF(1) => A_n_1_port, 
                           DIFF(0) => A_n_0_port, CO => n_1296);
   U80 : CLKBUF_X1 port map( A => PTMP_2_39_port, Z => n13);
   U81 : BUF_X1 port map( A => PTMP_5_45_port, Z => n14);
   U82 : BUF_X1 port map( A => PTMP_8_51_port, Z => n6);
   U83 : CLKBUF_X1 port map( A => PTMP_3_41_port, Z => n7);
   U84 : BUF_X1 port map( A => PTMP_13_61_port, Z => n9);
   U85 : BUF_X2 port map( A => A(1), Z => n8);
   U86 : CLKBUF_X1 port map( A => PTMP_9_53_port, Z => n10);
   U87 : CLKBUF_X1 port map( A => n6, Z => n11);
   U88 : CLKBUF_X1 port map( A => PTMP_4_43_port, Z => n12);
   U89 : CLKBUF_X1 port map( A => PTMP_10_55_port, Z => n15);
   U90 : CLKBUF_X1 port map( A => PTMP_7_49_port, Z => n16);
   U91 : CLKBUF_X1 port map( A => PTMP_6_47_port, Z => n17);
   U92 : CLKBUF_X1 port map( A => PTMP_11_57_port, Z => n18);
   U93 : BUF_X1 port map( A => SHIFT_3_37_port, Z => n19);

end SYN_BEHAVIOURAL;
