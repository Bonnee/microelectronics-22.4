
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_BOOTHMUL_NBIT32 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_BOOTHMUL_NBIT32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT64_DW01_add_0 is

   port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (63 downto 0);  CO : out std_logic);

end RCA_NBIT64_DW01_add_0;

architecture SYN_rpl of RCA_NBIT64_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_63_port, carry_62_port, carry_61_port, carry_60_port, 
      carry_59_port, carry_29_port, carry_28_port, carry_27_port, carry_26_port
      , carry_25_port, carry_24_port, carry_23_port, carry_22_port, 
      carry_21_port, carry_20_port, carry_19_port, carry_18_port, carry_17_port
      , carry_16_port, carry_15_port, carry_14_port, carry_13_port, 
      carry_12_port, carry_11_port, carry_10_port, carry_9_port, carry_8_port, 
      carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port, 
      carry_2_port, n1, net41892, net41964, net41962, net42392, net42403, 
      net42405, net43039, net43040, net42917, net44067, net44062, net44060, 
      net44055, net44024, net44094, net45334, net45410, net45412, net45417, 
      net45419, net45986, net47241, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, 
      n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27
      , n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, 
      n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56
      , n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, 
      n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85
      , n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, 
      n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, 
      n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, 
      n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, 
      n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, 
      n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, 
      n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, 
      n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, 
      n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, 
      n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, 
      n268 : std_logic;

begin
   
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : CLKBUF_X1 port map( A => n167, Z => n3);
   U3 : NOR2_X1 port map( A1 => n3, A2 => B(53), ZN => n4);
   U4 : CLKBUF_X1 port map( A => net45419, Z => n5);
   U5 : CLKBUF_X1 port map( A => A(34), Z => n6);
   U6 : CLKBUF_X1 port map( A => n233, Z => n7);
   U7 : CLKBUF_X1 port map( A => n217, Z => n8);
   U8 : CLKBUF_X1 port map( A => n235, Z => n9);
   U9 : CLKBUF_X1 port map( A => n216, Z => n10);
   U10 : NAND2_X1 port map( A1 => B(31), A2 => n225, ZN => n91);
   U11 : INV_X1 port map( A => A(30), ZN => n86);
   U12 : INV_X1 port map( A => A(35), ZN => n105);
   U13 : INV_X1 port map( A => A(36), ZN => n109);
   U14 : INV_X1 port map( A => A(39), ZN => n120);
   U15 : INV_X1 port map( A => A(43), ZN => n135);
   U16 : OAI21_X1 port map( B1 => n44, B2 => n45, A => n46, ZN => net44067);
   U17 : INV_X1 port map( A => n59, ZN => n44);
   U18 : NAND2_X1 port map( A1 => B(56), A2 => net44067, ZN => net44094);
   U19 : NAND2_X1 port map( A1 => n82, A2 => n83, ZN => n81);
   U20 : NAND2_X1 port map( A1 => B(29), A2 => A(29), ZN => n82);
   U21 : OAI21_X1 port map( B1 => A(29), B2 => B(29), A => carry_29_port, ZN =>
                           n83);
   U22 : NOR2_X1 port map( A1 => B(30), A2 => n81, ZN => n85);
   U23 : NAND2_X1 port map( A1 => B(30), A2 => n81, ZN => n87);
   U24 : XNOR2_X1 port map( A => A(29), B => n211, ZN => SUM(29));
   U25 : XNOR2_X1 port map( A => B(29), B => carry_29_port, ZN => n211);
   U26 : XNOR2_X1 port map( A => n210, B => n86, ZN => SUM(30));
   U27 : XNOR2_X1 port map( A => n81, B => n174, ZN => n210);
   U28 : INV_X1 port map( A => B(30), ZN => n174);
   U29 : XNOR2_X1 port map( A => n209, B => n90, ZN => SUM(31));
   U30 : XNOR2_X1 port map( A => n225, B => n175, ZN => n209);
   U31 : INV_X1 port map( A => B(31), ZN => n175);
   U32 : XNOR2_X1 port map( A => n208, B => n94, ZN => SUM(32));
   U33 : INV_X1 port map( A => B(32), ZN => n176);
   U34 : XNOR2_X1 port map( A => n63, B => n207, ZN => SUM(33));
   U35 : XNOR2_X1 port map( A => n205, B => n105, ZN => SUM(35));
   U36 : INV_X1 port map( A => B(35), ZN => n177);
   U37 : XNOR2_X1 port map( A => n204, B => n109, ZN => SUM(36));
   U38 : INV_X1 port map( A => B(36), ZN => n178);
   U39 : XNOR2_X1 port map( A => A(37), B => n203, ZN => SUM(37));
   U40 : XNOR2_X1 port map( A => B(37), B => n8, ZN => n203);
   U41 : XNOR2_X1 port map( A => n201, B => n120, ZN => SUM(39));
   U42 : INV_X1 port map( A => B(39), ZN => n179);
   U43 : INV_X1 port map( A => B(40), ZN => n180);
   U44 : XNOR2_X1 port map( A => B(41), B => n10, ZN => n199);
   U45 : XNOR2_X1 port map( A => n197, B => n135, ZN => SUM(43));
   U46 : INV_X1 port map( A => B(43), ZN => n181);
   U47 : XNOR2_X1 port map( A => n196, B => n139, ZN => SUM(44));
   U48 : INV_X1 port map( A => B(44), ZN => n182);
   U49 : XNOR2_X1 port map( A => B(45), B => n214, ZN => n195);
   U50 : XNOR2_X1 port map( A => n193, B => n150, ZN => SUM(47));
   U51 : INV_X1 port map( A => B(47), ZN => n183);
   U52 : INV_X1 port map( A => B(48), ZN => n184);
   U53 : XNOR2_X1 port map( A => B(49), B => n212, ZN => n191);
   U54 : XNOR2_X1 port map( A => net43040, B => n79, ZN => SUM(54));
   U55 : XNOR2_X1 port map( A => net44067, B => net44055, ZN => net41892);
   U56 : XNOR2_X1 port map( A => n78, B => n80, ZN => SUM(57));
   U57 : XNOR2_X1 port map( A => n200, B => n124, ZN => SUM(40));
   U58 : CLKBUF_X1 port map( A => n228, Z => n11);
   U59 : INV_X1 port map( A => A(44), ZN => n139);
   U60 : INV_X1 port map( A => B(56), ZN => net44055);
   U61 : CLKBUF_X1 port map( A => A(55), Z => n12);
   U62 : XNOR2_X1 port map( A => n253, B => n13, ZN => SUM(62));
   U63 : XNOR2_X1 port map( A => A(62), B => B(62), ZN => n13);
   U64 : XNOR2_X1 port map( A => n189, B => n165, ZN => SUM(51));
   U65 : INV_X1 port map( A => B(52), ZN => n186);
   U66 : INV_X1 port map( A => B(51), ZN => n185);
   U67 : INV_X1 port map( A => B(57), ZN => n52);
   U68 : OAI21_X1 port map( B1 => n98, B2 => n97, A => n99, ZN => n223);
   U69 : XNOR2_X1 port map( A => n192, B => n154, ZN => SUM(48));
   U70 : CLKBUF_X1 port map( A => n115, Z => n14);
   U71 : NOR2_X1 port map( A1 => B(47), A2 => n145, ZN => n15);
   U72 : NOR2_X1 port map( A1 => n107, A2 => B(37), ZN => n16);
   U73 : CLKBUF_X1 port map( A => n221, Z => n17);
   U74 : CLKBUF_X1 port map( A => A(42), Z => n18);
   U75 : NOR2_X1 port map( A1 => B(35), A2 => n100, ZN => n19);
   U76 : NOR2_X1 port map( A1 => B(32), A2 => n88, ZN => n20);
   U77 : CLKBUF_X1 port map( A => n231, Z => n21);
   U78 : INV_X1 port map( A => A(32), ZN => n94);
   U79 : CLKBUF_X1 port map( A => n222, Z => n22);
   U80 : NOR2_X1 port map( A1 => B(45), A2 => n137, ZN => n23);
   U81 : OAI21_X1 port map( B1 => n89, B2 => n90, A => n91, ZN => n24);
   U82 : CLKBUF_X1 port map( A => n155, Z => n25);
   U83 : XNOR2_X1 port map( A => n100, B => n177, ZN => n205);
   U84 : NOR2_X1 port map( A1 => B(31), A2 => n84, ZN => n89);
   U85 : INV_X1 port map( A => A(31), ZN => n90);
   U86 : CLKBUF_X1 port map( A => n56, Z => n39);
   U87 : CLKBUF_X1 port map( A => n234, Z => n26);
   U88 : NOR2_X1 port map( A1 => B(39), A2 => n115, ZN => n27);
   U89 : CLKBUF_X1 port map( A => n219, Z => n28);
   U90 : OAI21_X1 port map( B1 => B(54), B2 => net42917, A => A(54), ZN => n29)
                           ;
   U91 : CLKBUF_X1 port map( A => A(38), Z => n30);
   U92 : CLKBUF_X1 port map( A => n220, Z => n31);
   U93 : CLKBUF_X1 port map( A => A(50), Z => n32);
   U94 : OAI21_X1 port map( B1 => n169, B2 => n168, A => n170, ZN => n33);
   U95 : INV_X1 port map( A => A(40), ZN => n124);
   U96 : NOR2_X1 port map( A1 => B(49), A2 => n152, ZN => n34);
   U97 : INV_X1 port map( A => A(47), ZN => n150);
   U98 : XNOR2_X1 port map( A => n6, B => n206, ZN => SUM(34));
   U99 : INV_X1 port map( A => n172, ZN => n35);
   U100 : CLKBUF_X1 port map( A => n173, Z => n36);
   U101 : CLKBUF_X1 port map( A => n145, Z => n37);
   U102 : INV_X1 port map( A => A(48), ZN => n154);
   U103 : CLKBUF_X1 port map( A => n130, Z => n38);
   U104 : INV_X1 port map( A => A(37), ZN => n113);
   U105 : XNOR2_X1 port map( A => A(45), B => n195, ZN => SUM(45));
   U106 : XNOR2_X1 port map( A => n14, B => n179, ZN => n201);
   U107 : XNOR2_X1 port map( A => n30, B => n202, ZN => SUM(38));
   U108 : INV_X1 port map( A => A(51), ZN => n165);
   U109 : XNOR2_X1 port map( A => n188, B => n169, ZN => SUM(52));
   U110 : CLKBUF_X1 port map( A => n160, Z => n40);
   U111 : INV_X1 port map( A => A(53), ZN => n41);
   U112 : NAND2_X1 port map( A1 => n117, A2 => n116, ZN => n115);
   U113 : XNOR2_X1 port map( A => n18, B => n198, ZN => SUM(42));
   U114 : OAI21_X1 port map( B1 => B(55), B2 => net44024, A => A(55), ZN => n43
                           );
   U115 : AND2_X1 port map( A1 => net44024, A2 => B(55), ZN => n56);
   U116 : OAI211_X1 port map( C1 => net45419, C2 => n58, A => n50, B => n52, ZN
                           => n51);
   U117 : NAND2_X1 port map( A1 => n60, A2 => n43, ZN => net45412);
   U118 : AOI21_X1 port map( B1 => net45419, B2 => n47, A => n57, ZN => 
                           net44062);
   U119 : INV_X1 port map( A => n51, ZN => net47241);
   U120 : NAND2_X1 port map( A1 => n56, A2 => B(56), ZN => n55);
   U121 : NAND2_X1 port map( A1 => n53, A2 => n49, ZN => n54);
   U122 : AND2_X1 port map( A1 => n54, A2 => n55, ZN => n50);
   U123 : NAND2_X1 port map( A1 => net45986, A2 => B(55), ZN => n42);
   U124 : XNOR2_X1 port map( A => n61, B => B(55), ZN => net44060);
   U125 : AND2_X1 port map( A1 => n55, A2 => n54, ZN => n47);
   U126 : AND2_X1 port map( A1 => n48, A2 => n43, ZN => n57);
   U127 : OR2_X1 port map( A1 => net44024, A2 => B(55), ZN => n53);
   U128 : INV_X1 port map( A => A(56), ZN => net45419);
   U129 : AND2_X1 port map( A1 => n42, A2 => net44055, ZN => n48);
   U130 : INV_X1 port map( A => n39, ZN => n46);
   U131 : AND2_X1 port map( A1 => n48, A2 => n43, ZN => n58);
   U132 : CLKBUF_X1 port map( A => n53, Z => n59);
   U133 : CLKBUF_X1 port map( A => n42, Z => n60);
   U134 : CLKBUF_X1 port map( A => net45986, Z => n61);
   U135 : AND2_X1 port map( A1 => B(56), A2 => A(55), ZN => n49);
   U136 : INV_X1 port map( A => n12, ZN => n45);
   U137 : CLKBUF_X1 port map( A => A(54), Z => n62);
   U138 : INV_X1 port map( A => A(45), ZN => n143);
   U139 : OAI21_X1 port map( B1 => B(38), B2 => n111, A => A(38), ZN => n117);
   U140 : NAND2_X1 port map( A1 => B(37), A2 => n217, ZN => n114);
   U141 : XNOR2_X1 port map( A => A(49), B => n191, ZN => SUM(49));
   U142 : INV_X1 port map( A => A(49), ZN => n158);
   U143 : XNOR2_X1 port map( A => A(41), B => n199, ZN => SUM(41));
   U144 : INV_X1 port map( A => A(41), ZN => n128);
   U145 : NAND2_X1 port map( A1 => B(41), A2 => n216, ZN => n129);
   U146 : INV_X1 port map( A => n98, ZN => n63);
   U147 : INV_X1 port map( A => A(33), ZN => n98);
   U148 : XNOR2_X1 port map( A => n40, B => n185, ZN => n189);
   U149 : XNOR2_X1 port map( A => n38, B => n181, ZN => n197);
   U150 : NAND2_X1 port map( A1 => n74, A2 => n29, ZN => net45986);
   U151 : XNOR2_X1 port map( A => B(54), B => n62, ZN => n79);
   U152 : XNOR2_X1 port map( A => n32, B => n190, ZN => SUM(50));
   U153 : XNOR2_X1 port map( A => n37, B => n183, ZN => n193);
   U154 : NAND2_X1 port map( A1 => n213, A2 => B(49), ZN => n159);
   U155 : NAND2_X1 port map( A1 => B(45), A2 => n215, ZN => n144);
   U156 : CLKBUF_X1 port map( A => n77, Z => n64);
   U157 : XNOR2_X1 port map( A => n35, B => n187, ZN => SUM(53));
   U158 : INV_X1 port map( A => A(53), ZN => n172);
   U159 : OAI21_X1 port map( B1 => n141, B2 => B(46), A => A(46), ZN => n147);
   U160 : XNOR2_X1 port map( A => A(46), B => n194, ZN => SUM(46));
   U161 : CLKBUF_X1 port map( A => A(57), Z => n65);
   U162 : OAI21_X1 port map( B1 => net47241, B2 => n76, A => n77, ZN => n66);
   U163 : CLKBUF_X1 port map( A => net47241, Z => net45417);
   U164 : INV_X1 port map( A => n5, ZN => net45410);
   U165 : NAND2_X1 port map( A1 => net43039, A2 => B(54), ZN => n74);
   U166 : OAI21_X1 port map( B1 => n156, B2 => B(50), A => A(50), ZN => n162);
   U167 : INV_X1 port map( A => net45410, ZN => net45334);
   U168 : OAI21_X1 port map( B1 => B(42), B2 => n126, A => A(42), ZN => n132);
   U169 : CLKBUF_X1 port map( A => n267, Z => n67);
   U170 : NOR2_X1 port map( A1 => net45412, A2 => B(56), ZN => n68);
   U171 : CLKBUF_X1 port map( A => A(58), Z => n71);
   U172 : CLKBUF_X1 port map( A => A(59), Z => n69);
   U173 : CLKBUF_X1 port map( A => A(60), Z => n70);
   U174 : OAI21_X1 port map( B1 => net45417, B2 => n76, A => n64, ZN => n72);
   U175 : OAI21_X1 port map( B1 => n76, B2 => net47241, A => n77, ZN => 
                           net42392);
   U176 : INV_X1 port map( A => A(52), ZN => n169);
   U177 : NAND2_X1 port map( A1 => n146, A2 => n147, ZN => n145);
   U178 : NAND2_X1 port map( A1 => n162, A2 => n161, ZN => n160);
   U179 : CLKBUF_X1 port map( A => n251, Z => n73);
   U180 : OAI21_X1 port map( B1 => n68, B2 => net45334, A => net44094, ZN => 
                           n80);
   U181 : NAND2_X1 port map( A1 => A(58), A2 => net42392, ZN => net41962);
   U182 : NAND2_X1 port map( A1 => n66, A2 => B(58), ZN => net41964);
   U183 : OAI21_X1 port map( B1 => net42917, B2 => B(54), A => A(54), ZN => n75
                           );
   U184 : NAND2_X1 port map( A1 => n74, A2 => n75, ZN => net44024);
   U185 : XNOR2_X1 port map( A => n12, B => net44060, ZN => SUM(55));
   U186 : XNOR2_X1 port map( A => n65, B => B(57), ZN => n78);
   U187 : INV_X1 port map( A => A(57), ZN => n76);
   U188 : NAND2_X1 port map( A1 => net44062, A2 => B(57), ZN => n77);
   U189 : NOR2_X1 port map( A1 => n167, A2 => B(53), ZN => n171);
   U190 : OAI21_X1 port map( B1 => n171, B2 => n41, A => n173, ZN => net42917);
   U191 : OAI21_X1 port map( B1 => n4, B2 => n172, A => n36, ZN => net43040);
   U192 : OAI21_X1 port map( B1 => n226, B2 => n172, A => n173, ZN => net43039)
                           ;
   U193 : NOR2_X1 port map( A1 => B(48), A2 => n235, ZN => n153);
   U194 : OAI21_X1 port map( B1 => n153, B2 => n154, A => n155, ZN => n152);
   U195 : OAI21_X1 port map( B1 => n26, B2 => n154, A => n25, ZN => n212);
   U196 : OAI21_X1 port map( B1 => n234, B2 => n154, A => n155, ZN => n213);
   U197 : NOR2_X1 port map( A1 => B(44), A2 => n229, ZN => n138);
   U198 : OAI21_X1 port map( B1 => n138, B2 => n139, A => n140, ZN => n137);
   U199 : OAI21_X1 port map( B1 => n11, B2 => n139, A => n140, ZN => n214);
   U200 : OAI21_X1 port map( B1 => n228, B2 => n139, A => n140, ZN => n215);
   U201 : NOR2_X1 port map( A1 => B(40), A2 => n231, ZN => n123);
   U202 : OAI21_X1 port map( B1 => n123, B2 => n124, A => n125, ZN => n122);
   U203 : OAI21_X1 port map( B1 => n230, B2 => n124, A => n125, ZN => n216);
   U204 : NOR2_X1 port map( A1 => n233, A2 => B(36), ZN => n108);
   U205 : OAI21_X1 port map( B1 => n108, B2 => n109, A => n110, ZN => n107);
   U206 : OAI21_X1 port map( B1 => n232, B2 => n109, A => n110, ZN => n217);
   U207 : OAI21_X1 port map( B1 => n93, B2 => n94, A => n95, ZN => n92);
   U208 : NAND2_X1 port map( A1 => B(33), A2 => n218, ZN => n99);
   U209 : XNOR2_X1 port map( A => B(33), B => n218, ZN => n207);
   U210 : NOR2_X1 port map( A1 => B(33), A2 => n92, ZN => n97);
   U211 : NOR2_X1 port map( A1 => B(32), A2 => n88, ZN => n93);
   U212 : OAI21_X1 port map( B1 => n20, B2 => n94, A => n95, ZN => n218);
   U213 : NOR2_X1 port map( A1 => n152, A2 => B(49), ZN => n157);
   U214 : OAI21_X1 port map( B1 => n157, B2 => n158, A => n159, ZN => n156);
   U215 : OAI21_X1 port map( B1 => n34, B2 => n158, A => n159, ZN => n219);
   U216 : XNOR2_X1 port map( A => B(50), B => n28, ZN => n190);
   U217 : NAND2_X1 port map( A1 => B(50), A2 => n219, ZN => n161);
   U218 : NOR2_X1 port map( A1 => n137, A2 => B(45), ZN => n142);
   U219 : OAI21_X1 port map( B1 => n142, B2 => n143, A => n144, ZN => n141);
   U220 : OAI21_X1 port map( B1 => n23, B2 => n143, A => n144, ZN => n220);
   U221 : XNOR2_X1 port map( A => B(46), B => n31, ZN => n194);
   U222 : NAND2_X1 port map( A1 => B(46), A2 => n220, ZN => n146);
   U223 : NOR2_X1 port map( A1 => B(41), A2 => n122, ZN => n127);
   U224 : OAI21_X1 port map( B1 => n127, B2 => n128, A => n129, ZN => n126);
   U225 : OAI21_X1 port map( B1 => n127, B2 => n128, A => n129, ZN => n221);
   U226 : XNOR2_X1 port map( A => B(42), B => n17, ZN => n198);
   U227 : NAND2_X1 port map( A1 => B(42), A2 => n221, ZN => n131);
   U228 : NOR2_X1 port map( A1 => B(37), A2 => n107, ZN => n112);
   U229 : OAI21_X1 port map( B1 => n112, B2 => n113, A => n114, ZN => n111);
   U230 : OAI21_X1 port map( B1 => n16, B2 => n113, A => n114, ZN => n222);
   U231 : XNOR2_X1 port map( A => B(38), B => n22, ZN => n202);
   U232 : NAND2_X1 port map( A1 => B(38), A2 => n222, ZN => n116);
   U233 : OAI21_X1 port map( B1 => n97, B2 => n98, A => n99, ZN => n96);
   U234 : NAND2_X1 port map( A1 => B(34), A2 => n223, ZN => n101);
   U235 : OAI21_X1 port map( B1 => B(34), B2 => n96, A => A(34), ZN => n102);
   U236 : XNOR2_X1 port map( A => B(34), B => n223, ZN => n206);
   U237 : OAI21_X1 port map( B1 => n164, B2 => n165, A => n166, ZN => n163);
   U238 : XNOR2_X1 port map( A => n236, B => n186, ZN => n188);
   U239 : NAND2_X1 port map( A1 => B(52), A2 => n224, ZN => n170);
   U240 : NOR2_X1 port map( A1 => n163, A2 => B(52), ZN => n168);
   U241 : NOR2_X1 port map( A1 => n160, A2 => B(51), ZN => n164);
   U242 : OAI21_X1 port map( B1 => n164, B2 => n165, A => n166, ZN => n224);
   U243 : OAI21_X1 port map( B1 => n85, B2 => n86, A => n87, ZN => n84);
   U244 : OAI21_X1 port map( B1 => n85, B2 => n86, A => n87, ZN => n225);
   U245 : NOR2_X1 port map( A1 => B(53), A2 => n167, ZN => n226);
   U246 : OAI21_X1 port map( B1 => n168, B2 => n169, A => n170, ZN => n167);
   U247 : NAND2_X1 port map( A1 => n33, A2 => B(53), ZN => n173);
   U248 : XNOR2_X1 port map( A => B(53), B => n227, ZN => n187);
   U249 : CLKBUF_X1 port map( A => n33, Z => n227);
   U250 : NOR2_X1 port map( A1 => B(44), A2 => n133, ZN => n228);
   U251 : OAI21_X1 port map( B1 => n134, B2 => n135, A => n136, ZN => n133);
   U252 : XNOR2_X1 port map( A => n229, B => n182, ZN => n196);
   U253 : NAND2_X1 port map( A1 => n133, A2 => B(44), ZN => n140);
   U254 : NOR2_X1 port map( A1 => B(43), A2 => n130, ZN => n134);
   U255 : OAI21_X1 port map( B1 => n237, B2 => n135, A => n136, ZN => n229);
   U256 : NOR2_X1 port map( A1 => n118, A2 => B(40), ZN => n230);
   U257 : OAI21_X1 port map( B1 => n27, B2 => n120, A => n121, ZN => n118);
   U258 : XNOR2_X1 port map( A => n21, B => n180, ZN => n200);
   U259 : NAND2_X1 port map( A1 => n118, A2 => B(40), ZN => n125);
   U260 : NOR2_X1 port map( A1 => B(39), A2 => n115, ZN => n119);
   U261 : OAI21_X1 port map( B1 => n119, B2 => n120, A => n121, ZN => n231);
   U262 : NOR2_X1 port map( A1 => B(36), A2 => n103, ZN => n232);
   U263 : OAI21_X1 port map( B1 => n104, B2 => n105, A => n106, ZN => n103);
   U264 : XNOR2_X1 port map( A => n7, B => n178, ZN => n204);
   U265 : NAND2_X1 port map( A1 => n103, A2 => B(36), ZN => n110);
   U266 : NOR2_X1 port map( A1 => B(35), A2 => n100, ZN => n104);
   U267 : OAI21_X1 port map( B1 => n19, B2 => n105, A => n106, ZN => n233);
   U268 : NOR2_X1 port map( A1 => B(48), A2 => n148, ZN => n234);
   U269 : OAI21_X1 port map( B1 => n15, B2 => n150, A => n151, ZN => n148);
   U270 : XNOR2_X1 port map( A => n9, B => n184, ZN => n192);
   U271 : NAND2_X1 port map( A1 => n148, A2 => B(48), ZN => n155);
   U272 : NOR2_X1 port map( A1 => B(47), A2 => n145, ZN => n149);
   U273 : OAI21_X1 port map( B1 => n149, B2 => n150, A => n151, ZN => n235);
   U274 : OAI21_X1 port map( B1 => n89, B2 => n90, A => n91, ZN => n88);
   U275 : XNOR2_X1 port map( A => n24, B => n176, ZN => n208);
   U276 : NAND2_X1 port map( A1 => B(32), A2 => n24, ZN => n95);
   U277 : NAND2_X1 port map( A1 => n160, A2 => B(51), ZN => n166);
   U278 : CLKBUF_X1 port map( A => n224, Z => n236);
   U279 : NAND2_X1 port map( A1 => n101, A2 => n102, ZN => n100);
   U280 : NAND2_X1 port map( A1 => n145, A2 => B(47), ZN => n151);
   U281 : NAND2_X1 port map( A1 => n130, A2 => B(43), ZN => n136);
   U282 : NAND2_X1 port map( A1 => B(39), A2 => n115, ZN => n121);
   U283 : NAND2_X1 port map( A1 => B(35), A2 => n100, ZN => n106);
   U284 : NAND2_X1 port map( A1 => n132, A2 => n131, ZN => n130);
   U285 : NOR2_X1 port map( A1 => B(43), A2 => n130, ZN => n237);
   U286 : CLKBUF_X1 port map( A => n242, Z => n238);
   U287 : CLKBUF_X1 port map( A => n260, Z => n239);
   U288 : NAND3_X1 port map( A1 => n260, A2 => n259, A3 => n261, ZN => n240);
   U289 : CLKBUF_X1 port map( A => n266, Z => n241);
   U290 : NAND2_X1 port map( A1 => carry_59_port, A2 => B(59), ZN => n242);
   U291 : CLKBUF_X1 port map( A => net41964, Z => net42405);
   U292 : CLKBUF_X1 port map( A => net41962, Z => net42403);
   U293 : CLKBUF_X1 port map( A => n261, Z => n243);
   U294 : CLKBUF_X1 port map( A => n249, Z => n244);
   U295 : NAND3_X1 port map( A1 => n266, A2 => n268, A3 => n267, ZN => n245);
   U296 : NAND3_X1 port map( A1 => n241, A2 => n238, A3 => n67, ZN => n246);
   U297 : NAND3_X1 port map( A1 => net41964, A2 => n251, A3 => net41962, ZN => 
                           n247);
   U298 : NAND3_X1 port map( A1 => net42403, A2 => net42405, A3 => n73, ZN => 
                           n248);
   U299 : NAND3_X1 port map( A1 => n257, A2 => n256, A3 => n255, ZN => n249);
   U300 : XOR2_X1 port map( A => n72, B => B(58), Z => n250);
   U301 : XOR2_X1 port map( A => n250, B => n71, Z => SUM(58));
   U302 : NAND2_X1 port map( A1 => A(58), A2 => B(58), ZN => n251);
   U303 : NAND3_X1 port map( A1 => n251, A2 => net41964, A3 => net41962, ZN => 
                           carry_59_port);
   U304 : XNOR2_X1 port map( A => carry_63_port, B => n252, ZN => SUM(63));
   U305 : XNOR2_X1 port map( A => A(63), B => B(63), ZN => n252);
   U306 : XOR2_X1 port map( A => net45410, B => net41892, Z => SUM(56));
   U307 : NAND3_X1 port map( A1 => n239, A2 => n243, A3 => n259, ZN => n253);
   U308 : XOR2_X1 port map( A => n70, B => B(60), Z => n254);
   U309 : XOR2_X1 port map( A => n254, B => n246, Z => SUM(60));
   U310 : NAND2_X1 port map( A1 => A(60), A2 => B(60), ZN => n255);
   U311 : NAND2_X1 port map( A1 => n245, A2 => A(60), ZN => n256);
   U312 : NAND2_X1 port map( A1 => carry_60_port, A2 => B(60), ZN => n257);
   U313 : NAND3_X1 port map( A1 => n257, A2 => n256, A3 => n255, ZN => 
                           carry_61_port);
   U314 : XOR2_X1 port map( A => A(61), B => B(61), Z => n258);
   U315 : XOR2_X1 port map( A => n258, B => n244, Z => SUM(61));
   U316 : NAND2_X1 port map( A1 => A(61), A2 => B(61), ZN => n259);
   U317 : NAND2_X1 port map( A1 => n249, A2 => A(61), ZN => n260);
   U318 : NAND2_X1 port map( A1 => carry_61_port, A2 => B(61), ZN => n261);
   U319 : NAND3_X1 port map( A1 => n260, A2 => n259, A3 => n261, ZN => 
                           carry_62_port);
   U320 : NAND2_X1 port map( A1 => n240, A2 => A(62), ZN => n262);
   U321 : NAND2_X1 port map( A1 => carry_62_port, A2 => B(62), ZN => n263);
   U322 : NAND2_X1 port map( A1 => A(62), A2 => B(62), ZN => n264);
   U323 : NAND3_X1 port map( A1 => n263, A2 => n262, A3 => n264, ZN => 
                           carry_63_port);
   U324 : XOR2_X1 port map( A => n248, B => B(59), Z => n265);
   U325 : XOR2_X1 port map( A => n69, B => n265, Z => SUM(59));
   U326 : NAND2_X1 port map( A1 => n247, A2 => A(59), ZN => n266);
   U327 : NAND2_X1 port map( A1 => A(59), A2 => B(59), ZN => n267);
   U328 : NAND2_X1 port map( A1 => carry_59_port, A2 => B(59), ZN => n268);
   U329 : NAND3_X1 port map( A1 => n242, A2 => n266, A3 => n267, ZN => 
                           carry_60_port);
   U330 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n1);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT62_DW01_add_0 is

   port( A, B : in std_logic_vector (61 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (61 downto 0);  CO : out std_logic);

end RCA_NBIT62_DW01_add_0;

architecture SYN_rpl of RCA_NBIT62_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_61_port, carry_60_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, n1, net42064, net42063, 
      net42400, net45316, net45173, net45328, net46053, net45261, net73769, 
      net44091, net42091, net42090, carry_59_port, carry_58_port, carry_57_port
      , n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18
      , n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, 
      n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47
      , n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, 
      n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76
      , n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, 
      n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104
      , n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
      n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, 
      n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, 
      n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, 
      n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, 
      n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, 
      n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, 
      n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, 
      n201, n202, n203, n204 : std_logic;

begin
   
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1_57 : FA_X1 port map( A => A(57), B => B(57), CI => carry_57_port, CO => 
                           carry_58_port, S => SUM(57));
   U1_58 : FA_X1 port map( A => A(58), B => B(58), CI => carry_58_port, CO => 
                           carry_59_port, S => SUM(58));
   U1 : INV_X1 port map( A => n85, ZN => n3);
   U3 : CLKBUF_X1 port map( A => n69, Z => n4);
   U4 : NAND2_X1 port map( A1 => n42, A2 => n41, ZN => n5);
   U5 : OAI21_X1 port map( B1 => B(42), B2 => n83, A => A(42), ZN => n6);
   U6 : INV_X1 port map( A => n71, ZN => n7);
   U7 : OAI21_X1 port map( B1 => n55, B2 => B(34), A => A(34), ZN => n8);
   U8 : NAND2_X1 port map( A1 => n8, A2 => n60, ZN => n9);
   U9 : INV_X1 port map( A => B(31), ZN => n134);
   U10 : INV_X1 port map( A => B(30), ZN => n133);
   U11 : INV_X1 port map( A => B(32), ZN => n135);
   U12 : INV_X1 port map( A => B(35), ZN => n136);
   U13 : INV_X1 port map( A => B(36), ZN => n137);
   U14 : INV_X1 port map( A => B(40), ZN => n139);
   U15 : INV_X1 port map( A => B(44), ZN => n141);
   U16 : INV_X1 port map( A => B(47), ZN => n142);
   U17 : INV_X1 port map( A => A(36), ZN => n68);
   U18 : INV_X1 port map( A => B(51), ZN => n144);
   U19 : INV_X1 port map( A => B(52), ZN => n145);
   U20 : NOR2_X1 port map( A1 => n195, A2 => B(31), ZN => n10);
   U21 : INV_X1 port map( A => B(39), ZN => n138);
   U22 : INV_X1 port map( A => B(48), ZN => n143);
   U23 : INV_X1 port map( A => B(43), ZN => n140);
   U24 : OAI211_X1 port map( C1 => n80, C2 => n81, A => n82, B => n11, ZN => 
                           n12);
   U25 : INV_X1 port map( A => B(41), ZN => n11);
   U26 : INV_X1 port map( A => n12, ZN => n84);
   U27 : OAI21_X1 port map( B1 => n53, B2 => n52, A => n54, ZN => n196);
   U28 : OAI21_X1 port map( B1 => n56, B2 => n57, A => n58, ZN => n17);
   U29 : OAI21_X1 port map( B1 => B(38), B2 => n4, A => A(38), ZN => n13);
   U30 : CLKBUF_X1 port map( A => A(29), Z => n14);
   U31 : NOR2_X1 port map( A1 => n108, A2 => B(49), ZN => n15);
   U32 : CLKBUF_X1 port map( A => A(38), Z => n16);
   U33 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => n18);
   U34 : XNOR2_X1 port map( A => n168, B => n53, ZN => SUM(32));
   U35 : XNOR2_X1 port map( A => n165, B => n64, ZN => SUM(35));
   U36 : XNOR2_X1 port map( A => n9, B => n136, ZN => n165);
   U37 : NOR2_X1 port map( A1 => B(35), A2 => n9, ZN => n19);
   U38 : CLKBUF_X1 port map( A => A(34), Z => n20);
   U39 : INV_X1 port map( A => A(31), ZN => n49);
   U40 : XNOR2_X1 port map( A => carry_59_port, B => net45328, ZN => SUM(59));
   U41 : NAND2_X1 port map( A1 => carry_59_port, A2 => B(59), ZN => net42064);
   U42 : NAND2_X1 port map( A1 => carry_59_port, A2 => A(59), ZN => net42063);
   U43 : NAND3_X1 port map( A1 => n21, A2 => net42090, A3 => net42091, ZN => 
                           carry_57_port);
   U44 : NAND2_X1 port map( A1 => net44091, A2 => B(56), ZN => net42091);
   U45 : NAND2_X1 port map( A1 => A(56), A2 => B(56), ZN => n21);
   U46 : NAND2_X1 port map( A1 => A(56), A2 => net44091, ZN => net42090);
   U47 : NAND2_X1 port map( A1 => n23, A2 => n22, ZN => net44091);
   U48 : CLKBUF_X1 port map( A => net44091, Z => net46053);
   U49 : NAND2_X1 port map( A1 => net45316, A2 => B(55), ZN => n22);
   U50 : OAI21_X1 port map( B1 => net45316, B2 => B(55), A => A(55), ZN => n23)
                           ;
   U51 : XNOR2_X1 port map( A => A(56), B => B(56), ZN => net42400);
   U52 : XNOR2_X1 port map( A => net45173, B => B(55), ZN => net45261);
   U53 : CLKBUF_X1 port map( A => A(55), Z => net73769);
   U54 : CLKBUF_X1 port map( A => A(46), Z => n32);
   U55 : OAI21_X1 port map( B1 => n112, B2 => B(50), A => A(50), ZN => n24);
   U56 : NOR2_X1 port map( A1 => n94, A2 => B(45), ZN => n25);
   U57 : XNOR2_X1 port map( A => n170, B => n45, ZN => SUM(30));
   U58 : CLKBUF_X1 port map( A => A(50), Z => n36);
   U59 : NAND2_X1 port map( A1 => n117, A2 => n24, ZN => n26);
   U60 : NAND2_X1 port map( A1 => n88, A2 => n89, ZN => n27);
   U61 : CLKBUF_X1 port map( A => A(42), Z => n28);
   U62 : NAND2_X1 port map( A1 => n62, A2 => B(36), ZN => n29);
   U63 : NOR2_X1 port map( A1 => n47, A2 => B(32), ZN => n30);
   U64 : INV_X1 port map( A => A(44), ZN => n96);
   U65 : AND2_X1 port map( A1 => n13, A2 => n31, ZN => n77);
   U66 : AND2_X1 port map( A1 => n74, A2 => n138, ZN => n31);
   U67 : XNOR2_X1 port map( A => n164, B => n68, ZN => SUM(36));
   U68 : XNOR2_X1 port map( A => n161, B => n78, ZN => SUM(39));
   U69 : XNOR2_X1 port map( A => n73, B => n138, ZN => n161);
   U70 : XNOR2_X1 port map( A => n92, B => n157, ZN => SUM(43));
   U71 : XNOR2_X1 port map( A => net45261, B => net73769, ZN => SUM(55));
   U72 : XNOR2_X1 port map( A => n153, B => n106, ZN => SUM(47));
   U73 : INV_X1 port map( A => n99, ZN => n33);
   U74 : XNOR2_X1 port map( A => n27, B => n140, ZN => n157);
   U75 : XNOR2_X1 port map( A => n159, B => n3, ZN => SUM(41));
   U76 : INV_X1 port map( A => A(43), ZN => n92);
   U77 : NAND2_X1 port map( A1 => B(37), A2 => n178, ZN => n72);
   U78 : INV_X1 port map( A => A(35), ZN => n64);
   U79 : XNOR2_X1 port map( A => n160, B => n81, ZN => SUM(40));
   U80 : INV_X1 port map( A => A(39), ZN => n78);
   U81 : INV_X1 port map( A => A(30), ZN => n45);
   U82 : XNOR2_X1 port map( A => n169, B => n49, ZN => SUM(31));
   U83 : XNOR2_X1 port map( A => n149, B => n121, ZN => SUM(51));
   U84 : NOR2_X1 port map( A1 => B(51), A2 => n26, ZN => n34);
   U85 : INV_X1 port map( A => n114, ZN => n35);
   U86 : NOR2_X1 port map( A1 => B(47), A2 => n101, ZN => n37);
   U87 : OAI21_X1 port map( B1 => B(42), B2 => n83, A => A(42), ZN => n89);
   U88 : XNOR2_X1 port map( A => n156, B => n96, ZN => SUM(44));
   U89 : XNOR2_X1 port map( A => n152, B => n110, ZN => SUM(48));
   U90 : INV_X1 port map( A => A(48), ZN => n110);
   U91 : XNOR2_X1 port map( A => n7, B => n163, ZN => SUM(37));
   U92 : INV_X1 port map( A => A(37), ZN => n71);
   U93 : XNOR2_X1 port map( A => n116, B => n144, ZN => n149);
   U94 : CLKBUF_X1 port map( A => A(53), Z => n38);
   U95 : INV_X1 port map( A => A(51), ZN => n121);
   U96 : XNOR2_X1 port map( A => n33, B => n155, ZN => SUM(45));
   U97 : XNOR2_X1 port map( A => n18, B => n142, ZN => n153);
   U98 : NAND2_X1 port map( A1 => n103, A2 => n102, ZN => n101);
   U99 : NAND2_X1 port map( A1 => n6, A2 => n88, ZN => n87);
   U100 : NAND2_X1 port map( A1 => n75, A2 => n74, ZN => n73);
   U101 : INV_X1 port map( A => A(47), ZN => n106);
   U102 : NAND2_X1 port map( A1 => n173, A2 => B(54), ZN => n132);
   U103 : XNOR2_X1 port map( A => n148, B => n125, ZN => SUM(52));
   U104 : OAI21_X1 port map( B1 => n182, B2 => B(38), A => A(38), ZN => n75);
   U105 : NAND2_X1 port map( A1 => n176, A2 => B(41), ZN => n86);
   U106 : INV_X1 port map( A => A(41), ZN => n85);
   U107 : XNOR2_X1 port map( A => B(29), B => carry_29_port, ZN => n171);
   U108 : NAND2_X1 port map( A1 => n61, A2 => n60, ZN => n59);
   U109 : XNOR2_X1 port map( A => n199, B => n39, ZN => SUM(60));
   U110 : XNOR2_X1 port map( A => A(60), B => B(60), ZN => n39);
   U111 : OAI21_X1 port map( B1 => n98, B2 => B(46), A => A(46), ZN => n103);
   U112 : XNOR2_X1 port map( A => n35, B => n151, ZN => SUM(49));
   U113 : INV_X1 port map( A => A(54), ZN => n131);
   U114 : INV_X1 port map( A => A(52), ZN => n125);
   U115 : INV_X1 port map( A => A(53), ZN => n128);
   U116 : XNOR2_X1 port map( A => A(59), B => B(59), ZN => net45328);
   U117 : INV_X1 port map( A => A(40), ZN => n81);
   U118 : XNOR2_X1 port map( A => n176, B => B(41), ZN => n159);
   U119 : NOR2_X1 port map( A1 => B(53), A2 => n123, ZN => n127);
   U120 : OAI21_X1 port map( B1 => n127, B2 => n128, A => n129, ZN => n172);
   U121 : OAI21_X1 port map( B1 => n128, B2 => n185, A => n129, ZN => n173);
   U122 : NOR2_X1 port map( A1 => n194, A2 => B(48), ZN => n109);
   U123 : OAI21_X1 port map( B1 => n109, B2 => n110, A => n111, ZN => n108);
   U124 : OAI21_X1 port map( B1 => n193, B2 => n110, A => n111, ZN => n174);
   U125 : NOR2_X1 port map( A1 => n188, A2 => B(44), ZN => n95);
   U126 : OAI21_X1 port map( B1 => n95, B2 => n96, A => n97, ZN => n94);
   U127 : OAI21_X1 port map( B1 => n187, B2 => n96, A => n97, ZN => n175);
   U128 : NOR2_X1 port map( A1 => n190, A2 => B(40), ZN => n80);
   U129 : OAI21_X1 port map( B1 => n189, B2 => n81, A => n82, ZN => n176);
   U130 : OAI21_X1 port map( B1 => n67, B2 => n68, A => n29, ZN => n66);
   U131 : NOR2_X1 port map( A1 => B(36), A2 => n62, ZN => n67);
   U132 : OAI21_X1 port map( B1 => n191, B2 => n68, A => n29, ZN => n177);
   U133 : OAI21_X1 port map( B1 => n191, B2 => n68, A => n29, ZN => n178);
   U134 : NAND2_X1 port map( A1 => n196, A2 => B(33), ZN => n58);
   U135 : XNOR2_X1 port map( A => n196, B => B(33), ZN => n167);
   U136 : NOR2_X1 port map( A1 => n51, A2 => B(33), ZN => n56);
   U137 : NOR2_X1 port map( A1 => n108, A2 => B(49), ZN => n113);
   U138 : OAI21_X1 port map( B1 => n113, B2 => n114, A => n115, ZN => n112);
   U139 : OAI21_X1 port map( B1 => n15, B2 => n114, A => n115, ZN => n179);
   U140 : XNOR2_X1 port map( A => n179, B => B(50), ZN => n150);
   U141 : NAND2_X1 port map( A1 => n179, A2 => B(50), ZN => n117);
   U142 : OAI21_X1 port map( B1 => n25, B2 => n99, A => n100, ZN => n98);
   U143 : OAI21_X1 port map( B1 => n99, B2 => n25, A => n100, ZN => n180);
   U144 : XNOR2_X1 port map( A => B(46), B => n180, ZN => n154);
   U145 : NAND2_X1 port map( A1 => n98, A2 => B(46), ZN => n102);
   U146 : OAI21_X1 port map( B1 => n84, B2 => n85, A => n86, ZN => n83);
   U147 : OAI21_X1 port map( B1 => n85, B2 => n84, A => n86, ZN => n181);
   U148 : XNOR2_X1 port map( A => n181, B => B(42), ZN => n158);
   U149 : NAND2_X1 port map( A1 => n181, A2 => B(42), ZN => n88);
   U150 : NOR2_X1 port map( A1 => B(37), A2 => n66, ZN => n70);
   U151 : OAI21_X1 port map( B1 => n70, B2 => n71, A => n72, ZN => n69);
   U152 : OAI21_X1 port map( B1 => n71, B2 => n70, A => n72, ZN => n182);
   U153 : XNOR2_X1 port map( A => n182, B => B(38), ZN => n162);
   U154 : NAND2_X1 port map( A1 => n69, A2 => B(38), ZN => n74);
   U155 : OAI21_X1 port map( B1 => n56, B2 => n57, A => n58, ZN => n55);
   U156 : NAND2_X1 port map( A1 => n17, A2 => B(34), ZN => n60);
   U157 : OAI21_X1 port map( B1 => n17, B2 => B(34), A => A(34), ZN => n61);
   U158 : XNOR2_X1 port map( A => n55, B => B(34), ZN => n166);
   U159 : OAI21_X1 port map( B1 => n120, B2 => n121, A => n122, ZN => n119);
   U160 : XNOR2_X1 port map( A => n183, B => n145, ZN => n148);
   U161 : NAND2_X1 port map( A1 => n119, A2 => B(52), ZN => n126);
   U162 : NOR2_X1 port map( A1 => n119, A2 => B(52), ZN => n124);
   U163 : NOR2_X1 port map( A1 => n116, A2 => B(51), ZN => n120);
   U164 : OAI21_X1 port map( B1 => n34, B2 => n121, A => n122, ZN => n183);
   U165 : OAI21_X1 port map( B1 => n10, B2 => n49, A => n50, ZN => n47);
   U166 : XNOR2_X1 port map( A => n184, B => n135, ZN => n168);
   U167 : NAND2_X1 port map( A1 => n184, A2 => B(32), ZN => n54);
   U168 : NOR2_X1 port map( A1 => B(32), A2 => n47, ZN => n52);
   U169 : NOR2_X1 port map( A1 => B(31), A2 => n43, ZN => n48);
   U170 : OAI21_X1 port map( B1 => n48, B2 => n49, A => n50, ZN => n184);
   U171 : NOR2_X1 port map( A1 => n186, A2 => B(53), ZN => n185);
   U172 : OAI21_X1 port map( B1 => n124, B2 => n125, A => n126, ZN => n123);
   U173 : NAND2_X1 port map( A1 => n186, A2 => B(53), ZN => n129);
   U174 : XNOR2_X1 port map( A => n123, B => B(53), ZN => n147);
   U175 : OAI21_X1 port map( B1 => n124, B2 => n125, A => n126, ZN => n186);
   U176 : NOR2_X1 port map( A1 => n90, A2 => B(44), ZN => n187);
   U177 : OAI21_X1 port map( B1 => n91, B2 => n92, A => n93, ZN => n90);
   U178 : XNOR2_X1 port map( A => n188, B => n141, ZN => n156);
   U179 : NAND2_X1 port map( A1 => n90, A2 => B(44), ZN => n97);
   U180 : NOR2_X1 port map( A1 => B(43), A2 => n87, ZN => n91);
   U181 : OAI21_X1 port map( B1 => n197, B2 => n92, A => n93, ZN => n188);
   U182 : NOR2_X1 port map( A1 => n76, A2 => B(40), ZN => n189);
   U183 : OAI21_X1 port map( B1 => n77, B2 => n78, A => n79, ZN => n76);
   U184 : XNOR2_X1 port map( A => n190, B => n139, ZN => n160);
   U185 : NAND2_X1 port map( A1 => n76, A2 => B(40), ZN => n82);
   U186 : OAI21_X1 port map( B1 => n77, B2 => n78, A => n79, ZN => n190);
   U187 : NOR2_X1 port map( A1 => n192, A2 => B(36), ZN => n191);
   U188 : OAI21_X1 port map( B1 => n63, B2 => n64, A => n65, ZN => n62);
   U189 : XNOR2_X1 port map( A => n192, B => n137, ZN => n164);
   U190 : NOR2_X1 port map( A1 => B(35), A2 => n59, ZN => n63);
   U191 : OAI21_X1 port map( B1 => n19, B2 => n64, A => n65, ZN => n192);
   U192 : NOR2_X1 port map( A1 => n104, A2 => B(48), ZN => n193);
   U193 : OAI21_X1 port map( B1 => n37, B2 => n106, A => n107, ZN => n104);
   U194 : XNOR2_X1 port map( A => n104, B => n143, ZN => n152);
   U195 : NAND2_X1 port map( A1 => n194, A2 => B(48), ZN => n111);
   U196 : NOR2_X1 port map( A1 => B(47), A2 => n18, ZN => n105);
   U197 : OAI21_X1 port map( B1 => n105, B2 => n106, A => n107, ZN => n194);
   U198 : OAI21_X1 port map( B1 => n130, B2 => n131, A => n132, ZN => net45173)
                           ;
   U199 : NOR2_X1 port map( A1 => n173, A2 => B(54), ZN => n130);
   U200 : OAI21_X1 port map( B1 => n130, B2 => n131, A => n132, ZN => net45316)
                           ;
   U201 : XNOR2_X1 port map( A => n172, B => B(54), ZN => n146);
   U202 : OAI21_X1 port map( B1 => n44, B2 => n45, A => n46, ZN => n43);
   U203 : XNOR2_X1 port map( A => n195, B => n134, ZN => n169);
   U204 : NAND2_X1 port map( A1 => n43, A2 => B(31), ZN => n50);
   U205 : NOR2_X1 port map( A1 => B(30), A2 => n40, ZN => n44);
   U206 : OAI21_X1 port map( B1 => n44, B2 => n45, A => n46, ZN => n195);
   U207 : NAND2_X1 port map( A1 => B(29), A2 => A(29), ZN => n41);
   U208 : OAI21_X1 port map( B1 => A(29), B2 => B(29), A => carry_29_port, ZN 
                           => n42);
   U209 : XNOR2_X1 port map( A => n14, B => n171, ZN => SUM(29));
   U210 : XNOR2_X1 port map( A => n147, B => n38, ZN => SUM(53));
   U211 : XNOR2_X1 port map( A => n146, B => A(54), ZN => SUM(54));
   U212 : NAND2_X1 port map( A1 => n101, A2 => B(47), ZN => n107);
   U213 : NAND2_X1 port map( A1 => B(43), A2 => n87, ZN => n93);
   U214 : NAND2_X1 port map( A1 => B(39), A2 => n73, ZN => n79);
   U215 : XNOR2_X1 port map( A => n166, B => n20, ZN => SUM(34));
   U216 : NAND2_X1 port map( A1 => B(35), A2 => n59, ZN => n65);
   U217 : XNOR2_X1 port map( A => n174, B => B(49), ZN => n151);
   U218 : NAND2_X1 port map( A1 => n42, A2 => n41, ZN => n40);
   U219 : XNOR2_X1 port map( A => n5, B => n133, ZN => n170);
   U220 : NAND2_X1 port map( A1 => B(30), A2 => n5, ZN => n46);
   U221 : XNOR2_X1 port map( A => n198, B => n167, ZN => SUM(33));
   U222 : INV_X1 port map( A => A(33), ZN => n57);
   U223 : INV_X1 port map( A => A(32), ZN => n53);
   U224 : OAI21_X1 port map( B1 => n30, B2 => n53, A => n54, ZN => n51);
   U225 : NAND2_X1 port map( A1 => n26, A2 => B(51), ZN => n122);
   U226 : XNOR2_X1 port map( A => n150, B => n36, ZN => SUM(50));
   U227 : XNOR2_X1 port map( A => n175, B => B(45), ZN => n155);
   U228 : XNOR2_X1 port map( A => n154, B => n32, ZN => SUM(46));
   U229 : NOR2_X1 port map( A1 => B(43), A2 => n27, ZN => n197);
   U230 : INV_X1 port map( A => n57, ZN => n198);
   U231 : XNOR2_X1 port map( A => n162, B => n16, ZN => SUM(38));
   U232 : NAND2_X1 port map( A1 => n174, A2 => B(49), ZN => n115);
   U233 : INV_X1 port map( A => A(49), ZN => n114);
   U234 : XNOR2_X1 port map( A => n28, B => n158, ZN => SUM(42));
   U235 : NAND2_X1 port map( A1 => n175, A2 => B(45), ZN => n100);
   U236 : INV_X1 port map( A => A(45), ZN => n99);
   U237 : OAI21_X1 port map( B1 => n112, B2 => B(50), A => A(50), ZN => n118);
   U238 : NAND2_X1 port map( A1 => n118, A2 => n117, ZN => n116);
   U239 : XNOR2_X1 port map( A => B(37), B => n177, ZN => n163);
   U240 : NAND3_X1 port map( A1 => net42063, A2 => net42064, A3 => n200, ZN => 
                           n199);
   U241 : XNOR2_X1 port map( A => net42400, B => net46053, ZN => SUM(56));
   U242 : NAND2_X1 port map( A1 => A(59), A2 => B(59), ZN => n200);
   U243 : NAND3_X1 port map( A1 => net42063, A2 => net42064, A3 => n200, ZN => 
                           carry_60_port);
   U244 : NAND2_X1 port map( A1 => carry_60_port, A2 => A(60), ZN => n201);
   U245 : NAND2_X1 port map( A1 => carry_60_port, A2 => B(60), ZN => n202);
   U246 : NAND2_X1 port map( A1 => A(60), A2 => B(60), ZN => n203);
   U247 : NAND3_X1 port map( A1 => n201, A2 => n202, A3 => n203, ZN => 
                           carry_61_port);
   U248 : XOR2_X1 port map( A => A(61), B => B(61), Z => n204);
   U249 : XOR2_X1 port map( A => carry_61_port, B => n204, Z => SUM(61));
   U250 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n1);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT60_DW01_add_0 is

   port( A, B : in std_logic_vector (59 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (59 downto 0);  CO : out std_logic);

end RCA_NBIT60_DW01_add_0;

architecture SYN_rpl of RCA_NBIT60_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_59_port, carry_58_port, carry_30_port, carry_29_port, 
      carry_28_port, carry_27_port, carry_26_port, carry_25_port, carry_24_port
      , carry_23_port, carry_22_port, carry_21_port, carry_20_port, 
      carry_19_port, carry_18_port, carry_17_port, carry_16_port, carry_15_port
      , carry_14_port, carry_13_port, carry_12_port, carry_11_port, 
      carry_10_port, carry_9_port, carry_8_port, carry_7_port, carry_6_port, 
      carry_5_port, carry_4_port, carry_3_port, carry_2_port, n1, net41887, 
      net41886, net45414, net45945, net45910, net45909, net45888, net45887, 
      net45884, net45883, net45867, net45748, net46056, net46064, net47172, 
      net45886, net45885, net45778, net45877, net45776, net73713, net45922, 
      net45773, net45772, net45953, net45779, net45777, net45771, net73789, 
      net45928, net45889, net45767, net45765, net45761, net45974, net45931, 
      net45791, net45789, net45785, net45784, net45782, net45933, net45768, 
      net45766, net45921, net45882, net45911, net45797, net45796, net45794, 
      net45790, net45788, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, 
      n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29
      , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
      n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58
      , n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, 
      n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n167, n168, n169, n170 : std_logic;

begin
   
   U1_29 : FA_X1 port map( A => B(29), B => A(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => carry_27_port, B => B(27), CI => A(27), CO => 
                           carry_28_port, S => SUM(27));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : CLKBUF_X1 port map( A => n92, Z => n3);
   U3 : INV_X1 port map( A => n100, ZN => n4);
   U4 : AND2_X1 port map( A1 => n118, A2 => n50, ZN => n58);
   U5 : NOR2_X1 port map( A1 => n57, A2 => B(32), ZN => n5);
   U6 : INV_X1 port map( A => B(33), ZN => n120);
   U7 : INV_X1 port map( A => B(41), ZN => n124);
   U8 : INV_X1 port map( A => B(40), ZN => n123);
   U9 : INV_X1 port map( A => B(45), ZN => n126);
   U10 : XNOR2_X1 port map( A => carry_59_port, B => n166, ZN => SUM(59));
   U11 : NOR2_X1 port map( A1 => n80, A2 => B(38), ZN => n6);
   U12 : NOR2_X1 port map( A1 => B(36), A2 => n73, ZN => n7);
   U13 : OAI21_X1 port map( B1 => n98, B2 => B(43), A => A(43), ZN => n8);
   U14 : CLKBUF_X1 port map( A => A(48), Z => n9);
   U15 : INV_X1 port map( A => B(31), ZN => n118);
   U16 : NOR2_X1 port map( A1 => net45771, A2 => B(52), ZN => n10);
   U17 : INV_X1 port map( A => B(48), ZN => net45867);
   U18 : XNOR2_X1 port map( A => n144, B => n59, ZN => SUM(31));
   U19 : INV_X1 port map( A => B(37), ZN => n122);
   U20 : OAI21_X1 port map( B1 => n14, B2 => n15, A => n16, ZN => n11);
   U21 : INV_X1 port map( A => B(32), ZN => n119);
   U22 : INV_X1 port map( A => B(36), ZN => n121);
   U23 : INV_X1 port map( A => B(52), ZN => n27);
   U24 : INV_X1 port map( A => B(49), ZN => n20);
   U25 : CLKBUF_X1 port map( A => A(47), Z => n53);
   U26 : INV_X1 port map( A => B(44), ZN => n125);
   U27 : INV_X1 port map( A => B(53), ZN => net45877);
   U28 : OAI21_X1 port map( B1 => n25, B2 => n18, A => n19, ZN => n17);
   U29 : OAI21_X1 port map( B1 => n12, B2 => net45796, A => net45797, ZN => 
                           net45794);
   U30 : XNOR2_X1 port map( A => net45794, B => B(56), ZN => net45882);
   U31 : NOR2_X1 port map( A1 => net45788, A2 => B(55), ZN => n12);
   U32 : NAND2_X1 port map( A1 => net45911, A2 => B(55), ZN => net45797);
   U33 : OAI21_X1 port map( B1 => net45796, B2 => n13, A => net45797, ZN => 
                           net45921);
   U34 : BUF_X1 port map( A => A(55), Z => net46056);
   U35 : INV_X1 port map( A => A(55), ZN => net45796);
   U36 : OAI21_X1 port map( B1 => net45790, B2 => net45789, A => net45791, ZN 
                           => net45788);
   U37 : NOR2_X1 port map( A1 => B(55), A2 => net45788, ZN => n13);
   U38 : INV_X1 port map( A => A(54), ZN => net45790);
   U39 : OAI21_X1 port map( B1 => net45789, B2 => net45790, A => net45791, ZN 
                           => net45911);
   U40 : XNOR2_X1 port map( A => net45911, B => B(55), ZN => net45883);
   U41 : XNOR2_X1 port map( A => net45882, B => A(56), ZN => SUM(56));
   U42 : NAND2_X1 port map( A1 => B(56), A2 => net45921, ZN => net45910);
   U43 : OAI21_X1 port map( B1 => B(56), B2 => net45921, A => A(56), ZN => 
                           net45909);
   U44 : NOR2_X1 port map( A1 => n17, A2 => B(50), ZN => net45766);
   U45 : OAI21_X1 port map( B1 => net45766, B2 => net45767, A => net45768, ZN 
                           => net45922);
   U46 : OAI21_X1 port map( B1 => net45766, B2 => net45767, A => net45768, ZN 
                           => net45765);
   U47 : INV_X1 port map( A => A(49), ZN => n25);
   U48 : OAI21_X1 port map( B1 => n23, B2 => n25, A => n19, ZN => n22);
   U49 : NOR2_X1 port map( A1 => net45933, A2 => B(49), ZN => n18);
   U50 : NAND2_X1 port map( A1 => B(50), A2 => n21, ZN => net45768);
   U51 : XNOR2_X1 port map( A => n22, B => B(50), ZN => net45888);
   U52 : NAND2_X1 port map( A1 => n11, A2 => B(49), ZN => n19);
   U53 : OAI21_X1 port map( B1 => n23, B2 => net45761, A => n19, ZN => n21);
   U54 : INV_X1 port map( A => A(49), ZN => net45761);
   U55 : OAI21_X1 port map( B1 => n24, B2 => n15, A => n16, ZN => net45933);
   U56 : XNOR2_X1 port map( A => net45933, B => n20, ZN => net45889);
   U57 : INV_X1 port map( A => A(48), ZN => n15);
   U58 : NOR2_X1 port map( A1 => B(48), A2 => net45748, ZN => n24);
   U59 : NOR2_X1 port map( A1 => B(49), A2 => n11, ZN => n23);
   U60 : INV_X1 port map( A => n9, ZN => net73713);
   U61 : NOR2_X1 port map( A1 => net45945, A2 => B(48), ZN => n14);
   U62 : NAND2_X1 port map( A1 => net45748, A2 => B(48), ZN => n16);
   U63 : NOR2_X1 port map( A1 => net45782, A2 => B(54), ZN => net45789);
   U64 : OAI21_X1 port map( B1 => net45974, B2 => net45784, A => net45785, ZN 
                           => net45782);
   U65 : NAND2_X1 port map( A1 => net45782, A2 => B(54), ZN => net45791);
   U66 : INV_X1 port map( A => A(53), ZN => net45784);
   U67 : XNOR2_X1 port map( A => net45885, B => net45784, ZN => SUM(53));
   U68 : OAI21_X1 port map( B1 => net45784, B2 => n26, A => net45785, ZN => 
                           net45931);
   U69 : NOR2_X1 port map( A1 => net45928, A2 => B(53), ZN => net45974);
   U70 : XNOR2_X1 port map( A => net45931, B => B(54), ZN => net45884);
   U71 : NAND2_X1 port map( A1 => net45928, A2 => B(53), ZN => net45785);
   U72 : NOR2_X1 port map( A1 => B(53), A2 => net45776, ZN => n26);
   U73 : OAI21_X1 port map( B1 => net45765, B2 => B(51), A => A(51), ZN => 
                           net45773);
   U74 : NAND2_X1 port map( A1 => net45765, A2 => B(51), ZN => net45772);
   U75 : INV_X1 port map( A => A(50), ZN => net45767);
   U76 : XNOR2_X1 port map( A => net45889, B => net45761, ZN => SUM(49));
   U77 : CLKBUF_X1 port map( A => A(50), Z => net47172);
   U78 : OAI21_X1 port map( B1 => n10, B2 => net73789, A => net45779, ZN => 
                           net45928);
   U79 : INV_X1 port map( A => A(52), ZN => net73789);
   U80 : OAI21_X1 port map( B1 => net45778, B2 => net45777, A => net45779, ZN 
                           => net45776);
   U81 : INV_X1 port map( A => A(52), ZN => net45778);
   U82 : NOR2_X1 port map( A1 => net45771, A2 => B(52), ZN => net45777);
   U83 : NAND2_X1 port map( A1 => net45773, A2 => net45772, ZN => net45771);
   U84 : NAND2_X1 port map( A1 => net45953, A2 => B(52), ZN => net45779);
   U85 : NAND2_X1 port map( A1 => net45773, A2 => net45772, ZN => net45953);
   U86 : XNOR2_X1 port map( A => net45953, B => n27, ZN => net45886);
   U87 : XNOR2_X1 port map( A => net45922, B => B(51), ZN => net45887);
   U88 : CLKBUF_X1 port map( A => A(51), Z => net46064);
   U89 : CLKBUF_X1 port map( A => A(26), Z => n28);
   U90 : INV_X1 port map( A => A(37), ZN => n82);
   U91 : NOR2_X1 port map( A1 => B(34), A2 => n161, ZN => n29);
   U92 : NOR2_X1 port map( A1 => B(44), A2 => n102, ZN => n30);
   U93 : NOR2_X1 port map( A1 => B(40), A2 => n87, ZN => n31);
   U94 : XNOR2_X1 port map( A => n160, B => n118, ZN => n144);
   U95 : NOR2_X1 port map( A1 => n152, A2 => B(33), ZN => n32);
   U96 : INV_X1 port map( A => A(46), ZN => n33);
   U97 : CLKBUF_X1 port map( A => A(35), Z => n34);
   U98 : OAI21_X1 port map( B1 => n29, B2 => n71, A => n72, ZN => n35);
   U99 : OAI21_X1 port map( B1 => n70, B2 => n71, A => n72, ZN => n69);
   U100 : NOR2_X1 port map( A1 => n108, A2 => B(46), ZN => n36);
   U101 : XNOR2_X1 port map( A => n37, B => n165, ZN => SUM(58));
   U102 : XNOR2_X1 port map( A => A(58), B => B(58), ZN => n37);
   U103 : NAND2_X1 port map( A1 => n89, A2 => n88, ZN => n38);
   U104 : CLKBUF_X1 port map( A => A(30), Z => n39);
   U105 : NAND2_X1 port map( A1 => n148, A2 => B(42), ZN => n40);
   U106 : CLKBUF_X1 port map( A => A(38), Z => n41);
   U107 : NAND2_X1 port map( A1 => n158, A2 => B(37), ZN => n42);
   U108 : INV_X1 port map( A => A(45), ZN => n110);
   U109 : CLKBUF_X1 port map( A => A(39), Z => n43);
   U110 : INV_X1 port map( A => A(31), ZN => n59);
   U111 : XNOR2_X1 port map( A => n135, B => n3, ZN => SUM(40));
   U112 : XOR2_X1 port map( A => carry_26_port, B => B(26), Z => n44);
   U113 : XOR2_X1 port map( A => n28, B => n44, Z => SUM(26));
   U114 : NAND2_X1 port map( A1 => n28, A2 => carry_26_port, ZN => n45);
   U115 : NAND2_X1 port map( A1 => A(26), A2 => B(26), ZN => n46);
   U116 : NAND2_X1 port map( A1 => carry_26_port, A2 => B(26), ZN => n47);
   U117 : NAND3_X1 port map( A1 => n45, A2 => n46, A3 => n47, ZN => 
                           carry_27_port);
   U118 : INV_X1 port map( A => A(41), ZN => n96);
   U119 : NAND2_X1 port map( A1 => n75, A2 => n74, ZN => n48);
   U120 : NAND2_X1 port map( A1 => n8, A2 => n103, ZN => n49);
   U121 : XNOR2_X1 port map( A => net45776, B => net45877, ZN => net45885);
   U122 : XNOR2_X1 port map( A => net45886, B => net45778, ZN => SUM(52));
   U123 : AND2_X1 port map( A1 => n56, A2 => n55, ZN => n50);
   U124 : INV_X1 port map( A => A(33), ZN => n67);
   U125 : INV_X1 port map( A => A(36), ZN => n78);
   U126 : OAI21_X1 port map( B1 => A(30), B2 => B(30), A => carry_30_port, ZN 
                           => n56);
   U127 : XNOR2_X1 port map( A => n142, B => n67, ZN => SUM(33));
   U128 : CLKBUF_X1 port map( A => A(43), Z => n51);
   U129 : INV_X1 port map( A => n33, ZN => n52);
   U130 : INV_X1 port map( A => A(32), ZN => n63);
   U131 : XNOR2_X1 port map( A => n38, B => n123, ZN => n135);
   U132 : XNOR2_X1 port map( A => n130, B => n110, ZN => SUM(45));
   U133 : XNOR2_X1 port map( A => n139, B => n78, ZN => SUM(36));
   U134 : NAND2_X1 port map( A1 => n149, A2 => B(38), ZN => n86);
   U135 : INV_X1 port map( A => A(38), ZN => n85);
   U136 : CLKBUF_X1 port map( A => A(57), Z => n54);
   U137 : INV_X1 port map( A => A(40), ZN => n92);
   U138 : NAND2_X1 port map( A1 => n146, A2 => B(46), ZN => n114);
   U139 : INV_X1 port map( A => A(44), ZN => n106);
   U140 : XNOR2_X1 port map( A => n48, B => n121, ZN => n139);
   U141 : XNOR2_X1 port map( A => n127, B => net73713, ZN => SUM(48));
   U142 : XNOR2_X1 port map( A => net45945, B => net45867, ZN => n127);
   U143 : XNOR2_X1 port map( A => n131, B => n106, ZN => SUM(44));
   U144 : XNOR2_X1 port map( A => n49, B => n125, ZN => n131);
   U145 : XNOR2_X1 port map( A => net45414, B => n117, ZN => SUM(57));
   U146 : NAND2_X1 port map( A1 => n117, A2 => B(57), ZN => net41887);
   U147 : NAND2_X1 port map( A1 => n54, A2 => n117, ZN => net41886);
   U148 : NAND2_X1 port map( A1 => net45910, A2 => net45909, ZN => n117);
   U149 : XNOR2_X1 port map( A => n138, B => n82, ZN => SUM(37));
   U150 : NOR2_X1 port map( A1 => n154, A2 => B(45), ZN => n109);
   U151 : OAI21_X1 port map( B1 => n109, B2 => n110, A => n111, ZN => n108);
   U152 : OAI21_X1 port map( B1 => n153, B2 => n110, A => n111, ZN => n146);
   U153 : NOR2_X1 port map( A1 => B(41), A2 => n156, ZN => n95);
   U154 : OAI21_X1 port map( B1 => n95, B2 => n96, A => n97, ZN => n94);
   U155 : OAI21_X1 port map( B1 => n155, B2 => n96, A => n97, ZN => n147);
   U156 : OAI21_X1 port map( B1 => n155, B2 => n96, A => n97, ZN => n148);
   U157 : OAI21_X1 port map( B1 => n81, B2 => n82, A => n42, ZN => n80);
   U158 : NOR2_X1 port map( A1 => B(37), A2 => n158, ZN => n81);
   U159 : OAI21_X1 port map( B1 => n157, B2 => n82, A => n42, ZN => n149);
   U160 : NAND2_X1 port map( A1 => n65, A2 => B(34), ZN => n72);
   U161 : XNOR2_X1 port map( A => n65, B => B(34), ZN => n141);
   U162 : NOR2_X1 port map( A1 => n161, A2 => B(34), ZN => n70);
   U163 : OAI21_X1 port map( B1 => n33, B2 => n36, A => n114, ZN => n112);
   U164 : XNOR2_X1 port map( A => n112, B => B(47), ZN => n128);
   U165 : NAND2_X1 port map( A1 => n163, A2 => B(47), ZN => n115);
   U166 : NOR2_X1 port map( A1 => n94, A2 => B(42), ZN => n99);
   U167 : OAI21_X1 port map( B1 => n99, B2 => n100, A => n101, ZN => n98);
   U168 : OAI21_X1 port map( B1 => n100, B2 => n162, A => n40, ZN => n150);
   U169 : XNOR2_X1 port map( A => n164, B => B(43), ZN => n132);
   U170 : NAND2_X1 port map( A1 => B(43), A2 => n150, ZN => n103);
   U171 : NOR2_X1 port map( A1 => n80, A2 => B(38), ZN => n84);
   U172 : OAI21_X1 port map( B1 => n84, B2 => n85, A => n86, ZN => n83);
   U173 : OAI21_X1 port map( B1 => n85, B2 => n6, A => n86, ZN => n151);
   U174 : XNOR2_X1 port map( A => n151, B => B(39), ZN => n136);
   U175 : NAND2_X1 port map( A1 => n151, A2 => B(39), ZN => n88);
   U176 : NAND2_X1 port map( A1 => n69, A2 => B(35), ZN => n74);
   U177 : OAI21_X1 port map( B1 => n69, B2 => B(35), A => A(35), ZN => n75);
   U178 : XNOR2_X1 port map( A => n35, B => B(35), ZN => n140);
   U179 : OAI21_X1 port map( B1 => n62, B2 => n63, A => n64, ZN => n61);
   U180 : XNOR2_X1 port map( A => n152, B => n120, ZN => n142);
   U181 : NAND2_X1 port map( A1 => n61, A2 => B(33), ZN => n68);
   U182 : NOR2_X1 port map( A1 => n61, A2 => B(33), ZN => n66);
   U183 : NOR2_X1 port map( A1 => n57, A2 => B(32), ZN => n62);
   U184 : OAI21_X1 port map( B1 => n5, B2 => n63, A => n64, ZN => n152);
   U185 : NOR2_X1 port map( A1 => B(45), A2 => n104, ZN => n153);
   U186 : OAI21_X1 port map( B1 => n105, B2 => n106, A => n107, ZN => n104);
   U187 : XNOR2_X1 port map( A => n154, B => n126, ZN => n130);
   U188 : NAND2_X1 port map( A1 => n104, A2 => B(45), ZN => n111);
   U189 : NOR2_X1 port map( A1 => B(44), A2 => n102, ZN => n105);
   U190 : OAI21_X1 port map( B1 => n30, B2 => n106, A => n107, ZN => n154);
   U191 : NOR2_X1 port map( A1 => n90, A2 => B(41), ZN => n155);
   U192 : OAI21_X1 port map( B1 => n91, B2 => n92, A => n93, ZN => n90);
   U193 : XNOR2_X1 port map( A => n156, B => n124, ZN => n134);
   U194 : NAND2_X1 port map( A1 => n90, A2 => B(41), ZN => n97);
   U195 : NOR2_X1 port map( A1 => B(40), A2 => n87, ZN => n91);
   U196 : OAI21_X1 port map( B1 => n31, B2 => n92, A => n93, ZN => n156);
   U197 : NOR2_X1 port map( A1 => n76, A2 => B(37), ZN => n157);
   U198 : OAI21_X1 port map( B1 => n77, B2 => n78, A => n79, ZN => n76);
   U199 : XNOR2_X1 port map( A => n76, B => n122, ZN => n138);
   U200 : NOR2_X1 port map( A1 => B(36), A2 => n73, ZN => n77);
   U201 : OAI21_X1 port map( B1 => n7, B2 => n78, A => n79, ZN => n158);
   U202 : XNOR2_X1 port map( A => net45884, B => A(54), ZN => SUM(54));
   U203 : XNOR2_X1 port map( A => net45888, B => net47172, ZN => SUM(50));
   U204 : XNOR2_X1 port map( A => net45883, B => net46056, ZN => SUM(55));
   U205 : OAI21_X1 port map( B1 => n58, B2 => n59, A => n60, ZN => n57);
   U206 : XNOR2_X1 port map( A => n159, B => n119, ZN => n143);
   U207 : NAND2_X1 port map( A1 => n159, A2 => B(32), ZN => n64);
   U208 : OAI21_X1 port map( B1 => n59, B2 => n58, A => n60, ZN => n159);
   U209 : XNOR2_X1 port map( A => n146, B => B(46), ZN => n129);
   U210 : XNOR2_X1 port map( A => net45887, B => net46064, ZN => SUM(51));
   U211 : NAND2_X1 port map( A1 => n49, A2 => B(44), ZN => n107);
   U212 : NAND2_X1 port map( A1 => n38, A2 => B(40), ZN => n93);
   U213 : NAND2_X1 port map( A1 => n48, A2 => B(36), ZN => n79);
   U214 : XNOR2_X1 port map( A => n140, B => n34, ZN => SUM(35));
   U215 : NAND2_X1 port map( A1 => n75, A2 => n74, ZN => n73);
   U216 : NAND2_X1 port map( A1 => n116, A2 => n115, ZN => net45748);
   U217 : NAND2_X1 port map( A1 => n56, A2 => n55, ZN => n160);
   U218 : XNOR2_X1 port map( A => n149, B => B(38), ZN => n137);
   U219 : XNOR2_X1 port map( A => n141, B => A(34), ZN => SUM(34));
   U220 : INV_X1 port map( A => A(34), ZN => n71);
   U221 : XNOR2_X1 port map( A => B(42), B => n147, ZN => n133);
   U222 : XNOR2_X1 port map( A => carry_30_port, B => B(30), ZN => n145);
   U223 : XNOR2_X1 port map( A => n39, B => n145, ZN => SUM(30));
   U224 : XNOR2_X1 port map( A => n129, B => n52, ZN => SUM(46));
   U225 : OAI21_X1 port map( B1 => n163, B2 => B(47), A => A(47), ZN => n116);
   U226 : NAND2_X1 port map( A1 => n116, A2 => n115, ZN => net45945);
   U227 : OAI21_X1 port map( B1 => n66, B2 => n67, A => n68, ZN => n65);
   U228 : OAI21_X1 port map( B1 => n32, B2 => n67, A => n68, ZN => n161);
   U229 : XNOR2_X1 port map( A => n128, B => n53, ZN => SUM(47));
   U230 : XNOR2_X1 port map( A => n132, B => n51, ZN => SUM(43));
   U231 : XNOR2_X1 port map( A => n133, B => n4, ZN => SUM(42));
   U232 : NAND2_X1 port map( A1 => n148, A2 => B(42), ZN => n101);
   U233 : NOR2_X1 port map( A1 => n94, A2 => B(42), ZN => n162);
   U234 : XNOR2_X1 port map( A => n136, B => n43, ZN => SUM(39));
   U235 : NAND2_X1 port map( A1 => B(31), A2 => n160, ZN => n60);
   U236 : XNOR2_X1 port map( A => n143, B => n63, ZN => SUM(32));
   U237 : NAND2_X1 port map( A1 => n8, A2 => n103, ZN => n102);
   U238 : NAND2_X1 port map( A1 => A(30), A2 => B(30), ZN => n55);
   U239 : INV_X1 port map( A => A(46), ZN => n113);
   U240 : OAI21_X1 port map( B1 => n36, B2 => n113, A => n114, ZN => n163);
   U241 : XNOR2_X1 port map( A => n134, B => n96, ZN => SUM(41));
   U242 : XNOR2_X1 port map( A => n41, B => n137, ZN => SUM(38));
   U243 : OAI21_X1 port map( B1 => n83, B2 => B(39), A => A(39), ZN => n89);
   U244 : NAND2_X1 port map( A1 => n89, A2 => n88, ZN => n87);
   U245 : INV_X1 port map( A => A(42), ZN => n100);
   U246 : OAI21_X1 port map( B1 => n162, B2 => n100, A => n40, ZN => n164);
   U247 : NAND3_X1 port map( A1 => n167, A2 => net41886, A3 => net41887, ZN => 
                           n165);
   U248 : XNOR2_X1 port map( A => A(57), B => B(57), ZN => net45414);
   U249 : XNOR2_X1 port map( A => A(59), B => B(59), ZN => n166);
   U250 : NAND2_X1 port map( A1 => n54, A2 => B(57), ZN => n167);
   U251 : NAND3_X1 port map( A1 => n167, A2 => net41886, A3 => net41887, ZN => 
                           carry_58_port);
   U252 : NAND2_X1 port map( A1 => A(58), A2 => B(58), ZN => n168);
   U253 : NAND2_X1 port map( A1 => A(58), A2 => carry_58_port, ZN => n169);
   U254 : NAND2_X1 port map( A1 => B(58), A2 => carry_58_port, ZN => n170);
   U255 : NAND3_X1 port map( A1 => n168, A2 => n169, A3 => n170, ZN => 
                           carry_59_port);
   U256 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n1);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT58_DW01_add_0 is

   port( A, B : in std_logic_vector (57 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (57 downto 0);  CO : out std_logic);

end RCA_NBIT58_DW01_add_0;

architecture SYN_rpl of RCA_NBIT58_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_57_port, carry_56_port, carry_55_port, carry_54_port, 
      carry_26_port, carry_25_port, carry_24_port, carry_23_port, carry_22_port
      , carry_21_port, carry_20_port, carry_19_port, carry_18_port, 
      carry_17_port, carry_16_port, carry_15_port, carry_14_port, carry_13_port
      , carry_12_port, carry_11_port, carry_10_port, carry_9_port, carry_8_port
      , carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port, 
      carry_2_port, n1, net42004, net42003, net45975, net47117, net47106, 
      net47082, net47059, net47058, net47057, net47056, net47054, net47038, 
      net46924, net47190, net47079, net47050, net46972, net51391, net47084, 
      net47081, net47080, net47052, net46971, net46959, net73644, net73650, 
      net73661, net73751, net46930, net46944, net46943, net46936, net47198, 
      net47097, net47053, net47185, net47113, net47096, net47086, net46962, 
      net46960, net46956, net46955, net46954, net46942, net51392, net47114, 
      net47055, net47045, net46947, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, 
      n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27
      , n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, 
      n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56
      , n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, 
      n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85
      , n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, 
      n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, 
      n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, 
      n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, 
      n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, 
      n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, 
      n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, 
      n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194 : 
      std_logic;

begin
   
   U1_56 : FA_X1 port map( A => A(56), B => B(56), CI => carry_56_port, CO => 
                           carry_57_port, S => SUM(56));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : OAI21_X1 port map( B1 => n123, B2 => n122, A => n124, ZN => n3);
   U3 : NOR2_X1 port map( A1 => B(34), A2 => n102, ZN => n4);
   U4 : OAI21_X1 port map( B1 => n45, B2 => n41, A => n43, ZN => n5);
   U5 : NAND3_X1 port map( A1 => n66, A2 => n67, A3 => n68, ZN => n6);
   U6 : NAND3_X1 port map( A1 => n62, A2 => n63, A3 => n64, ZN => n7);
   U7 : NAND3_X1 port map( A1 => n62, A2 => n63, A3 => n64, ZN => n8);
   U8 : CLKBUF_X1 port map( A => n104, Z => n9);
   U9 : NOR2_X1 port map( A1 => B(34), A2 => n102, ZN => n107);
   U10 : OAI21_X1 port map( B1 => n92, B2 => B(31), A => A(31), ZN => n10);
   U11 : CLKBUF_X1 port map( A => n100, Z => n11);
   U12 : OAI21_X1 port map( B1 => n44, B2 => n42, A => n43, ZN => n12);
   U13 : NOR2_X1 port map( A1 => n15, A2 => n14, ZN => n13);
   U14 : NOR2_X1 port map( A1 => n15, A2 => n14, ZN => n99);
   U15 : INV_X32 port map( A => n147, ZN => n14);
   U16 : NAND2_X1 port map( A1 => n10, A2 => n96, ZN => n15);
   U17 : INV_X1 port map( A => A(34), ZN => n16);
   U18 : INV_X1 port map( A => A(28), ZN => n17);
   U19 : OAI21_X1 port map( B1 => n44, B2 => n42, A => n43, ZN => n18);
   U20 : NOR2_X1 port map( A1 => n117, A2 => B(38), ZN => n19);
   U21 : CLKBUF_X1 port map( A => A(43), Z => n70);
   U22 : INV_X1 port map( A => B(33), ZN => n148);
   U23 : INV_X1 port map( A => B(44), ZN => n153);
   U24 : INV_X1 port map( A => B(52), ZN => net46971);
   U25 : INV_X1 port map( A => B(28), ZN => n145);
   U26 : INV_X1 port map( A => B(29), ZN => n146);
   U27 : INV_X1 port map( A => A(29), ZN => n20);
   U28 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => n21);
   U29 : INV_X1 port map( A => B(27), ZN => n144);
   U30 : CLKBUF_X1 port map( A => A(47), Z => net73751);
   U31 : INV_X1 port map( A => B(37), ZN => n150);
   U32 : INV_X1 port map( A => B(40), ZN => n151);
   U33 : INV_X1 port map( A => B(49), ZN => net47045);
   U34 : INV_X1 port map( A => B(41), ZN => n152);
   U35 : INV_X1 port map( A => B(45), ZN => net47038);
   U36 : INV_X1 port map( A => B(36), ZN => n149);
   U37 : INV_X1 port map( A => B(32), ZN => n147);
   U38 : OAI211_X1 port map( C1 => n132, C2 => n133, A => n134, B => n22, ZN =>
                           n23);
   U39 : INV_X1 port map( A => B(42), ZN => n22);
   U40 : INV_X1 port map( A => n23, ZN => n49);
   U41 : OAI21_X1 port map( B1 => n86, B2 => n85, A => n87, ZN => n179);
   U42 : XNOR2_X1 port map( A => net47114, B => net47045, ZN => net47055);
   U43 : XNOR2_X1 port map( A => net47055, B => net51392, ZN => SUM(49));
   U44 : OAI21_X1 port map( B1 => n24, B2 => n25, A => n26, ZN => net47114);
   U45 : NOR2_X1 port map( A1 => B(49), A2 => net47114, ZN => net46954);
   U46 : INV_X1 port map( A => A(48), ZN => n25);
   U47 : XNOR2_X1 port map( A => net47056, B => n25, ZN => SUM(48));
   U48 : OAI21_X1 port map( B1 => n27, B2 => n25, A => n26, ZN => net46947);
   U49 : NOR2_X1 port map( A1 => net46942, A2 => B(48), ZN => n24);
   U50 : NOR2_X1 port map( A1 => B(49), A2 => net46947, ZN => net47113);
   U51 : NAND2_X1 port map( A1 => net46947, A2 => B(49), ZN => net46956);
   U52 : NAND2_X1 port map( A1 => net46942, A2 => B(48), ZN => n26);
   U53 : NOR2_X1 port map( A1 => net46942, A2 => B(48), ZN => n27);
   U54 : INV_X1 port map( A => A(49), ZN => net51392);
   U55 : OAI21_X1 port map( B1 => net51392, B2 => net47113, A => net46956, ZN 
                           => net47086);
   U56 : INV_X1 port map( A => A(49), ZN => net46955);
   U57 : NAND2_X1 port map( A1 => net46944, A2 => net46943, ZN => net46942);
   U58 : AND2_X1 port map( A1 => net46944, A2 => net46943, ZN => net73661);
   U59 : OAI21_X1 port map( B1 => net46960, B2 => net47185, A => net46962, ZN 
                           => net47096);
   U60 : XNOR2_X1 port map( A => net47096, B => B(51), ZN => net47053);
   U61 : INV_X1 port map( A => A(50), ZN => net47185);
   U62 : NOR2_X1 port map( A1 => n28, A2 => B(50), ZN => net46960);
   U63 : OAI21_X1 port map( B1 => n29, B2 => net46960, A => net46962, ZN => 
                           net46959);
   U64 : OAI21_X1 port map( B1 => n29, B2 => net46960, A => net46962, ZN => 
                           net47097);
   U65 : OAI21_X1 port map( B1 => net46955, B2 => net46954, A => net46956, ZN 
                           => n28);
   U66 : OAI21_X1 port map( B1 => net46955, B2 => net47113, A => net46956, ZN 
                           => n30);
   U67 : NAND2_X1 port map( A1 => net47086, A2 => B(50), ZN => net46962);
   U68 : CLKBUF_X1 port map( A => A(50), Z => net73644);
   U69 : INV_X1 port map( A => A(50), ZN => n29);
   U70 : XNOR2_X1 port map( A => n30, B => B(50), ZN => net47054);
   U71 : XNOR2_X1 port map( A => net47053, B => net47198, ZN => SUM(51));
   U72 : OAI21_X1 port map( B1 => B(51), B2 => net73650, A => net47198, ZN => 
                           net47117);
   U73 : NAND2_X1 port map( A1 => B(51), A2 => net47097, ZN => net47080);
   U74 : OAI21_X1 port map( B1 => net46959, B2 => B(51), A => A(51), ZN => 
                           net47081);
   U75 : CLKBUF_X1 port map( A => A(51), Z => net47198);
   U76 : OAI21_X1 port map( B1 => n189, B2 => B(35), A => A(35), ZN => n31);
   U77 : NAND2_X1 port map( A1 => n97, A2 => n96, ZN => n32);
   U78 : NOR2_X1 port map( A1 => B(29), A2 => n84, ZN => n33);
   U79 : NOR2_X1 port map( A1 => B(28), A2 => n186, ZN => n34);
   U80 : INV_X1 port map( A => A(46), ZN => n35);
   U81 : OAI21_X1 port map( B1 => n39, B2 => B(47), A => A(47), ZN => net46944)
                           ;
   U82 : OAI21_X1 port map( B1 => n35, B2 => n36, A => n38, ZN => n39);
   U83 : NAND2_X1 port map( A1 => n39, A2 => B(47), ZN => net46943);
   U84 : INV_X1 port map( A => A(46), ZN => n37);
   U85 : INV_X1 port map( A => n37, ZN => net47190);
   U86 : OAI21_X1 port map( B1 => n37, B2 => n40, A => n38, ZN => net46936);
   U87 : NOR2_X1 port map( A1 => net46930, A2 => B(46), ZN => n36);
   U88 : XNOR2_X1 port map( A => net46936, B => B(47), ZN => net47057);
   U89 : NOR2_X1 port map( A1 => B(46), A2 => n5, ZN => n40);
   U90 : XNOR2_X1 port map( A => n12, B => B(46), ZN => net47058);
   U91 : NAND2_X1 port map( A1 => n18, A2 => B(46), ZN => n38);
   U92 : INV_X1 port map( A => A(45), ZN => n42);
   U93 : OAI21_X1 port map( B1 => n45, B2 => n41, A => n43, ZN => net46930);
   U94 : NOR2_X1 port map( A1 => net46924, A2 => B(45), ZN => n41);
   U95 : INV_X1 port map( A => A(45), ZN => n45);
   U96 : XNOR2_X1 port map( A => net47059, B => n45, ZN => SUM(45));
   U97 : NOR2_X1 port map( A1 => net46924, A2 => B(45), ZN => n44);
   U98 : NAND2_X1 port map( A1 => net47106, A2 => B(45), ZN => n43);
   U99 : AND2_X1 port map( A1 => n46, A2 => n79, ZN => n81);
   U100 : AND2_X1 port map( A1 => n78, A2 => n144, ZN => n46);
   U101 : INV_X1 port map( A => A(37), ZN => n47);
   U102 : INV_X1 port map( A => n136, ZN => n48);
   U103 : XNOR2_X1 port map( A => n165, B => n9, ZN => SUM(33));
   U104 : INV_X1 port map( A => A(27), ZN => n82);
   U105 : CLKBUF_X1 port map( A => net46959, Z => net73650);
   U106 : BUF_X1 port map( A => A(53), Z => n51);
   U107 : CLKBUF_X1 port map( A => A(26), Z => n50);
   U108 : NOR2_X1 port map( A1 => B(44), A2 => n138, ZN => n52);
   U109 : INV_X1 port map( A => A(44), ZN => n53);
   U110 : XNOR2_X1 port map( A => net73661, B => B(48), ZN => net47056);
   U111 : NAND2_X1 port map( A1 => net47080, A2 => net46971, ZN => net47079);
   U112 : XNOR2_X1 port map( A => carry_54_port, B => n54, ZN => SUM(54));
   U113 : XNOR2_X1 port map( A => A(54), B => B(54), ZN => n54);
   U114 : NAND2_X1 port map( A1 => carry_54_port, A2 => A(54), ZN => n55);
   U115 : NAND2_X1 port map( A1 => carry_54_port, A2 => B(54), ZN => n56);
   U116 : NAND2_X1 port map( A1 => A(54), A2 => B(54), ZN => n57);
   U117 : NAND3_X1 port map( A1 => n55, A2 => n56, A3 => n57, ZN => 
                           carry_55_port);
   U118 : OAI21_X1 port map( B1 => n182, B2 => n119, A => n120, ZN => n58);
   U119 : INV_X1 port map( A => A(33), ZN => n104);
   U120 : OAI21_X1 port map( B1 => n93, B2 => n94, A => n95, ZN => n59);
   U121 : INV_X1 port map( A => n16, ZN => n60);
   U122 : XOR2_X1 port map( A => A(24), B => B(24), Z => n61);
   U123 : XOR2_X1 port map( A => n61, B => carry_24_port, Z => SUM(24));
   U124 : NAND2_X1 port map( A1 => A(24), A2 => B(24), ZN => n62);
   U125 : NAND2_X1 port map( A1 => A(24), A2 => carry_24_port, ZN => n63);
   U126 : NAND2_X1 port map( A1 => B(24), A2 => carry_24_port, ZN => n64);
   U127 : NAND3_X1 port map( A1 => n62, A2 => n63, A3 => n64, ZN => 
                           carry_25_port);
   U128 : XOR2_X1 port map( A => A(25), B => B(25), Z => n65);
   U129 : XOR2_X1 port map( A => n65, B => n8, Z => SUM(25));
   U130 : NAND2_X1 port map( A1 => A(25), A2 => B(25), ZN => n66);
   U131 : NAND2_X1 port map( A1 => A(25), A2 => n7, ZN => n67);
   U132 : NAND2_X1 port map( A1 => B(25), A2 => carry_25_port, ZN => n68);
   U133 : NAND3_X1 port map( A1 => n66, A2 => n67, A3 => n68, ZN => 
                           carry_26_port);
   U134 : XNOR2_X1 port map( A => n171, B => n82, ZN => SUM(27));
   U135 : INV_X1 port map( A => A(41), ZN => n133);
   U136 : XNOR2_X1 port map( A => n162, B => n115, ZN => SUM(36));
   U137 : XNOR2_X1 port map( A => n161, B => n47, ZN => SUM(37));
   U138 : XNOR2_X1 port map( A => n191, B => n153, ZN => n154);
   U139 : NAND2_X1 port map( A1 => n31, A2 => n111, ZN => n69);
   U140 : NAND2_X1 port map( A1 => n175, A2 => B(38), ZN => n124);
   U141 : OAI21_X1 port map( B1 => net51391, B2 => net46971, A => net46972, ZN 
                           => net45975);
   U142 : XNOR2_X1 port map( A => net47084, B => net46971, ZN => net47052);
   U143 : XNOR2_X1 port map( A => net47052, B => net47050, ZN => SUM(52));
   U144 : NAND2_X1 port map( A1 => net47081, A2 => net47080, ZN => net47084);
   U145 : AND2_X1 port map( A1 => net47117, A2 => net47080, ZN => net51391);
   U146 : INV_X1 port map( A => A(52), ZN => net47050);
   U147 : OAI21_X1 port map( B1 => net47082, B2 => net47079, A => A(52), ZN => 
                           net46972);
   U148 : OAI21_X1 port map( B1 => n93, B2 => n94, A => n95, ZN => n92);
   U149 : XNOR2_X1 port map( A => n169, B => n90, ZN => SUM(29));
   U150 : XOR2_X1 port map( A => A(55), B => B(55), Z => n71);
   U151 : XOR2_X1 port map( A => carry_55_port, B => n71, Z => SUM(55));
   U152 : NAND2_X1 port map( A1 => carry_55_port, A2 => A(55), ZN => n72);
   U153 : NAND2_X1 port map( A1 => carry_55_port, A2 => B(55), ZN => n73);
   U154 : NAND2_X1 port map( A1 => A(55), A2 => B(55), ZN => n74);
   U155 : NAND3_X1 port map( A1 => n72, A2 => n73, A3 => n74, ZN => 
                           carry_56_port);
   U156 : NAND2_X1 port map( A1 => net45975, A2 => n51, ZN => net42003);
   U157 : NAND2_X1 port map( A1 => net45975, A2 => B(53), ZN => net42004);
   U158 : OAI21_X1 port map( B1 => B(43), B2 => n135, A => A(43), ZN => n75);
   U159 : XNOR2_X1 port map( A => n154, B => n53, ZN => SUM(44));
   U160 : XNOR2_X1 port map( A => n157, B => n133, ZN => SUM(41));
   U161 : XNOR2_X1 port map( A => n166, B => n11, ZN => SUM(32));
   U162 : NAND2_X1 port map( A1 => n176, A2 => B(34), ZN => n109);
   U163 : INV_X1 port map( A => A(37), ZN => n119);
   U164 : XNOR2_X1 port map( A => n158, B => n130, ZN => SUM(40));
   U165 : XNOR2_X1 port map( A => n21, B => n151, ZN => n158);
   U166 : XNOR2_X1 port map( A => n170, B => n17, ZN => SUM(28));
   U167 : OAI21_X1 port map( B1 => n52, B2 => n142, A => n143, ZN => n76);
   U168 : NOR2_X1 port map( A1 => B(41), A2 => n128, ZN => n132);
   U169 : OAI21_X1 port map( B1 => n133, B2 => n180, A => n134, ZN => n173);
   U170 : OAI21_X1 port map( B1 => n180, B2 => n133, A => n134, ZN => n174);
   U171 : OAI21_X1 port map( B1 => n118, B2 => n119, A => n120, ZN => n117);
   U172 : NOR2_X1 port map( A1 => n113, A2 => B(37), ZN => n118);
   U173 : OAI21_X1 port map( B1 => n182, B2 => n47, A => n120, ZN => n175);
   U174 : OAI21_X1 port map( B1 => n103, B2 => n104, A => n105, ZN => n102);
   U175 : NOR2_X1 port map( A1 => n185, A2 => B(33), ZN => n103);
   U176 : OAI21_X1 port map( B1 => n184, B2 => n104, A => n105, ZN => n176);
   U177 : NAND2_X1 port map( A1 => n88, A2 => B(30), ZN => n95);
   U178 : XNOR2_X1 port map( A => n187, B => B(30), ZN => n168);
   U179 : NOR2_X1 port map( A1 => n88, A2 => B(30), ZN => n93);
   U180 : OAI21_X1 port map( B1 => n49, B2 => n136, A => n137, ZN => n135);
   U181 : OAI21_X1 port map( B1 => n49, B2 => n136, A => n137, ZN => n177);
   U182 : XNOR2_X1 port map( A => n135, B => B(43), ZN => n155);
   U183 : NAND2_X1 port map( A1 => n177, A2 => B(43), ZN => n139);
   U184 : NOR2_X1 port map( A1 => n117, A2 => B(38), ZN => n122);
   U185 : OAI21_X1 port map( B1 => n19, B2 => n123, A => n124, ZN => n121);
   U186 : XNOR2_X1 port map( A => n3, B => B(39), ZN => n159);
   U187 : NAND2_X1 port map( A1 => n190, A2 => B(39), ZN => n126);
   U188 : OAI21_X1 port map( B1 => n4, B2 => n108, A => n109, ZN => n106);
   U189 : OAI21_X1 port map( B1 => n4, B2 => n16, A => n109, ZN => n178);
   U190 : XNOR2_X1 port map( A => B(35), B => n178, ZN => n163);
   U191 : NAND2_X1 port map( A1 => B(35), A2 => n106, ZN => n111);
   U192 : NAND2_X1 port map( A1 => n59, A2 => B(31), ZN => n96);
   U193 : OAI21_X1 port map( B1 => n92, B2 => B(31), A => A(31), ZN => n97);
   U194 : XNOR2_X1 port map( A => n59, B => B(31), ZN => n167);
   U195 : OAI21_X1 port map( B1 => n34, B2 => n17, A => n87, ZN => n84);
   U196 : XNOR2_X1 port map( A => n179, B => n146, ZN => n169);
   U197 : NAND2_X1 port map( A1 => n179, A2 => B(29), ZN => n91);
   U198 : NOR2_X1 port map( A1 => B(29), A2 => n84, ZN => n89);
   U199 : NOR2_X1 port map( A1 => B(28), A2 => n186, ZN => n85);
   U200 : OAI21_X1 port map( B1 => n141, B2 => n142, A => n143, ZN => net46924)
                           ;
   U201 : XNOR2_X1 port map( A => n76, B => net47038, ZN => net47059);
   U202 : NOR2_X1 port map( A1 => n138, A2 => B(44), ZN => n141);
   U203 : OAI21_X1 port map( B1 => n53, B2 => n141, A => n143, ZN => net47106);
   U204 : NOR2_X1 port map( A1 => B(41), A2 => n181, ZN => n180);
   U205 : OAI21_X1 port map( B1 => n129, B2 => n130, A => n131, ZN => n128);
   U206 : XNOR2_X1 port map( A => n128, B => n152, ZN => n157);
   U207 : NAND2_X1 port map( A1 => n181, A2 => B(41), ZN => n134);
   U208 : NOR2_X1 port map( A1 => n125, A2 => B(40), ZN => n129);
   U209 : OAI21_X1 port map( B1 => n129, B2 => n130, A => n131, ZN => n181);
   U210 : NOR2_X1 port map( A1 => n183, A2 => B(37), ZN => n182);
   U211 : OAI21_X1 port map( B1 => n114, B2 => n115, A => n116, ZN => n113);
   U212 : XNOR2_X1 port map( A => n113, B => n150, ZN => n161);
   U213 : NAND2_X1 port map( A1 => n183, A2 => B(37), ZN => n120);
   U214 : NOR2_X1 port map( A1 => B(36), A2 => n110, ZN => n114);
   U215 : OAI21_X1 port map( B1 => n114, B2 => n115, A => n116, ZN => n183);
   U216 : NOR2_X1 port map( A1 => n98, A2 => B(33), ZN => n184);
   U217 : OAI21_X1 port map( B1 => n13, B2 => n100, A => n101, ZN => n98);
   U218 : XNOR2_X1 port map( A => n185, B => n148, ZN => n165);
   U219 : NAND2_X1 port map( A1 => n98, A2 => B(33), ZN => n105);
   U220 : OAI21_X1 port map( B1 => n99, B2 => n100, A => n101, ZN => n185);
   U221 : OAI21_X1 port map( B1 => n81, B2 => n82, A => n83, ZN => n80);
   U222 : XNOR2_X1 port map( A => n80, B => n145, ZN => n170);
   U223 : NAND2_X1 port map( A1 => n80, A2 => B(28), ZN => n87);
   U224 : OAI21_X1 port map( B1 => n81, B2 => n82, A => n83, ZN => n186);
   U225 : NAND2_X1 port map( A1 => A(26), A2 => B(26), ZN => n78);
   U226 : OAI21_X1 port map( B1 => A(26), B2 => B(26), A => n6, ZN => n79);
   U227 : XNOR2_X1 port map( A => n172, B => n50, ZN => SUM(26));
   U228 : INV_X1 port map( A => net47081, ZN => net47082);
   U229 : XNOR2_X1 port map( A => net47054, B => net73644, ZN => SUM(50));
   U230 : NAND2_X1 port map( A1 => n138, A2 => B(44), ZN => n143);
   U231 : NAND2_X1 port map( A1 => n21, A2 => B(40), ZN => n131);
   U232 : NAND2_X1 port map( A1 => B(36), A2 => n69, ZN => n116);
   U233 : XNOR2_X1 port map( A => n167, B => A(31), ZN => SUM(31));
   U234 : NAND2_X1 port map( A1 => B(32), A2 => n32, ZN => n101);
   U235 : NAND2_X1 port map( A1 => n78, A2 => n79, ZN => n77);
   U236 : XNOR2_X1 port map( A => n168, B => n188, ZN => SUM(30));
   U237 : INV_X1 port map( A => A(30), ZN => n94);
   U238 : XNOR2_X1 port map( A => n77, B => n144, ZN => n171);
   U239 : NAND2_X1 port map( A1 => n77, A2 => B(27), ZN => n83);
   U240 : OAI21_X1 port map( B1 => n89, B2 => n20, A => n91, ZN => n88);
   U241 : OAI21_X1 port map( B1 => n33, B2 => n90, A => n91, ZN => n187);
   U242 : XNOR2_X1 port map( A => net47057, B => net73751, ZN => SUM(47));
   U243 : XNOR2_X1 port map( A => B(38), B => n58, ZN => n160);
   U244 : NAND2_X1 port map( A1 => n140, A2 => n139, ZN => n138);
   U245 : XNOR2_X1 port map( A => n176, B => B(34), ZN => n164);
   U246 : INV_X1 port map( A => n94, ZN => n188);
   U247 : XNOR2_X1 port map( A => n155, B => n70, ZN => SUM(43));
   U248 : INV_X1 port map( A => A(29), ZN => n90);
   U249 : XNOR2_X1 port map( A => n173, B => B(42), ZN => n156);
   U250 : XNOR2_X1 port map( A => A(35), B => n163, ZN => SUM(35));
   U251 : XNOR2_X1 port map( A => carry_26_port, B => B(26), ZN => n172);
   U252 : XNOR2_X1 port map( A => n159, B => A(39), ZN => SUM(39));
   U253 : OAI21_X1 port map( B1 => n177, B2 => B(43), A => A(43), ZN => n140);
   U254 : INV_X1 port map( A => A(34), ZN => n108);
   U255 : OAI21_X1 port map( B1 => n107, B2 => n108, A => n109, ZN => n189);
   U256 : OAI21_X1 port map( B1 => n189, B2 => B(35), A => A(35), ZN => n112);
   U257 : NAND2_X1 port map( A1 => n112, A2 => n111, ZN => n110);
   U258 : NAND2_X1 port map( A1 => n174, A2 => B(42), ZN => n137);
   U259 : INV_X1 port map( A => A(42), ZN => n136);
   U260 : INV_X1 port map( A => A(32), ZN => n100);
   U261 : INV_X1 port map( A => A(38), ZN => n123);
   U262 : OAI21_X1 port map( B1 => n123, B2 => n122, A => n124, ZN => n190);
   U263 : INV_X1 port map( A => A(44), ZN => n142);
   U264 : OAI21_X1 port map( B1 => n121, B2 => B(39), A => A(39), ZN => n127);
   U265 : NAND2_X1 port map( A1 => n127, A2 => n126, ZN => n125);
   U266 : XNOR2_X1 port map( A => n164, B => n60, ZN => SUM(34));
   U267 : XNOR2_X1 port map( A => A(38), B => n160, ZN => SUM(38));
   U268 : XNOR2_X1 port map( A => n32, B => n147, ZN => n166);
   U269 : NAND2_X1 port map( A1 => n139, A2 => n75, ZN => n191);
   U270 : XNOR2_X1 port map( A => net47058, B => net47190, ZN => SUM(46));
   U271 : INV_X1 port map( A => A(40), ZN => n130);
   U272 : XNOR2_X1 port map( A => n156, B => n48, ZN => SUM(42));
   U273 : XNOR2_X1 port map( A => n69, B => n149, ZN => n162);
   U274 : INV_X1 port map( A => A(36), ZN => n115);
   U275 : INV_X1 port map( A => A(28), ZN => n86);
   U276 : XNOR2_X1 port map( A => net45975, B => n192, ZN => SUM(53));
   U277 : XNOR2_X1 port map( A => A(53), B => B(53), ZN => n192);
   U278 : XNOR2_X1 port map( A => carry_57_port, B => n193, ZN => SUM(57));
   U279 : XNOR2_X1 port map( A => A(57), B => B(57), ZN => n193);
   U280 : NAND2_X1 port map( A1 => n51, A2 => B(53), ZN => n194);
   U281 : NAND3_X1 port map( A1 => net42003, A2 => net42004, A3 => n194, ZN => 
                           carry_54_port);
   U282 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n1);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT56_DW01_add_0 is

   port( A, B : in std_logic_vector (55 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (55 downto 0);  CO : out std_logic);

end RCA_NBIT56_DW01_add_0;

architecture SYN_rpl of RCA_NBIT56_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_55_port, carry_54_port, carry_53_port, carry_25_port, 
      carry_24_port, carry_23_port, carry_22_port, carry_21_port, carry_20_port
      , carry_19_port, carry_18_port, carry_17_port, carry_16_port, 
      carry_15_port, carry_14_port, carry_13_port, carry_12_port, carry_11_port
      , carry_10_port, carry_9_port, carry_8_port, carry_7_port, carry_6_port, 
      carry_5_port, carry_4_port, carry_3_port, carry_2_port, n1, net46026, 
      net46025, net73431, net73429, net73384, net73382, net73380, net73363, 
      net73286, net73264, net73259, net73253, net73248, net73246, net73576, 
      net73776, net73381, net79778, net73668, net73642, net73289, net73287, 
      net73409, net73408, net73378, net73377, net73282, net73280, net73527, 
      net73428, net73283, net73281, net73277, net73276, net73275, net73260, 
      net73258, net73245, net73699, net73465, net73418, net73265, net73762, 
      net73424, net73379, net73370, net73691, net73687, net73271, net73269, 
      net73268, net73263, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, 
      n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29
      , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
      n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58
      , n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, 
      n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, 
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186 : std_logic;

begin
   
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : CLKBUF_X1 port map( A => A(23), Z => n3);
   U3 : OAI21_X1 port map( B1 => n50, B2 => B(30), A => A(30), ZN => n4);
   U4 : CLKBUF_X1 port map( A => A(22), Z => n5);
   U5 : OAI21_X1 port map( B1 => n65, B2 => n66, A => n67, ZN => n6);
   U6 : NOR2_X1 port map( A1 => B(26), A2 => n51, ZN => n7);
   U7 : CLKBUF_X1 port map( A => A(34), Z => n8);
   U8 : INV_X1 port map( A => A(32), ZN => n9);
   U9 : CLKBUF_X1 port map( A => n63, Z => n10);
   U10 : OAI21_X1 port map( B1 => n56, B2 => n7, A => n57, ZN => n11);
   U11 : NOR2_X1 port map( A1 => B(29), A2 => n61, ZN => n12);
   U12 : NOR2_X1 port map( A1 => n90, A2 => B(37), ZN => n13);
   U13 : INV_X1 port map( A => A(41), ZN => n14);
   U14 : BUF_X1 port map( A => A(38), Z => n15);
   U15 : CLKBUF_X1 port map( A => A(53), Z => n16);
   U16 : XNOR2_X1 port map( A => n142, B => n59, ZN => SUM(27));
   U17 : INV_X1 port map( A => B(28), ZN => n117);
   U18 : NAND2_X1 port map( A1 => n146, A2 => n145, ZN => n114);
   U19 : NAND2_X1 port map( A1 => n114, A2 => B(52), ZN => net46026);
   U20 : INV_X1 port map( A => B(44), ZN => net73363);
   U21 : INV_X1 port map( A => B(48), ZN => net73370);
   U22 : INV_X1 port map( A => B(32), ZN => n119);
   U23 : INV_X1 port map( A => B(36), ZN => n121);
   U24 : INV_X1 port map( A => B(39), ZN => n122);
   U25 : INV_X1 port map( A => B(40), ZN => n123);
   U26 : OAI21_X1 port map( B1 => n79, B2 => B(34), A => A(34), ZN => n17);
   U27 : INV_X1 port map( A => B(31), ZN => n118);
   U28 : INV_X1 port map( A => B(35), ZN => n120);
   U29 : INV_X1 port map( A => B(47), ZN => n19);
   U30 : INV_X1 port map( A => B(43), ZN => n124);
   U31 : OAI21_X1 port map( B1 => B(38), B2 => n94, A => A(38), ZN => n18);
   U32 : INV_X1 port map( A => B(27), ZN => n116);
   U33 : AND3_X1 port map( A1 => n84, A2 => n85, A3 => n120, ZN => n87);
   U34 : AND3_X1 port map( A1 => n113, A2 => n112, A3 => n124, ZN => net73246);
   U35 : OAI21_X1 port map( B1 => n77, B2 => n76, A => n78, ZN => n75);
   U36 : OAI21_X1 port map( B1 => net73687, B2 => net73269, A => net73271, ZN 
                           => net73268);
   U37 : XNOR2_X1 port map( A => net73268, B => net73370, ZN => net73379);
   U38 : INV_X1 port map( A => A(47), ZN => net73687);
   U39 : OAI21_X1 port map( B1 => net73687, B2 => net73269, A => net73271, ZN 
                           => net73762);
   U40 : AND2_X1 port map( A1 => net73265, A2 => net73691, ZN => net73269);
   U41 : OAI21_X1 port map( B1 => net73687, B2 => net73269, A => net73271, ZN 
                           => net73424);
   U42 : AND2_X1 port map( A1 => net73264, A2 => n19, ZN => net73691);
   U43 : NAND2_X1 port map( A1 => net73263, A2 => B(47), ZN => net73271);
   U44 : NAND2_X1 port map( A1 => net73265, A2 => net73264, ZN => net73263);
   U45 : XNOR2_X1 port map( A => net73263, B => n19, ZN => net73380);
   U46 : XNOR2_X1 port map( A => net73276, B => net73379, ZN => SUM(48));
   U47 : NAND2_X1 port map( A1 => net73424, A2 => B(48), ZN => net73277);
   U48 : NOR2_X1 port map( A1 => B(48), A2 => net73762, ZN => net73527);
   U49 : NOR2_X1 port map( A1 => net73424, A2 => B(48), ZN => net73275);
   U50 : OAI21_X1 port map( B1 => net73465, B2 => B(46), A => A(46), ZN => 
                           net73265);
   U51 : OAI21_X1 port map( B1 => net73258, B2 => net73699, A => net73260, ZN 
                           => net73465);
   U52 : XNOR2_X1 port map( A => net73465, B => B(46), ZN => net73381);
   U53 : INV_X1 port map( A => A(45), ZN => net73699);
   U54 : NAND2_X1 port map( A1 => net73418, A2 => B(46), ZN => net73264);
   U55 : CLKBUF_X1 port map( A => A(46), Z => net73776);
   U56 : OAI21_X1 port map( B1 => net73259, B2 => net73258, A => net73260, ZN 
                           => net73418);
   U57 : INV_X1 port map( A => A(45), ZN => net73259);
   U58 : NOR2_X1 port map( A1 => n21, A2 => B(45), ZN => net73258);
   U59 : OAI21_X1 port map( B1 => n27, B2 => n22, A => n23, ZN => n21);
   U60 : NOR2_X1 port map( A1 => B(44), A2 => net73431, ZN => n22);
   U61 : INV_X1 port map( A => A(44), ZN => n27);
   U62 : OAI21_X1 port map( B1 => n26, B2 => n27, A => n23, ZN => n24);
   U63 : NAND2_X1 port map( A1 => n24, A2 => B(45), ZN => net73260);
   U64 : XNOR2_X1 port map( A => n25, B => B(45), ZN => net73382);
   U65 : NAND2_X1 port map( A1 => net73245, A2 => B(44), ZN => n23);
   U66 : OAI21_X1 port map( B1 => net73253, B2 => n26, A => n23, ZN => n25);
   U67 : NOR2_X1 port map( A1 => net73245, A2 => B(44), ZN => n26);
   U68 : OAI21_X1 port map( B1 => net73246, B2 => n20, A => net73248, ZN => 
                           net73245);
   U69 : INV_X1 port map( A => A(43), ZN => n20);
   U70 : XNOR2_X1 port map( A => net73384, B => n20, ZN => SUM(43));
   U71 : OAI21_X1 port map( B1 => n20, B2 => net73246, A => net73248, ZN => 
                           net73431);
   U72 : INV_X1 port map( A => A(44), ZN => net73253);
   U73 : NAND2_X1 port map( A1 => n28, A2 => B(49), ZN => net73283);
   U74 : OAI21_X1 port map( B1 => net73281, B2 => net73282, A => net73283, ZN 
                           => net73280);
   U75 : OAI21_X1 port map( B1 => n29, B2 => net73282, A => net73283, ZN => 
                           net73409);
   U76 : OAI21_X1 port map( B1 => net73281, B2 => net73282, A => net73283, ZN 
                           => net73408);
   U77 : OAI21_X1 port map( B1 => net73276, B2 => net73527, A => net73277, ZN 
                           => n28);
   U78 : NOR2_X1 port map( A1 => B(49), A2 => n28, ZN => net73281);
   U79 : INV_X1 port map( A => A(48), ZN => net73276);
   U80 : OAI21_X1 port map( B1 => net73276, B2 => net73275, A => net73277, ZN 
                           => net73428);
   U81 : XNOR2_X1 port map( A => net73428, B => B(49), ZN => net73378);
   U82 : NOR2_X1 port map( A1 => B(49), A2 => net73428, ZN => n29);
   U83 : XNOR2_X1 port map( A => net73409, B => B(50), ZN => net73377);
   U84 : XNOR2_X1 port map( A => net73377, B => net73668, ZN => SUM(50));
   U85 : INV_X1 port map( A => A(49), ZN => net73282);
   U86 : NAND2_X1 port map( A1 => B(50), A2 => net73408, ZN => net73289);
   U87 : NOR2_X1 port map( A1 => B(50), A2 => net73280, ZN => net73642);
   U88 : NOR2_X1 port map( A1 => net73280, A2 => B(50), ZN => net73287);
   U89 : XNOR2_X1 port map( A => net73378, B => A(49), ZN => SUM(49));
   U90 : INV_X1 port map( A => net79778, ZN => net73668);
   U91 : INV_X1 port map( A => A(50), ZN => net79778);
   U92 : OAI21_X1 port map( B1 => net73642, B2 => net79778, A => net73289, ZN 
                           => net73429);
   U93 : OAI21_X1 port map( B1 => net73287, B2 => net79778, A => net73289, ZN 
                           => net73286);
   U94 : NOR2_X1 port map( A1 => B(26), A2 => n51, ZN => n30);
   U95 : NAND2_X1 port map( A1 => n112, A2 => n113, ZN => n31);
   U96 : NOR2_X1 port map( A1 => B(28), A2 => n58, ZN => n32);
   U97 : OAI21_X1 port map( B1 => n34, B2 => n81, A => n82, ZN => n33);
   U98 : NOR2_X1 port map( A1 => B(33), A2 => n75, ZN => n34);
   U99 : NOR2_X1 port map( A1 => B(41), A2 => n105, ZN => n35);
   U100 : XOR2_X1 port map( A => carry_23_port, B => B(23), Z => n36);
   U101 : XOR2_X1 port map( A => n3, B => n36, Z => SUM(23));
   U102 : NAND2_X1 port map( A1 => A(23), A2 => carry_23_port, ZN => n37);
   U103 : NAND2_X1 port map( A1 => A(23), A2 => B(23), ZN => n38);
   U104 : NAND2_X1 port map( A1 => carry_23_port, A2 => B(23), ZN => n39);
   U105 : NAND3_X1 port map( A1 => n37, A2 => n38, A3 => n39, ZN => 
                           carry_24_port);
   U106 : XNOR2_X1 port map( A => net73381, B => net73776, ZN => SUM(46));
   U107 : CLKBUF_X1 port map( A => A(33), Z => n40);
   U108 : NAND2_X1 port map( A1 => n153, A2 => B(33), ZN => n82);
   U109 : NOR2_X1 port map( A1 => B(29), A2 => n61, ZN => n65);
   U110 : CLKBUF_X1 port map( A => A(42), Z => n43);
   U111 : AND2_X1 port map( A1 => n41, A2 => n4, ZN => n72);
   U112 : AND2_X1 port map( A1 => n69, A2 => n118, ZN => n41);
   U113 : NAND2_X1 port map( A1 => n18, A2 => n99, ZN => n42);
   U114 : XNOR2_X1 port map( A => n83, B => n120, ZN => n134);
   U115 : XNOR2_X1 port map( A => n177, B => n44, ZN => SUM(54));
   U116 : XNOR2_X1 port map( A => A(54), B => B(54), ZN => n44);
   U117 : NAND2_X1 port map( A1 => n114, A2 => A(52), ZN => net46025);
   U118 : NOR2_X1 port map( A1 => n54, A2 => B(27), ZN => n45);
   U119 : NAND2_X1 port map( A1 => n165, A2 => B(26), ZN => n57);
   U120 : XNOR2_X1 port map( A => n138, B => n73, ZN => SUM(31));
   U121 : XNOR2_X1 port map( A => n42, B => n122, ZN => n130);
   U122 : INV_X1 port map( A => A(40), ZN => n46);
   U123 : XNOR2_X1 port map( A => A(52), B => B(52), ZN => n48);
   U124 : XNOR2_X1 port map( A => carry_53_port, B => n47, ZN => SUM(53));
   U125 : XNOR2_X1 port map( A => A(53), B => B(53), ZN => n47);
   U126 : XNOR2_X1 port map( A => n48, B => n114, ZN => SUM(52));
   U127 : INV_X1 port map( A => net73259, ZN => net73576);
   U128 : XNOR2_X1 port map( A => net73380, B => net73687, ZN => SUM(47));
   U129 : XNOR2_X1 port map( A => n134, B => n88, ZN => SUM(35));
   U130 : XNOR2_X1 port map( A => n143, B => n56, ZN => SUM(26));
   U131 : XNOR2_X1 port map( A => n165, B => n115, ZN => n143);
   U132 : OAI21_X1 port map( B1 => n65, B2 => n66, A => n67, ZN => n49);
   U133 : OAI21_X1 port map( B1 => n12, B2 => n66, A => n67, ZN => n50);
   U134 : INV_X1 port map( A => A(32), ZN => n77);
   U135 : NAND2_X1 port map( A1 => n17, A2 => n84, ZN => n83);
   U136 : XNOR2_X1 port map( A => n130, B => n103, ZN => SUM(39));
   U137 : INV_X1 port map( A => A(31), ZN => n73);
   U138 : NAND2_X1 port map( A1 => B(41), A2 => n149, ZN => n111);
   U139 : XNOR2_X1 port map( A => n141, B => n10, ZN => SUM(28));
   U140 : NAND2_X1 port map( A1 => n100, A2 => n99, ZN => n98);
   U141 : XNOR2_X1 port map( A => n31, B => n124, ZN => net73384);
   U142 : INV_X1 port map( A => A(40), ZN => n107);
   U143 : XNOR2_X1 port map( A => n126, B => net73253, ZN => SUM(44));
   U144 : INV_X2 port map( A => B(26), ZN => n115);
   U145 : NAND2_X1 port map( A1 => A(25), A2 => B(25), ZN => n52);
   U146 : OAI21_X1 port map( B1 => A(25), B2 => B(25), A => carry_25_port, ZN 
                           => n53);
   U147 : XNOR2_X1 port map( A => n144, B => n147, ZN => SUM(25));
   U148 : CLKBUF_X1 port map( A => A(25), Z => n147);
   U149 : NOR2_X1 port map( A1 => B(40), A2 => n160, ZN => n106);
   U150 : OAI21_X1 port map( B1 => n107, B2 => n106, A => n108, ZN => n105);
   U151 : OAI21_X1 port map( B1 => n159, B2 => n107, A => n108, ZN => n148);
   U152 : OAI21_X1 port map( B1 => n159, B2 => n46, A => n108, ZN => n149);
   U153 : OAI21_X1 port map( B1 => n92, B2 => n91, A => n93, ZN => n90);
   U154 : NOR2_X1 port map( A1 => B(36), A2 => n86, ZN => n91);
   U155 : OAI21_X1 port map( B1 => n92, B2 => n161, A => n93, ZN => n150);
   U156 : OAI21_X1 port map( B1 => n161, B2 => n92, A => n93, ZN => n151);
   U157 : NOR2_X1 port map( A1 => B(32), A2 => n71, ZN => n76);
   U158 : OAI21_X1 port map( B1 => n163, B2 => n77, A => n78, ZN => n152);
   U159 : OAI21_X1 port map( B1 => n163, B2 => n9, A => n78, ZN => n153);
   U160 : NAND2_X1 port map( A1 => n166, A2 => B(29), ZN => n67);
   U161 : XNOR2_X1 port map( A => n166, B => B(29), ZN => n140);
   U162 : NAND2_X1 port map( A1 => B(51), A2 => net73429, ZN => n146);
   U163 : OAI21_X1 port map( B1 => B(51), B2 => net73429, A => A(51), ZN => 
                           n145);
   U164 : XNOR2_X1 port map( A => net73286, B => B(51), ZN => n125);
   U165 : OAI21_X1 port map( B1 => n110, B2 => n35, A => n111, ZN => n109);
   U166 : OAI21_X1 port map( B1 => n35, B2 => n14, A => n111, ZN => n154);
   U167 : XNOR2_X1 port map( A => n109, B => B(42), ZN => n127);
   U168 : NAND2_X1 port map( A1 => n154, A2 => B(42), ZN => n112);
   U169 : OAI21_X1 port map( B1 => n95, B2 => n96, A => n97, ZN => n94);
   U170 : NOR2_X1 port map( A1 => n90, A2 => B(37), ZN => n95);
   U171 : OAI21_X1 port map( B1 => n13, B2 => n96, A => n97, ZN => n155);
   U172 : XNOR2_X1 port map( A => n155, B => B(38), ZN => n131);
   U173 : NAND2_X1 port map( A1 => n155, A2 => B(38), ZN => n99);
   U174 : OAI21_X1 port map( B1 => n80, B2 => n81, A => n82, ZN => n79);
   U175 : NOR2_X1 port map( A1 => n75, A2 => B(33), ZN => n80);
   U176 : OAI21_X1 port map( B1 => n81, B2 => n34, A => n82, ZN => n156);
   U177 : XNOR2_X1 port map( A => B(34), B => n33, ZN => n135);
   U178 : NAND2_X1 port map( A1 => n156, A2 => B(34), ZN => n84);
   U179 : NAND2_X1 port map( A1 => n49, A2 => B(30), ZN => n69);
   U180 : OAI21_X1 port map( B1 => n50, B2 => B(30), A => A(30), ZN => n70);
   U181 : XNOR2_X1 port map( A => n6, B => B(30), ZN => n139);
   U182 : OAI21_X1 port map( B1 => n55, B2 => n56, A => n57, ZN => n54);
   U183 : XNOR2_X1 port map( A => n157, B => n116, ZN => n142);
   U184 : NAND2_X1 port map( A1 => n11, A2 => B(27), ZN => n60);
   U185 : NOR2_X1 port map( A1 => B(26), A2 => n51, ZN => n55);
   U186 : OAI21_X1 port map( B1 => n30, B2 => n56, A => n57, ZN => n157);
   U187 : OAI21_X1 port map( B1 => n45, B2 => n59, A => n60, ZN => n58);
   U188 : XNOR2_X1 port map( A => n158, B => n117, ZN => n141);
   U189 : NAND2_X1 port map( A1 => n158, A2 => B(28), ZN => n64);
   U190 : NOR2_X1 port map( A1 => n58, A2 => B(28), ZN => n62);
   U191 : OAI21_X1 port map( B1 => n59, B2 => n45, A => n60, ZN => n158);
   U192 : XNOR2_X1 port map( A => net73431, B => net73363, ZN => n126);
   U193 : NOR2_X1 port map( A1 => B(40), A2 => n101, ZN => n159);
   U194 : OAI21_X1 port map( B1 => n102, B2 => n103, A => n104, ZN => n101);
   U195 : XNOR2_X1 port map( A => n101, B => n123, ZN => n129);
   U196 : NAND2_X1 port map( A1 => n160, A2 => B(40), ZN => n108);
   U197 : NOR2_X1 port map( A1 => B(39), A2 => n98, ZN => n102);
   U198 : OAI21_X1 port map( B1 => n102, B2 => n103, A => n104, ZN => n160);
   U199 : NOR2_X1 port map( A1 => n162, A2 => B(36), ZN => n161);
   U200 : OAI21_X1 port map( B1 => n87, B2 => n88, A => n89, ZN => n86);
   U201 : XNOR2_X1 port map( A => n86, B => n121, ZN => n133);
   U202 : NAND2_X1 port map( A1 => n162, A2 => B(36), ZN => n93);
   U203 : OAI21_X1 port map( B1 => n87, B2 => n88, A => n89, ZN => n162);
   U204 : NOR2_X1 port map( A1 => n164, A2 => B(32), ZN => n163);
   U205 : OAI21_X1 port map( B1 => n72, B2 => n73, A => n74, ZN => n71);
   U206 : XNOR2_X1 port map( A => n71, B => n119, ZN => n137);
   U207 : NAND2_X1 port map( A1 => n164, A2 => B(32), ZN => n78);
   U208 : OAI21_X1 port map( B1 => n72, B2 => n73, A => n74, ZN => n164);
   U209 : INV_X1 port map( A => A(29), ZN => n66);
   U210 : XNOR2_X1 port map( A => n125, B => A(51), ZN => SUM(51));
   U211 : NAND2_X1 port map( A1 => n31, A2 => B(43), ZN => net73248);
   U212 : NAND2_X1 port map( A1 => B(39), A2 => n42, ZN => n104);
   U213 : XNOR2_X1 port map( A => n139, B => n169, ZN => SUM(30));
   U214 : NAND2_X1 port map( A1 => B(35), A2 => n83, ZN => n89);
   U215 : NAND2_X1 port map( A1 => B(31), A2 => n68, ZN => n74);
   U216 : INV_X1 port map( A => A(28), ZN => n63);
   U217 : NAND2_X1 port map( A1 => n53, A2 => n52, ZN => n51);
   U218 : NAND2_X1 port map( A1 => n53, A2 => n52, ZN => n165);
   U219 : OAI21_X1 port map( B1 => n32, B2 => n63, A => n64, ZN => n61);
   U220 : OAI21_X1 port map( B1 => n62, B2 => n63, A => n64, ZN => n166);
   U221 : CLKBUF_X1 port map( A => A(29), Z => n167);
   U222 : OAI21_X1 port map( B1 => B(34), B2 => n79, A => A(34), ZN => n85);
   U223 : XNOR2_X1 port map( A => n135, B => n8, ZN => SUM(34));
   U224 : XNOR2_X1 port map( A => n170, B => n132, ZN => SUM(37));
   U225 : INV_X1 port map( A => A(37), ZN => n96);
   U226 : OAI21_X1 port map( B1 => n94, B2 => B(38), A => A(38), ZN => n100);
   U227 : XNOR2_X1 port map( A => n131, B => n15, ZN => SUM(38));
   U228 : XNOR2_X1 port map( A => n148, B => B(41), ZN => n128);
   U229 : INV_X1 port map( A => A(41), ZN => n110);
   U230 : INV_X1 port map( A => n110, ZN => n168);
   U231 : XNOR2_X1 port map( A => n152, B => B(33), ZN => n136);
   U232 : XNOR2_X1 port map( A => net73382, B => net73576, ZN => SUM(45));
   U233 : XNOR2_X1 port map( A => B(37), B => n150, ZN => n132);
   U234 : XNOR2_X1 port map( A => carry_25_port, B => B(25), ZN => n144);
   U235 : XNOR2_X1 port map( A => n136, B => n40, ZN => SUM(33));
   U236 : INV_X1 port map( A => A(33), ZN => n81);
   U237 : XNOR2_X1 port map( A => n43, B => n127, ZN => SUM(42));
   U238 : INV_X1 port map( A => A(35), ZN => n88);
   U239 : XNOR2_X1 port map( A => n128, B => n168, ZN => SUM(41));
   U240 : INV_X1 port map( A => A(39), ZN => n103);
   U241 : CLKBUF_X1 port map( A => A(30), Z => n169);
   U242 : XNOR2_X1 port map( A => n140, B => n167, ZN => SUM(29));
   U243 : NAND2_X1 port map( A1 => B(37), A2 => n151, ZN => n97);
   U244 : INV_X1 port map( A => A(26), ZN => n56);
   U245 : XNOR2_X1 port map( A => n137, B => n9, ZN => SUM(32));
   U246 : NAND2_X1 port map( A1 => n70, A2 => n69, ZN => n68);
   U247 : INV_X1 port map( A => n96, ZN => n170);
   U248 : XNOR2_X1 port map( A => n133, B => n92, ZN => SUM(36));
   U249 : OAI21_X1 port map( B1 => n154, B2 => B(42), A => A(42), ZN => n113);
   U250 : XNOR2_X1 port map( A => n129, B => n46, ZN => SUM(40));
   U251 : INV_X1 port map( A => A(27), ZN => n59);
   U252 : XNOR2_X1 port map( A => n68, B => n118, ZN => n138);
   U253 : INV_X1 port map( A => A(36), ZN => n92);
   U254 : XOR2_X1 port map( A => n5, B => B(22), Z => n171);
   U255 : XOR2_X1 port map( A => carry_22_port, B => n171, Z => SUM(22));
   U256 : NAND2_X1 port map( A1 => carry_22_port, A2 => n5, ZN => n172);
   U257 : NAND2_X1 port map( A1 => carry_22_port, A2 => B(22), ZN => n173);
   U258 : NAND2_X1 port map( A1 => A(22), A2 => B(22), ZN => n174);
   U259 : NAND3_X1 port map( A1 => n172, A2 => n173, A3 => n174, ZN => 
                           carry_23_port);
   U260 : XOR2_X1 port map( A => A(55), B => B(55), Z => n175);
   U261 : XOR2_X1 port map( A => carry_55_port, B => n175, Z => SUM(55));
   U262 : NAND2_X1 port map( A1 => carry_53_port, A2 => B(53), ZN => n176);
   U263 : NAND3_X1 port map( A1 => n184, A2 => n176, A3 => n186, ZN => n177);
   U264 : NAND3_X1 port map( A1 => n176, A2 => n184, A3 => n186, ZN => n178);
   U265 : NAND2_X1 port map( A1 => n178, A2 => A(54), ZN => n179);
   U266 : NAND2_X1 port map( A1 => carry_54_port, A2 => B(54), ZN => n180);
   U267 : NAND2_X1 port map( A1 => A(54), A2 => B(54), ZN => n181);
   U268 : NAND3_X1 port map( A1 => n179, A2 => n180, A3 => n181, ZN => 
                           carry_55_port);
   U269 : NAND3_X1 port map( A1 => net46025, A2 => net46026, A3 => n183, ZN => 
                           n182);
   U270 : NAND2_X1 port map( A1 => A(52), A2 => B(52), ZN => n183);
   U271 : NAND3_X1 port map( A1 => net46026, A2 => net46025, A3 => n183, ZN => 
                           carry_53_port);
   U272 : NAND2_X1 port map( A1 => n182, A2 => n16, ZN => n184);
   U273 : NAND2_X1 port map( A1 => carry_53_port, A2 => B(53), ZN => n185);
   U274 : NAND2_X1 port map( A1 => A(53), A2 => B(53), ZN => n186);
   U275 : NAND3_X1 port map( A1 => n184, A2 => n185, A3 => n186, ZN => 
                           carry_54_port);
   U276 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n1);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT54_DW01_add_0 is

   port( A, B : in std_logic_vector (53 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (53 downto 0);  CO : out std_logic);

end RCA_NBIT54_DW01_add_0;

architecture SYN_rpl of RCA_NBIT54_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_53_port, carry_52_port, carry_51_port, carry_50_port, 
      carry_16_port, carry_15_port, carry_14_port, carry_13_port, carry_12_port
      , carry_11_port, carry_10_port, carry_9_port, carry_8_port, carry_7_port,
      carry_6_port, carry_5_port, carry_4_port, carry_3_port, carry_2_port, n1,
      net44085, net44084, net47540, carry_49_port, carry_48_port, net65737, 
      net65698, net65682, net65671, net65600, net65599, net65525, net65524, 
      net65505, net65710, net65678, carry_47_port, carry_46_port, net65743, 
      net65520, net65519, net65518, net65718, net65717, net65511, net65697, 
      net79733, net65598, net76626, net73574, net65679, net65675, net65674, 
      net73529, net65681, net65606, net65604, net65603, n3, n4, n5, n6, n7, n8,
      n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
      n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67
      , n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, 
      n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96
      , n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180 : 
      std_logic;

begin
   
   U1_52 : FA_X1 port map( A => A(52), B => B(52), CI => carry_52_port, CO => 
                           carry_53_port, S => SUM(52));
   U1_50 : FA_X1 port map( A => A(50), B => B(50), CI => carry_50_port, CO => 
                           carry_51_port, S => SUM(50));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1_48 : FA_X1 port map( A => A(48), B => B(48), CI => carry_48_port, CO => 
                           carry_49_port, S => SUM(48));
   U1_47 : FA_X1 port map( A => A(47), B => B(47), CI => carry_47_port, CO => 
                           carry_48_port, S => SUM(47));
   U1_46 : FA_X1 port map( A => A(46), B => B(46), CI => carry_46_port, CO => 
                           carry_47_port, S => SUM(46));
   U1 : CLKBUF_X1 port map( A => A(21), Z => n3);
   U3 : CLKBUF_X1 port map( A => n31, Z => n6);
   U4 : CLKBUF_X1 port map( A => A(20), Z => n4);
   U5 : CLKBUF_X1 port map( A => A(24), Z => n32);
   U6 : XNOR2_X1 port map( A => carry_53_port, B => n5, ZN => SUM(53));
   U7 : XNOR2_X1 port map( A => A(53), B => B(53), ZN => n5);
   U8 : CLKBUF_X1 port map( A => n151, Z => n8);
   U9 : BUF_X1 port map( A => A(26), Z => n28);
   U10 : NOR2_X1 port map( A1 => B(38), A2 => n105, ZN => n7);
   U11 : CLKBUF_X1 port map( A => n77, Z => n9);
   U12 : INV_X1 port map( A => B(39), ZN => n124);
   U13 : INV_X1 port map( A => B(43), ZN => net65671);
   U14 : NAND2_X1 port map( A1 => B(20), A2 => n48, ZN => n55);
   U15 : XNOR2_X1 port map( A => B(16), B => carry_16_port, ZN => n148);
   U16 : XNOR2_X1 port map( A => B(17), B => A(17), ZN => n147);
   U17 : NAND2_X1 port map( A1 => n38, A2 => n39, ZN => n37);
   U18 : NAND2_X1 port map( A1 => B(16), A2 => A(16), ZN => n38);
   U19 : OAI21_X1 port map( B1 => A(16), B2 => B(16), A => carry_16_port, ZN =>
                           n39);
   U20 : XNOR2_X1 port map( A => B(18), B => A(18), ZN => n146);
   U21 : OAI21_X1 port map( B1 => n41, B2 => n42, A => n43, ZN => n40);
   U22 : INV_X1 port map( A => A(17), ZN => n42);
   U23 : NAND2_X1 port map( A1 => B(17), A2 => n37, ZN => n43);
   U24 : NOR2_X1 port map( A1 => B(17), A2 => n37, ZN => n41);
   U25 : XNOR2_X1 port map( A => B(19), B => A(19), ZN => n145);
   U26 : OAI21_X1 port map( B1 => n45, B2 => n46, A => n47, ZN => n44);
   U27 : INV_X1 port map( A => A(18), ZN => n46);
   U28 : NAND2_X1 port map( A1 => B(18), A2 => n40, ZN => n47);
   U29 : NOR2_X1 port map( A1 => B(18), A2 => n40, ZN => n45);
   U30 : OAI21_X1 port map( B1 => n49, B2 => n50, A => n51, ZN => n48);
   U31 : INV_X1 port map( A => A(19), ZN => n50);
   U32 : NAND2_X1 port map( A1 => B(19), A2 => n44, ZN => n51);
   U33 : NOR2_X1 port map( A1 => B(19), A2 => n44, ZN => n49);
   U34 : XNOR2_X1 port map( A => B(21), B => n3, ZN => n143);
   U35 : INV_X1 port map( A => B(38), ZN => n123);
   U36 : XNOR2_X1 port map( A => A(16), B => n148, ZN => SUM(16));
   U37 : XNOR2_X1 port map( A => n147, B => n37, ZN => SUM(17));
   U38 : XNOR2_X1 port map( A => n146, B => n40, ZN => SUM(18));
   U39 : XNOR2_X1 port map( A => n145, B => n44, ZN => SUM(19));
   U40 : XNOR2_X1 port map( A => n144, B => n48, ZN => SUM(20));
   U41 : CLKBUF_X1 port map( A => n153, Z => n14);
   U42 : NOR2_X1 port map( A1 => n116, A2 => B(41), ZN => n10);
   U43 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => n56);
   U44 : XNOR2_X1 port map( A => B(20), B => n4, ZN => n144);
   U45 : INV_X1 port map( A => A(20), ZN => n54);
   U46 : NAND2_X1 port map( A1 => B(24), A2 => n156, ZN => n70);
   U47 : CLKBUF_X1 port map( A => carry_49_port, Z => net47540);
   U48 : AND3_X1 port map( A1 => n92, A2 => n91, A3 => n11, ZN => n94);
   U49 : INV_X1 port map( A => B(34), ZN => n11);
   U50 : XNOR2_X1 port map( A => net65603, B => B(44), ZN => net65681);
   U51 : XNOR2_X1 port map( A => net65681, B => net73574, ZN => SUM(44));
   U52 : OAI21_X1 port map( B1 => net65604, B2 => n12, A => net65606, ZN => 
                           net65603);
   U53 : NOR2_X1 port map( A1 => B(44), A2 => net65603, ZN => net65674);
   U54 : INV_X1 port map( A => A(43), ZN => n12);
   U55 : XNOR2_X1 port map( A => n12, B => net65682, ZN => SUM(43));
   U56 : OAI21_X1 port map( B1 => n13, B2 => n12, A => net65606, ZN => net73529
                           );
   U57 : NOR2_X1 port map( A1 => net65598, A2 => B(43), ZN => net65604);
   U58 : NAND2_X1 port map( A1 => net73529, A2 => B(44), ZN => net65679);
   U59 : NOR2_X1 port map( A1 => net73529, A2 => B(44), ZN => net76626);
   U60 : NOR2_X1 port map( A1 => B(43), A2 => net65598, ZN => n13);
   U61 : NAND2_X1 port map( A1 => net65598, A2 => B(43), ZN => net65606);
   U62 : INV_X1 port map( A => net65675, ZN => net73574);
   U63 : INV_X1 port map( A => A(44), ZN => net65675);
   U64 : OAI21_X1 port map( B1 => net65675, B2 => net65674, A => net65679, ZN 
                           => net65710);
   U65 : OAI21_X1 port map( B1 => net76626, B2 => net65675, A => net65679, ZN 
                           => net65678);
   U66 : NAND2_X1 port map( A1 => net65600, A2 => net65599, ZN => net65598);
   U67 : NAND2_X1 port map( A1 => net65600, A2 => net65599, ZN => net79733);
   U68 : NOR2_X1 port map( A1 => B(30), A2 => n77, ZN => n15);
   U69 : NAND2_X1 port map( A1 => B(28), A2 => net65717, ZN => net65520);
   U70 : CLKBUF_X1 port map( A => n158, Z => n16);
   U71 : CLKBUF_X1 port map( A => n159, Z => n17);
   U72 : NAND2_X1 port map( A1 => B(36), A2 => n152, ZN => n104);
   U73 : NAND2_X1 port map( A1 => n154, A2 => B(32), ZN => n89);
   U74 : XNOR2_X1 port map( A => n143, B => n161, ZN => SUM(21));
   U75 : NAND2_X1 port map( A1 => B(21), A2 => n161, ZN => n57);
   U76 : CLKBUF_X1 port map( A => A(42), Z => n18);
   U77 : INV_X1 port map( A => n118, ZN => n19);
   U78 : NAND2_X1 port map( A1 => n164, A2 => B(40), ZN => n20);
   U79 : BUF_X1 port map( A => A(45), Z => n21);
   U80 : NAND2_X1 port map( A1 => net65525, A2 => net65524, ZN => n77);
   U81 : NAND2_X1 port map( A1 => n91, A2 => n92, ZN => n90);
   U82 : NAND2_X1 port map( A1 => n72, A2 => n73, ZN => n71);
   U83 : OAI21_X1 port map( B1 => B(21), B2 => n52, A => A(21), ZN => n58);
   U84 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => n22);
   U85 : CLKBUF_X1 port map( A => A(41), Z => n23);
   U86 : INV_X1 port map( A => A(40), ZN => n118);
   U87 : INV_X1 port map( A => A(38), ZN => n110);
   U88 : XNOR2_X1 port map( A => A(28), B => B(28), ZN => net65697);
   U89 : XNOR2_X1 port map( A => net65697, B => net65511, ZN => SUM(28));
   U90 : NOR2_X1 port map( A1 => B(28), A2 => net65718, ZN => net65743);
   U91 : NOR2_X1 port map( A1 => net65511, A2 => B(28), ZN => net65518);
   U92 : OAI21_X1 port map( B1 => n25, B2 => n24, A => n26, ZN => net65718);
   U93 : INV_X1 port map( A => A(27), ZN => n25);
   U94 : OAI21_X1 port map( B1 => n27, B2 => n25, A => n26, ZN => net65717);
   U95 : OAI21_X1 port map( B1 => n24, B2 => n25, A => n26, ZN => net65511);
   U96 : NOR2_X1 port map( A1 => net65505, A2 => B(27), ZN => n24);
   U97 : NAND2_X1 port map( A1 => net65505, A2 => B(27), ZN => n26);
   U98 : XNOR2_X1 port map( A => A(27), B => B(27), ZN => net65698);
   U99 : NOR2_X1 port map( A1 => B(27), A2 => net65737, ZN => n27);
   U100 : XNOR2_X1 port map( A => n30, B => n6, ZN => SUM(29));
   U101 : XNOR2_X1 port map( A => A(29), B => B(29), ZN => n30);
   U102 : OAI21_X1 port map( B1 => net65743, B2 => net65519, A => net65520, ZN 
                           => n31);
   U103 : NAND2_X1 port map( A1 => n31, A2 => B(29), ZN => net65524);
   U104 : INV_X1 port map( A => A(28), ZN => net65519);
   U105 : OAI21_X1 port map( B1 => net65518, B2 => net65519, A => net65520, ZN 
                           => n29);
   U106 : OAI21_X1 port map( B1 => B(29), B2 => n29, A => A(29), ZN => net65525
                           );
   U107 : INV_X1 port map( A => A(45), ZN => n33);
   U108 : XNOR2_X1 port map( A => net79733, B => net65671, ZN => net65682);
   U109 : OAI21_X1 port map( B1 => n34, B2 => n33, A => n35, ZN => 
                           carry_46_port);
   U110 : NAND2_X1 port map( A1 => net65678, A2 => B(45), ZN => n35);
   U111 : NOR2_X1 port map( A1 => net65678, A2 => B(45), ZN => n34);
   U112 : XNOR2_X1 port map( A => net65710, B => B(45), ZN => n36);
   U113 : XNOR2_X1 port map( A => n36, B => n21, ZN => SUM(45));
   U114 : XNOR2_X1 port map( A => n129, B => n110, ZN => SUM(38));
   U115 : XNOR2_X1 port map( A => n114, B => n128, ZN => SUM(39));
   U116 : NOR2_X1 port map( A1 => n112, A2 => B(40), ZN => n117);
   U117 : OAI21_X1 port map( B1 => n117, B2 => n118, A => n20, ZN => n116);
   U118 : OAI21_X1 port map( B1 => n118, B2 => n117, A => n20, ZN => n149);
   U119 : OAI21_X1 port map( B1 => n163, B2 => n118, A => n20, ZN => n150);
   U120 : NOR2_X1 port map( A1 => n93, A2 => B(35), ZN => n98);
   U121 : OAI21_X1 port map( B1 => n98, B2 => n99, A => n100, ZN => n97);
   U122 : OAI21_X1 port map( B1 => n98, B2 => n99, A => n100, ZN => n151);
   U123 : OAI21_X1 port map( B1 => n165, B2 => n99, A => n100, ZN => n152);
   U124 : NOR2_X1 port map( A1 => n78, A2 => B(31), ZN => n83);
   U125 : OAI21_X1 port map( B1 => n83, B2 => n84, A => n85, ZN => n82);
   U126 : OAI21_X1 port map( B1 => n83, B2 => n84, A => n85, ZN => n153);
   U127 : OAI21_X1 port map( B1 => n167, B2 => n84, A => n85, ZN => n154);
   U128 : NOR2_X1 port map( A1 => n59, A2 => B(23), ZN => n64);
   U129 : OAI21_X1 port map( B1 => n64, B2 => n65, A => n66, ZN => n63);
   U130 : OAI21_X1 port map( B1 => n64, B2 => n65, A => n66, ZN => n155);
   U131 : OAI21_X1 port map( B1 => n169, B2 => n65, A => n66, ZN => n156);
   U132 : NOR2_X1 port map( A1 => B(41), A2 => n116, ZN => n120);
   U133 : OAI21_X1 port map( B1 => n120, B2 => n121, A => n122, ZN => n119);
   U134 : NOR2_X1 port map( A1 => n97, A2 => B(36), ZN => n102);
   U135 : OAI21_X1 port map( B1 => n102, B2 => n103, A => n104, ZN => n101);
   U136 : OAI21_X1 port map( B1 => n171, B2 => n103, A => n104, ZN => n158);
   U137 : XNOR2_X1 port map( A => n130, B => n16, ZN => SUM(37));
   U138 : NAND2_X1 port map( A1 => n158, A2 => B(37), ZN => n106);
   U139 : NOR2_X1 port map( A1 => n82, A2 => B(32), ZN => n87);
   U140 : OAI21_X1 port map( B1 => n87, B2 => n88, A => n89, ZN => n86);
   U141 : OAI21_X1 port map( B1 => n172, B2 => n88, A => n89, ZN => n159);
   U142 : XNOR2_X1 port map( A => n134, B => n17, ZN => SUM(33));
   U143 : NAND2_X1 port map( A1 => n159, A2 => B(33), ZN => n91);
   U144 : NOR2_X1 port map( A1 => n63, A2 => B(24), ZN => n68);
   U145 : OAI21_X1 port map( B1 => n68, B2 => n69, A => n70, ZN => n67);
   U146 : OAI21_X1 port map( B1 => n173, B2 => n69, A => n70, ZN => n160);
   U147 : XNOR2_X1 port map( A => n139, B => n160, ZN => SUM(25));
   U148 : NAND2_X1 port map( A1 => n160, A2 => B(25), ZN => n72);
   U149 : NOR2_X1 port map( A1 => B(20), A2 => n48, ZN => n53);
   U150 : OAI21_X1 port map( B1 => n53, B2 => n54, A => n55, ZN => n52);
   U151 : OAI21_X1 port map( B1 => n53, B2 => n54, A => n55, ZN => n161);
   U152 : OAI21_X1 port map( B1 => n109, B2 => n110, A => n111, ZN => n108);
   U153 : XNOR2_X1 port map( A => n162, B => n124, ZN => n128);
   U154 : NAND2_X1 port map( A1 => n108, A2 => B(39), ZN => n115);
   U155 : NOR2_X1 port map( A1 => n108, A2 => B(39), ZN => n113);
   U156 : NOR2_X1 port map( A1 => n22, A2 => B(38), ZN => n109);
   U157 : OAI21_X1 port map( B1 => n110, B2 => n7, A => n111, ZN => n162);
   U158 : NOR2_X1 port map( A1 => B(40), A2 => n164, ZN => n163);
   U159 : OAI21_X1 port map( B1 => n113, B2 => n114, A => n115, ZN => n112);
   U160 : XNOR2_X1 port map( A => n112, B => B(40), ZN => n127);
   U161 : OAI21_X1 port map( B1 => n174, B2 => n114, A => n115, ZN => n164);
   U162 : NOR2_X1 port map( A1 => B(35), A2 => n166, ZN => n165);
   U163 : OAI21_X1 port map( B1 => n94, B2 => n95, A => n96, ZN => n93);
   U164 : OAI21_X1 port map( B1 => n94, B2 => n95, A => n96, ZN => n166);
   U165 : NAND2_X1 port map( A1 => n93, A2 => B(35), ZN => n100);
   U166 : NOR2_X1 port map( A1 => B(31), A2 => n168, ZN => n167);
   U167 : NOR2_X1 port map( A1 => n77, A2 => B(30), ZN => n79);
   U168 : OAI21_X1 port map( B1 => n79, B2 => n80, A => n81, ZN => n78);
   U169 : OAI21_X1 port map( B1 => n15, B2 => n80, A => n81, ZN => n168);
   U170 : NAND2_X1 port map( A1 => n78, A2 => B(31), ZN => n85);
   U171 : NOR2_X1 port map( A1 => n71, A2 => B(26), ZN => n74);
   U172 : OAI21_X1 port map( B1 => n74, B2 => n75, A => n76, ZN => net65505);
   U173 : OAI21_X1 port map( B1 => n75, B2 => n74, A => n76, ZN => net65737);
   U174 : NOR2_X1 port map( A1 => B(23), A2 => n170, ZN => n169);
   U175 : NOR2_X1 port map( A1 => B(22), A2 => n56, ZN => n60);
   U176 : OAI21_X1 port map( B1 => n60, B2 => n61, A => n62, ZN => n59);
   U177 : OAI21_X1 port map( B1 => n60, B2 => n61, A => n62, ZN => n170);
   U178 : NAND2_X1 port map( A1 => n59, A2 => B(23), ZN => n66);
   U179 : XNOR2_X1 port map( A => n127, B => n19, ZN => SUM(40));
   U180 : NAND2_X1 port map( A1 => B(34), A2 => n90, ZN => n96);
   U181 : NAND2_X1 port map( A1 => n77, A2 => B(30), ZN => n81);
   U182 : NAND2_X1 port map( A1 => n71, A2 => B(26), ZN => n76);
   U183 : NAND2_X1 port map( A1 => B(22), A2 => n56, ZN => n62);
   U184 : NOR2_X1 port map( A1 => n151, A2 => B(36), ZN => n171);
   U185 : XNOR2_X1 port map( A => n132, B => n166, ZN => SUM(35));
   U186 : NOR2_X1 port map( A1 => n153, A2 => B(32), ZN => n172);
   U187 : XNOR2_X1 port map( A => n136, B => n168, ZN => SUM(31));
   U188 : XNOR2_X1 port map( A => net65698, B => net65737, ZN => SUM(27));
   U189 : NOR2_X1 port map( A1 => B(24), A2 => n63, ZN => n173);
   U190 : XNOR2_X1 port map( A => n141, B => n170, ZN => SUM(23));
   U191 : NAND2_X1 port map( A1 => n107, A2 => n106, ZN => n105);
   U192 : XNOR2_X1 port map( A => n105, B => n123, ZN => n129);
   U193 : NAND2_X1 port map( A1 => n22, A2 => B(38), ZN => n111);
   U194 : OAI21_X1 port map( B1 => n10, B2 => n121, A => n122, ZN => n157);
   U195 : XNOR2_X1 port map( A => n119, B => B(42), ZN => n125);
   U196 : NAND2_X1 port map( A1 => n157, A2 => B(42), ZN => net65599);
   U197 : NOR2_X1 port map( A1 => B(39), A2 => n108, ZN => n174);
   U198 : XNOR2_X1 port map( A => n149, B => B(41), ZN => n126);
   U199 : XNOR2_X1 port map( A => A(37), B => B(37), ZN => n130);
   U200 : OAI21_X1 port map( B1 => n101, B2 => B(37), A => A(37), ZN => n107);
   U201 : XNOR2_X1 port map( A => A(36), B => B(36), ZN => n131);
   U202 : INV_X1 port map( A => A(36), ZN => n103);
   U203 : XNOR2_X1 port map( A => A(32), B => B(32), ZN => n135);
   U204 : INV_X1 port map( A => A(32), ZN => n88);
   U205 : XNOR2_X1 port map( A => A(24), B => B(24), ZN => n140);
   U206 : INV_X1 port map( A => n32, ZN => n69);
   U207 : XNOR2_X1 port map( A => A(34), B => B(34), ZN => n133);
   U208 : INV_X1 port map( A => A(34), ZN => n95);
   U209 : XNOR2_X1 port map( A => A(30), B => B(30), ZN => n137);
   U210 : INV_X1 port map( A => A(30), ZN => n80);
   U211 : XNOR2_X1 port map( A => A(26), B => B(26), ZN => n138);
   U212 : INV_X1 port map( A => n28, ZN => n75);
   U213 : XNOR2_X1 port map( A => n125, B => n18, ZN => SUM(42));
   U214 : XNOR2_X1 port map( A => B(22), B => A(22), ZN => n142);
   U215 : INV_X1 port map( A => A(22), ZN => n61);
   U216 : XNOR2_X1 port map( A => A(35), B => B(35), ZN => n132);
   U217 : XNOR2_X1 port map( A => A(31), B => B(31), ZN => n136);
   U218 : XNOR2_X1 port map( A => A(23), B => B(23), ZN => n141);
   U219 : XNOR2_X1 port map( A => A(33), B => B(33), ZN => n134);
   U220 : XNOR2_X1 port map( A => A(25), B => B(25), ZN => n139);
   U221 : INV_X1 port map( A => A(39), ZN => n114);
   U222 : OAI21_X1 port map( B1 => n157, B2 => B(42), A => A(42), ZN => 
                           net65600);
   U223 : XNOR2_X1 port map( A => n126, B => n23, ZN => SUM(41));
   U224 : XNOR2_X1 port map( A => n131, B => n8, ZN => SUM(36));
   U225 : XNOR2_X1 port map( A => n135, B => n14, ZN => SUM(32));
   U226 : XNOR2_X1 port map( A => n140, B => n155, ZN => SUM(24));
   U227 : XNOR2_X1 port map( A => n133, B => n90, ZN => SUM(34));
   U228 : XNOR2_X1 port map( A => n137, B => n9, ZN => SUM(30));
   U229 : XNOR2_X1 port map( A => n138, B => n71, ZN => SUM(26));
   U230 : INV_X1 port map( A => A(41), ZN => n121);
   U231 : XNOR2_X1 port map( A => n142, B => n56, ZN => SUM(22));
   U232 : INV_X1 port map( A => A(35), ZN => n99);
   U233 : INV_X1 port map( A => A(31), ZN => n84);
   U234 : INV_X1 port map( A => A(23), ZN => n65);
   U235 : OAI21_X1 port map( B1 => n86, B2 => B(33), A => A(33), ZN => n92);
   U236 : OAI21_X1 port map( B1 => B(25), B2 => n67, A => A(25), ZN => n73);
   U237 : NAND2_X1 port map( A1 => B(41), A2 => n150, ZN => n122);
   U238 : NAND2_X1 port map( A1 => carry_49_port, A2 => B(49), ZN => net44085);
   U239 : NAND2_X1 port map( A1 => carry_49_port, A2 => A(49), ZN => net44084);
   U240 : XOR2_X1 port map( A => A(49), B => B(49), Z => n175);
   U241 : XOR2_X1 port map( A => net47540, B => n175, Z => SUM(49));
   U242 : NAND2_X1 port map( A1 => A(49), A2 => B(49), ZN => n176);
   U243 : NAND3_X1 port map( A1 => net44084, A2 => net44085, A3 => n176, ZN => 
                           carry_50_port);
   U244 : XOR2_X1 port map( A => A(51), B => B(51), Z => n177);
   U245 : XOR2_X1 port map( A => carry_51_port, B => n177, Z => SUM(51));
   U246 : NAND2_X1 port map( A1 => carry_51_port, A2 => A(51), ZN => n178);
   U247 : NAND2_X1 port map( A1 => carry_51_port, A2 => B(51), ZN => n179);
   U248 : NAND2_X1 port map( A1 => A(51), A2 => B(51), ZN => n180);
   U249 : NAND3_X1 port map( A1 => n178, A2 => n179, A3 => n180, ZN => 
                           carry_52_port);
   U250 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n1);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT52_DW01_add_0 is

   port( A, B : in std_logic_vector (51 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (51 downto 0);  CO : out std_logic);

end RCA_NBIT52_DW01_add_0;

architecture SYN_rpl of RCA_NBIT52_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_51_port, carry_50_port, carry_19_port, carry_18_port, 
      carry_17_port, carry_16_port, carry_15_port, carry_14_port, carry_13_port
      , carry_12_port, carry_11_port, carry_10_port, carry_9_port, carry_8_port
      , carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port, 
      carry_2_port, n1, net42107, net42106, carry_49_port, carry_48_port, 
      net63168, net63167, net69343, net69305, net69304, net69278, net69277, 
      net69276, net69176, net69104, net69103, net69084, net69414, net69331, 
      net69312, net69311, net69098, net69097, net69096, net69095, net69332, 
      net69089, net69293, net73628, net73640, net79647, net69336, net69181, 
      net69275, net69193, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, 
      n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29
      , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
      n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58
      , n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, 
      n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, 
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, 
      n198, n199, n200, n201, n202, n203, n204 : std_logic;

begin
   
   U1_50 : FA_X1 port map( A => A(50), B => B(50), CI => carry_50_port, CO => 
                           carry_51_port, S => SUM(50));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1_48 : FA_X1 port map( A => A(48), B => B(48), CI => carry_48_port, CO => 
                           carry_49_port, S => SUM(48));
   U1 : NOR2_X1 port map( A1 => B(23), A2 => n77, ZN => n3);
   U3 : CLKBUF_X1 port map( A => n181, Z => n4);
   U4 : NOR2_X1 port map( A1 => B(21), A2 => n70, ZN => n5);
   U5 : CLKBUF_X1 port map( A => n113, Z => n6);
   U6 : CLKBUF_X1 port map( A => A(30), Z => n7);
   U7 : CLKBUF_X1 port map( A => n77, Z => n8);
   U8 : NOR2_X1 port map( A1 => n176, A2 => B(37), ZN => n9);
   U9 : NAND2_X1 port map( A1 => n110, A2 => n109, ZN => n10);
   U10 : INV_X1 port map( A => n103, ZN => n11);
   U11 : INV_X1 port map( A => B(19), ZN => n68);
   U12 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => n30);
   U13 : NOR2_X1 port map( A1 => B(45), A2 => B(44), ZN => n26);
   U14 : INV_X1 port map( A => B(40), ZN => n145);
   U15 : INV_X1 port map( A => B(43), ZN => n36);
   U16 : INV_X1 port map( A => B(47), ZN => n147);
   U17 : INV_X1 port map( A => B(31), ZN => n141);
   U18 : INV_X1 port map( A => B(35), ZN => n142);
   U19 : INV_X1 port map( A => B(36), ZN => n143);
   U20 : INV_X1 port map( A => B(39), ZN => n144);
   U21 : CLKBUF_X1 port map( A => net69084, Z => n12);
   U22 : NOR2_X1 port map( A1 => n176, A2 => B(37), ZN => n13);
   U23 : CLKBUF_X1 port map( A => n87, Z => n14);
   U24 : CLKBUF_X1 port map( A => n180, Z => n15);
   U25 : OAI21_X1 port map( B1 => n126, B2 => n50, A => n127, ZN => n16);
   U26 : INV_X1 port map( A => A(44), ZN => n17);
   U27 : NAND2_X1 port map( A1 => B(21), A2 => n70, ZN => n76);
   U28 : NAND3_X1 port map( A1 => n30, A2 => n29, A3 => A(45), ZN => n20);
   U29 : NAND2_X1 port map( A1 => n31, A2 => net73640, ZN => n28);
   U30 : NAND2_X1 port map( A1 => n25, A2 => n31, ZN => n29);
   U31 : OAI211_X1 port map( C1 => n17, C2 => n32, A => n31, B => n22, ZN => 
                           n19);
   U32 : NAND2_X1 port map( A1 => n20, A2 => n18, ZN => n23);
   U33 : XNOR2_X1 port map( A => n23, B => B(46), ZN => net69275);
   U34 : INV_X1 port map( A => net69336, ZN => n27);
   U35 : NAND2_X1 port map( A1 => n24, A2 => n28, ZN => n18);
   U36 : NAND2_X1 port map( A1 => n18, A2 => n20, ZN => net69193);
   U37 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => net69276);
   U38 : INV_X1 port map( A => B(45), ZN => n22);
   U39 : INV_X1 port map( A => B(44), ZN => n21);
   U40 : XNOR2_X1 port map( A => net69336, B => n21, ZN => net69277);
   U41 : NAND2_X1 port map( A1 => net69181, A2 => B(44), ZN => n31);
   U42 : NOR2_X1 port map( A1 => A(44), A2 => B(45), ZN => n25);
   U43 : INV_X1 port map( A => A(44), ZN => net73640);
   U44 : NOR2_X1 port map( A1 => net69181, A2 => B(44), ZN => n32);
   U45 : NOR2_X1 port map( A1 => n32, A2 => n22, ZN => n24);
   U46 : XNOR2_X1 port map( A => net69275, B => net79647, ZN => SUM(46));
   U47 : NAND2_X1 port map( A1 => net69193, A2 => B(46), ZN => net69305);
   U48 : OAI21_X1 port map( B1 => B(46), B2 => net69193, A => A(46), ZN => 
                           net69304);
   U49 : OAI21_X1 port map( B1 => n37, B2 => n34, A => n35, ZN => net69336);
   U50 : INV_X1 port map( A => A(43), ZN => n34);
   U51 : BUF_X1 port map( A => n34, Z => net73628);
   U52 : OAI21_X1 port map( B1 => n33, B2 => n34, A => n35, ZN => net69181);
   U53 : NOR2_X1 port map( A1 => B(43), A2 => net69414, ZN => n37);
   U54 : NOR2_X1 port map( A1 => B(43), A2 => net69176, ZN => n33);
   U55 : NAND2_X1 port map( A1 => net69176, A2 => B(43), ZN => n35);
   U56 : XNOR2_X1 port map( A => net69414, B => n36, ZN => net69278);
   U57 : BUF_X1 port map( A => A(46), Z => net79647);
   U58 : NOR2_X1 port map( A1 => net69095, A2 => B(29), ZN => n38);
   U59 : NOR2_X1 port map( A1 => B(29), A2 => net69095, ZN => net69343);
   U60 : XNOR2_X1 port map( A => n167, B => n190, ZN => SUM(21));
   U61 : NOR2_X1 port map( A1 => B(36), A2 => n189, ZN => n39);
   U62 : CLKBUF_X1 port map( A => n85, Z => n40);
   U63 : INV_X1 port map( A => n69, ZN => n41);
   U64 : CLKBUF_X1 port map( A => A(19), Z => n42);
   U65 : NOR2_X1 port map( A1 => n94, A2 => B(31), ZN => n43);
   U66 : NAND2_X1 port map( A1 => B(25), A2 => n173, ZN => n91);
   U67 : NOR2_X1 port map( A1 => n195, A2 => B(35), ZN => n44);
   U68 : INV_X1 port map( A => n107, ZN => n45);
   U69 : NAND2_X1 port map( A1 => n124, A2 => n123, ZN => n46);
   U70 : BUF_X1 port map( A => A(38), Z => n53);
   U71 : XNOR2_X1 port map( A => n196, B => n141, ZN => n160);
   U72 : INV_X1 port map( A => A(36), ZN => n47);
   U73 : INV_X1 port map( A => n62, ZN => n48);
   U74 : NOR2_X1 port map( A1 => B(33), A2 => n101, ZN => n49);
   U75 : NAND2_X1 port map( A1 => n78, A2 => n79, ZN => n77);
   U76 : INV_X1 port map( A => A(21), ZN => n75);
   U77 : NOR2_X1 port map( A1 => B(39), A2 => n46, ZN => n50);
   U78 : XNOR2_X1 port map( A => n10, B => n142, ZN => n156);
   U79 : NAND2_X1 port map( A1 => A(47), A2 => B(47), ZN => n139);
   U80 : INV_X1 port map( A => A(47), ZN => n146);
   U81 : OAI21_X1 port map( B1 => n177, B2 => B(42), A => A(42), ZN => n51);
   U82 : NAND2_X1 port map( A1 => n92, A2 => n93, ZN => net69084);
   U83 : XNOR2_X1 port map( A => B(21), B => A(21), ZN => n167);
   U84 : CLKBUF_X1 port map( A => A(42), Z => n52);
   U85 : NAND2_X1 port map( A1 => net69304, A2 => net69305, ZN => n54);
   U86 : INV_X1 port map( A => A(39), ZN => n55);
   U87 : NOR2_X1 port map( A1 => n128, A2 => B(41), ZN => n56);
   U88 : NOR2_X1 port map( A1 => B(41), A2 => n128, ZN => n133);
   U89 : XNOR2_X1 port map( A => A(28), B => B(28), ZN => net69293);
   U90 : XNOR2_X1 port map( A => net69293, B => net69332, ZN => SUM(28));
   U91 : INV_X1 port map( A => A(28), ZN => net69097);
   U92 : NOR2_X1 port map( A1 => B(28), A2 => net69332, ZN => net69331);
   U93 : NOR2_X1 port map( A1 => net69089, A2 => B(28), ZN => net69096);
   U94 : NAND2_X1 port map( A1 => net69089, A2 => B(28), ZN => net69098);
   U95 : OAI21_X1 port map( B1 => n61, B2 => n58, A => n59, ZN => net69332);
   U96 : INV_X1 port map( A => A(27), ZN => n58);
   U97 : OAI21_X1 port map( B1 => n57, B2 => n58, A => n59, ZN => net69089);
   U98 : NOR2_X1 port map( A1 => B(27), A2 => net69084, ZN => n61);
   U99 : XNOR2_X1 port map( A => A(27), B => B(27), ZN => n60);
   U100 : NOR2_X1 port map( A1 => net69084, A2 => B(27), ZN => n57);
   U101 : NAND2_X1 port map( A1 => net69084, A2 => B(27), ZN => n59);
   U102 : XNOR2_X1 port map( A => n60, B => n12, ZN => SUM(27));
   U103 : XNOR2_X1 port map( A => n156, B => n6, ZN => SUM(35));
   U104 : NAND2_X1 port map( A1 => B(29), A2 => net69311, ZN => net69104);
   U105 : INV_X1 port map( A => A(41), ZN => n62);
   U106 : XNOR2_X1 port map( A => net69312, B => B(29), ZN => n63);
   U107 : XNOR2_X1 port map( A => n63, B => n64, ZN => SUM(29));
   U108 : INV_X1 port map( A => A(29), ZN => net69103);
   U109 : INV_X1 port map( A => net69103, ZN => n64);
   U110 : OAI21_X1 port map( B1 => net69097, B2 => net69096, A => net69098, ZN 
                           => net69312);
   U111 : OAI21_X1 port map( B1 => net69331, B2 => net69097, A => net69098, ZN 
                           => net69311);
   U112 : OAI21_X1 port map( B1 => net69096, B2 => net69097, A => net69098, ZN 
                           => net69095);
   U113 : XNOR2_X1 port map( A => n151, B => n130, ZN => SUM(40));
   U114 : XNOR2_X1 port map( A => n160, B => n99, ZN => SUM(31));
   U115 : XNOR2_X1 port map( A => carry_49_port, B => n65, ZN => SUM(49));
   U116 : XNOR2_X1 port map( A => A(49), B => B(49), ZN => n65);
   U117 : OAI21_X1 port map( B1 => n126, B2 => n125, A => n127, ZN => n66);
   U118 : XNOR2_X1 port map( A => net69277, B => n17, ZN => SUM(44));
   U119 : NAND2_X1 port map( A1 => n136, A2 => n51, ZN => net69414);
   U120 : XNOR2_X1 port map( A => n152, B => n55, ZN => SUM(39));
   U121 : INV_X1 port map( A => A(35), ZN => n113);
   U122 : INV_X1 port map( A => A(32), ZN => n103);
   U123 : NAND3_X1 port map( A1 => n138, A2 => n139, A3 => n140, ZN => 
                           carry_48_port);
   U124 : NOR2_X1 port map( A1 => n97, A2 => B(32), ZN => n102);
   U125 : OAI21_X1 port map( B1 => n102, B2 => n103, A => n104, ZN => n101);
   U126 : OAI21_X1 port map( B1 => n103, B2 => n102, A => n104, ZN => n170);
   U127 : OAI21_X1 port map( B1 => n184, B2 => n103, A => n104, ZN => n171);
   U128 : NOR2_X1 port map( A1 => n80, A2 => B(24), ZN => n85);
   U129 : OAI21_X1 port map( B1 => n85, B2 => n86, A => n87, ZN => n84);
   U130 : OAI21_X1 port map( B1 => n40, B2 => n86, A => n14, ZN => n172);
   U131 : OAI21_X1 port map( B1 => n186, B2 => n86, A => n87, ZN => n173);
   U132 : OAI21_X1 port map( B1 => n129, B2 => n130, A => n131, ZN => n128);
   U133 : NOR2_X1 port map( A1 => B(40), A2 => n16, ZN => n129);
   U134 : OAI21_X1 port map( B1 => n188, B2 => n130, A => n131, ZN => n174);
   U135 : OAI21_X1 port map( B1 => n188, B2 => n130, A => n131, ZN => n175);
   U136 : OAI21_X1 port map( B1 => n47, B2 => n116, A => n118, ZN => n115);
   U137 : NAND2_X1 port map( A1 => n115, A2 => B(37), ZN => n121);
   U138 : XNOR2_X1 port map( A => n115, B => B(37), ZN => n154);
   U139 : NOR2_X1 port map( A1 => n189, A2 => B(36), ZN => n116);
   U140 : OAI21_X1 port map( B1 => n117, B2 => n39, A => n118, ZN => n176);
   U141 : OAI21_X1 port map( B1 => n56, B2 => n62, A => n135, ZN => n132);
   U142 : OAI21_X1 port map( B1 => n133, B2 => n134, A => n135, ZN => n177);
   U143 : XNOR2_X1 port map( A => n132, B => B(42), ZN => n149);
   U144 : NAND2_X1 port map( A1 => B(42), A2 => n192, ZN => n136);
   U145 : NOR2_X1 port map( A1 => n101, A2 => B(33), ZN => n106);
   U146 : OAI21_X1 port map( B1 => n49, B2 => n107, A => n108, ZN => n105);
   U147 : OAI21_X1 port map( B1 => n106, B2 => n107, A => n108, ZN => n178);
   U148 : XNOR2_X1 port map( A => n105, B => B(34), ZN => n157);
   U149 : NAND2_X1 port map( A1 => n178, A2 => B(34), ZN => n109);
   U150 : OAI21_X1 port map( B1 => n38, B2 => net69103, A => net69104, ZN => 
                           n179);
   U151 : XNOR2_X1 port map( A => B(30), B => n194, ZN => n161);
   U152 : NAND2_X1 port map( A1 => n179, A2 => B(30), ZN => n95);
   U153 : NOR2_X1 port map( A1 => n84, A2 => B(25), ZN => n89);
   U154 : OAI21_X1 port map( B1 => n89, B2 => n90, A => n91, ZN => n88);
   U155 : OAI21_X1 port map( B1 => n191, B2 => n90, A => n91, ZN => n180);
   U156 : XNOR2_X1 port map( A => n162, B => n15, ZN => SUM(26));
   U157 : NAND2_X1 port map( A1 => B(26), A2 => n180, ZN => n92);
   U158 : NOR2_X1 port map( A1 => B(21), A2 => n70, ZN => n74);
   U159 : OAI21_X1 port map( B1 => n74, B2 => n75, A => n76, ZN => n73);
   U160 : OAI21_X1 port map( B1 => n75, B2 => n5, A => n76, ZN => n181);
   U161 : XNOR2_X1 port map( A => n166, B => n4, ZN => SUM(22));
   U162 : NAND2_X1 port map( A1 => B(22), A2 => n181, ZN => n78);
   U163 : OAI21_X1 port map( B1 => n120, B2 => n13, A => n121, ZN => n119);
   U164 : NAND2_X1 port map( A1 => n182, A2 => B(38), ZN => n123);
   U165 : OAI21_X1 port map( B1 => n182, B2 => B(38), A => A(38), ZN => n124);
   U166 : XNOR2_X1 port map( A => n119, B => B(38), ZN => n153);
   U167 : OAI21_X1 port map( B1 => n9, B2 => n120, A => n121, ZN => n182);
   U168 : INV_X1 port map( A => carry_19_port, ZN => n69);
   U169 : OAI211_X1 port map( C1 => n68, C2 => n69, A => net63167, B => 
                           net63168, ZN => n67);
   U170 : OAI211_X1 port map( C1 => n68, C2 => n69, A => net63168, B => 
                           net63167, ZN => n183);
   U171 : NOR2_X1 port map( A1 => n185, A2 => B(32), ZN => n184);
   U172 : NOR2_X1 port map( A1 => B(31), A2 => n196, ZN => n98);
   U173 : OAI21_X1 port map( B1 => n43, B2 => n99, A => n100, ZN => n97);
   U174 : OAI21_X1 port map( B1 => n98, B2 => n99, A => n100, ZN => n185);
   U175 : NAND2_X1 port map( A1 => n97, A2 => B(32), ZN => n104);
   U176 : NOR2_X1 port map( A1 => B(24), A2 => n187, ZN => n186);
   U177 : NOR2_X1 port map( A1 => B(23), A2 => n77, ZN => n81);
   U178 : OAI21_X1 port map( B1 => n81, B2 => n82, A => n83, ZN => n80);
   U179 : OAI21_X1 port map( B1 => n82, B2 => n3, A => n83, ZN => n187);
   U180 : NAND2_X1 port map( A1 => n80, A2 => B(24), ZN => n87);
   U181 : NOR2_X1 port map( A1 => n16, A2 => B(40), ZN => n188);
   U182 : XNOR2_X1 port map( A => n66, B => n145, ZN => n151);
   U183 : NAND2_X1 port map( A1 => B(40), A2 => n193, ZN => n131);
   U184 : NOR2_X1 port map( A1 => B(39), A2 => n122, ZN => n125);
   U185 : OAI21_X1 port map( B1 => n112, B2 => n113, A => n114, ZN => n111);
   U186 : XNOR2_X1 port map( A => n111, B => n143, ZN => n155);
   U187 : NAND2_X1 port map( A1 => n111, A2 => B(36), ZN => n118);
   U188 : NOR2_X1 port map( A1 => n10, A2 => B(35), ZN => n112);
   U189 : OAI21_X1 port map( B1 => n44, B2 => n113, A => n114, ZN => n189);
   U190 : OAI21_X1 port map( B1 => B(20), B2 => n67, A => A(20), ZN => n72);
   U191 : NAND2_X1 port map( A1 => B(20), A2 => n183, ZN => n71);
   U192 : NAND2_X1 port map( A1 => n72, A2 => n71, ZN => n70);
   U193 : CLKBUF_X1 port map( A => n70, Z => n190);
   U194 : NAND2_X1 port map( A1 => net69305, A2 => net69304, ZN => n168);
   U195 : XNOR2_X1 port map( A => n168, B => n147, ZN => n148);
   U196 : NAND2_X1 port map( A1 => B(47), A2 => n54, ZN => n140);
   U197 : NAND2_X1 port map( A1 => A(47), A2 => n54, ZN => n138);
   U198 : XNOR2_X1 port map( A => n185, B => B(32), ZN => n159);
   U199 : XNOR2_X1 port map( A => n175, B => B(41), ZN => n150);
   U200 : XNOR2_X1 port map( A => n154, B => A(37), ZN => SUM(37));
   U201 : XNOR2_X1 port map( A => n148, B => n146, ZN => SUM(47));
   U202 : XNOR2_X1 port map( A => A(45), B => net69276, ZN => SUM(45));
   U203 : XNOR2_X1 port map( A => n149, B => n52, ZN => SUM(42));
   U204 : NAND2_X1 port map( A1 => n124, A2 => n123, ZN => n122);
   U205 : XNOR2_X1 port map( A => n170, B => B(33), ZN => n158);
   U206 : XNOR2_X1 port map( A => n159, B => n11, ZN => SUM(32));
   U207 : NAND2_X1 port map( A1 => n195, A2 => B(35), ZN => n114);
   U208 : XNOR2_X1 port map( A => A(34), B => n157, ZN => SUM(34));
   U209 : NAND2_X1 port map( A1 => B(23), A2 => n77, ZN => n83);
   U210 : XNOR2_X1 port map( A => n155, B => n117, ZN => SUM(36));
   U211 : NAND2_X1 port map( A1 => n94, A2 => B(31), ZN => n100);
   U212 : NOR2_X1 port map( A1 => n84, A2 => B(25), ZN => n191);
   U213 : XNOR2_X1 port map( A => n164, B => n187, ZN => SUM(24));
   U214 : OAI21_X1 port map( B1 => n177, B2 => B(42), A => A(42), ZN => n137);
   U215 : XNOR2_X1 port map( A => A(20), B => B(20), ZN => n169);
   U216 : XNOR2_X1 port map( A => n7, B => n161, ZN => SUM(30));
   U217 : XNOR2_X1 port map( A => A(25), B => B(25), ZN => n163);
   U218 : INV_X1 port map( A => A(25), ZN => n90);
   U219 : NAND2_X1 port map( A1 => n174, A2 => B(41), ZN => n135);
   U220 : INV_X1 port map( A => A(41), ZN => n134);
   U221 : XNOR2_X1 port map( A => A(23), B => B(23), ZN => n165);
   U222 : INV_X1 port map( A => A(23), ZN => n82);
   U223 : XNOR2_X1 port map( A => A(26), B => B(26), ZN => n162);
   U224 : XNOR2_X1 port map( A => n153, B => n53, ZN => SUM(38));
   U225 : NAND2_X1 port map( A1 => n137, A2 => n136, ZN => net69176);
   U226 : XNOR2_X1 port map( A => A(24), B => B(24), ZN => n164);
   U227 : XNOR2_X1 port map( A => n150, B => n48, ZN => SUM(41));
   U228 : XNOR2_X1 port map( A => A(22), B => B(22), ZN => n166);
   U229 : INV_X1 port map( A => A(33), ZN => n107);
   U230 : INV_X1 port map( A => A(37), ZN => n120);
   U231 : OAI21_X1 port map( B1 => n178, B2 => B(34), A => A(34), ZN => n110);
   U232 : OAI21_X1 port map( B1 => n179, B2 => B(30), A => A(30), ZN => n96);
   U233 : NAND2_X1 port map( A1 => n96, A2 => n95, ZN => n94);
   U234 : INV_X1 port map( A => A(39), ZN => n126);
   U235 : XNOR2_X1 port map( A => n158, B => n45, ZN => SUM(33));
   U236 : XNOR2_X1 port map( A => n46, B => n144, ZN => n152);
   U237 : NAND2_X1 port map( A1 => B(39), A2 => n122, ZN => n127);
   U238 : XNOR2_X1 port map( A => n163, B => n172, ZN => SUM(25));
   U239 : OAI21_X1 port map( B1 => n134, B2 => n56, A => n135, ZN => n192);
   U240 : INV_X1 port map( A => A(31), ZN => n99);
   U241 : OAI21_X1 port map( B1 => B(26), B2 => n88, A => A(26), ZN => n93);
   U242 : XNOR2_X1 port map( A => net69278, B => net73628, ZN => SUM(43));
   U243 : OAI21_X1 port map( B1 => n125, B2 => n55, A => n127, ZN => n193);
   U244 : INV_X1 port map( A => A(36), ZN => n117);
   U245 : INV_X1 port map( A => A(24), ZN => n86);
   U246 : XNOR2_X1 port map( A => n165, B => n8, ZN => SUM(23));
   U247 : XNOR2_X1 port map( A => n183, B => n169, ZN => SUM(20));
   U248 : OAI21_X1 port map( B1 => net69343, B2 => net69103, A => net69104, ZN 
                           => n194);
   U249 : NAND2_X1 port map( A1 => B(33), A2 => n171, ZN => n108);
   U250 : OAI21_X1 port map( B1 => B(22), B2 => n73, A => A(22), ZN => n79);
   U251 : NAND2_X1 port map( A1 => n110, A2 => n109, ZN => n195);
   U252 : NAND2_X1 port map( A1 => n96, A2 => n95, ZN => n196);
   U253 : INV_X1 port map( A => A(40), ZN => n130);
   U254 : CLKBUF_X1 port map( A => A(18), Z => n197);
   U255 : XOR2_X1 port map( A => n41, B => B(19), Z => n198);
   U256 : XOR2_X1 port map( A => n42, B => n198, Z => SUM(19));
   U257 : NAND2_X1 port map( A1 => A(19), A2 => carry_19_port, ZN => net63167);
   U258 : NAND2_X1 port map( A1 => A(19), A2 => B(19), ZN => net63168);
   U259 : XOR2_X1 port map( A => n197, B => B(18), Z => n199);
   U260 : XOR2_X1 port map( A => carry_18_port, B => n199, Z => SUM(18));
   U261 : NAND2_X1 port map( A1 => carry_18_port, A2 => n197, ZN => n200);
   U262 : NAND2_X1 port map( A1 => carry_18_port, A2 => B(18), ZN => n201);
   U263 : NAND2_X1 port map( A1 => A(18), A2 => B(18), ZN => n202);
   U264 : NAND3_X1 port map( A1 => n200, A2 => n201, A3 => n202, ZN => 
                           carry_19_port);
   U265 : NAND2_X1 port map( A1 => carry_49_port, A2 => B(49), ZN => net42107);
   U266 : NAND2_X1 port map( A1 => carry_49_port, A2 => A(49), ZN => net42106);
   U267 : NAND2_X1 port map( A1 => A(49), A2 => B(49), ZN => n203);
   U268 : NAND3_X1 port map( A1 => net42106, A2 => net42107, A3 => n203, ZN => 
                           carry_50_port);
   U269 : XOR2_X2 port map( A => carry_51_port, B => n204, Z => SUM(51));
   U270 : XOR2_X1 port map( A => A(51), B => B(51), Z => n204);
   U271 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n1);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT50_DW01_add_0 is

   port( A, B : in std_logic_vector (49 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (49 downto 0);  CO : out std_logic);

end RCA_NBIT50_DW01_add_0;

architecture SYN_rpl of RCA_NBIT50_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_49_port, carry_48_port, carry_46_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_10_port
      , carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, n1, carry_44_port, 
      carry_16_port, net52609, net52608, net52676, net55502, carry_43_port, 
      carry_42_port, carry_41_port, net63222, net70828, net73512, net73510, 
      net73508, net73507, net73573, net73746, net73785, net52611, net52610, n3,
      n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
      n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92
      , n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, 
      n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, 
      n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, 
      n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, 
      n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
      n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, 
      n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, 
      n178, n179, n180, n181, n182, n183, n184, n185 : std_logic;

begin
   
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_44 : FA_X1 port map( A => A(44), B => B(44), CI => carry_44_port, CO => 
                           net70828, S => SUM(44));
   U1_41 : FA_X1 port map( A => A(41), B => B(41), CI => carry_41_port, CO => 
                           carry_42_port, S => SUM(41));
   U1_43 : FA_X1 port map( A => A(43), B => B(43), CI => carry_43_port, CO => 
                           carry_44_port, S => SUM(43));
   U1_42 : FA_X1 port map( A => A(42), B => B(42), CI => carry_42_port, CO => 
                           carry_43_port, S => SUM(42));
   U1 : CLKBUF_X1 port map( A => n147, Z => n3);
   U3 : NOR2_X1 port map( A1 => n46, A2 => B(23), ZN => n4);
   U4 : CLKBUF_X1 port map( A => A(35), Z => n5);
   U5 : NOR2_X1 port map( A1 => n35, A2 => B(20), ZN => n6);
   U6 : NAND2_X1 port map( A1 => n77, A2 => n78, ZN => n7);
   U7 : AND2_X1 port map( A1 => n8, A2 => n9, ZN => n32);
   U8 : NOR2_X1 port map( A1 => B(18), A2 => n113, ZN => n8);
   U9 : NAND2_X1 port map( A1 => net55502, A2 => n172, ZN => n9);
   U10 : OR2_X2 port map( A1 => n166, A2 => n113, ZN => n30);
   U11 : OAI21_X1 port map( B1 => n84, B2 => n85, A => n86, ZN => n10);
   U12 : OAI21_X1 port map( B1 => n69, B2 => n70, A => n71, ZN => n11);
   U13 : BUF_X1 port map( A => n165, Z => n12);
   U14 : NOR2_X1 port map( A1 => B(27), A2 => n62, ZN => n13);
   U15 : NAND2_X1 port map( A1 => B(18), A2 => n30, ZN => n14);
   U16 : XOR2_X1 port map( A => A(48), B => B(48), Z => n15);
   U17 : XOR2_X1 port map( A => carry_48_port, B => n15, Z => SUM(48));
   U18 : NAND2_X1 port map( A1 => carry_48_port, A2 => A(48), ZN => n16);
   U19 : NAND2_X1 port map( A1 => carry_48_port, A2 => B(48), ZN => n17);
   U20 : NAND2_X1 port map( A1 => A(48), A2 => B(48), ZN => n18);
   U21 : NAND3_X1 port map( A1 => n16, A2 => n17, A3 => n18, ZN => 
                           carry_49_port);
   U22 : INV_X1 port map( A => B(17), ZN => n112);
   U23 : NAND2_X1 port map( A1 => n173, A2 => n176, ZN => n175);
   U24 : INV_X1 port map( A => B(40), ZN => n29);
   U25 : INV_X1 port map( A => B(22), ZN => n48);
   U26 : XNOR2_X1 port map( A => carry_49_port, B => n178, ZN => SUM(49));
   U27 : CLKBUF_X1 port map( A => n43, Z => n167);
   U28 : BUF_X1 port map( A => A(27), Z => n169);
   U29 : BUF_X1 port map( A => n108, Z => n25);
   U30 : BUF_X1 port map( A => n148, Z => n26);
   U31 : NAND2_X1 port map( A1 => B(25), A2 => n146, ZN => n61);
   U32 : NAND2_X1 port map( A1 => B(29), A2 => n144, ZN => n75);
   U33 : INV_X1 port map( A => B(46), ZN => n176);
   U34 : NAND2_X1 port map( A1 => n20, A2 => net70828, ZN => n19);
   U35 : OR2_X1 port map( A1 => A(45), A2 => B(45), ZN => n20);
   U36 : OAI211_X1 port map( C1 => n98, C2 => n99, A => n100, B => n21, ZN => 
                           n22);
   U37 : INV_X1 port map( A => B(37), ZN => n21);
   U38 : INV_X1 port map( A => n22, ZN => n102);
   U39 : CLKBUF_X1 port map( A => A(19), Z => n23);
   U40 : CLKBUF_X1 port map( A => n105, Z => n24);
   U41 : BUF_X1 port map( A => A(31), Z => n168);
   U42 : BUF_X1 port map( A => A(17), Z => n172);
   U43 : OAI21_X1 port map( B1 => n109, B2 => n110, A => n111, ZN => n108);
   U44 : OAI21_X1 port map( B1 => n4, B2 => n52, A => n53, ZN => n27);
   U45 : OAI21_X1 port map( B1 => n89, B2 => n162, A => n90, ZN => n28);
   U46 : INV_X1 port map( A => carry_46_port, ZN => net73785);
   U47 : XNOR2_X1 port map( A => n136, B => n30, ZN => SUM(18));
   U48 : XNOR2_X1 port map( A => B(21), B => A(21), ZN => n133);
   U49 : XNOR2_X1 port map( A => A(22), B => B(22), ZN => n132);
   U50 : NAND2_X1 port map( A1 => n106, A2 => n107, ZN => n105);
   U51 : BUF_X1 port map( A => n50, Z => n157);
   U52 : NAND2_X1 port map( A1 => B(33), A2 => n142, ZN => n90);
   U53 : XNOR2_X1 port map( A => A(46), B => n176, ZN => net73510);
   U54 : XNOR2_X1 port map( A => n129, B => n145, ZN => SUM(25));
   U55 : XNOR2_X1 port map( A => A(40), B => n29, ZN => n179);
   U56 : XNOR2_X1 port map( A => n134, B => n138, ZN => SUM(20));
   U57 : XNOR2_X1 port map( A => n115, B => n24, ZN => SUM(39));
   U58 : XNOR2_X1 port map( A => n117, B => n140, ZN => SUM(37));
   U59 : XNOR2_X1 port map( A => n11, B => n125, ZN => SUM(29));
   U60 : XNOR2_X1 port map( A => n10, B => n121, ZN => SUM(33));
   U61 : XNOR2_X1 port map( A => n127, B => n62, ZN => SUM(27));
   U62 : XNOR2_X1 port map( A => n123, B => n7, ZN => SUM(31));
   U63 : NOR2_X1 port map( A1 => n31, A2 => B(19), ZN => n36);
   U64 : OAI21_X1 port map( B1 => n36, B2 => n37, A => n38, ZN => n35);
   U65 : OAI21_X1 port map( B1 => n37, B2 => n36, A => n38, ZN => n138);
   U66 : OAI21_X1 port map( B1 => n160, B2 => n37, A => n38, ZN => n139);
   U67 : NOR2_X1 port map( A1 => n94, A2 => B(36), ZN => n98);
   U68 : OAI21_X1 port map( B1 => n98, B2 => n99, A => n100, ZN => n140);
   U69 : OAI21_X1 port map( B1 => n158, B2 => n99, A => n100, ZN => n141);
   U70 : NOR2_X1 port map( A1 => n79, A2 => B(32), ZN => n84);
   U71 : OAI21_X1 port map( B1 => n84, B2 => n85, A => n86, ZN => n83);
   U72 : OAI21_X1 port map( B1 => n152, B2 => n85, A => n86, ZN => n142);
   U73 : NOR2_X1 port map( A1 => n65, A2 => B(28), ZN => n69);
   U74 : OAI21_X1 port map( B1 => n69, B2 => n70, A => n71, ZN => n143);
   U75 : OAI21_X1 port map( B1 => n154, B2 => n70, A => n71, ZN => n144);
   U76 : NOR2_X1 port map( A1 => n27, A2 => B(24), ZN => n55);
   U77 : OAI21_X1 port map( B1 => n55, B2 => n56, A => n57, ZN => n54);
   U78 : OAI21_X1 port map( B1 => n55, B2 => n56, A => n57, ZN => n145);
   U79 : OAI21_X1 port map( B1 => n156, B2 => n56, A => n57, ZN => n146);
   U80 : NAND2_X1 port map( A1 => n165, A2 => B(23), ZN => n53);
   U81 : XNOR2_X1 port map( A => n12, B => n131, ZN => SUM(23));
   U82 : NOR2_X1 port map( A1 => n46, A2 => B(23), ZN => n51);
   U83 : NOR2_X1 port map( A1 => n35, A2 => B(20), ZN => n40);
   U84 : OAI21_X1 port map( B1 => n6, B2 => n41, A => n42, ZN => n39);
   U85 : OAI21_X1 port map( B1 => n41, B2 => n40, A => n42, ZN => n147);
   U86 : XNOR2_X1 port map( A => n3, B => n133, ZN => SUM(21));
   U87 : NAND2_X1 port map( A1 => n147, A2 => B(21), ZN => n44);
   U88 : OAI21_X1 port map( B1 => n102, B2 => n103, A => n104, ZN => n101);
   U89 : OAI21_X1 port map( B1 => n102, B2 => n103, A => n104, ZN => n148);
   U90 : XNOR2_X1 port map( A => n116, B => n26, ZN => SUM(38));
   U91 : NAND2_X1 port map( A1 => n148, A2 => B(38), ZN => n106);
   U92 : NOR2_X1 port map( A1 => n83, A2 => B(33), ZN => n88);
   U93 : OAI21_X1 port map( B1 => n88, B2 => n89, A => n90, ZN => n87);
   U94 : OAI21_X1 port map( B1 => n162, B2 => n89, A => n90, ZN => n149);
   U95 : XNOR2_X1 port map( A => n120, B => n28, ZN => SUM(34));
   U96 : NAND2_X1 port map( A1 => B(34), A2 => n149, ZN => n92);
   U97 : NOR2_X1 port map( A1 => n143, A2 => B(29), ZN => n73);
   U98 : OAI21_X1 port map( B1 => n73, B2 => n74, A => n75, ZN => n72);
   U99 : OAI21_X1 port map( B1 => n163, B2 => n74, A => n75, ZN => n150);
   U100 : XNOR2_X1 port map( A => n124, B => n150, ZN => SUM(30));
   U101 : NAND2_X1 port map( A1 => n150, A2 => B(30), ZN => n77);
   U102 : NOR2_X1 port map( A1 => n54, A2 => B(25), ZN => n59);
   U103 : OAI21_X1 port map( B1 => n59, B2 => n60, A => n61, ZN => n58);
   U104 : OAI21_X1 port map( B1 => n164, B2 => n60, A => n61, ZN => n151);
   U105 : XNOR2_X1 port map( A => n128, B => n151, ZN => SUM(26));
   U106 : NAND2_X1 port map( A1 => n151, A2 => B(26), ZN => n63);
   U107 : NOR2_X1 port map( A1 => n153, A2 => B(32), ZN => n152);
   U108 : NOR2_X1 port map( A1 => n76, A2 => B(31), ZN => n80);
   U109 : OAI21_X1 port map( B1 => n80, B2 => n81, A => n82, ZN => n79);
   U110 : OAI21_X1 port map( B1 => n81, B2 => n80, A => n82, ZN => n153);
   U111 : NAND2_X1 port map( A1 => n79, A2 => B(32), ZN => n86);
   U112 : NOR2_X1 port map( A1 => n155, A2 => B(28), ZN => n154);
   U113 : NOR2_X1 port map( A1 => B(27), A2 => n62, ZN => n66);
   U114 : OAI21_X1 port map( B1 => n66, B2 => n67, A => n68, ZN => n65);
   U115 : OAI21_X1 port map( B1 => n67, B2 => n13, A => n68, ZN => n155);
   U116 : NAND2_X1 port map( A1 => n65, A2 => B(28), ZN => n71);
   U117 : NOR2_X1 port map( A1 => B(24), A2 => n27, ZN => n156);
   U118 : OAI21_X1 port map( B1 => n51, B2 => n52, A => n53, ZN => n50);
   U119 : NAND2_X1 port map( A1 => n50, A2 => B(24), ZN => n57);
   U120 : XNOR2_X1 port map( A => n130, B => n157, ZN => SUM(24));
   U121 : NOR2_X1 port map( A1 => B(36), A2 => n159, ZN => n158);
   U122 : OAI21_X1 port map( B1 => n95, B2 => n96, A => n97, ZN => n94);
   U123 : NOR2_X1 port map( A1 => n91, A2 => B(35), ZN => n95);
   U124 : OAI21_X1 port map( B1 => n96, B2 => n95, A => n97, ZN => n159);
   U125 : NAND2_X1 port map( A1 => n94, A2 => B(36), ZN => n100);
   U126 : NOR2_X1 port map( A1 => B(19), A2 => n161, ZN => n160);
   U127 : OAI21_X1 port map( B1 => n32, B2 => n33, A => n34, ZN => n31);
   U128 : OAI21_X1 port map( B1 => n33, B2 => n32, A => n14, ZN => n161);
   U129 : NAND2_X1 port map( A1 => n31, A2 => B(19), ZN => n38);
   U130 : NAND2_X1 port map( A1 => n108, A2 => B(40), ZN => net73508);
   U131 : NAND2_X1 port map( A1 => n171, A2 => n108, ZN => net73507);
   U132 : NOR2_X1 port map( A1 => B(39), A2 => n105, ZN => n109);
   U133 : NAND2_X1 port map( A1 => B(39), A2 => n105, ZN => n111);
   U134 : NAND2_X1 port map( A1 => B(18), A2 => n30, ZN => n34);
   U135 : XNOR2_X1 port map( A => n118, B => n159, ZN => SUM(36));
   U136 : NAND2_X1 port map( A1 => n91, A2 => B(35), ZN => n97);
   U137 : NAND2_X1 port map( A1 => B(31), A2 => n7, ZN => n82);
   U138 : XNOR2_X1 port map( A => n126, B => n155, ZN => SUM(28));
   U139 : NAND2_X1 port map( A1 => B(27), A2 => n62, ZN => n68);
   U140 : NOR2_X1 port map( A1 => n10, A2 => B(33), ZN => n162);
   U141 : XNOR2_X1 port map( A => n122, B => n153, ZN => SUM(32));
   U142 : NOR2_X1 port map( A1 => n11, A2 => B(29), ZN => n163);
   U143 : XNOR2_X1 port map( A => n135, B => n161, ZN => SUM(19));
   U144 : NOR2_X1 port map( A1 => B(25), A2 => n54, ZN => n164);
   U145 : NAND2_X1 port map( A1 => n77, A2 => n78, ZN => n76);
   U146 : NAND2_X1 port map( A1 => n63, A2 => n64, ZN => n62);
   U147 : NAND2_X1 port map( A1 => n92, A2 => n93, ZN => n91);
   U148 : NAND2_X1 port map( A1 => B(20), A2 => n139, ZN => n42);
   U149 : NAND2_X1 port map( A1 => B(37), A2 => n141, ZN => n104);
   U150 : OAI21_X1 port map( B1 => n39, B2 => B(21), A => A(21), ZN => n45);
   U151 : NAND2_X1 port map( A1 => n45, A2 => n44, ZN => n43);
   U152 : NAND2_X1 port map( A1 => A(22), A2 => n43, ZN => n49);
   U153 : XNOR2_X1 port map( A => n132, B => n167, ZN => SUM(22));
   U154 : NOR2_X1 port map( A1 => n43, A2 => A(22), ZN => n47);
   U155 : OAI21_X1 port map( B1 => n47, B2 => n48, A => n49, ZN => n46);
   U156 : OAI21_X1 port map( B1 => n48, B2 => n47, A => n49, ZN => n165);
   U157 : AOI21_X1 port map( B1 => n114, B2 => net52609, A => n112, ZN => n113)
                           ;
   U158 : AND2_X1 port map( A1 => n172, A2 => net55502, ZN => n166);
   U159 : NAND2_X1 port map( A1 => net52610, A2 => net52611, ZN => n137);
   U160 : NOR2_X1 port map( A1 => A(17), A2 => n137, ZN => n114);
   U161 : XNOR2_X1 port map( A => A(35), B => B(35), ZN => n119);
   U162 : INV_X1 port map( A => n5, ZN => n96);
   U163 : XNOR2_X1 port map( A => A(31), B => B(31), ZN => n123);
   U164 : INV_X1 port map( A => n168, ZN => n81);
   U165 : XNOR2_X1 port map( A => A(27), B => B(27), ZN => n127);
   U166 : INV_X1 port map( A => n169, ZN => n67);
   U167 : XNOR2_X1 port map( A => A(25), B => B(25), ZN => n129);
   U168 : INV_X1 port map( A => n170, ZN => n60);
   U169 : XNOR2_X1 port map( A => A(32), B => B(32), ZN => n122);
   U170 : INV_X1 port map( A => A(32), ZN => n85);
   U171 : XNOR2_X1 port map( A => A(18), B => B(18), ZN => n136);
   U172 : INV_X1 port map( A => A(18), ZN => n33);
   U173 : XNOR2_X1 port map( A => A(33), B => B(33), ZN => n121);
   U174 : INV_X1 port map( A => A(33), ZN => n89);
   U175 : XNOR2_X1 port map( A => A(29), B => B(29), ZN => n125);
   U176 : INV_X1 port map( A => A(29), ZN => n74);
   U177 : XNOR2_X1 port map( A => A(36), B => B(36), ZN => n118);
   U178 : INV_X1 port map( A => A(36), ZN => n99);
   U179 : XNOR2_X1 port map( A => A(34), B => B(34), ZN => n120);
   U180 : OAI21_X1 port map( B1 => B(34), B2 => n87, A => A(34), ZN => n93);
   U181 : XNOR2_X1 port map( A => A(30), B => B(30), ZN => n124);
   U182 : OAI21_X1 port map( B1 => B(30), B2 => n72, A => A(30), ZN => n78);
   U183 : XNOR2_X1 port map( A => A(23), B => B(23), ZN => n131);
   U184 : INV_X1 port map( A => A(23), ZN => n52);
   U185 : XNOR2_X1 port map( A => A(20), B => B(20), ZN => n134);
   U186 : INV_X1 port map( A => A(20), ZN => n41);
   U187 : XNOR2_X1 port map( A => A(26), B => B(26), ZN => n128);
   U188 : OAI21_X1 port map( B1 => B(26), B2 => n58, A => A(26), ZN => n64);
   U189 : XNOR2_X1 port map( A => A(28), B => B(28), ZN => n126);
   U190 : INV_X1 port map( A => A(28), ZN => n70);
   U191 : XNOR2_X1 port map( A => A(39), B => B(39), ZN => n115);
   U192 : INV_X1 port map( A => A(39), ZN => n110);
   U193 : XNOR2_X1 port map( A => A(24), B => B(24), ZN => n130);
   U194 : INV_X1 port map( A => A(24), ZN => n56);
   U195 : XNOR2_X1 port map( A => A(19), B => B(19), ZN => n135);
   U196 : INV_X1 port map( A => n23, ZN => n37);
   U197 : XNOR2_X1 port map( A => B(37), B => A(37), ZN => n117);
   U198 : INV_X1 port map( A => A(37), ZN => n103);
   U199 : XNOR2_X1 port map( A => A(38), B => B(38), ZN => n116);
   U200 : OAI21_X1 port map( B1 => B(38), B2 => n101, A => A(38), ZN => n107);
   U201 : XNOR2_X1 port map( A => n119, B => n91, ZN => SUM(35));
   U202 : BUF_X1 port map( A => A(40), Z => n171);
   U203 : CLKBUF_X1 port map( A => A(25), Z => n170);
   U204 : NAND2_X1 port map( A1 => A(16), A2 => B(16), ZN => net52611);
   U205 : NAND3_X1 port map( A1 => net52609, A2 => net52610, A3 => net52611, ZN
                           => net55502);
   U206 : CLKBUF_X1 port map( A => A(16), Z => net52676);
   U207 : XOR2_X1 port map( A => net52676, B => B(16), Z => net52608);
   U208 : NAND2_X1 port map( A1 => carry_16_port, A2 => B(16), ZN => net52610);
   U209 : INV_X1 port map( A => n19, ZN => n177);
   U210 : NAND2_X1 port map( A1 => n19, A2 => n173, ZN => carry_46_port);
   U211 : OAI21_X1 port map( B1 => n177, B2 => n175, A => A(46), ZN => n174);
   U212 : NAND2_X1 port map( A1 => net73512, A2 => n174, ZN => net73573);
   U213 : NAND2_X1 port map( A1 => B(45), A2 => A(45), ZN => n173);
   U214 : XNOR2_X1 port map( A => B(45), B => A(45), ZN => net73746);
   U215 : XNOR2_X1 port map( A => net73785, B => net73510, ZN => SUM(46));
   U216 : XNOR2_X1 port map( A => net70828, B => net73746, ZN => SUM(45));
   U217 : XNOR2_X1 port map( A => A(49), B => B(49), ZN => n178);
   U218 : XOR2_X1 port map( A => n25, B => n179, Z => SUM(40));
   U219 : NAND2_X1 port map( A1 => n171, A2 => B(40), ZN => n180);
   U220 : NAND3_X1 port map( A1 => n180, A2 => net73507, A3 => net73508, ZN => 
                           carry_41_port);
   U221 : NAND2_X1 port map( A1 => carry_46_port, A2 => B(46), ZN => net73512);
   U222 : CLKBUF_X1 port map( A => n172, Z => net63222);
   U223 : XOR2_X1 port map( A => net63222, B => B(17), Z => n181);
   U224 : XOR2_X1 port map( A => net55502, B => n181, Z => SUM(17));
   U225 : XOR2_X1 port map( A => carry_16_port, B => net52608, Z => SUM(16));
   U226 : NAND2_X1 port map( A1 => carry_16_port, A2 => net52676, ZN => 
                           net52609);
   U227 : XOR2_X1 port map( A => A(47), B => B(47), Z => n182);
   U228 : XOR2_X1 port map( A => net73573, B => n182, Z => SUM(47));
   U229 : NAND2_X1 port map( A1 => net73573, A2 => A(47), ZN => n183);
   U230 : NAND2_X1 port map( A1 => net73573, A2 => B(47), ZN => n184);
   U231 : NAND2_X1 port map( A1 => A(47), A2 => B(47), ZN => n185);
   U232 : NAND3_X1 port map( A1 => n183, A2 => n184, A3 => n185, ZN => 
                           carry_48_port);
   U233 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n1);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT48_DW01_add_0 is

   port( A, B : in std_logic_vector (47 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (47 downto 0);  CO : out std_logic);

end RCA_NBIT48_DW01_add_0;

architecture SYN_rpl of RCA_NBIT48_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_47_port, carry_46_port, carry_45_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_10_port
      , carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, n1, net42193, net42192, 
      net42190, carry_44_port, net52615, net52614, net52656, net52655, net52654
      , net62366, net62347, net62331, net62320, net62271, net62270, net62254, 
      net62234, net62232, net62184, net62183, net62178, net62164, net62081, 
      net62080, net62079, net62067, net62058, net62057, net62056, net63145, 
      net63135, net63127, net63126, net63123, net62326, net62072, net63180, 
      net62050, net62356, net62269, net62176, n3, n4, n5, n6, n7, n8, n9, n10, 
      n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25
      , n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, 
      n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54
      , n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, 
      n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83
      , n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, 
      n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, 
      n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
      n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, 
      n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, 
      n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, 
      n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, 
      n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, 
      n182, n183 : std_logic;

begin
   
   U1_46 : FA_X1 port map( A => A(46), B => B(46), CI => carry_46_port, CO => 
                           carry_47_port, S => SUM(46));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : CLKBUF_X1 port map( A => A(15), Z => n3);
   U3 : OAI21_X1 port map( B1 => n68, B2 => n69, A => n70, ZN => n4);
   U4 : NOR2_X1 port map( A1 => B(25), A2 => n71, ZN => n5);
   U5 : CLKBUF_X1 port map( A => A(36), Z => n6);
   U6 : AND2_X1 port map( A1 => n117, A2 => n34, ZN => n7);
   U7 : AND2_X1 port map( A1 => n117, A2 => n34, ZN => n119);
   U8 : INV_X1 port map( A => A(34), ZN => n8);
   U9 : BUF_X1 port map( A => n4, Z => n166);
   U10 : CLKBUF_X1 port map( A => n101, Z => n9);
   U11 : NOR2_X1 port map( A1 => B(26), A2 => n74, ZN => n10);
   U12 : BUF_X1 port map( A => n86, Z => n11);
   U13 : NOR2_X1 port map( A1 => B(41), A2 => n36, ZN => n12);
   U14 : OR2_X1 port map( A1 => net62232, A2 => net62234, ZN => net63180);
   U15 : BUF_X1 port map( A => n159, Z => n13);
   U16 : INV_X1 port map( A => B(41), ZN => n131);
   U17 : INV_X1 port map( A => B(34), ZN => n129);
   U18 : INV_X1 port map( A => B(38), ZN => net62254);
   U19 : INV_X1 port map( A => B(42), ZN => n132);
   U20 : XNOR2_X1 port map( A => n3, B => n55, ZN => SUM(15));
   U21 : CLKBUF_X1 port map( A => n31, Z => n161);
   U22 : INV_X1 port map( A => B(17), ZN => n171);
   U23 : INV_X1 port map( A => B(37), ZN => n130);
   U24 : AND3_X1 port map( A1 => n102, A2 => n103, A3 => n14, ZN => n105);
   U25 : INV_X1 port map( A => B(33), ZN => n14);
   U26 : OAI21_X1 port map( B1 => n8, B2 => n109, A => n111, ZN => n172);
   U27 : OAI21_X1 port map( B1 => n24, B2 => n19, A => n20, ZN => n22);
   U28 : XNOR2_X1 port map( A => n22, B => B(40), ZN => net62269);
   U29 : INV_X1 port map( A => A(39), ZN => n24);
   U30 : NOR2_X1 port map( A1 => n15, A2 => B(39), ZN => n19);
   U31 : OAI21_X1 port map( B1 => net62178, B2 => n19, A => n20, ZN => net62176
                           );
   U32 : OAI21_X1 port map( B1 => n16, B2 => n17, A => n18, ZN => n15);
   U33 : INV_X1 port map( A => A(38), ZN => n17);
   U34 : XNOR2_X1 port map( A => net62271, B => n17, ZN => SUM(38));
   U35 : NOR2_X1 port map( A1 => net62164, A2 => B(38), ZN => n16);
   U36 : NAND2_X1 port map( A1 => n21, A2 => B(39), ZN => n20);
   U37 : INV_X1 port map( A => A(39), ZN => net62178);
   U38 : XNOR2_X1 port map( A => n21, B => B(39), ZN => net62270);
   U39 : OAI21_X1 port map( B1 => n25, B2 => n23, A => n18, ZN => n21);
   U40 : INV_X1 port map( A => A(38), ZN => n23);
   U41 : NAND2_X1 port map( A1 => net62320, A2 => B(38), ZN => n18);
   U42 : NOR2_X1 port map( A1 => B(38), A2 => net62164, ZN => n25);
   U43 : XNOR2_X1 port map( A => net62269, B => net62356, ZN => SUM(40));
   U44 : OAI21_X1 port map( B1 => net62176, B2 => B(40), A => A(40), ZN => 
                           net62184);
   U45 : NAND2_X1 port map( A1 => net62176, A2 => B(40), ZN => net62183);
   U46 : BUF_X1 port map( A => A(40), Z => net62356);
   U47 : NOR2_X1 port map( A1 => B(21), A2 => net62067, ZN => n26);
   U48 : CLKBUF_X1 port map( A => n157, Z => n27);
   U49 : OAI21_X1 port map( B1 => n169, B2 => n91, A => n92, ZN => n157);
   U50 : NOR2_X1 port map( A1 => net62326, A2 => B(22), ZN => n28);
   U51 : NAND2_X1 port map( A1 => n65, A2 => n64, ZN => n29);
   U52 : NOR2_X1 port map( A1 => B(33), A2 => n101, ZN => n30);
   U53 : OAI21_X1 port map( B1 => n28, B2 => net62080, A => net62081, ZN => n31
                           );
   U54 : CLKBUF_X1 port map( A => A(14), Z => n32);
   U55 : OAI21_X1 port map( B1 => n105, B2 => n106, A => n107, ZN => n33);
   U56 : AND2_X1 port map( A1 => n118, A2 => n130, ZN => n34);
   U57 : NOR2_X1 port map( A1 => n104, A2 => B(34), ZN => n35);
   U58 : NAND2_X1 port map( A1 => B(28), A2 => n164, ZN => n87);
   U59 : NOR2_X1 port map( A1 => B(30), A2 => n89, ZN => n94);
   U60 : NAND2_X1 port map( A1 => n87, A2 => n88, ZN => n86);
   U61 : NAND2_X1 port map( A1 => net62184, A2 => net62183, ZN => n36);
   U62 : BUF_X1 port map( A => A(18), Z => net62366);
   U63 : XOR2_X1 port map( A => carry_47_port, B => n183, Z => SUM(47));
   U64 : INV_X1 port map( A => A(37), ZN => n37);
   U65 : NAND2_X1 port map( A1 => n102, A2 => n103, ZN => n101);
   U66 : XNOR2_X1 port map( A => A(43), B => B(43), ZN => n38);
   U67 : NAND3_X1 port map( A1 => net52614, A2 => net52615, A3 => n174, ZN => 
                           n39);
   U68 : XNOR2_X1 port map( A => n40, B => carry_45_port, ZN => SUM(45));
   U69 : XNOR2_X1 port map( A => A(45), B => B(45), ZN => n40);
   U70 : XNOR2_X1 port map( A => n116, B => n130, ZN => n137);
   U71 : CLKBUF_X1 port map( A => n126, Z => n41);
   U72 : XNOR2_X1 port map( A => A(16), B => n42, ZN => n43);
   U73 : NAND2_X1 port map( A1 => n43, A2 => net63135, ZN => net63127);
   U74 : INV_X1 port map( A => B(16), ZN => n42);
   U75 : NAND2_X1 port map( A1 => net63123, A2 => n42, ZN => n44);
   U76 : MUX2_X1 port map( A => n44, B => net52656, S => A(16), Z => net63126);
   U77 : NAND2_X1 port map( A1 => A(16), A2 => net63145, ZN => net52655);
   U78 : NAND2_X1 port map( A1 => A(16), A2 => B(16), ZN => net52654);
   U79 : NAND2_X1 port map( A1 => net63123, A2 => B(16), ZN => net52656);
   U80 : XNOR2_X1 port map( A => A(18), B => B(18), ZN => n45);
   U81 : XNOR2_X1 port map( A => n45, B => net63180, ZN => SUM(18));
   U82 : NAND2_X1 port map( A1 => B(18), A2 => net62050, ZN => net62058);
   U83 : NOR2_X1 port map( A1 => B(18), A2 => net62050, ZN => net62056);
   U84 : NOR2_X1 port map( A1 => B(18), A2 => net63180, ZN => net62331);
   U85 : OR2_X1 port map( A1 => net62232, A2 => net62234, ZN => net62050);
   U86 : OAI21_X1 port map( B1 => n133, B2 => n134, A => n154, ZN => n126);
   U87 : INV_X1 port map( A => A(42), ZN => n134);
   U88 : NAND2_X1 port map( A1 => B(42), A2 => n167, ZN => n154);
   U89 : NOR2_X1 port map( A1 => B(42), A2 => n167, ZN => n133);
   U90 : NAND2_X1 port map( A1 => n126, A2 => A(43), ZN => net52614);
   U91 : NAND2_X1 port map( A1 => n126, A2 => B(43), ZN => net52615);
   U92 : BUF_X1 port map( A => A(21), Z => n51);
   U93 : XNOR2_X1 port map( A => A(22), B => B(22), ZN => n46);
   U94 : XNOR2_X1 port map( A => n46, B => net62326, ZN => SUM(22));
   U95 : INV_X1 port map( A => A(22), ZN => net62080);
   U96 : NAND2_X1 port map( A1 => net62072, A2 => B(22), ZN => net62081);
   U97 : NOR2_X1 port map( A1 => net62072, A2 => B(22), ZN => net62079);
   U98 : OAI21_X1 port map( B1 => n50, B2 => n47, A => n48, ZN => net62326);
   U99 : INV_X1 port map( A => n51, ZN => n47);
   U100 : OAI21_X1 port map( B1 => n26, B2 => n47, A => n48, ZN => net62072);
   U101 : XNOR2_X1 port map( A => A(21), B => B(21), ZN => n49);
   U102 : NAND2_X1 port map( A1 => n29, A2 => B(21), ZN => n48);
   U103 : NOR2_X1 port map( A1 => B(21), A2 => net62067, ZN => n50);
   U104 : XNOR2_X1 port map( A => n49, B => n29, ZN => SUM(21));
   U105 : NOR2_X1 port map( A1 => n59, A2 => B(19), ZN => n52);
   U106 : XNOR2_X1 port map( A => carry_15_port, B => B(15), ZN => n55);
   U107 : NAND2_X1 port map( A1 => carry_15_port, A2 => B(15), ZN => n53);
   U108 : OAI21_X1 port map( B1 => B(15), B2 => carry_15_port, A => A(15), ZN 
                           => n54);
   U109 : NAND2_X1 port map( A1 => n53, A2 => n54, ZN => net63123);
   U110 : INV_X1 port map( A => net63145, ZN => net63135);
   U111 : NAND2_X1 port map( A1 => net63127, A2 => net63126, ZN => SUM(16));
   U112 : NAND2_X1 port map( A1 => n53, A2 => n56, ZN => net63145);
   U113 : OAI21_X1 port map( B1 => B(15), B2 => carry_15_port, A => A(15), ZN 
                           => n56);
   U114 : CLKBUF_X1 port map( A => A(19), Z => n57);
   U115 : XNOR2_X1 port map( A => n136, B => n124, ZN => SUM(41));
   U116 : XNOR2_X1 port map( A => n41, B => n38, ZN => SUM(43));
   U117 : XNOR2_X1 port map( A => n122, B => n132, ZN => n135);
   U118 : XNOR2_X1 port map( A => n135, B => n134, ZN => SUM(42));
   U119 : XNOR2_X1 port map( A => n137, B => n37, ZN => SUM(37));
   U120 : NAND3_X1 port map( A1 => net52656, A2 => net52655, A3 => net52654, ZN
                           => n58);
   U121 : INV_X1 port map( A => A(17), ZN => n127);
   U122 : OAI21_X1 port map( B1 => net62331, B2 => net62057, A => net62058, ZN 
                           => n59);
   U123 : NOR2_X1 port map( A1 => B(29), A2 => n86, ZN => n90);
   U124 : OAI21_X1 port map( B1 => n90, B2 => n91, A => n92, ZN => n89);
   U125 : NOR2_X1 port map( A1 => B(25), A2 => n71, ZN => n75);
   U126 : OAI21_X1 port map( B1 => n5, B2 => n76, A => n77, ZN => n74);
   U127 : NAND2_X1 port map( A1 => B(30), A2 => n157, ZN => n96);
   U128 : OAI21_X1 port map( B1 => n94, B2 => n95, A => n96, ZN => n93);
   U129 : OAI21_X1 port map( B1 => n94, B2 => n95, A => n96, ZN => n159);
   U130 : XNOR2_X1 port map( A => n143, B => n13, ZN => SUM(31));
   U131 : NAND2_X1 port map( A1 => B(31), A2 => n159, ZN => n100);
   U132 : NAND2_X1 port map( A1 => B(26), A2 => n158, ZN => n81);
   U133 : OAI21_X1 port map( B1 => n79, B2 => n80, A => n81, ZN => n78);
   U134 : OAI21_X1 port map( B1 => n10, B2 => n80, A => n81, ZN => n160);
   U135 : XNOR2_X1 port map( A => n147, B => n160, ZN => SUM(27));
   U136 : NAND2_X1 port map( A1 => B(27), A2 => n160, ZN => n85);
   U137 : OAI21_X1 port map( B1 => n35, B2 => n110, A => n111, ZN => n108);
   U138 : NAND2_X1 port map( A1 => n172, A2 => B(35), ZN => n115);
   U139 : XNOR2_X1 port map( A => n108, B => B(35), ZN => n139);
   U140 : NOR2_X1 port map( A1 => n172, A2 => B(35), ZN => n113);
   U141 : NOR2_X1 port map( A1 => B(34), A2 => n33, ZN => n109);
   U142 : OAI21_X1 port map( B1 => net62079, B2 => net62080, A => net62081, ZN 
                           => n66);
   U143 : NAND2_X1 port map( A1 => n31, A2 => B(23), ZN => n70);
   U144 : XNOR2_X1 port map( A => n151, B => n161, ZN => SUM(23));
   U145 : NOR2_X1 port map( A1 => n66, A2 => B(23), ZN => n68);
   U146 : OAI21_X1 port map( B1 => n113, B2 => n114, A => n115, ZN => n112);
   U147 : NAND2_X1 port map( A1 => n162, A2 => B(36), ZN => n117);
   U148 : OAI21_X1 port map( B1 => n112, B2 => B(36), A => A(36), ZN => n118);
   U149 : XNOR2_X1 port map( A => n162, B => B(36), ZN => n138);
   U150 : OAI21_X1 port map( B1 => n113, B2 => n114, A => n115, ZN => n162);
   U151 : NOR2_X1 port map( A1 => n93, A2 => B(31), ZN => n98);
   U152 : OAI21_X1 port map( B1 => n98, B2 => n99, A => n100, ZN => n97);
   U153 : OAI21_X1 port map( B1 => n99, B2 => n98, A => n100, ZN => n163);
   U154 : NOR2_X1 port map( A1 => B(27), A2 => n78, ZN => n83);
   U155 : OAI21_X1 port map( B1 => n83, B2 => n84, A => n85, ZN => n82);
   U156 : OAI21_X1 port map( B1 => n83, B2 => n84, A => n85, ZN => n164);
   U157 : OAI21_X1 port map( B1 => n52, B2 => n62, A => n63, ZN => n60);
   U158 : NAND2_X1 port map( A1 => n156, A2 => B(19), ZN => n63);
   U159 : OAI21_X1 port map( B1 => n61, B2 => n62, A => n63, ZN => n165);
   U160 : OAI21_X1 port map( B1 => n68, B2 => n69, A => n70, ZN => n67);
   U161 : NAND2_X1 port map( A1 => n4, A2 => B(24), ZN => n72);
   U162 : OAI21_X1 port map( B1 => n67, B2 => B(24), A => A(24), ZN => n73);
   U163 : XNOR2_X1 port map( A => n150, B => n166, ZN => SUM(24));
   U164 : OAI21_X1 port map( B1 => n12, B2 => n124, A => n125, ZN => n122);
   U165 : NOR2_X1 port map( A1 => B(41), A2 => n36, ZN => n123);
   U166 : OAI21_X1 port map( B1 => n124, B2 => n123, A => n125, ZN => n167);
   U167 : XNOR2_X1 port map( A => net62347, B => net62270, ZN => SUM(39));
   U168 : OAI21_X1 port map( B1 => n7, B2 => n37, A => n120, ZN => net62164);
   U169 : XNOR2_X1 port map( A => net62320, B => net62254, ZN => net62271);
   U170 : OAI21_X1 port map( B1 => n119, B2 => n37, A => n120, ZN => net62320);
   U171 : XNOR2_X1 port map( A => n139, B => n173, ZN => SUM(35));
   U172 : XNOR2_X1 port map( A => n138, B => n6, ZN => SUM(36));
   U173 : OAI21_X1 port map( B1 => n105, B2 => n106, A => n107, ZN => n104);
   U174 : XNOR2_X1 port map( A => n168, B => n129, ZN => n140);
   U175 : NAND2_X1 port map( A1 => n104, A2 => B(34), ZN => n111);
   U176 : OAI21_X1 port map( B1 => n30, B2 => n106, A => n107, ZN => n168);
   U177 : NOR2_X1 port map( A1 => B(29), A2 => n86, ZN => n169);
   U178 : OAI21_X1 port map( B1 => n75, B2 => n76, A => n77, ZN => n158);
   U179 : NOR2_X1 port map( A1 => B(19), A2 => n59, ZN => n61);
   U180 : OAI21_X1 port map( B1 => net62056, B2 => net62057, A => net62058, ZN 
                           => n156);
   U181 : XNOR2_X1 port map( A => n152, B => n165, ZN => SUM(20));
   U182 : NAND2_X1 port map( A1 => B(20), A2 => n165, ZN => n64);
   U183 : XNOR2_X1 port map( A => n153, B => n156, ZN => SUM(19));
   U184 : NAND2_X1 port map( A1 => B(33), A2 => n101, ZN => n107);
   U185 : XNOR2_X1 port map( A => n140, B => n110, ZN => SUM(34));
   U186 : NAND2_X1 port map( A1 => B(37), A2 => n116, ZN => n120);
   U187 : NAND2_X1 port map( A1 => n73, A2 => n72, ZN => n71);
   U188 : CLKBUF_X1 port map( A => n71, Z => n170);
   U189 : NAND2_X1 port map( A1 => n118, A2 => n117, ZN => n116);
   U190 : INV_X1 port map( A => n58, ZN => n128);
   U191 : XNOR2_X1 port map( A => n155, B => n58, ZN => SUM(17));
   U192 : NAND2_X1 port map( A1 => B(25), A2 => n71, ZN => n77);
   U193 : NOR2_X1 port map( A1 => B(26), A2 => n74, ZN => n79);
   U194 : XNOR2_X1 port map( A => n148, B => n158, ZN => SUM(26));
   U195 : NAND2_X1 port map( A1 => B(29), A2 => n86, ZN => n92);
   U196 : OAI21_X1 port map( B1 => n97, B2 => B(32), A => A(32), ZN => n103);
   U197 : XNOR2_X1 port map( A => n142, B => n163, ZN => SUM(32));
   U198 : NAND2_X1 port map( A1 => B(32), A2 => n163, ZN => n102);
   U199 : OAI21_X1 port map( B1 => n60, B2 => B(20), A => A(20), ZN => n65);
   U200 : NAND2_X1 port map( A1 => n65, A2 => n64, ZN => net62067);
   U201 : AOI21_X1 port map( B1 => n128, B2 => n171, A => n127, ZN => net62232)
                           ;
   U202 : XNOR2_X1 port map( A => A(28), B => B(28), ZN => n146);
   U203 : OAI21_X1 port map( B1 => B(28), B2 => n82, A => A(28), ZN => n88);
   U204 : XNOR2_X1 port map( A => A(29), B => B(29), ZN => n145);
   U205 : INV_X1 port map( A => A(29), ZN => n91);
   U206 : NOR2_X1 port map( A1 => n171, A2 => n128, ZN => net62234);
   U207 : XNOR2_X1 port map( A => A(25), B => B(25), ZN => n149);
   U208 : INV_X1 port map( A => A(25), ZN => n76);
   U209 : XNOR2_X1 port map( A => A(17), B => B(17), ZN => n155);
   U210 : XNOR2_X1 port map( A => A(31), B => B(31), ZN => n143);
   U211 : INV_X1 port map( A => A(31), ZN => n99);
   U212 : XNOR2_X1 port map( A => A(27), B => B(27), ZN => n147);
   U213 : INV_X1 port map( A => A(27), ZN => n84);
   U214 : XNOR2_X1 port map( A => A(30), B => B(30), ZN => n144);
   U215 : INV_X1 port map( A => A(30), ZN => n95);
   U216 : XNOR2_X1 port map( A => A(33), B => B(33), ZN => n141);
   U217 : INV_X1 port map( A => A(33), ZN => n106);
   U218 : INV_X1 port map( A => net62366, ZN => net62057);
   U219 : XNOR2_X1 port map( A => A(19), B => B(19), ZN => n153);
   U220 : INV_X1 port map( A => n57, ZN => n62);
   U221 : XNOR2_X1 port map( A => A(23), B => B(23), ZN => n151);
   U222 : INV_X1 port map( A => A(23), ZN => n69);
   U223 : XNOR2_X1 port map( A => A(24), B => B(24), ZN => n150);
   U224 : XNOR2_X1 port map( A => A(26), B => B(26), ZN => n148);
   U225 : INV_X1 port map( A => A(26), ZN => n80);
   U226 : INV_X1 port map( A => net62178, ZN => net62347);
   U227 : INV_X1 port map( A => A(34), ZN => n110);
   U228 : XNOR2_X1 port map( A => A(20), B => B(20), ZN => n152);
   U229 : INV_X1 port map( A => A(35), ZN => n114);
   U230 : INV_X1 port map( A => n114, ZN => n173);
   U231 : XNOR2_X1 port map( A => A(32), B => B(32), ZN => n142);
   U232 : XNOR2_X1 port map( A => n146, B => n164, ZN => SUM(28));
   U233 : XNOR2_X1 port map( A => n145, B => n11, ZN => SUM(29));
   U234 : INV_X1 port map( A => A(41), ZN => n124);
   U235 : NAND2_X1 port map( A1 => net62184, A2 => net62183, ZN => n121);
   U236 : XNOR2_X1 port map( A => n149, B => n170, ZN => SUM(25));
   U237 : XNOR2_X1 port map( A => n144, B => n27, ZN => SUM(30));
   U238 : XNOR2_X1 port map( A => n141, B => n9, ZN => SUM(33));
   U239 : XNOR2_X1 port map( A => n121, B => n131, ZN => n136);
   U240 : NAND2_X1 port map( A1 => n36, A2 => B(41), ZN => n125);
   U241 : NAND2_X1 port map( A1 => A(43), A2 => B(43), ZN => n174);
   U242 : NAND3_X1 port map( A1 => net52614, A2 => net52615, A3 => n174, ZN => 
                           carry_44_port);
   U243 : XOR2_X1 port map( A => n32, B => B(14), Z => n175);
   U244 : XOR2_X1 port map( A => carry_14_port, B => n175, Z => SUM(14));
   U245 : NAND2_X1 port map( A1 => carry_14_port, A2 => n32, ZN => n176);
   U246 : NAND2_X1 port map( A1 => carry_14_port, A2 => B(14), ZN => n177);
   U247 : NAND2_X1 port map( A1 => A(14), A2 => B(14), ZN => n178);
   U248 : NAND3_X1 port map( A1 => n176, A2 => n177, A3 => n178, ZN => 
                           carry_15_port);
   U249 : NAND2_X1 port map( A1 => B(44), A2 => carry_44_port, ZN => net42193);
   U250 : NAND2_X1 port map( A1 => A(44), A2 => n39, ZN => net42192);
   U251 : XOR2_X1 port map( A => net42190, B => carry_44_port, Z => SUM(44));
   U252 : XOR2_X1 port map( A => A(44), B => B(44), Z => net42190);
   U253 : NAND2_X1 port map( A1 => A(44), A2 => B(44), ZN => n179);
   U254 : NAND3_X1 port map( A1 => n179, A2 => net42192, A3 => net42193, ZN => 
                           carry_45_port);
   U255 : NAND2_X1 port map( A1 => A(45), A2 => B(45), ZN => n180);
   U256 : NAND2_X1 port map( A1 => A(45), A2 => carry_45_port, ZN => n181);
   U257 : NAND2_X1 port map( A1 => B(45), A2 => carry_45_port, ZN => n182);
   U258 : NAND3_X1 port map( A1 => n180, A2 => n181, A3 => n182, ZN => 
                           carry_46_port);
   U259 : XOR2_X1 port map( A => A(47), B => B(47), Z => n183);
   U260 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n1);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT46_DW01_add_0 is

   port( A, B : in std_logic_vector (45 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (45 downto 0);  CO : out std_logic);

end RCA_NBIT46_DW01_add_0;

architecture SYN_rpl of RCA_NBIT46_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_45_port, carry_44_port, carry_43_port, carry_42_port, 
      carry_12_port, carry_11_port, carry_10_port, carry_9_port, carry_8_port, 
      carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port, 
      carry_2_port, n1, net51366, net51324, net51309, net51303, net51302, 
      net51301, net51297, net51296, net51295, net51278, net51247, net51233, 
      net51226, net51177, net51169, net51167, net51117, net51116, net51115, 
      net51105, net51104, net51103, net51102, net51080, net51079, net51075, 
      net51056, net51035, net51021, net51380, net52606, net52803, net52807, 
      net55239, net55370, net51479, net51312, net51288, net51108, net52687, 
      net51299, net51082, net51081, net51340, net51353, net62443, net51321, 
      net51076, net51071, net51069, net51065, net51064, net51063, net51062, 
      net51074, net51325, net51223, net51030, net51028, net51027, net55374, 
      net51322, net51053, net51052, net51045, net52617, net51059, net51058, 
      net51057, net51048, net51046, net51482, net51298, net51230, net51051, 
      net51300, net51039, net55358, net52805, net52589, net51315, net51041, 
      net51040, net51036, net51034, net51316, net51166, net87441, net51180, 
      net51179, net51178, net79782, net51364, n3, n4, n5, n6, n7, n8, n9, n10, 
      n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25
      , n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, 
      n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54
      , n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, 
      n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83
      , n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, 
      n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, 
      n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
      n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, 
      n134, n135, n136 : std_logic;

begin
   
   U1_42 : FA_X1 port map( A => carry_42_port, B => B(42), CI => A(42), CO => 
                           carry_43_port, S => SUM(42));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : OAI21_X1 port map( B1 => n28, B2 => net51028, A => net51030, ZN => n3);
   U3 : OAI21_X1 port map( B1 => n28, B2 => net51028, A => net51030, ZN => 
                           net51325);
   U4 : INV_X1 port map( A => A(19), ZN => n4);
   U5 : CLKBUF_X1 port map( A => A(37), Z => n5);
   U6 : NAND2_X1 port map( A1 => n66, A2 => n65, ZN => n6);
   U7 : BUF_X1 port map( A => A(38), Z => net52606);
   U8 : AND2_X1 port map( A1 => n7, A2 => n62, ZN => net51103);
   U9 : AND2_X1 port map( A1 => n61, A2 => n8, ZN => n7);
   U10 : INV_X1 port map( A => B(26), ZN => n8);
   U11 : INV_X1 port map( A => B(15), ZN => net51226);
   U12 : INV_X1 port map( A => B(39), ZN => n13);
   U13 : NAND2_X1 port map( A1 => net79782, A2 => B(39), ZN => net51180);
   U14 : INV_X1 port map( A => B(18), ZN => net51230);
   U15 : XNOR2_X1 port map( A => B(12), B => carry_12_port, ZN => n118);
   U16 : INV_X1 port map( A => B(14), ZN => net51223);
   U17 : INV_X1 port map( A => B(13), ZN => n27);
   U18 : INV_X1 port map( A => B(19), ZN => net51233);
   U19 : INV_X1 port map( A => B(31), ZN => n95);
   U20 : INV_X1 port map( A => B(30), ZN => n94);
   U21 : INV_X1 port map( A => B(35), ZN => n97);
   U22 : INV_X1 port map( A => B(23), ZN => n92);
   U23 : CLKBUF_X1 port map( A => A(16), Z => n9);
   U24 : BUF_X1 port map( A => A(33), Z => n45);
   U25 : AND2_X1 port map( A1 => A(41), A2 => B(41), ZN => n10);
   U26 : INV_X1 port map( A => B(22), ZN => n30);
   U27 : INV_X1 port map( A => B(34), ZN => n96);
   U28 : INV_X1 port map( A => B(26), ZN => n93);
   U29 : INV_X1 port map( A => B(27), ZN => net51247);
   U30 : XNOR2_X1 port map( A => A(43), B => B(43), ZN => n18);
   U31 : OAI21_X1 port map( B1 => n82, B2 => n81, A => n83, ZN => n49);
   U32 : XNOR2_X1 port map( A => net51364, B => n13, ZN => n14);
   U33 : XNOR2_X1 port map( A => n14, B => net51179, ZN => SUM(39));
   U34 : NAND2_X1 port map( A1 => n12, A2 => n11, ZN => net51364);
   U35 : NOR2_X1 port map( A1 => B(39), A2 => net79782, ZN => net51178);
   U36 : NOR2_X1 port map( A1 => B(39), A2 => net79782, ZN => net87441);
   U37 : OAI21_X1 port map( B1 => net51316, B2 => B(38), A => A(38), ZN => n12)
                           ;
   U38 : NAND2_X1 port map( A1 => n12, A2 => n11, ZN => net79782);
   U39 : NAND2_X1 port map( A1 => net51316, A2 => B(38), ZN => n11);
   U40 : XNOR2_X1 port map( A => net51166, B => B(38), ZN => net51278);
   U41 : INV_X1 port map( A => A(39), ZN => net51179);
   U42 : OAI21_X1 port map( B1 => net87441, B2 => net51179, A => net51180, ZN 
                           => net51309);
   U43 : OAI21_X1 port map( B1 => net51179, B2 => net51178, A => net51180, ZN 
                           => net51177);
   U44 : OAI21_X1 port map( B1 => net51167, B2 => n15, A => net51169, ZN => 
                           net51316);
   U45 : INV_X1 port map( A => A(37), ZN => n15);
   U46 : OAI21_X1 port map( B1 => net51167, B2 => n15, A => net51169, ZN => 
                           net51166);
   U47 : NOR2_X1 port map( A1 => B(32), A2 => n71, ZN => n16);
   U48 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => n17);
   U49 : OAI21_X1 port map( B1 => net51064, B2 => net51063, A => net51065, ZN 
                           => net51062);
   U50 : XNOR2_X1 port map( A => carry_43_port, B => n18, ZN => SUM(43));
   U51 : XNOR2_X1 port map( A => carry_44_port, B => n19, ZN => SUM(44));
   U52 : XNOR2_X1 port map( A => A(44), B => B(44), ZN => n19);
   U53 : CLKBUF_X1 port map( A => n17, Z => n20);
   U54 : BUF_X1 port map( A => A(12), Z => n47);
   U55 : AND2_X1 port map( A1 => n21, A2 => n80, ZN => n81);
   U56 : AND2_X1 port map( A1 => n79, A2 => n96, ZN => n21);
   U57 : NAND2_X1 port map( A1 => n128, A2 => B(34), ZN => n83);
   U58 : OAI21_X1 port map( B1 => net51041, B2 => net52589, A => n22, ZN => 
                           net51315);
   U59 : XNOR2_X1 port map( A => net51315, B => B(16), ZN => net51300);
   U60 : NOR2_X1 port map( A1 => B(15), A2 => net52805, ZN => net52589);
   U61 : INV_X1 port map( A => A(15), ZN => net51041);
   U62 : XNOR2_X1 port map( A => net51041, B => net51301, ZN => SUM(15));
   U63 : NAND2_X1 port map( A1 => net55358, A2 => B(15), ZN => n22);
   U64 : OAI21_X1 port map( B1 => net51040, B2 => n24, A => n22, ZN => net51039
                           );
   U65 : OAI21_X1 port map( B1 => n25, B2 => n23, A => net51036, ZN => net55358
                           );
   U66 : INV_X1 port map( A => A(14), ZN => n23);
   U67 : OAI21_X1 port map( B1 => n23, B2 => net51034, A => net51036, ZN => 
                           net52805);
   U68 : NOR2_X1 port map( A1 => net52805, A2 => B(15), ZN => net51040);
   U69 : NOR2_X1 port map( A1 => net51027, A2 => B(14), ZN => net51034);
   U70 : INV_X1 port map( A => A(15), ZN => n24);
   U71 : OAI21_X1 port map( B1 => net51035, B2 => n25, A => net51036, ZN => 
                           net51366);
   U72 : INV_X1 port map( A => A(14), ZN => net51035);
   U73 : NOR2_X1 port map( A1 => net51027, A2 => B(14), ZN => n25);
   U74 : NAND2_X1 port map( A1 => net51325, A2 => B(14), ZN => net51036);
   U75 : XNOR2_X1 port map( A => net51300, B => n9, ZN => SUM(16));
   U76 : NAND2_X1 port map( A1 => net51039, A2 => B(16), ZN => net51048);
   U77 : NOR2_X1 port map( A1 => net51039, A2 => B(16), ZN => net51046);
   U78 : INV_X1 port map( A => A(16), ZN => net55374);
   U79 : XNOR2_X1 port map( A => net51482, B => net51230, ZN => net51298);
   U80 : XNOR2_X1 port map( A => net51298, B => net51058, ZN => SUM(18));
   U81 : NAND2_X1 port map( A1 => net51053, A2 => net51052, ZN => net51482);
   U82 : NOR2_X1 port map( A1 => B(18), A2 => net51482, ZN => net52617);
   U83 : NOR2_X1 port map( A1 => net51051, A2 => B(18), ZN => net51057);
   U84 : NAND2_X1 port map( A1 => net51051, A2 => B(18), ZN => net51059);
   U85 : NAND2_X1 port map( A1 => net51053, A2 => net51052, ZN => net51051);
   U86 : OAI21_X1 port map( B1 => net51046, B2 => net55374, A => net51048, ZN 
                           => net51045);
   U87 : OAI21_X1 port map( B1 => net51046, B2 => net55374, A => net51048, ZN 
                           => net51322);
   U88 : INV_X1 port map( A => A(18), ZN => net51058);
   U89 : OAI21_X1 port map( B1 => net51058, B2 => net52617, A => net51059, ZN 
                           => net51056);
   U90 : OAI21_X1 port map( B1 => net51057, B2 => net51058, A => net51059, ZN 
                           => net51340);
   U91 : OAI21_X1 port map( B1 => net51045, B2 => B(17), A => A(17), ZN => 
                           net51053);
   U92 : NAND2_X1 port map( A1 => net51045, A2 => B(17), ZN => net51052);
   U93 : XNOR2_X1 port map( A => net51322, B => B(17), ZN => net51299);
   U94 : CLKBUF_X1 port map( A => A(17), Z => net52687);
   U95 : OAI21_X1 port map( B1 => n26, B2 => n29, A => net51030, ZN => net51027
                           );
   U96 : NOR2_X1 port map( A1 => net51021, A2 => B(13), ZN => n29);
   U97 : INV_X1 port map( A => A(13), ZN => n26);
   U98 : CLKBUF_X1 port map( A => n26, Z => net55370);
   U99 : XNOR2_X1 port map( A => n3, B => net51223, ZN => net51302);
   U100 : NOR2_X1 port map( A1 => n17, A2 => B(13), ZN => net51028);
   U101 : NAND2_X1 port map( A1 => B(13), A2 => net51021, ZN => net51030);
   U102 : XNOR2_X1 port map( A => n20, B => n27, ZN => net51303);
   U103 : INV_X1 port map( A => A(13), ZN => n28);
   U104 : XNOR2_X1 port map( A => net51074, B => n30, ZN => n31);
   U105 : XNOR2_X1 port map( A => n31, B => net51081, ZN => SUM(22));
   U106 : NAND2_X1 port map( A1 => net51075, A2 => net51076, ZN => net51074);
   U107 : NAND2_X1 port map( A1 => net51074, A2 => B(22), ZN => net51082);
   U108 : AND2_X1 port map( A1 => net51075, A2 => n30, ZN => net51380);
   U109 : NOR2_X1 port map( A1 => B(20), A2 => net51062, ZN => net51069);
   U110 : NOR2_X1 port map( A1 => net51353, A2 => B(20), ZN => net62443);
   U111 : NAND2_X1 port map( A1 => net51353, A2 => B(20), ZN => net51071);
   U112 : INV_X1 port map( A => A(19), ZN => net51064);
   U113 : XNOR2_X1 port map( A => net51064, B => net51297, ZN => SUM(19));
   U114 : OAI21_X1 port map( B1 => net51063, B2 => n4, A => net51065, ZN => 
                           net51353);
   U115 : NOR2_X1 port map( A1 => net51340, A2 => B(19), ZN => net51063);
   U116 : NAND2_X1 port map( A1 => net51340, A2 => B(19), ZN => net51065);
   U117 : OAI21_X1 port map( B1 => B(21), B2 => n32, A => A(21), ZN => net51076
                           );
   U118 : OAI21_X1 port map( B1 => net62443, B2 => n33, A => net51071, ZN => 
                           n32);
   U119 : NAND2_X1 port map( A1 => n32, A2 => B(21), ZN => net51075);
   U120 : INV_X1 port map( A => A(20), ZN => n33);
   U121 : OAI21_X1 port map( B1 => net51069, B2 => n33, A => net51071, ZN => 
                           net51321);
   U122 : XNOR2_X1 port map( A => net51321, B => B(21), ZN => net51295);
   U123 : CLKBUF_X1 port map( A => A(21), Z => net52803);
   U124 : CLKBUF_X1 port map( A => A(20), Z => net52807);
   U125 : XNOR2_X1 port map( A => net51062, B => B(20), ZN => net51296);
   U126 : INV_X1 port map( A => A(22), ZN => net51081);
   U127 : OAI21_X1 port map( B1 => net51081, B2 => net51080, A => net51082, ZN 
                           => net51324);
   U128 : OAI21_X1 port map( B1 => net51080, B2 => net51081, A => net51082, ZN 
                           => net51079);
   U129 : XNOR2_X1 port map( A => net51299, B => net52687, ZN => SUM(17));
   U130 : OAI21_X1 port map( B1 => n38, B2 => n35, A => n36, ZN => n37);
   U131 : XNOR2_X1 port map( A => n37, B => B(28), ZN => net51288);
   U132 : INV_X1 port map( A => A(27), ZN => n35);
   U133 : OAI21_X1 port map( B1 => n34, B2 => n35, A => n36, ZN => net51108);
   U134 : NOR2_X1 port map( A1 => n39, A2 => B(27), ZN => n38);
   U135 : OAI21_X1 port map( B1 => n38, B2 => n35, A => n36, ZN => net51312);
   U136 : NAND2_X1 port map( A1 => net51102, A2 => B(27), ZN => n36);
   U137 : OAI21_X1 port map( B1 => net51104, B2 => net51103, A => net51105, ZN 
                           => n39);
   U138 : NOR2_X1 port map( A1 => B(27), A2 => n39, ZN => n34);
   U139 : OAI21_X1 port map( B1 => net51103, B2 => net51104, A => net51105, ZN 
                           => net51102);
   U140 : INV_X1 port map( A => A(26), ZN => net51104);
   U141 : XNOR2_X1 port map( A => net51288, B => net51479, ZN => SUM(28));
   U142 : NAND2_X1 port map( A1 => B(28), A2 => net51312, ZN => net51117);
   U143 : NOR2_X1 port map( A1 => net51108, A2 => B(28), ZN => net51115);
   U144 : NOR2_X1 port map( A1 => B(28), A2 => net51108, ZN => net55239);
   U145 : CLKBUF_X1 port map( A => A(28), Z => net51479);
   U146 : INV_X1 port map( A => A(28), ZN => net51116);
   U147 : CLKBUF_X1 port map( A => A(32), Z => n40);
   U148 : OAI21_X1 port map( B1 => n48, B2 => n84, A => n85, ZN => n41);
   U149 : XNOR2_X1 port map( A => net51303, B => net55370, ZN => SUM(13));
   U150 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => net51021);
   U151 : CLKBUF_X1 port map( A => A(29), Z => n42);
   U152 : CLKBUF_X1 port map( A => A(36), Z => n43);
   U153 : CLKBUF_X1 port map( A => n100, Z => n44);
   U154 : XNOR2_X1 port map( A => n117, B => n55, ZN => SUM(23));
   U155 : NAND2_X1 port map( A1 => n61, A2 => n62, ZN => n46);
   U156 : INV_X1 port map( A => A(35), ZN => n48);
   U157 : NOR2_X1 port map( A1 => n91, A2 => n90, ZN => carry_42_port);
   U158 : XNOR2_X1 port map( A => n106, B => n48, ZN => SUM(35));
   U159 : INV_X1 port map( A => A(31), ZN => n50);
   U160 : XNOR2_X1 port map( A => n114, B => net51104, ZN => SUM(26));
   U161 : INV_X1 port map( A => A(40), ZN => n99);
   U162 : NAND2_X1 port map( A1 => B(40), A2 => net51309, ZN => n101);
   U163 : OAI21_X1 port map( B1 => n59, B2 => n58, A => n60, ZN => n51);
   U164 : AND2_X1 port map( A1 => net51380, A2 => net51076, ZN => net51080);
   U165 : XNOR2_X1 port map( A => net51302, B => net51035, ZN => SUM(14));
   U166 : OAI21_X1 port map( B1 => n88, B2 => n87, A => n89, ZN => n86);
   U167 : NOR2_X1 port map( A1 => n125, A2 => B(36), ZN => n87);
   U168 : OAI21_X1 port map( B1 => n87, B2 => n88, A => n89, ZN => n119);
   U169 : NOR2_X1 port map( A1 => n67, A2 => B(31), ZN => n72);
   U170 : OAI21_X1 port map( B1 => n72, B2 => n73, A => n74, ZN => n71);
   U171 : OAI21_X1 port map( B1 => n50, B2 => n123, A => n74, ZN => n120);
   U172 : NAND2_X1 port map( A1 => n129, A2 => B(24), ZN => n60);
   U173 : XNOR2_X1 port map( A => n126, B => B(24), ZN => n116);
   U174 : NOR2_X1 port map( A1 => n129, A2 => B(24), ZN => n58);
   U175 : NOR2_X1 port map( A1 => n119, A2 => B(37), ZN => net51167);
   U176 : NOR2_X1 port map( A1 => n71, A2 => B(32), ZN => n76);
   U177 : OAI21_X1 port map( B1 => n16, B2 => n77, A => n78, ZN => n75);
   U178 : OAI21_X1 port map( B1 => n76, B2 => n77, A => n78, ZN => n121);
   U179 : OAI21_X1 port map( B1 => net51116, B2 => net55239, A => net51117, ZN 
                           => n63);
   U180 : OAI21_X1 port map( B1 => n58, B2 => n59, A => n60, ZN => n57);
   U181 : NAND2_X1 port map( A1 => n57, A2 => B(25), ZN => n61);
   U182 : OAI21_X1 port map( B1 => n57, B2 => B(25), A => A(25), ZN => n62);
   U183 : XNOR2_X1 port map( A => n51, B => B(25), ZN => n115);
   U184 : XNOR2_X1 port map( A => n122, B => n97, ZN => n106);
   U185 : NAND2_X1 port map( A1 => n49, A2 => B(35), ZN => n85);
   U186 : NOR2_X1 port map( A1 => n49, A2 => B(35), ZN => n84);
   U187 : OAI21_X1 port map( B1 => n82, B2 => n81, A => n83, ZN => n122);
   U188 : XNOR2_X1 port map( A => net51324, B => n92, ZN => n117);
   U189 : NAND2_X1 port map( A1 => net51079, A2 => B(23), ZN => n56);
   U190 : NOR2_X1 port map( A1 => net51079, A2 => B(23), ZN => n54);
   U191 : NAND2_X1 port map( A1 => n125, A2 => B(36), ZN => n89);
   U192 : XNOR2_X1 port map( A => n41, B => B(36), ZN => n105);
   U193 : NOR2_X1 port map( A1 => n124, A2 => B(31), ZN => n123);
   U194 : OAI21_X1 port map( B1 => n69, B2 => n68, A => n70, ZN => n67);
   U195 : XNOR2_X1 port map( A => n67, B => n95, ZN => n110);
   U196 : NAND2_X1 port map( A1 => n124, A2 => B(31), ZN => n74);
   U197 : NOR2_X1 port map( A1 => n64, A2 => B(30), ZN => n68);
   U198 : OAI21_X1 port map( B1 => n69, B2 => n68, A => n70, ZN => n124);
   U199 : XNOR2_X1 port map( A => net51102, B => net51247, ZN => n113);
   U200 : NAND2_X1 port map( A1 => n119, A2 => B(37), ZN => net51169);
   U201 : XNOR2_X1 port map( A => n86, B => B(37), ZN => n104);
   U202 : OAI21_X1 port map( B1 => n84, B2 => n48, A => n85, ZN => n125);
   U203 : XNOR2_X1 port map( A => net51177, B => B(40), ZN => n103);
   U204 : NAND2_X1 port map( A1 => n120, A2 => B(32), ZN => n78);
   U205 : XNOR2_X1 port map( A => n115, B => A(25), ZN => SUM(25));
   U206 : XNOR2_X1 port map( A => n75, B => B(33), ZN => n108);
   U207 : NAND2_X1 port map( A1 => n121, A2 => B(33), ZN => n79);
   U208 : XNOR2_X1 port map( A => B(29), B => n63, ZN => n112);
   U209 : NAND2_X1 port map( A1 => n127, A2 => B(29), ZN => n65);
   U210 : XNOR2_X1 port map( A => n120, B => B(32), ZN => n109);
   U211 : XNOR2_X1 port map( A => n103, B => A(40), ZN => SUM(40));
   U212 : XNOR2_X1 port map( A => net51056, B => net51233, ZN => net51297);
   U213 : INV_X1 port map( A => A(24), ZN => n59);
   U214 : OAI21_X1 port map( B1 => n55, B2 => n54, A => n56, ZN => n126);
   U215 : XNOR2_X1 port map( A => n105, B => n43, ZN => SUM(36));
   U216 : XNOR2_X1 port map( A => net51366, B => net51226, ZN => net51301);
   U217 : XNOR2_X1 port map( A => net51295, B => net52803, ZN => SUM(21));
   U218 : XNOR2_X1 port map( A => net51278, B => net52606, ZN => SUM(38));
   U219 : XNOR2_X1 port map( A => n108, B => n45, ZN => SUM(33));
   U220 : XNOR2_X1 port map( A => n42, B => n112, ZN => SUM(29));
   U221 : XNOR2_X1 port map( A => n104, B => n5, ZN => SUM(37));
   U222 : INV_X1 port map( A => A(23), ZN => n55);
   U223 : XNOR2_X1 port map( A => net51296, B => net52807, ZN => SUM(20));
   U224 : XNOR2_X1 port map( A => n109, B => n40, ZN => SUM(32));
   U225 : XNOR2_X1 port map( A => n128, B => n96, ZN => n107);
   U226 : XNOR2_X1 port map( A => n6, B => n94, ZN => n111);
   U227 : XNOR2_X1 port map( A => n69, B => n111, ZN => SUM(30));
   U228 : XNOR2_X1 port map( A => n116, B => A(24), ZN => SUM(24));
   U229 : XNOR2_X1 port map( A => A(41), B => B(41), ZN => n102);
   U230 : NOR2_X1 port map( A1 => A(41), A2 => B(41), ZN => n90);
   U231 : OAI21_X1 port map( B1 => n98, B2 => n99, A => n101, ZN => n100);
   U232 : XNOR2_X1 port map( A => n102, B => n44, ZN => SUM(41));
   U233 : NOR2_X1 port map( A1 => n100, A2 => n10, ZN => n91);
   U234 : NAND2_X1 port map( A1 => B(12), A2 => A(12), ZN => n52);
   U235 : OAI21_X1 port map( B1 => n47, B2 => B(12), A => carry_12_port, ZN => 
                           n53);
   U236 : XNOR2_X1 port map( A => n47, B => n118, ZN => SUM(12));
   U237 : INV_X1 port map( A => A(32), ZN => n77);
   U238 : INV_X1 port map( A => A(36), ZN => n88);
   U239 : INV_X1 port map( A => A(31), ZN => n73);
   U240 : INV_X1 port map( A => A(34), ZN => n82);
   U241 : XNOR2_X1 port map( A => n46, B => n93, ZN => n114);
   U242 : NAND2_X1 port map( A1 => n46, A2 => B(26), ZN => net51105);
   U243 : XNOR2_X1 port map( A => n107, B => n82, ZN => SUM(34));
   U244 : NAND2_X1 port map( A1 => n6, A2 => B(30), ZN => n70);
   U245 : INV_X1 port map( A => A(30), ZN => n69);
   U246 : XNOR2_X1 port map( A => n110, B => n73, ZN => SUM(31));
   U247 : OAI21_X1 port map( B1 => net51115, B2 => net51116, A => net51117, ZN 
                           => n127);
   U248 : XNOR2_X1 port map( A => n113, B => n35, ZN => SUM(27));
   U249 : OAI21_X1 port map( B1 => n121, B2 => B(33), A => A(33), ZN => n80);
   U250 : NAND2_X1 port map( A1 => n80, A2 => n79, ZN => n128);
   U251 : NAND2_X1 port map( A1 => n66, A2 => n65, ZN => n64);
   U252 : NOR2_X1 port map( A1 => B(40), A2 => net51309, ZN => n98);
   U253 : OAI21_X1 port map( B1 => n54, B2 => n55, A => n56, ZN => n129);
   U254 : OAI21_X1 port map( B1 => n127, B2 => B(29), A => A(29), ZN => n66);
   U255 : NAND2_X1 port map( A1 => carry_43_port, A2 => A(43), ZN => n130);
   U256 : NAND2_X1 port map( A1 => carry_43_port, A2 => B(43), ZN => n131);
   U257 : NAND2_X1 port map( A1 => A(43), A2 => B(43), ZN => n132);
   U258 : NAND3_X1 port map( A1 => n130, A2 => n131, A3 => n132, ZN => 
                           carry_44_port);
   U259 : NAND2_X1 port map( A1 => carry_44_port, A2 => A(44), ZN => n133);
   U260 : NAND2_X1 port map( A1 => carry_44_port, A2 => B(44), ZN => n134);
   U261 : NAND2_X1 port map( A1 => A(44), A2 => B(44), ZN => n135);
   U262 : NAND3_X1 port map( A1 => n133, A2 => n134, A3 => n135, ZN => 
                           carry_45_port);
   U263 : XOR2_X1 port map( A => A(45), B => B(45), Z => n136);
   U264 : XOR2_X1 port map( A => carry_45_port, B => n136, Z => SUM(45));
   U265 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n1);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT44_DW01_add_0 is

   port( A, B : in std_logic_vector (43 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (43 downto 0);  CO : out std_logic);

end RCA_NBIT44_DW01_add_0;

architecture SYN_rpl of RCA_NBIT44_DW01_add_0 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_43_port, carry_42_port, net45992, net45991, net51441, net52575,
      net52564, net52506, net52420, net52419, net52418, net52413, net52405, 
      net52356, net52355, net52342, net52287, net52285, net52284, net52280, 
      net52279, net52706, net52524, net52348, net52685, n1, carry_9_port, 
      carry_8_port, carry_7_port, carry_6_port, carry_5_port, carry_4_port, 
      carry_3_port, carry_2_port, carry_14_port, carry_13_port, carry_12_port, 
      carry_11_port, carry_10_port, net52605, net52286, net52414, net52412, 
      net79780, net52558, net52513, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, 
      n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27
      , n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, 
      n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56
      , n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, 
      n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85
      , n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, 
      n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, 
      n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, 
      n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, 
      n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, 
      n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, 
      n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n174, n175, n176, n177, n178, n179, n180 : std_logic;

begin
   
   U1_42 : FA_X1 port map( A => A(42), B => B(42), CI => carry_42_port, CO => 
                           carry_43_port, S => SUM(42));
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_13 : FA_X1 port map( A => B(13), B => A(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1 : NAND2_X1 port map( A1 => n62, A2 => n61, ZN => n3);
   U3 : OAI21_X1 port map( B1 => n80, B2 => n79, A => n81, ZN => n4);
   U4 : INV_X1 port map( A => B(17), ZN => n124);
   U5 : INV_X1 port map( A => B(36), ZN => n133);
   U6 : INV_X1 port map( A => B(37), ZN => net52506);
   U7 : XNOR2_X1 port map( A => B(40), B => A(40), ZN => n134);
   U8 : INV_X1 port map( A => B(16), ZN => n123);
   U9 : INV_X1 port map( A => B(15), ZN => n25);
   U10 : INV_X1 port map( A => B(20), ZN => n125);
   U11 : INV_X1 port map( A => B(21), ZN => n126);
   U12 : INV_X1 port map( A => B(25), ZN => n128);
   U13 : INV_X1 port map( A => B(29), ZN => n130);
   U14 : INV_X1 port map( A => B(33), ZN => n132);
   U15 : INV_X1 port map( A => B(28), ZN => n129);
   U16 : INV_X1 port map( A => B(32), ZN => n131);
   U17 : INV_X1 port map( A => B(24), ZN => n127);
   U18 : XOR2_X1 port map( A => A(10), B => B(10), Z => n5);
   U19 : XOR2_X1 port map( A => carry_10_port, B => n5, Z => SUM(10));
   U20 : NAND2_X1 port map( A1 => carry_10_port, A2 => A(10), ZN => n6);
   U21 : NAND2_X1 port map( A1 => carry_10_port, A2 => B(10), ZN => n7);
   U22 : NAND2_X1 port map( A1 => A(10), A2 => B(10), ZN => n8);
   U23 : NAND3_X1 port map( A1 => n6, A2 => n7, A3 => n8, ZN => carry_11_port);
   U24 : OAI211_X1 port map( C1 => n89, C2 => n90, A => n91, B => n9, ZN => n10
                           );
   U25 : INV_X1 port map( A => B(30), ZN => n9);
   U26 : INV_X1 port map( A => n10, ZN => n93);
   U27 : XNOR2_X1 port map( A => n11, B => B(38), ZN => net52513);
   U28 : XNOR2_X1 port map( A => net52513, B => net79780, ZN => SUM(38));
   U29 : OAI21_X1 port map( B1 => n12, B2 => net52412, A => net52414, ZN => n11
                           );
   U30 : NAND2_X1 port map( A1 => n11, A2 => B(38), ZN => net52420);
   U31 : INV_X1 port map( A => A(37), ZN => n12);
   U32 : NOR2_X1 port map( A1 => net52558, A2 => B(38), ZN => net52564);
   U33 : NOR2_X1 port map( A1 => B(38), A2 => net52558, ZN => net52418);
   U34 : OAI21_X1 port map( B1 => net52413, B2 => net52412, A => net52414, ZN 
                           => net52558);
   U35 : INV_X1 port map( A => A(37), ZN => net52413);
   U36 : CLKBUF_X1 port map( A => A(38), Z => net79780);
   U37 : INV_X1 port map( A => A(38), ZN => net52419);
   U38 : NOR2_X1 port map( A1 => net52405, A2 => B(37), ZN => net52412);
   U39 : NAND2_X1 port map( A1 => net52405, A2 => B(37), ZN => net52414);
   U40 : CLKBUF_X1 port map( A => carry_11_port, Z => n13);
   U41 : XNOR2_X1 port map( A => carry_43_port, B => n45, ZN => SUM(43));
   U42 : CLKBUF_X1 port map( A => A(26), Z => n35);
   U43 : INV_X1 port map( A => A(32), ZN => n14);
   U44 : CLKBUF_X1 port map( A => A(11), Z => n15);
   U45 : NAND2_X1 port map( A1 => B(33), A2 => n173, ZN => n16);
   U46 : NOR2_X1 port map( A1 => n60, A2 => B(20), ZN => n17);
   U47 : NOR2_X1 port map( A1 => n178, A2 => B(16), ZN => n18);
   U48 : OAI21_X1 port map( B1 => n100, B2 => n101, A => n102, ZN => n19);
   U49 : CLKBUF_X1 port map( A => A(31), Z => n21);
   U50 : CLKBUF_X1 port map( A => A(35), Z => n20);
   U51 : NOR2_X1 port map( A1 => n41, A2 => B(28), ZN => n22);
   U52 : AND2_X1 port map( A1 => n77, A2 => n23, ZN => n79);
   U53 : AND2_X1 port map( A1 => n76, A2 => n127, ZN => n23);
   U54 : XNOR2_X1 port map( A => n27, B => n25, ZN => n26);
   U55 : XNOR2_X1 port map( A => n26, B => net52286, ZN => SUM(15));
   U56 : NAND2_X1 port map( A1 => net52280, A2 => net52279, ZN => n27);
   U57 : NOR2_X1 port map( A1 => B(15), A2 => n27, ZN => net52605);
   U58 : NAND2_X1 port map( A1 => n24, A2 => B(15), ZN => net52287);
   U59 : NOR2_X1 port map( A1 => n24, A2 => B(15), ZN => net52285);
   U60 : NAND2_X1 port map( A1 => net52280, A2 => net52279, ZN => n24);
   U61 : INV_X1 port map( A => A(15), ZN => net52286);
   U62 : OAI21_X1 port map( B1 => net52605, B2 => net52286, A => net52287, ZN 
                           => net52284);
   U63 : INV_X1 port map( A => A(15), ZN => net52706);
   U64 : XOR2_X1 port map( A => n15, B => B(11), Z => n28);
   U65 : XOR2_X1 port map( A => n13, B => n28, Z => SUM(11));
   U66 : NAND2_X1 port map( A1 => A(11), A2 => carry_11_port, ZN => n29);
   U67 : NAND2_X1 port map( A1 => carry_11_port, A2 => B(11), ZN => n30);
   U68 : NAND2_X1 port map( A1 => A(11), A2 => B(11), ZN => n31);
   U69 : NAND3_X1 port map( A1 => n29, A2 => n31, A3 => n30, ZN => 
                           carry_12_port);
   U70 : XNOR2_X1 port map( A => carry_14_port, B => B(14), ZN => n32);
   U71 : XNOR2_X1 port map( A => n32, B => net52685, ZN => SUM(14));
   U72 : OAI21_X1 port map( B1 => A(14), B2 => B(14), A => carry_14_port, ZN =>
                           net52280);
   U73 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n1);
   U74 : NAND2_X1 port map( A1 => A(14), A2 => B(14), ZN => net52279);
   U75 : CLKBUF_X1 port map( A => A(14), Z => net52685);
   U76 : NOR2_X1 port map( A1 => n48, A2 => B(17), ZN => n33);
   U77 : CLKBUF_X1 port map( A => A(22), Z => n34);
   U78 : AND2_X2 port map( A1 => n97, A2 => n42, ZN => n100);
   U79 : NAND2_X1 port map( A1 => n157, A2 => n156, ZN => n122);
   U80 : NAND2_X1 port map( A1 => B(39), A2 => n159, ZN => n121);
   U81 : XNOR2_X1 port map( A => B(27), B => n40, ZN => net52524);
   U82 : XNOR2_X1 port map( A => net52524, B => A(27), ZN => SUM(27));
   U83 : OAI21_X1 port map( B1 => n37, B2 => n36, A => n38, ZN => n40);
   U84 : INV_X1 port map( A => A(26), ZN => n37);
   U85 : OAI21_X1 port map( B1 => n37, B2 => n36, A => n38, ZN => net52348);
   U86 : OAI21_X1 port map( B1 => net52348, B2 => B(27), A => A(27), ZN => 
                           net52356);
   U87 : NAND2_X1 port map( A1 => net52348, A2 => B(27), ZN => net52355);
   U88 : NOR2_X1 port map( A1 => net52575, A2 => B(26), ZN => n36);
   U89 : NAND2_X1 port map( A1 => net52342, A2 => B(26), ZN => n38);
   U90 : XNOR2_X1 port map( A => n35, B => n39, ZN => SUM(26));
   U91 : XNOR2_X1 port map( A => net52342, B => B(26), ZN => n39);
   U92 : NAND2_X1 port map( A1 => net52356, A2 => net52355, ZN => n41);
   U93 : AND2_X1 port map( A1 => n98, A2 => n131, ZN => n42);
   U94 : NAND2_X1 port map( A1 => B(36), A2 => n111, ZN => n116);
   U95 : NOR2_X1 port map( A1 => n176, A2 => B(21), ZN => n43);
   U96 : NOR2_X1 port map( A1 => B(22), A2 => n67, ZN => n44);
   U97 : XNOR2_X1 port map( A => A(43), B => B(43), ZN => n45);
   U98 : OAI21_X1 port map( B1 => n100, B2 => n14, A => n102, ZN => n46);
   U99 : XNOR2_X1 port map( A => n147, B => n80, ZN => SUM(24));
   U100 : OAI21_X1 port map( B1 => n172, B2 => n105, A => n16, ZN => n47);
   U101 : NAND2_X1 port map( A1 => n113, A2 => n112, ZN => n111);
   U102 : XNOR2_X1 port map( A => n141, B => n14, ZN => SUM(32));
   U103 : INV_X1 port map( A => A(29), ZN => n90);
   U104 : XNOR2_X1 port map( A => n145, B => n87, ZN => SUM(28));
   U105 : INV_X1 port map( A => A(16), ZN => n50);
   U106 : XNOR2_X1 port map( A => n150, B => n69, ZN => SUM(21));
   U107 : XNOR2_X1 port map( A => n151, B => n65, ZN => SUM(20));
   U108 : XNOR2_X1 port map( A => net51441, B => n122, ZN => SUM(41));
   U109 : NAND2_X1 port map( A1 => n122, A2 => n179, ZN => net45991);
   U110 : NAND2_X1 port map( A1 => n122, A2 => B(41), ZN => net45992);
   U111 : NAND2_X1 port map( A1 => B(24), A2 => n75, ZN => n81);
   U112 : XNOR2_X1 port map( A => n75, B => n127, ZN => n147);
   U113 : NAND2_X1 port map( A1 => n77, A2 => n76, ZN => n75);
   U114 : INV_X1 port map( A => A(36), ZN => n115);
   U115 : XNOR2_X1 port map( A => n146, B => n83, ZN => SUM(25));
   U116 : INV_X1 port map( A => A(32), ZN => n101);
   U117 : XNOR2_X1 port map( A => n144, B => n90, ZN => SUM(29));
   U118 : INV_X1 port map( A => A(21), ZN => n69);
   U119 : INV_X1 port map( A => A(17), ZN => n54);
   U120 : XNOR2_X1 port map( A => n136, B => net52413, ZN => SUM(37));
   U121 : OAI21_X1 port map( B1 => B(35), B2 => n166, A => A(35), ZN => n113);
   U122 : XNOR2_X1 port map( A => n155, B => n50, ZN => SUM(16));
   U123 : OAI21_X1 port map( B1 => net52418, B2 => net52419, A => net52420, ZN 
                           => n117);
   U124 : OAI21_X1 port map( B1 => net52419, B2 => net52418, A => net52420, ZN 
                           => n158);
   U125 : OAI21_X1 port map( B1 => net52564, B2 => net52419, A => net52420, ZN 
                           => n159);
   U126 : NOR2_X1 port map( A1 => B(33), A2 => n46, ZN => n104);
   U127 : OAI21_X1 port map( B1 => n104, B2 => n105, A => n106, ZN => n103);
   U128 : OAI21_X1 port map( B1 => n172, B2 => n105, A => n16, ZN => n160);
   U129 : NOR2_X1 port map( A1 => n175, A2 => B(29), ZN => n89);
   U130 : OAI21_X1 port map( B1 => n90, B2 => n174, A => n91, ZN => n161);
   U131 : OAI21_X1 port map( B1 => n174, B2 => n90, A => n91, ZN => n162);
   U132 : OAI21_X1 port map( B1 => n43, B2 => n69, A => n70, ZN => n67);
   U133 : NAND2_X1 port map( A1 => n163, A2 => B(22), ZN => n74);
   U134 : XNOR2_X1 port map( A => n163, B => B(22), ZN => n149);
   U135 : NOR2_X1 port map( A1 => n67, A2 => B(22), ZN => n72);
   U136 : NOR2_X1 port map( A1 => n63, A2 => B(21), ZN => n68);
   U137 : OAI21_X1 port map( B1 => n69, B2 => n68, A => n70, ZN => n163);
   U138 : OAI21_X1 port map( B1 => n54, B2 => n53, A => n55, ZN => n52);
   U139 : NAND2_X1 port map( A1 => n164, A2 => B(18), ZN => n59);
   U140 : XNOR2_X1 port map( A => n52, B => B(18), ZN => n153);
   U141 : NOR2_X1 port map( A1 => n164, A2 => B(18), ZN => n57);
   U142 : NOR2_X1 port map( A1 => B(17), A2 => n48, ZN => n53);
   U143 : OAI21_X1 port map( B1 => n33, B2 => n54, A => n55, ZN => n164);
   U144 : OAI21_X1 port map( B1 => n119, B2 => n120, A => n121, ZN => n118);
   U145 : NOR2_X1 port map( A1 => B(39), A2 => n117, ZN => n119);
   U146 : OAI21_X1 port map( B1 => n119, B2 => n120, A => n121, ZN => n165);
   U147 : NOR2_X1 port map( A1 => n103, A2 => B(34), ZN => n108);
   U148 : OAI21_X1 port map( B1 => n108, B2 => n109, A => n110, ZN => n107);
   U149 : OAI21_X1 port map( B1 => n108, B2 => n109, A => n110, ZN => n166);
   U150 : OAI21_X1 port map( B1 => n93, B2 => n94, A => n95, ZN => n92);
   U151 : OAI21_X1 port map( B1 => n93, B2 => n94, A => n95, ZN => n167);
   U152 : OAI21_X1 port map( B1 => n44, B2 => n73, A => n74, ZN => n71);
   U153 : NAND2_X1 port map( A1 => B(23), A2 => n168, ZN => n76);
   U154 : OAI21_X1 port map( B1 => B(23), B2 => n168, A => A(23), ZN => n77);
   U155 : XNOR2_X1 port map( A => n71, B => B(23), ZN => n148);
   U156 : OAI21_X1 port map( B1 => n72, B2 => n73, A => n74, ZN => n168);
   U157 : OAI21_X1 port map( B1 => n58, B2 => n57, A => n59, ZN => n56);
   U158 : NAND2_X1 port map( A1 => n169, A2 => B(19), ZN => n61);
   U159 : OAI21_X1 port map( B1 => n56, B2 => B(19), A => A(19), ZN => n62);
   U160 : XNOR2_X1 port map( A => n169, B => B(19), ZN => n152);
   U161 : OAI21_X1 port map( B1 => n57, B2 => n58, A => n59, ZN => n169);
   U162 : OAI21_X1 port map( B1 => n115, B2 => n114, A => n116, ZN => net52405)
                           ;
   U163 : XNOR2_X1 port map( A => n170, B => net52506, ZN => n136);
   U164 : NOR2_X1 port map( A1 => B(36), A2 => n111, ZN => n114);
   U165 : OAI21_X1 port map( B1 => n115, B2 => n114, A => n116, ZN => n170);
   U166 : OAI21_X1 port map( B1 => n79, B2 => n80, A => n81, ZN => n78);
   U167 : XNOR2_X1 port map( A => n78, B => n128, ZN => n146);
   U168 : NAND2_X1 port map( A1 => n171, A2 => B(25), ZN => n84);
   U169 : NOR2_X1 port map( A1 => n4, A2 => B(25), ZN => n82);
   U170 : OAI21_X1 port map( B1 => n80, B2 => n79, A => n81, ZN => n171);
   U171 : XNOR2_X1 port map( A => net52284, B => n123, ZN => n155);
   U172 : NAND2_X1 port map( A1 => n178, A2 => B(16), ZN => n51);
   U173 : NOR2_X1 port map( A1 => n178, A2 => B(16), ZN => n49);
   U174 : NOR2_X1 port map( A1 => n99, A2 => B(33), ZN => n172);
   U175 : OAI21_X1 port map( B1 => n14, B2 => n100, A => n102, ZN => n99);
   U176 : XNOR2_X1 port map( A => n19, B => n132, ZN => n140);
   U177 : NAND2_X1 port map( A1 => B(33), A2 => n173, ZN => n106);
   U178 : OAI21_X1 port map( B1 => n100, B2 => n101, A => n102, ZN => n173);
   U179 : NOR2_X1 port map( A1 => n85, A2 => B(29), ZN => n174);
   U180 : OAI21_X1 port map( B1 => n87, B2 => n22, A => n88, ZN => n85);
   U181 : XNOR2_X1 port map( A => n175, B => n130, ZN => n144);
   U182 : NAND2_X1 port map( A1 => n85, A2 => B(29), ZN => n91);
   U183 : NOR2_X1 port map( A1 => n41, A2 => B(28), ZN => n86);
   U184 : OAI21_X1 port map( B1 => n87, B2 => n86, A => n88, ZN => n175);
   U185 : NAND2_X1 port map( A1 => B(34), A2 => n160, ZN => n110);
   U186 : NAND2_X1 port map( A1 => B(30), A2 => n162, ZN => n95);
   U187 : INV_X1 port map( A => A(30), ZN => n94);
   U188 : XNOR2_X1 port map( A => n92, B => B(31), ZN => n142);
   U189 : NAND2_X1 port map( A1 => n167, A2 => B(31), ZN => n97);
   U190 : XNOR2_X1 port map( A => n107, B => B(35), ZN => n138);
   U191 : NAND2_X1 port map( A1 => n166, A2 => B(35), ZN => n112);
   U192 : OAI21_X1 port map( B1 => n17, B2 => n65, A => n66, ZN => n63);
   U193 : XNOR2_X1 port map( A => n176, B => n126, ZN => n150);
   U194 : NAND2_X1 port map( A1 => n63, A2 => B(21), ZN => n70);
   U195 : NOR2_X1 port map( A1 => n3, A2 => B(20), ZN => n64);
   U196 : OAI21_X1 port map( B1 => n65, B2 => n64, A => n66, ZN => n176);
   U197 : OAI21_X1 port map( B1 => n50, B2 => n18, A => n51, ZN => n48);
   U198 : XNOR2_X1 port map( A => n177, B => n124, ZN => n154);
   U199 : NAND2_X1 port map( A1 => n177, A2 => B(17), ZN => n55);
   U200 : OAI21_X1 port map( B1 => n49, B2 => n50, A => n51, ZN => n177);
   U201 : XNOR2_X1 port map( A => n47, B => B(34), ZN => n139);
   U202 : XNOR2_X1 port map( A => n134, B => n165, ZN => SUM(40));
   U203 : NAND2_X1 port map( A1 => B(40), A2 => n165, ZN => n157);
   U204 : XNOR2_X1 port map( A => n158, B => B(39), ZN => n135);
   U205 : XNOR2_X1 port map( A => n152, B => A(19), ZN => SUM(19));
   U206 : XNOR2_X1 port map( A => n138, B => n20, ZN => SUM(35));
   U207 : XNOR2_X1 port map( A => n148, B => A(23), ZN => SUM(23));
   U208 : XNOR2_X1 port map( A => n161, B => B(30), ZN => n143);
   U209 : XNOR2_X1 port map( A => n139, B => A(34), ZN => SUM(34));
   U210 : OAI21_X1 port map( B1 => n167, B2 => B(31), A => A(31), ZN => n98);
   U211 : XNOR2_X1 port map( A => n142, B => n21, ZN => SUM(31));
   U212 : XNOR2_X1 port map( A => n135, B => A(39), ZN => SUM(39));
   U213 : XNOR2_X1 port map( A => n153, B => A(18), ZN => SUM(18));
   U214 : XNOR2_X1 port map( A => n149, B => n34, ZN => SUM(22));
   U215 : XNOR2_X1 port map( A => n111, B => n133, ZN => n137);
   U216 : XNOR2_X1 port map( A => n115, B => n137, ZN => SUM(36));
   U217 : OAI21_X1 port map( B1 => B(40), B2 => n118, A => A(40), ZN => n156);
   U218 : OAI21_X1 port map( B1 => net52285, B2 => net52706, A => net52287, ZN 
                           => n178);
   U219 : INV_X1 port map( A => A(34), ZN => n109);
   U220 : INV_X1 port map( A => A(18), ZN => n58);
   U221 : XNOR2_X1 port map( A => n143, B => A(30), ZN => SUM(30));
   U222 : XNOR2_X1 port map( A => n140, B => n105, ZN => SUM(33));
   U223 : OAI21_X1 port map( B1 => n82, B2 => n83, A => n84, ZN => net52342);
   U224 : OAI21_X1 port map( B1 => n83, B2 => n82, A => n84, ZN => net52575);
   U225 : INV_X1 port map( A => A(22), ZN => n73);
   U226 : INV_X1 port map( A => A(39), ZN => n120);
   U227 : CLKBUF_X1 port map( A => A(41), Z => n179);
   U228 : INV_X1 port map( A => A(28), ZN => n87);
   U229 : INV_X1 port map( A => A(24), ZN => n80);
   U230 : XNOR2_X1 port map( A => n41, B => n129, ZN => n145);
   U231 : NAND2_X1 port map( A1 => B(28), A2 => n41, ZN => n88);
   U232 : XNOR2_X1 port map( A => n154, B => n54, ZN => SUM(17));
   U233 : INV_X1 port map( A => A(33), ZN => n105);
   U234 : NAND2_X1 port map( A1 => n62, A2 => n61, ZN => n60);
   U235 : NAND2_X1 port map( A1 => n98, A2 => n97, ZN => n96);
   U236 : INV_X1 port map( A => A(25), ZN => n83);
   U237 : INV_X1 port map( A => A(20), ZN => n65);
   U238 : XNOR2_X1 port map( A => n3, B => n125, ZN => n151);
   U239 : NAND2_X1 port map( A1 => n60, A2 => B(20), ZN => n66);
   U240 : XNOR2_X1 port map( A => n96, B => n131, ZN => n141);
   U241 : NAND2_X1 port map( A1 => n96, A2 => B(32), ZN => n102);
   U242 : XNOR2_X1 port map( A => A(41), B => B(41), ZN => net51441);
   U243 : NAND2_X1 port map( A1 => A(41), A2 => B(41), ZN => n180);
   U244 : NAND3_X1 port map( A1 => net45991, A2 => net45992, A3 => n180, ZN => 
                           carry_42_port);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT42_DW01_add_0 is

   port( A, B : in std_logic_vector (41 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (41 downto 0);  CO : out std_logic);

end RCA_NBIT42_DW01_add_0;

architecture SYN_rpl of RCA_NBIT42_DW01_add_0 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_41_port, carry_40_port, carry_39_port, carry_38_port, 
      carry_37_port, carry_36_port, carry_35_port, carry_34_port, carry_33_port
      , net55500, net58080, net58075, net58076, net58048, net58044, net57936, 
      net57935, net57934, net73543, net73542, net73541, net73568, net62414, 
      net52672, carry_32_port, carry_31_port, carry_30_port, carry_29_port, 
      carry_28_port, carry_27_port, carry_26_port, carry_25_port, carry_24_port
      , carry_23_port, carry_22_port, carry_21_port, carry_20_port, 
      carry_19_port, carry_18_port, net58099, net58043, net57939, net58042, 
      net57944, net52674, net52673, net62406, net58087, net58083, net58041, 
      net57959, net57957, net57953, net57951, net57950, net52797, n3, n4, n5, 
      n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, 
      n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35
      , n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, 
      n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64
      , n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
      n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, 
      n119, n120, n121, n122, n123 : std_logic;

begin
   
   U1_38 : FA_X1 port map( A => A(38), B => B(38), CI => carry_38_port, CO => 
                           carry_39_port, S => SUM(38));
   U1_37 : FA_X1 port map( A => A(37), B => B(37), CI => carry_37_port, CO => 
                           carry_38_port, S => SUM(37));
   U1_36 : FA_X1 port map( A => A(36), B => B(36), CI => carry_36_port, CO => 
                           carry_37_port, S => SUM(36));
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => carry_35_port, CO => 
                           carry_36_port, S => SUM(35));
   U1_34 : FA_X1 port map( A => A(34), B => B(34), CI => carry_34_port, CO => 
                           carry_35_port, S => SUM(34));
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U1 : CLKBUF_X1 port map( A => n14, Z => n3);
   U2 : NAND3_X1 port map( A1 => n15, A2 => n14, A3 => n16, ZN => n4);
   U3 : BUF_X1 port map( A => A(10), Z => n67);
   U4 : CLKBUF_X1 port map( A => carry_24_port, Z => n5);
   U5 : NAND3_X1 port map( A1 => n29, A2 => n30, A3 => n31, ZN => n6);
   U6 : CLKBUF_X1 port map( A => A(13), Z => n45);
   U7 : XOR2_X1 port map( A => A(24), B => B(24), Z => n7);
   U8 : XOR2_X1 port map( A => n5, B => n7, Z => SUM(24));
   U9 : NAND2_X1 port map( A1 => carry_24_port, A2 => A(24), ZN => n8);
   U10 : NAND2_X1 port map( A1 => carry_24_port, A2 => B(24), ZN => n9);
   U11 : NAND2_X1 port map( A1 => A(24), A2 => B(24), ZN => n10);
   U12 : NAND3_X1 port map( A1 => n8, A2 => n9, A3 => n10, ZN => carry_25_port)
                           ;
   U13 : NAND3_X1 port map( A1 => n15, A2 => n14, A3 => n16, ZN => n11);
   U14 : NAND3_X1 port map( A1 => n30, A2 => n31, A3 => n29, ZN => n12);
   U15 : INV_X1 port map( A => B(32), ZN => net73568);
   U16 : INV_X1 port map( A => B(8), ZN => n79);
   U17 : NAND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n82);
   U18 : NAND2_X1 port map( A1 => n82, A2 => n81, ZN => n109);
   U19 : INV_X1 port map( A => B(1), ZN => n81);
   U20 : INV_X1 port map( A => A(7), ZN => n93);
   U21 : INV_X1 port map( A => A(1), ZN => n83);
   U22 : XNOR2_X1 port map( A => B(1), B => n82, ZN => n107);
   U23 : XNOR2_X1 port map( A => A(0), B => n80, ZN => SUM(0));
   U24 : INV_X1 port map( A => B(0), ZN => n80);
   U25 : XNOR2_X1 port map( A => B(2), B => A(2), ZN => n105);
   U26 : NAND2_X1 port map( A1 => n111, A2 => n110, ZN => n106);
   U27 : NAND2_X1 port map( A1 => n108, A2 => B(1), ZN => n111);
   U28 : NAND2_X1 port map( A1 => A(1), A2 => n109, ZN => n110);
   U29 : INV_X1 port map( A => n82, ZN => n108);
   U30 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n103);
   U31 : OAI222_X1 port map( A1 => n112, A2 => n84, B1 => n112, B2 => n85, C1 
                           => n85, C2 => n84, ZN => n104);
   U32 : INV_X1 port map( A => n106, ZN => n112);
   U33 : INV_X1 port map( A => B(2), ZN => n84);
   U34 : INV_X1 port map( A => A(2), ZN => n85);
   U35 : XNOR2_X1 port map( A => B(4), B => A(4), ZN => n101);
   U36 : OAI222_X1 port map( A1 => n113, A2 => n86, B1 => n113, B2 => n87, C1 
                           => n87, C2 => n86, ZN => n102);
   U37 : INV_X1 port map( A => B(3), ZN => n86);
   U38 : INV_X1 port map( A => A(3), ZN => n87);
   U39 : INV_X1 port map( A => n104, ZN => n113);
   U40 : XNOR2_X1 port map( A => B(5), B => A(5), ZN => n99);
   U41 : OAI222_X1 port map( A1 => n114, A2 => n88, B1 => n114, B2 => n89, C1 
                           => n89, C2 => n88, ZN => n100);
   U42 : INV_X1 port map( A => B(4), ZN => n88);
   U43 : INV_X1 port map( A => A(4), ZN => n89);
   U44 : INV_X1 port map( A => n102, ZN => n114);
   U45 : XNOR2_X1 port map( A => B(6), B => A(6), ZN => n98);
   U46 : OAI222_X1 port map( A1 => n74, A2 => n75, B1 => n74, B2 => n76, C1 => 
                           n76, C2 => n75, ZN => n73);
   U47 : INV_X1 port map( A => B(5), ZN => n75);
   U48 : INV_X1 port map( A => A(5), ZN => n76);
   U49 : INV_X1 port map( A => n100, ZN => n74);
   U50 : XNOR2_X1 port map( A => B(7), B => A(7), ZN => n96);
   U51 : OAI21_X1 port map( B1 => n90, B2 => n91, A => n115, ZN => n97);
   U52 : INV_X1 port map( A => A(6), ZN => n91);
   U53 : NAND2_X1 port map( A1 => B(6), A2 => n73, ZN => n115);
   U54 : NOR2_X1 port map( A1 => B(6), A2 => n73, ZN => n90);
   U55 : OAI221_X1 port map( B1 => n116, B2 => n93, C1 => n116, C2 => n92, A =>
                           n117, ZN => n95);
   U56 : INV_X1 port map( A => B(7), ZN => n92);
   U57 : INV_X1 port map( A => n97, ZN => n116);
   U58 : NAND2_X1 port map( A1 => B(7), A2 => A(7), ZN => n117);
   U59 : INV_X1 port map( A => B(17), ZN => net62414);
   U60 : XNOR2_X1 port map( A => n107, B => n83, ZN => SUM(1));
   U61 : XNOR2_X1 port map( A => n105, B => n106, ZN => SUM(2));
   U62 : XNOR2_X1 port map( A => n103, B => n104, ZN => SUM(3));
   U63 : XNOR2_X1 port map( A => n101, B => n102, ZN => SUM(4));
   U64 : XNOR2_X1 port map( A => n99, B => n100, ZN => SUM(5));
   U65 : XNOR2_X1 port map( A => n98, B => n73, ZN => SUM(6));
   U66 : XNOR2_X1 port map( A => n96, B => n97, ZN => SUM(7));
   U67 : XNOR2_X1 port map( A => n94, B => n95, ZN => SUM(8));
   U68 : AND3_X1 port map( A1 => n68, A2 => n69, A3 => n70, ZN => net58080);
   U69 : XOR2_X1 port map( A => A(19), B => B(19), Z => n13);
   U70 : XOR2_X1 port map( A => n6, B => n13, Z => SUM(19));
   U71 : NAND2_X1 port map( A1 => n12, A2 => A(19), ZN => n14);
   U72 : NAND2_X1 port map( A1 => carry_19_port, A2 => B(19), ZN => n15);
   U73 : NAND2_X1 port map( A1 => A(19), A2 => B(19), ZN => n16);
   U74 : NAND3_X1 port map( A1 => n3, A2 => n15, A3 => n16, ZN => carry_20_port
                           );
   U75 : INV_X1 port map( A => B(11), ZN => net57935);
   U76 : XOR2_X1 port map( A => B(9), B => n58, Z => n17);
   U77 : OAI21_X1 port map( B1 => n41, B2 => n42, A => n43, ZN => n18);
   U78 : INV_X1 port map( A => n32, ZN => n19);
   U79 : XOR2_X1 port map( A => A(20), B => B(20), Z => n20);
   U80 : XOR2_X1 port map( A => carry_20_port, B => n20, Z => SUM(20));
   U81 : NAND2_X1 port map( A1 => n4, A2 => A(20), ZN => n21);
   U82 : NAND2_X1 port map( A1 => n11, A2 => B(20), ZN => n22);
   U83 : NAND2_X1 port map( A1 => A(20), A2 => B(20), ZN => n23);
   U84 : NAND3_X1 port map( A1 => n21, A2 => n22, A3 => n23, ZN => 
                           carry_21_port);
   U85 : AND3_X2 port map( A1 => n69, A2 => n68, A3 => n70, ZN => n24);
   U86 : NAND3_X1 port map( A1 => net52674, A2 => n40, A3 => net52673, ZN => 
                           n25);
   U87 : NAND3_X1 port map( A1 => net52673, A2 => net52674, A3 => n40, ZN => 
                           n26);
   U88 : NAND2_X1 port map( A1 => B(13), A2 => net58099, ZN => n27);
   U89 : XOR2_X1 port map( A => A(18), B => B(18), Z => n28);
   U90 : XOR2_X1 port map( A => n26, B => n28, Z => SUM(18));
   U91 : NAND2_X1 port map( A1 => n25, A2 => A(18), ZN => n29);
   U92 : NAND2_X1 port map( A1 => carry_18_port, A2 => B(18), ZN => n30);
   U93 : NAND2_X1 port map( A1 => A(18), A2 => B(18), ZN => n31);
   U94 : NAND3_X1 port map( A1 => n29, A2 => n30, A3 => n31, ZN => 
                           carry_19_port);
   U95 : INV_X1 port map( A => A(8), ZN => n32);
   U96 : NAND2_X1 port map( A1 => n36, A2 => n35, ZN => net52797);
   U97 : XOR2_X1 port map( A => net52797, B => net52672, Z => SUM(17));
   U98 : NAND2_X1 port map( A1 => net52797, A2 => A(17), ZN => net52673);
   U99 : NAND2_X1 port map( A1 => net52797, A2 => B(17), ZN => net52674);
   U100 : NAND2_X1 port map( A1 => net58087, A2 => B(16), ZN => n35);
   U101 : OAI21_X1 port map( B1 => n33, B2 => B(16), A => A(16), ZN => n36);
   U102 : OAI21_X1 port map( B1 => net57957, B2 => n34, A => net57959, ZN => 
                           n33);
   U103 : INV_X1 port map( A => A(15), ZN => n34);
   U104 : OAI21_X1 port map( B1 => net62406, B2 => n34, A => net57959, ZN => 
                           net58087);
   U105 : NOR2_X1 port map( A1 => net58083, A2 => B(15), ZN => net57957);
   U106 : XNOR2_X1 port map( A => net58087, B => n37, ZN => SUM(16));
   U107 : NOR2_X1 port map( A1 => net57950, A2 => B(15), ZN => net62406);
   U108 : XNOR2_X1 port map( A => B(16), B => A(16), ZN => n37);
   U109 : NAND2_X1 port map( A1 => net58083, A2 => B(15), ZN => net57959);
   U110 : XNOR2_X1 port map( A => A(15), B => B(15), ZN => net58041);
   U111 : OAI21_X1 port map( B1 => net57951, B2 => n38, A => net57953, ZN => 
                           net58083);
   U112 : INV_X1 port map( A => A(14), ZN => n38);
   U113 : OAI21_X1 port map( B1 => n39, B2 => n38, A => net57953, ZN => 
                           net57950);
   U114 : NOR2_X1 port map( A1 => net57944, A2 => B(14), ZN => net57951);
   U115 : XNOR2_X1 port map( A => net57950, B => net58041, ZN => SUM(15));
   U116 : XNOR2_X1 port map( A => A(14), B => B(14), ZN => net58042);
   U117 : NOR2_X1 port map( A1 => net57944, A2 => B(14), ZN => n39);
   U118 : NAND2_X1 port map( A1 => n18, A2 => B(14), ZN => net57953);
   U119 : NAND3_X1 port map( A1 => net52673, A2 => net52674, A3 => n40, ZN => 
                           carry_18_port);
   U120 : NAND2_X1 port map( A1 => A(17), A2 => B(17), ZN => n40);
   U121 : OAI21_X1 port map( B1 => n44, B2 => n42, A => n27, ZN => net57944);
   U122 : INV_X1 port map( A => n45, ZN => n42);
   U123 : NOR2_X1 port map( A1 => net57939, A2 => B(13), ZN => n44);
   U124 : XNOR2_X1 port map( A => n18, B => net58042, ZN => SUM(14));
   U125 : XNOR2_X1 port map( A => A(13), B => B(13), ZN => net58043);
   U126 : NOR2_X1 port map( A1 => net57939, A2 => B(13), ZN => n41);
   U127 : NAND2_X1 port map( A1 => net58099, A2 => B(13), ZN => n43);
   U128 : NAND2_X1 port map( A1 => n49, A2 => n46, ZN => net57939);
   U129 : OAI21_X1 port map( B1 => B(12), B2 => net58075, A => n48, ZN => n49);
   U130 : BUF_X1 port map( A => A(12), Z => n48);
   U131 : OAI21_X1 port map( B1 => net58075, B2 => B(12), A => n48, ZN => n47);
   U132 : XNOR2_X1 port map( A => net58043, B => net58099, ZN => SUM(13));
   U133 : NAND2_X1 port map( A1 => n47, A2 => n46, ZN => net58099);
   U134 : XNOR2_X1 port map( A => A(12), B => B(12), ZN => net58044);
   U135 : NAND2_X1 port map( A1 => B(12), A2 => net58076, ZN => n46);
   U136 : CLKBUF_X1 port map( A => net55500, Z => n50);
   U137 : CLKBUF_X1 port map( A => carry_32_port, Z => n51);
   U138 : CLKBUF_X1 port map( A => carry_26_port, Z => n52);
   U139 : XOR2_X1 port map( A => A(26), B => B(26), Z => n53);
   U140 : XOR2_X1 port map( A => n52, B => n53, Z => SUM(26));
   U141 : NAND2_X1 port map( A1 => carry_26_port, A2 => A(26), ZN => n54);
   U142 : NAND2_X1 port map( A1 => carry_26_port, A2 => B(26), ZN => n55);
   U143 : NAND2_X1 port map( A1 => A(26), A2 => B(26), ZN => n56);
   U144 : NAND3_X1 port map( A1 => n54, A2 => n55, A3 => n56, ZN => 
                           carry_27_port);
   U145 : XNOR2_X1 port map( A => n59, B => n57, ZN => SUM(39));
   U146 : XNOR2_X1 port map( A => A(39), B => B(39), ZN => n57);
   U147 : CLKBUF_X1 port map( A => A(9), Z => n58);
   U148 : NAND2_X1 port map( A1 => carry_32_port, A2 => B(32), ZN => net73543);
   U149 : NAND2_X1 port map( A1 => carry_32_port, A2 => A(32), ZN => net73542);
   U150 : XOR2_X1 port map( A => n51, B => net73541, Z => SUM(32));
   U151 : XNOR2_X1 port map( A => A(17), B => net62414, ZN => net52672);
   U152 : CLKBUF_X1 port map( A => carry_39_port, Z => n59);
   U153 : NAND3_X1 port map( A1 => n61, A2 => n62, A3 => n63, ZN => n60);
   U154 : NAND2_X1 port map( A1 => carry_39_port, A2 => A(39), ZN => n61);
   U155 : NAND2_X1 port map( A1 => carry_39_port, A2 => B(39), ZN => n62);
   U156 : NAND2_X1 port map( A1 => A(39), A2 => B(39), ZN => n63);
   U157 : NAND3_X1 port map( A1 => n61, A2 => n62, A3 => n63, ZN => 
                           carry_40_port);
   U158 : XNOR2_X1 port map( A => A(11), B => net57935, ZN => n64);
   U159 : XNOR2_X1 port map( A => n24, B => n64, ZN => SUM(11));
   U160 : NAND2_X1 port map( A1 => A(11), A2 => B(11), ZN => net57936);
   U161 : INV_X1 port map( A => A(11), ZN => net57934);
   U162 : INV_X1 port map( A => n66, ZN => n70);
   U163 : AND2_X1 port map( A1 => A(10), A2 => B(10), ZN => n66);
   U164 : NAND2_X1 port map( A1 => net58048, A2 => B(10), ZN => n69);
   U165 : NAND2_X1 port map( A1 => net58048, A2 => n67, ZN => n68);
   U166 : XNOR2_X1 port map( A => A(10), B => B(10), ZN => n65);
   U167 : XNOR2_X1 port map( A => net58048, B => n65, ZN => SUM(10));
   U168 : XNOR2_X1 port map( A => carry_41_port, B => n71, ZN => SUM(41));
   U169 : XNOR2_X1 port map( A => A(41), B => B(41), ZN => n71);
   U170 : XNOR2_X1 port map( A => A(32), B => net73568, ZN => net73541);
   U171 : NAND2_X1 port map( A1 => A(32), A2 => B(32), ZN => n72);
   U172 : NAND3_X1 port map( A1 => net73542, A2 => net73543, A3 => n72, ZN => 
                           carry_33_port);
   U173 : XNOR2_X1 port map( A => B(8), B => n19, ZN => n94);
   U174 : OAI221_X1 port map( B1 => net58080, B2 => net57934, C1 => n24, C2 => 
                           net57935, A => net57936, ZN => net58076);
   U175 : OAI221_X1 port map( B1 => net58080, B2 => net57934, C1 => n24, C2 => 
                           net57935, A => net57936, ZN => net58075);
   U176 : INV_X1 port map( A => n95, ZN => n78);
   U177 : OAI222_X1 port map( A1 => n78, A2 => n79, B1 => n78, B2 => n32, C1 =>
                           n32, C2 => n79, ZN => n77);
   U178 : OAI222_X1 port map( A1 => n78, A2 => n79, B1 => n78, B2 => n32, C1 =>
                           n32, C2 => n79, ZN => net55500);
   U179 : NAND2_X1 port map( A1 => B(9), A2 => net55500, ZN => n119);
   U180 : NAND2_X1 port map( A1 => n119, A2 => n118, ZN => net58048);
   U181 : OAI21_X1 port map( B1 => n77, B2 => B(9), A => A(9), ZN => n118);
   U182 : XNOR2_X1 port map( A => net58076, B => net58044, ZN => SUM(12));
   U183 : XOR2_X1 port map( A => n50, B => n17, Z => SUM(9));
   U184 : XOR2_X1 port map( A => A(40), B => B(40), Z => n120);
   U185 : XOR2_X1 port map( A => carry_40_port, B => n120, Z => SUM(40));
   U186 : NAND2_X1 port map( A1 => n60, A2 => A(40), ZN => n121);
   U187 : NAND2_X1 port map( A1 => n60, A2 => B(40), ZN => n122);
   U188 : NAND2_X1 port map( A1 => A(40), A2 => B(40), ZN => n123);
   U189 : NAND3_X1 port map( A1 => n121, A2 => n122, A3 => n123, ZN => 
                           carry_41_port);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT40_DW01_add_0 is

   port( A, B : in std_logic_vector (39 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (39 downto 0);  CO : out std_logic);

end RCA_NBIT40_DW01_add_0;

architecture SYN_rpl of RCA_NBIT40_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_39_port, carry_38_port, carry_37_port, carry_36_port, 
      carry_35_port, carry_34_port, carry_33_port, carry_32_port, carry_31_port
      , carry_30_port, carry_29_port, carry_28_port, carry_27_port, 
      carry_26_port, carry_25_port, carry_24_port, carry_23_port, carry_22_port
      , carry_21_port, carry_20_port, carry_19_port, carry_18_port, 
      carry_17_port, carry_16_port, carry_6_port, carry_5_port, carry_4_port, 
      carry_3_port, carry_2_port, n1, net43092, net52752, net52751, net55496, 
      net62409, net42117, net42116, net42115, net79905, net82393, net82360, 
      net82357, net82309, net82308, net82307, net82293, net82477, net82495, 
      net82392, net82303, net82301, net82300, n3, n4, n5, n6, n7, n8, n9, n10, 
      n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25
      , n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, 
      n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54
      , n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, 
      n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83
      , n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, 
      n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, 
      n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, 
      n122, n123, n124, n125, n126, n127, n128 : std_logic;

begin
   
   U1_38 : FA_X1 port map( A => A(38), B => B(38), CI => carry_38_port, CO => 
                           carry_39_port, S => SUM(38));
   U1_37 : FA_X1 port map( A => A(37), B => B(37), CI => carry_37_port, CO => 
                           carry_38_port, S => SUM(37));
   U1_36 : FA_X1 port map( A => A(36), B => B(36), CI => carry_36_port, CO => 
                           carry_37_port, S => SUM(36));
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => carry_35_port, CO => 
                           carry_36_port, S => SUM(35));
   U1_34 : FA_X1 port map( A => A(34), B => B(34), CI => carry_34_port, CO => 
                           carry_35_port, S => SUM(34));
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => carry_32_port, CO => 
                           carry_33_port, S => SUM(32));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : XNOR2_X1 port map( A => carry_30_port, B => n3, ZN => SUM(30));
   U3 : XOR2_X1 port map( A => A(30), B => n53, Z => n3);
   U4 : CLKBUF_X1 port map( A => carry_20_port, Z => n4);
   U5 : CLKBUF_X1 port map( A => n118, Z => n5);
   U6 : CLKBUF_X1 port map( A => n51, Z => n6);
   U7 : CLKBUF_X1 port map( A => n60, Z => n25);
   U8 : NAND2_X1 port map( A1 => n96, A2 => B(17), ZN => n7);
   U9 : CLKBUF_X1 port map( A => n41, Z => n8);
   U10 : NAND2_X1 port map( A1 => net82393, A2 => B(10), ZN => n9);
   U11 : CLKBUF_X1 port map( A => n77, Z => n19);
   U12 : CLKBUF_X1 port map( A => n81, Z => n10);
   U13 : CLKBUF_X1 port map( A => A(8), Z => n11);
   U14 : CLKBUF_X1 port map( A => n114, Z => n12);
   U15 : XNOR2_X1 port map( A => n4, B => n13, ZN => SUM(20));
   U16 : XNOR2_X1 port map( A => A(20), B => B(20), ZN => n13);
   U17 : NAND2_X1 port map( A1 => carry_20_port, A2 => A(20), ZN => n14);
   U18 : NAND2_X1 port map( A1 => carry_20_port, A2 => B(20), ZN => n15);
   U19 : NAND2_X1 port map( A1 => A(20), A2 => B(20), ZN => n16);
   U20 : NAND3_X1 port map( A1 => n14, A2 => n15, A3 => n16, ZN => 
                           carry_21_port);
   U21 : INV_X1 port map( A => B(12), ZN => n27);
   U22 : OR2_X1 port map( A1 => A(11), A2 => B(11), ZN => n39);
   U23 : NOR2_X1 port map( A1 => n37, A2 => n28, ZN => net82301);
   U24 : INV_X1 port map( A => B(8), ZN => n56);
   U25 : INV_X1 port map( A => B(25), ZN => n52);
   U26 : INV_X1 port map( A => B(31), ZN => n54);
   U27 : INV_X1 port map( A => B(30), ZN => n53);
   U28 : INV_X1 port map( A => B(22), ZN => n82);
   U29 : INV_X1 port map( A => B(23), ZN => n99);
   U30 : CLKBUF_X1 port map( A => A(8), Z => n17);
   U31 : XNOR2_X1 port map( A => carry_17_port, B => n18, ZN => SUM(17));
   U32 : XNOR2_X1 port map( A => A(17), B => B(17), ZN => n18);
   U33 : BUF_X1 port map( A => A(9), Z => n80);
   U34 : NAND2_X1 port map( A1 => n26, A2 => B(12), ZN => n20);
   U35 : NAND2_X1 port map( A1 => n38, A2 => n40, ZN => n21);
   U36 : BUF_X1 port map( A => n76, Z => n22);
   U37 : OAI211_X1 port map( C1 => n48, C2 => n56, A => n77, B => n58, ZN => 
                           n23);
   U38 : BUF_X1 port map( A => A(12), Z => n45);
   U39 : NOR2_X1 port map( A1 => net82300, A2 => B(13), ZN => n24);
   U40 : CLKBUF_X1 port map( A => A(7), Z => net55496);
   U41 : BUF_X1 port map( A => A(15), Z => n50);
   U42 : XNOR2_X1 port map( A => n64, B => n61, ZN => net43092);
   U43 : NAND3_X1 port map( A1 => n9, A2 => n33, A3 => net82477, ZN => n32);
   U44 : NAND3_X1 port map( A1 => n35, A2 => n33, A3 => net82477, ZN => n34);
   U45 : NAND2_X1 port map( A1 => net82393, A2 => B(10), ZN => n35);
   U46 : NAND2_X1 port map( A1 => n36, A2 => B(11), ZN => n30);
   U47 : NAND2_X1 port map( A1 => n39, A2 => n32, ZN => n29);
   U48 : NAND2_X1 port map( A1 => n38, A2 => n40, ZN => n26);
   U49 : NAND2_X1 port map( A1 => n29, A2 => n40, ZN => net82293);
   U50 : CLKBUF_X1 port map( A => A(11), Z => n36);
   U51 : NAND2_X1 port map( A1 => B(10), A2 => A(10), ZN => n33);
   U52 : XNOR2_X1 port map( A => B(10), B => A(10), ZN => net82360);
   U53 : AND2_X1 port map( A1 => n34, A2 => n39, ZN => n37);
   U54 : XNOR2_X1 port map( A => n31, B => n32, ZN => SUM(11));
   U55 : XNOR2_X1 port map( A => A(11), B => B(11), ZN => n31);
   U56 : NAND2_X1 port map( A1 => n30, A2 => n27, ZN => n28);
   U57 : NAND2_X1 port map( A1 => n39, A2 => n34, ZN => n38);
   U58 : NAND2_X1 port map( A1 => n36, A2 => B(11), ZN => n40);
   U59 : NAND2_X1 port map( A1 => n26, A2 => B(12), ZN => net82303);
   U60 : NAND3_X1 port map( A1 => n110, A2 => n109, A3 => n108, ZN => n41);
   U61 : CLKBUF_X1 port map( A => A(6), Z => n94);
   U62 : XNOR2_X1 port map( A => A(13), B => B(13), ZN => n42);
   U63 : XNOR2_X1 port map( A => n42, B => net82495, ZN => SUM(13));
   U64 : INV_X1 port map( A => A(13), ZN => net82308);
   U65 : NAND2_X1 port map( A1 => net82392, A2 => B(13), ZN => net82309);
   U66 : NOR2_X1 port map( A1 => net82300, A2 => B(13), ZN => net82307);
   U67 : BUF_X1 port map( A => net82392, Z => net82495);
   U68 : OAI21_X1 port map( B1 => net82301, B2 => n43, A => n20, ZN => net82392
                           );
   U69 : INV_X1 port map( A => n45, ZN => n43);
   U70 : OAI21_X1 port map( B1 => n44, B2 => n43, A => net82303, ZN => net82300
                           );
   U71 : XNOR2_X1 port map( A => A(12), B => B(12), ZN => net82357);
   U72 : NOR2_X1 port map( A1 => net82293, A2 => B(12), ZN => n44);
   U73 : OAI211_X1 port map( C1 => n48, C2 => n56, A => n57, B => n58, ZN => 
                           n46);
   U74 : OR2_X1 port map( A1 => A(7), A2 => B(7), ZN => n69);
   U75 : INV_X1 port map( A => B(7), ZN => n61);
   U76 : OAI21_X1 port map( B1 => n46, B2 => B(9), A => n80, ZN => n47);
   U77 : XNOR2_X1 port map( A => n75, B => n74, ZN => SUM(9));
   U78 : AND2_X1 port map( A1 => n70, A2 => n71, ZN => n48);
   U79 : CLKBUF_X1 port map( A => net52752, Z => n49);
   U80 : NAND2_X1 port map( A1 => net55496, A2 => B(7), ZN => n71);
   U81 : NAND2_X1 port map( A1 => n68, A2 => A(10), ZN => net82477);
   U82 : NAND3_X1 port map( A1 => n123, A2 => n122, A3 => n121, ZN => n51);
   U83 : XNOR2_X1 port map( A => A(25), B => n52, ZN => n89);
   U84 : XNOR2_X1 port map( A => n65, B => n78, ZN => SUM(8));
   U85 : XNOR2_X1 port map( A => A(31), B => n54, ZN => n124);
   U86 : NAND3_X1 port map( A1 => net42116, A2 => net42117, A3 => net42115, ZN 
                           => n64);
   U87 : XNOR2_X1 port map( A => net82357, B => n21, ZN => SUM(12));
   U88 : NAND2_X1 port map( A1 => n72, A2 => n47, ZN => n68);
   U89 : OAI21_X1 port map( B1 => n24, B2 => net82308, A => net82309, ZN => n59
                           );
   U90 : NAND2_X1 port map( A1 => n76, A2 => B(14), ZN => n73);
   U91 : XNOR2_X1 port map( A => n67, B => n22, ZN => SUM(14));
   U92 : NOR2_X1 port map( A1 => n59, A2 => B(14), ZN => n62);
   U93 : NAND2_X1 port map( A1 => n66, A2 => n11, ZN => n57);
   U94 : OAI211_X1 port map( C1 => n48, C2 => n56, A => n57, B => n58, ZN => 
                           n55);
   U95 : OAI211_X1 port map( C1 => n48, C2 => n56, A => n19, B => n58, ZN => 
                           n75);
   U96 : OAI21_X1 port map( B1 => net82307, B2 => net82308, A => net82309, ZN 
                           => n76);
   U97 : OAI21_X1 port map( B1 => n62, B2 => n63, A => n73, ZN => n60);
   U98 : XNOR2_X1 port map( A => n25, B => net62409, ZN => SUM(15));
   U99 : NAND2_X1 port map( A1 => n60, A2 => n50, ZN => net52751);
   U100 : NAND2_X1 port map( A1 => n60, A2 => B(15), ZN => net52752);
   U101 : NAND2_X1 port map( A1 => n72, A2 => n79, ZN => net82393);
   U102 : NAND2_X1 port map( A1 => n78, A2 => n17, ZN => n77);
   U103 : NAND2_X1 port map( A1 => n69, A2 => n64, ZN => n70);
   U104 : NAND2_X1 port map( A1 => n70, A2 => n71, ZN => n66);
   U105 : NAND2_X1 port map( A1 => n70, A2 => n71, ZN => n78);
   U106 : XNOR2_X1 port map( A => net82393, B => net82360, ZN => SUM(10));
   U107 : OAI21_X1 port map( B1 => n55, B2 => B(9), A => n80, ZN => n79);
   U108 : NAND2_X1 port map( A1 => n23, A2 => B(9), ZN => n72);
   U109 : XNOR2_X1 port map( A => A(9), B => B(9), ZN => n74);
   U110 : XNOR2_X1 port map( A => A(8), B => B(8), ZN => n65);
   U111 : NAND2_X1 port map( A1 => A(8), A2 => B(8), ZN => n58);
   U112 : XNOR2_X1 port map( A => A(14), B => B(14), ZN => n67);
   U113 : INV_X1 port map( A => A(14), ZN => n63);
   U114 : NAND2_X1 port map( A1 => n97, A2 => A(16), ZN => n81);
   U115 : XNOR2_X1 port map( A => A(22), B => n82, ZN => n103);
   U116 : CLKBUF_X1 port map( A => net52751, Z => net79905);
   U117 : NAND2_X1 port map( A1 => A(15), A2 => B(15), ZN => n111);
   U118 : NAND3_X1 port map( A1 => n81, A2 => n114, A3 => n112, ZN => n83);
   U119 : NAND3_X1 port map( A1 => n86, A2 => n87, A3 => n88, ZN => n84);
   U120 : XOR2_X1 port map( A => A(24), B => B(24), Z => n85);
   U121 : XOR2_X1 port map( A => n85, B => n8, Z => SUM(24));
   U122 : NAND2_X1 port map( A1 => A(24), A2 => B(24), ZN => n86);
   U123 : NAND2_X1 port map( A1 => A(24), A2 => n41, ZN => n87);
   U124 : NAND2_X1 port map( A1 => B(24), A2 => carry_24_port, ZN => n88);
   U125 : NAND3_X1 port map( A1 => n86, A2 => n87, A3 => n88, ZN => 
                           carry_25_port);
   U126 : XOR2_X1 port map( A => n89, B => n84, Z => SUM(25));
   U127 : NAND2_X1 port map( A1 => A(25), A2 => B(25), ZN => n90);
   U128 : NAND2_X1 port map( A1 => A(25), A2 => carry_25_port, ZN => n91);
   U129 : NAND2_X1 port map( A1 => B(25), A2 => carry_25_port, ZN => n92);
   U130 : NAND3_X1 port map( A1 => n92, A2 => n91, A3 => n90, ZN => 
                           carry_26_port);
   U131 : NAND2_X1 port map( A1 => carry_6_port, A2 => n94, ZN => net42115);
   U132 : XOR2_X1 port map( A => n94, B => B(6), Z => n93);
   U133 : NAND2_X1 port map( A1 => carry_6_port, A2 => B(6), ZN => net42116);
   U134 : NAND2_X1 port map( A1 => A(6), A2 => B(6), ZN => net42117);
   U135 : XOR2_X1 port map( A => carry_6_port, B => n93, Z => SUM(6));
   U136 : XNOR2_X1 port map( A => n100, B => n95, ZN => SUM(18));
   U137 : NAND3_X1 port map( A1 => n5, A2 => n7, A3 => n120, ZN => n95);
   U138 : XNOR2_X1 port map( A => A(15), B => B(15), ZN => net62409);
   U139 : NAND3_X1 port map( A1 => n114, A2 => n113, A3 => n112, ZN => n96);
   U140 : NAND3_X1 port map( A1 => net52752, A2 => net52751, A3 => n111, ZN => 
                           n97);
   U141 : NAND3_X1 port map( A1 => net79905, A2 => n49, A3 => n111, ZN => n98);
   U142 : XNOR2_X1 port map( A => A(23), B => n99, ZN => n107);
   U143 : XNOR2_X1 port map( A => A(18), B => B(18), ZN => n100);
   U144 : XNOR2_X1 port map( A => n101, B => n98, ZN => SUM(16));
   U145 : XNOR2_X1 port map( A => A(16), B => B(16), ZN => n101);
   U146 : NAND3_X1 port map( A1 => n7, A2 => n118, A3 => n120, ZN => n102);
   U147 : XOR2_X1 port map( A => n103, B => carry_22_port, Z => SUM(22));
   U148 : NAND2_X1 port map( A1 => A(22), A2 => B(22), ZN => n104);
   U149 : NAND2_X1 port map( A1 => A(22), A2 => carry_22_port, ZN => n105);
   U150 : NAND2_X1 port map( A1 => carry_22_port, A2 => B(22), ZN => n106);
   U151 : NAND3_X1 port map( A1 => n104, A2 => n105, A3 => n106, ZN => 
                           carry_23_port);
   U152 : XOR2_X1 port map( A => n107, B => carry_23_port, Z => SUM(23));
   U153 : NAND2_X1 port map( A1 => A(23), A2 => B(23), ZN => n108);
   U154 : NAND2_X1 port map( A1 => carry_23_port, A2 => A(23), ZN => n109);
   U155 : NAND2_X1 port map( A1 => B(23), A2 => carry_23_port, ZN => n110);
   U156 : NAND3_X1 port map( A1 => n110, A2 => n109, A3 => n108, ZN => 
                           carry_24_port);
   U157 : NAND3_X1 port map( A1 => net52751, A2 => net52752, A3 => n111, ZN => 
                           carry_16_port);
   U158 : NAND2_X1 port map( A1 => A(16), A2 => B(16), ZN => n112);
   U159 : NAND2_X1 port map( A1 => n97, A2 => A(16), ZN => n113);
   U160 : NAND2_X1 port map( A1 => carry_16_port, A2 => B(16), ZN => n114);
   U161 : NAND3_X1 port map( A1 => n12, A2 => n10, A3 => n112, ZN => 
                           carry_17_port);
   U162 : NAND2_X1 port map( A1 => n102, A2 => A(18), ZN => n115);
   U163 : NAND2_X1 port map( A1 => carry_18_port, A2 => B(18), ZN => n116);
   U164 : NAND2_X1 port map( A1 => A(18), A2 => B(18), ZN => n117);
   U165 : NAND3_X1 port map( A1 => n115, A2 => n116, A3 => n117, ZN => 
                           carry_19_port);
   U166 : XOR2_X1 port map( A => net55496, B => net43092, Z => SUM(7));
   U167 : NAND2_X1 port map( A1 => n83, A2 => A(17), ZN => n118);
   U168 : NAND2_X1 port map( A1 => n96, A2 => B(17), ZN => n119);
   U169 : NAND2_X1 port map( A1 => A(17), A2 => B(17), ZN => n120);
   U170 : NAND3_X1 port map( A1 => n118, A2 => n120, A3 => n119, ZN => 
                           carry_18_port);
   U171 : NAND2_X1 port map( A1 => A(30), A2 => B(30), ZN => n121);
   U172 : NAND2_X1 port map( A1 => carry_30_port, A2 => A(30), ZN => n122);
   U173 : NAND2_X1 port map( A1 => B(30), A2 => carry_30_port, ZN => n123);
   U174 : NAND3_X1 port map( A1 => n123, A2 => n122, A3 => n121, ZN => 
                           carry_31_port);
   U175 : XOR2_X1 port map( A => n124, B => n6, Z => SUM(31));
   U176 : NAND2_X1 port map( A1 => A(31), A2 => B(31), ZN => n125);
   U177 : NAND2_X1 port map( A1 => A(31), A2 => n51, ZN => n126);
   U178 : NAND2_X1 port map( A1 => B(31), A2 => carry_31_port, ZN => n127);
   U179 : NAND3_X1 port map( A1 => n125, A2 => n126, A3 => n127, ZN => 
                           carry_32_port);
   U180 : XOR2_X2 port map( A => carry_39_port, B => n128, Z => SUM(39));
   U181 : XOR2_X1 port map( A => A(39), B => B(39), Z => n128);
   U182 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n1);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT38_DW01_add_0 is

   port( A, B : in std_logic_vector (37 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (37 downto 0);  CO : out std_logic);

end RCA_NBIT38_DW01_add_0;

architecture SYN_rpl of RCA_NBIT38_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_37_port, carry_36_port, carry_35_port, carry_34_port, 
      carry_33_port, carry_32_port, carry_31_port, carry_30_port, carry_29_port
      , carry_28_port, carry_27_port, carry_26_port, carry_25_port, 
      carry_23_port, carry_22_port, carry_21_port, carry_20_port, carry_19_port
      , carry_17_port, carry_13_port, carry_12_port, carry_11_port, 
      carry_5_port, carry_4_port, carry_3_port, carry_2_port, n1, net42046, 
      net42045, net42044, net42178, net42177, net43100, net41814, carry_6_port,
      net52801, net55136, net55123, net55122, net55117, net55092, net55291, 
      net58111, net65826, net52799, net43194, net43182, net42127, net42102, 
      net82557, net87234, net87250, net87249, net87580, net55091, carry_10_port
      , n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18
      , n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, 
      n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47
      , n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, 
      n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76
      , n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, 
      n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104
      , n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
      n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, 
      n129, n130, n131, n132, n133, n134, n135, n136, n137 : std_logic;

begin
   
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => carry_35_port, CO => 
                           carry_36_port, S => SUM(35));
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => carry_32_port, CO => 
                           carry_33_port, S => SUM(32));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           net58111, S => SUM(13));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : CLKBUF_X1 port map( A => A(25), Z => n3);
   U3 : XNOR2_X1 port map( A => A(19), B => n4, ZN => n98);
   U4 : INV_X32 port map( A => B(19), ZN => n4);
   U5 : NAND3_X1 port map( A1 => n18, A2 => n19, A3 => n20, ZN => n5);
   U6 : NAND3_X1 port map( A1 => n18, A2 => n19, A3 => n20, ZN => n6);
   U7 : NAND2_X1 port map( A1 => net82557, A2 => n8, ZN => n7);
   U8 : CLKBUF_X1 port map( A => A(15), Z => n8);
   U9 : XNOR2_X1 port map( A => n90, B => n9, ZN => SUM(12));
   U10 : XOR2_X1 port map( A => A(12), B => B(12), Z => n9);
   U11 : NAND2_X1 port map( A1 => n88, A2 => B(16), ZN => n10);
   U12 : XOR2_X1 port map( A => A(25), B => B(25), Z => n11);
   U13 : XOR2_X1 port map( A => carry_25_port, B => n11, Z => SUM(25));
   U14 : NAND2_X1 port map( A1 => carry_25_port, A2 => n3, ZN => n12);
   U15 : NAND2_X1 port map( A1 => carry_25_port, A2 => B(25), ZN => n13);
   U16 : NAND2_X1 port map( A1 => A(25), A2 => B(25), ZN => n14);
   U17 : NAND3_X1 port map( A1 => n12, A2 => n13, A3 => n14, ZN => 
                           carry_26_port);
   U18 : BUF_X1 port map( A => A(23), Z => n15);
   U19 : XOR2_X2 port map( A => carry_37_port, B => n137, Z => SUM(37));
   U20 : CLKBUF_X1 port map( A => A(21), Z => n16);
   U21 : XOR2_X1 port map( A => A(26), B => B(26), Z => n17);
   U22 : XOR2_X1 port map( A => n17, B => carry_26_port, Z => SUM(26));
   U23 : NAND2_X1 port map( A1 => A(26), A2 => B(26), ZN => n18);
   U24 : NAND2_X1 port map( A1 => A(26), A2 => carry_26_port, ZN => n19);
   U25 : NAND2_X1 port map( A1 => B(26), A2 => carry_26_port, ZN => n20);
   U26 : NAND3_X1 port map( A1 => n18, A2 => n19, A3 => n20, ZN => 
                           carry_27_port);
   U27 : XOR2_X1 port map( A => A(27), B => B(27), Z => n21);
   U28 : XOR2_X1 port map( A => n21, B => n6, Z => SUM(27));
   U29 : NAND2_X1 port map( A1 => A(27), A2 => B(27), ZN => n22);
   U30 : NAND2_X1 port map( A1 => A(27), A2 => n5, ZN => n23);
   U31 : NAND2_X1 port map( A1 => B(27), A2 => carry_27_port, ZN => n24);
   U32 : NAND3_X1 port map( A1 => n22, A2 => n23, A3 => n24, ZN => 
                           carry_28_port);
   U33 : NAND3_X1 port map( A1 => n64, A2 => n65, A3 => n66, ZN => n25);
   U34 : NAND3_X1 port map( A1 => n64, A2 => n65, A3 => n66, ZN => 
                           carry_21_port);
   U35 : BUF_X1 port map( A => A(17), Z => n59);
   U36 : XOR2_X1 port map( A => A(34), B => B(34), Z => n26);
   U37 : XOR2_X1 port map( A => carry_34_port, B => n26, Z => SUM(34));
   U38 : NAND2_X1 port map( A1 => carry_34_port, A2 => A(34), ZN => n27);
   U39 : NAND2_X1 port map( A1 => carry_34_port, A2 => B(34), ZN => n28);
   U40 : NAND2_X1 port map( A1 => A(34), A2 => B(34), ZN => n29);
   U41 : NAND3_X1 port map( A1 => n27, A2 => n28, A3 => n29, ZN => 
                           carry_35_port);
   U42 : XOR2_X1 port map( A => A(36), B => B(36), Z => n30);
   U43 : XOR2_X1 port map( A => carry_36_port, B => n30, Z => SUM(36));
   U44 : NAND2_X1 port map( A1 => carry_36_port, A2 => A(36), ZN => n31);
   U45 : NAND2_X1 port map( A1 => carry_36_port, A2 => B(36), ZN => n32);
   U46 : NAND2_X1 port map( A1 => A(36), A2 => B(36), ZN => n33);
   U47 : NAND3_X1 port map( A1 => n31, A2 => n32, A3 => n33, ZN => 
                           carry_37_port);
   U48 : XNOR2_X1 port map( A => n34, B => n79, ZN => SUM(24));
   U49 : XNOR2_X1 port map( A => A(24), B => B(24), ZN => n34);
   U50 : XNOR2_X1 port map( A => A(20), B => n35, ZN => n63);
   U51 : INV_X32 port map( A => B(20), ZN => n35);
   U52 : XNOR2_X1 port map( A => A(23), B => n36, ZN => n81);
   U53 : INV_X32 port map( A => B(23), ZN => n36);
   U54 : XOR2_X1 port map( A => A(21), B => B(21), Z => n37);
   U55 : XOR2_X1 port map( A => n25, B => n37, Z => SUM(21));
   U56 : NAND2_X1 port map( A1 => n25, A2 => n16, ZN => n38);
   U57 : NAND2_X1 port map( A1 => carry_21_port, A2 => B(21), ZN => n39);
   U58 : NAND2_X1 port map( A1 => n16, A2 => B(21), ZN => n40);
   U59 : NAND3_X1 port map( A1 => n38, A2 => n39, A3 => n40, ZN => 
                           carry_22_port);
   U60 : NAND2_X1 port map( A1 => B(6), A2 => net43100, ZN => net52799);
   U61 : XNOR2_X1 port map( A => net87249, B => net87250, ZN => SUM(9));
   U62 : XNOR2_X1 port map( A => n71, B => n67, ZN => SUM(16));
   U63 : INV_X1 port map( A => B(28), ZN => n62);
   U64 : XNOR2_X1 port map( A => net55117, B => net55136, ZN => SUM(8));
   U65 : NAND2_X1 port map( A1 => n41, A2 => n42, ZN => n43);
   U66 : NAND2_X1 port map( A1 => n43, A2 => net58111, ZN => n45);
   U67 : INV_X4 port map( A => B(14), ZN => n41);
   U68 : INV_X1 port map( A => A(14), ZN => n42);
   U69 : INV_X1 port map( A => B(9), ZN => n50);
   U70 : BUF_X1 port map( A => A(10), Z => net52801);
   U71 : NAND2_X1 port map( A1 => B(14), A2 => n47, ZN => n44);
   U72 : CLKBUF_X1 port map( A => A(14), Z => n47);
   U73 : XOR2_X1 port map( A => A(14), B => B(14), Z => net55291);
   U74 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => n46);
   U75 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => net82557);
   U76 : NAND2_X1 port map( A1 => n46, A2 => n8, ZN => net87580);
   U77 : NAND2_X1 port map( A1 => n46, A2 => B(15), ZN => net65826);
   U78 : NOR2_X1 port map( A1 => n55, A2 => n56, ZN => carry_10_port);
   U79 : NAND2_X1 port map( A1 => carry_10_port, A2 => B(10), ZN => net42178);
   U80 : NAND2_X1 port map( A1 => carry_10_port, A2 => net52801, ZN => net42177
                           );
   U81 : AND3_X1 port map( A1 => n53, A2 => n51, A3 => n52, ZN => n55);
   U82 : AND2_X1 port map( A1 => n49, A2 => n50, ZN => n56);
   U83 : NOR2_X1 port map( A1 => n56, A2 => n57, ZN => net87234);
   U84 : INV_X1 port map( A => A(9), ZN => n49);
   U85 : NAND2_X1 port map( A1 => A(9), A2 => B(9), ZN => n53);
   U86 : AND3_X1 port map( A1 => n53, A2 => n51, A3 => n52, ZN => n57);
   U87 : OAI21_X1 port map( B1 => n54, B2 => B(8), A => net55091, ZN => n51);
   U88 : NAND2_X1 port map( A1 => n51, A2 => n52, ZN => net87250);
   U89 : NAND2_X1 port map( A1 => n48, A2 => net55092, ZN => net55091);
   U90 : NAND2_X1 port map( A1 => net55123, A2 => net55122, ZN => n48);
   U91 : BUF_X1 port map( A => A(8), Z => n54);
   U92 : NAND2_X1 port map( A1 => n54, A2 => B(8), ZN => n52);
   U93 : XNOR2_X1 port map( A => A(9), B => B(9), ZN => net87249);
   U94 : XNOR2_X1 port map( A => A(8), B => B(8), ZN => net55117);
   U95 : NAND2_X1 port map( A1 => net55092, A2 => n48, ZN => net55136);
   U96 : NAND2_X1 port map( A1 => net82557, A2 => B(15), ZN => n58);
   U97 : BUF_X1 port map( A => A(20), Z => n61);
   U98 : NAND3_X1 port map( A1 => n99, A2 => n100, A3 => n101, ZN => n60);
   U99 : CLKBUF_X1 port map( A => carry_28_port, Z => n102);
   U100 : XNOR2_X1 port map( A => A(28), B => n62, ZN => n127);
   U101 : BUF_X1 port map( A => A(11), Z => n68);
   U102 : XOR2_X1 port map( A => n60, B => n63, Z => SUM(20));
   U103 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => n64);
   U104 : NAND2_X1 port map( A1 => carry_20_port, A2 => B(20), ZN => n65);
   U105 : NAND2_X1 port map( A1 => n61, A2 => B(20), ZN => n66);
   U106 : XNOR2_X1 port map( A => A(16), B => B(16), ZN => n67);
   U107 : XNOR2_X1 port map( A => n46, B => n69, ZN => SUM(15));
   U108 : XNOR2_X1 port map( A => A(15), B => B(15), ZN => n69);
   U109 : NAND2_X1 port map( A1 => carry_11_port, A2 => B(11), ZN => n70);
   U110 : OR2_X1 port map( A1 => A(7), A2 => B(7), ZN => net55123);
   U111 : NAND3_X1 port map( A1 => n7, A2 => n58, A3 => n91, ZN => n71);
   U112 : NAND2_X1 port map( A1 => carry_17_port, A2 => B(17), ZN => n72);
   U113 : NAND3_X1 port map( A1 => n72, A2 => n131, A3 => n133, ZN => n73);
   U114 : NAND3_X1 port map( A1 => n119, A2 => n10, A3 => n121, ZN => n74);
   U115 : CLKBUF_X1 port map( A => A(19), Z => n75);
   U116 : NAND3_X1 port map( A1 => n134, A2 => n135, A3 => n136, ZN => n76);
   U117 : NAND3_X1 port map( A1 => n119, A2 => n120, A3 => n121, ZN => n77);
   U118 : NAND3_X1 port map( A1 => n84, A2 => n83, A3 => n82, ZN => n78);
   U119 : NAND3_X1 port map( A1 => n84, A2 => n83, A3 => n82, ZN => n79);
   U120 : XNOR2_X1 port map( A => A(7), B => B(7), ZN => net42102);
   U121 : XNOR2_X1 port map( A => net42102, B => net42127, ZN => SUM(7));
   U122 : CLKBUF_X1 port map( A => A(7), Z => n80);
   U123 : NAND2_X1 port map( A1 => n80, A2 => B(7), ZN => net55092);
   U124 : NAND3_X1 port map( A1 => net43182, A2 => net52799, A3 => net43194, ZN
                           => net42127);
   U125 : NAND2_X1 port map( A1 => A(6), A2 => net43100, ZN => net43182);
   U126 : NAND3_X1 port map( A1 => net43182, A2 => net52799, A3 => net43194, ZN
                           => net55122);
   U127 : NAND2_X1 port map( A1 => A(6), A2 => B(6), ZN => net43194);
   U128 : XNOR2_X1 port map( A => A(6), B => B(6), ZN => net41814);
   U129 : BUF_X1 port map( A => A(28), Z => n94);
   U130 : XOR2_X1 port map( A => carry_23_port, B => n81, Z => SUM(23));
   U131 : NAND2_X1 port map( A1 => A(23), A2 => B(23), ZN => n82);
   U132 : NAND2_X1 port map( A1 => n15, A2 => carry_23_port, ZN => n83);
   U133 : NAND2_X1 port map( A1 => B(23), A2 => carry_23_port, ZN => n84);
   U134 : NAND2_X1 port map( A1 => A(24), A2 => B(24), ZN => n85);
   U135 : NAND2_X1 port map( A1 => A(24), A2 => n78, ZN => n86);
   U136 : NAND2_X1 port map( A1 => B(24), A2 => n78, ZN => n87);
   U137 : NAND3_X1 port map( A1 => n85, A2 => n86, A3 => n87, ZN => 
                           carry_25_port);
   U138 : NAND3_X1 port map( A1 => n7, A2 => net65826, A3 => n91, ZN => n88);
   U139 : NAND3_X1 port map( A1 => net87580, A2 => n58, A3 => n91, ZN => n89);
   U140 : AND3_X1 port map( A1 => n116, A2 => n70, A3 => n115, ZN => n90);
   U141 : NAND2_X1 port map( A1 => A(15), A2 => B(15), ZN => n91);
   U142 : BUF_X1 port map( A => A(18), Z => n93);
   U143 : XNOR2_X1 port map( A => n74, B => n92, ZN => SUM(17));
   U144 : XNOR2_X1 port map( A => A(17), B => B(17), ZN => n92);
   U145 : NAND3_X1 port map( A1 => n70, A2 => n116, A3 => n115, ZN => n95);
   U146 : XNOR2_X1 port map( A => net87234, B => n96, ZN => SUM(10));
   U147 : XNOR2_X1 port map( A => A(10), B => B(10), ZN => n96);
   U148 : XNOR2_X1 port map( A => n105, B => n97, ZN => SUM(11));
   U149 : XOR2_X1 port map( A => A(11), B => B(11), Z => n97);
   U150 : XOR2_X1 port map( A => net58111, B => net55291, Z => SUM(14));
   U151 : XOR2_X1 port map( A => n76, B => n98, Z => SUM(19));
   U152 : NAND2_X1 port map( A1 => n76, A2 => n75, ZN => n99);
   U153 : NAND2_X1 port map( A1 => carry_19_port, A2 => B(19), ZN => n100);
   U154 : NAND2_X1 port map( A1 => n75, A2 => B(19), ZN => n101);
   U155 : NAND3_X1 port map( A1 => n99, A2 => n100, A3 => n101, ZN => 
                           carry_20_port);
   U156 : NAND3_X1 port map( A1 => n131, A2 => n132, A3 => n133, ZN => n103);
   U157 : NAND3_X1 port map( A1 => n131, A2 => n72, A3 => n133, ZN => n104);
   U158 : AND3_X1 port map( A1 => net42177, A2 => net42178, A3 => n114, ZN => 
                           n105);
   U159 : XNOR2_X1 port map( A => n106, B => n104, ZN => SUM(18));
   U160 : XNOR2_X1 port map( A => A(18), B => B(18), ZN => n106);
   U161 : NAND2_X1 port map( A1 => n95, A2 => A(12), ZN => n107);
   U162 : NAND2_X1 port map( A1 => carry_12_port, A2 => B(12), ZN => n108);
   U163 : NAND2_X1 port map( A1 => A(12), A2 => B(12), ZN => n109);
   U164 : NAND3_X1 port map( A1 => n107, A2 => n108, A3 => n109, ZN => 
                           carry_13_port);
   U165 : NAND3_X1 port map( A1 => net42178, A2 => net42177, A3 => n114, ZN => 
                           n110);
   U166 : NAND3_X1 port map( A1 => net42044, A2 => net42045, A3 => net42046, ZN
                           => carry_6_port);
   U167 : XNOR2_X1 port map( A => net41814, B => carry_6_port, ZN => SUM(6));
   U168 : NAND3_X1 port map( A1 => net42044, A2 => net42045, A3 => net42046, ZN
                           => net43100);
   U169 : CLKBUF_X1 port map( A => A(5), Z => n111);
   U170 : NAND3_X1 port map( A1 => n124, A2 => n125, A3 => n126, ZN => n112);
   U171 : NAND3_X1 port map( A1 => n124, A2 => n125, A3 => n126, ZN => n113);
   U172 : NAND2_X1 port map( A1 => net52801, A2 => B(10), ZN => n114);
   U173 : NAND3_X1 port map( A1 => net42177, A2 => net42178, A3 => n114, ZN => 
                           carry_11_port);
   U174 : NAND2_X1 port map( A1 => n68, A2 => B(11), ZN => n115);
   U175 : NAND2_X1 port map( A1 => n110, A2 => n68, ZN => n116);
   U176 : NAND2_X1 port map( A1 => carry_11_port, A2 => B(11), ZN => n117);
   U177 : NAND3_X1 port map( A1 => n116, A2 => n117, A3 => n115, ZN => 
                           carry_12_port);
   U178 : CLKBUF_X1 port map( A => A(4), Z => n118);
   U179 : NAND2_X1 port map( A1 => n89, A2 => A(16), ZN => n119);
   U180 : NAND2_X1 port map( A1 => n88, A2 => B(16), ZN => n120);
   U181 : NAND2_X1 port map( A1 => A(16), A2 => B(16), ZN => n121);
   U182 : NAND3_X1 port map( A1 => n10, A2 => n119, A3 => n121, ZN => 
                           carry_17_port);
   U183 : XOR2_X1 port map( A => n113, B => B(5), Z => n122);
   U184 : XOR2_X1 port map( A => n111, B => n122, Z => SUM(5));
   U185 : NAND2_X1 port map( A1 => A(5), A2 => n112, ZN => net42044);
   U186 : NAND2_X1 port map( A1 => A(5), A2 => B(5), ZN => net42045);
   U187 : NAND2_X1 port map( A1 => carry_5_port, A2 => B(5), ZN => net42046);
   U188 : XOR2_X1 port map( A => n118, B => B(4), Z => n123);
   U189 : XOR2_X1 port map( A => carry_4_port, B => n123, Z => SUM(4));
   U190 : NAND2_X1 port map( A1 => carry_4_port, A2 => n118, ZN => n124);
   U191 : NAND2_X1 port map( A1 => carry_4_port, A2 => B(4), ZN => n125);
   U192 : NAND2_X1 port map( A1 => A(4), A2 => B(4), ZN => n126);
   U193 : NAND3_X1 port map( A1 => n124, A2 => n125, A3 => n126, ZN => 
                           carry_5_port);
   U194 : XOR2_X1 port map( A => n102, B => n127, Z => SUM(28));
   U195 : NAND2_X1 port map( A1 => n94, A2 => carry_28_port, ZN => n128);
   U196 : NAND2_X1 port map( A1 => carry_28_port, A2 => B(28), ZN => n129);
   U197 : NAND2_X1 port map( A1 => n94, A2 => B(28), ZN => n130);
   U198 : NAND3_X1 port map( A1 => n128, A2 => n129, A3 => n130, ZN => 
                           carry_29_port);
   U199 : NAND2_X1 port map( A1 => n77, A2 => n59, ZN => n131);
   U200 : NAND2_X1 port map( A1 => carry_17_port, A2 => B(17), ZN => n132);
   U201 : NAND2_X1 port map( A1 => n59, A2 => B(17), ZN => n133);
   U202 : NAND2_X1 port map( A1 => n73, A2 => n93, ZN => n134);
   U203 : NAND2_X1 port map( A1 => n103, A2 => B(18), ZN => n135);
   U204 : NAND2_X1 port map( A1 => n93, A2 => B(18), ZN => n136);
   U205 : NAND3_X1 port map( A1 => n135, A2 => n134, A3 => n136, ZN => 
                           carry_19_port);
   U206 : XOR2_X1 port map( A => A(37), B => B(37), Z => n137);
   U207 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n1);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT36_DW01_add_0 is

   port( A, B : in std_logic_vector (35 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (35 downto 0);  CO : out std_logic);

end RCA_NBIT36_DW01_add_0;

architecture SYN_rpl of RCA_NBIT36_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_35_port, carry_34_port, carry_33_port, carry_32_port, 
      carry_31_port, carry_30_port, carry_29_port, carry_28_port, carry_27_port
      , carry_26_port, carry_25_port, carry_24_port, carry_23_port, 
      carry_22_port, carry_21_port, carry_20_port, carry_19_port, carry_18_port
      , carry_15_port, carry_14_port, carry_13_port, carry_12_port, 
      carry_11_port, carry_10_port, carry_2_port, n1, net41723, net41782, 
      net41781, net41777, net41795, net42000, net42031, net42075, net42087, 
      net42085, net42095, net42103, net42248, net43189, net42093, net41972, 
      net41797, net41784, net41783, carry_5_port, net51473, net43087, net41728,
      net55627, net55615, net55614, net55610, net55598, net55590, net42083, 
      net41945, net41778, carry_3_port, net43114, net42242, net42173, net41837,
      carry_7_port, net42058, net42021, net42008, net41983, net41982, net41780,
      net41779, net41984, net42059, net41730, net41729, n3, n4, n5, n6, n7, n8,
      n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
      n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67
      , n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, 
      n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96
      , n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n_1030 : std_logic;

begin
   
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => carry_35_port, CO => 
                           n_1030, S => SUM(35));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => carry_32_port, CO => 
                           carry_33_port, S => SUM(32));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : NAND3_X1 port map( A1 => n81, A2 => n82, A3 => n83, ZN => n3);
   U3 : NAND3_X1 port map( A1 => n81, A2 => n82, A3 => n83, ZN => n4);
   U4 : NAND3_X1 port map( A1 => n20, A2 => n21, A3 => n22, ZN => n5);
   U5 : NAND2_X1 port map( A1 => net55590, A2 => B(9), ZN => n6);
   U6 : CLKBUF_X1 port map( A => n78, Z => n7);
   U7 : XOR2_X1 port map( A => B(31), B => A(31), Z => n8);
   U8 : XOR2_X1 port map( A => carry_31_port, B => n8, Z => SUM(31));
   U9 : NAND2_X1 port map( A1 => carry_31_port, A2 => B(31), ZN => n9);
   U10 : NAND2_X1 port map( A1 => carry_31_port, A2 => A(31), ZN => n10);
   U11 : NAND2_X1 port map( A1 => B(31), A2 => A(31), ZN => n11);
   U12 : NAND3_X1 port map( A1 => n9, A2 => n10, A3 => n11, ZN => carry_32_port
                           );
   U13 : NAND3_X1 port map( A1 => n71, A2 => n72, A3 => n73, ZN => n12);
   U14 : NAND3_X1 port map( A1 => n71, A2 => n72, A3 => n73, ZN => n13);
   U15 : NAND3_X1 port map( A1 => n94, A2 => n95, A3 => n96, ZN => n14);
   U16 : NAND3_X1 port map( A1 => n20, A2 => n21, A3 => n22, ZN => n15);
   U17 : XNOR2_X1 port map( A => n16, B => n138, ZN => SUM(17));
   U18 : AND3_X1 port map( A1 => n135, A2 => n136, A3 => n137, ZN => n16);
   U19 : NAND2_X1 port map( A1 => n75, A2 => B(17), ZN => n17);
   U20 : XNOR2_X1 port map( A => n98, B => n18, ZN => SUM(14));
   U21 : XNOR2_X1 port map( A => B(14), B => A(14), ZN => n18);
   U22 : XOR2_X1 port map( A => B(25), B => A(25), Z => n19);
   U23 : XOR2_X1 port map( A => n14, B => n19, Z => SUM(25));
   U24 : NAND2_X1 port map( A1 => n14, A2 => B(25), ZN => n20);
   U25 : NAND2_X1 port map( A1 => carry_25_port, A2 => A(25), ZN => n21);
   U26 : NAND2_X1 port map( A1 => B(25), A2 => A(25), ZN => n22);
   U27 : NAND3_X1 port map( A1 => n20, A2 => n21, A3 => n22, ZN => 
                           carry_26_port);
   U28 : NAND3_X1 port map( A1 => n63, A2 => n64, A3 => n65, ZN => n23);
   U29 : NAND3_X1 port map( A1 => n28, A2 => n27, A3 => n29, ZN => n24);
   U30 : XNOR2_X1 port map( A => n47, B => n25, ZN => SUM(20));
   U31 : XNOR2_X1 port map( A => B(20), B => A(20), ZN => n25);
   U32 : XNOR2_X1 port map( A => n4, B => n26, ZN => SUM(21));
   U33 : XNOR2_X1 port map( A => B(21), B => A(21), ZN => n26);
   U34 : NAND2_X1 port map( A1 => n3, A2 => B(21), ZN => n27);
   U35 : NAND2_X1 port map( A1 => carry_21_port, A2 => A(21), ZN => n28);
   U36 : NAND2_X1 port map( A1 => B(21), A2 => A(21), ZN => n29);
   U37 : NAND3_X1 port map( A1 => n27, A2 => n28, A3 => n29, ZN => 
                           carry_22_port);
   U38 : INV_X1 port map( A => n37, ZN => n40);
   U39 : NAND2_X1 port map( A1 => n38, A2 => A(9), ZN => net55615);
   U40 : NAND2_X1 port map( A1 => n99, A2 => net55598, ZN => n100);
   U41 : BUF_X1 port map( A => A(4), Z => net42093);
   U42 : INV_X1 port map( A => A(8), ZN => n35);
   U43 : XOR2_X1 port map( A => B(7), B => A(7), Z => n30);
   U44 : AND2_X1 port map( A1 => n37, A2 => A(9), ZN => n31);
   U45 : XOR2_X1 port map( A => A(8), B => B(8), Z => n32);
   U46 : NAND2_X1 port map( A1 => net42059, A2 => n31, ZN => net55614);
   U47 : NAND2_X1 port map( A1 => n35, A2 => n34, ZN => n37);
   U48 : NAND3_X1 port map( A1 => n107, A2 => n106, A3 => n108, ZN => n33);
   U49 : INV_X1 port map( A => n39, ZN => n38);
   U50 : NAND3_X1 port map( A1 => net41778, A2 => net41779, A3 => net41780, ZN 
                           => net42083);
   U51 : XOR2_X1 port map( A => A(9), B => B(9), Z => net55627);
   U52 : AOI21_X1 port map( B1 => net42059, B2 => n37, A => n38, ZN => n36);
   U53 : MUX2_X1 port map( A => net55610, B => net55627, S => n36, Z => SUM(9))
                           ;
   U54 : NAND3_X1 port map( A1 => net41728, A2 => n42, A3 => net41730, ZN => 
                           net42059);
   U55 : NAND2_X1 port map( A1 => net43114, A2 => A(7), ZN => n42);
   U56 : INV_X1 port map( A => B(8), ZN => n34);
   U57 : NAND2_X1 port map( A1 => A(8), A2 => B(8), ZN => n39);
   U58 : OAI21_X1 port map( B1 => n41, B2 => n40, A => n39, ZN => net55590);
   U59 : AND3_X1 port map( A1 => net41729, A2 => net41728, A3 => net41730, ZN 
                           => n41);
   U60 : AND3_X1 port map( A1 => net41729, A2 => net41728, A3 => net41730, ZN 
                           => net43087);
   U61 : NAND2_X1 port map( A1 => net43114, A2 => A(7), ZN => net41729);
   U62 : NAND2_X1 port map( A1 => B(7), A2 => A(7), ZN => net41730);
   U63 : AND2_X1 port map( A1 => net55614, A2 => net55615, ZN => n43);
   U64 : AND2_X1 port map( A1 => net55614, A2 => net55615, ZN => n44);
   U65 : AND2_X1 port map( A1 => net55614, A2 => net55615, ZN => n84);
   U66 : CLKBUF_X1 port map( A => net41782, Z => n45);
   U67 : NAND3_X1 port map( A1 => n86, A2 => n87, A3 => n88, ZN => n46);
   U68 : NAND3_X1 port map( A1 => n86, A2 => n87, A3 => n88, ZN => n47);
   U69 : XNOR2_X1 port map( A => n80, B => n48, ZN => SUM(15));
   U70 : XNOR2_X1 port map( A => B(15), B => A(15), ZN => n48);
   U71 : NAND3_X1 port map( A1 => n17, A2 => n139, A3 => n140, ZN => n49);
   U72 : NAND3_X1 port map( A1 => n17, A2 => n139, A3 => n140, ZN => n50);
   U73 : NAND3_X1 port map( A1 => n53, A2 => n54, A3 => n55, ZN => n51);
   U74 : XOR2_X1 port map( A => B(18), B => A(18), Z => n52);
   U75 : XOR2_X1 port map( A => n50, B => n52, Z => SUM(18));
   U76 : NAND2_X1 port map( A1 => n49, A2 => B(18), ZN => n53);
   U77 : NAND2_X1 port map( A1 => carry_18_port, A2 => A(18), ZN => n54);
   U78 : NAND2_X1 port map( A1 => B(18), A2 => A(18), ZN => n55);
   U79 : NAND3_X1 port map( A1 => n54, A2 => n53, A3 => n55, ZN => 
                           carry_19_port);
   U80 : NAND2_X1 port map( A1 => B(2), A2 => A(2), ZN => net41984);
   U81 : NAND3_X1 port map( A1 => net41982, A2 => net41983, A3 => net41984, ZN 
                           => carry_3_port);
   U82 : NAND3_X1 port map( A1 => net41982, A2 => net41983, A3 => net41984, ZN 
                           => net42008);
   U83 : NAND3_X1 port map( A1 => net41982, A2 => net41983, A3 => net41984, ZN 
                           => net42248);
   U84 : CLKBUF_X1 port map( A => B(2), Z => net42058);
   U85 : CLKBUF_X1 port map( A => A(2), Z => net42021);
   U86 : NAND2_X1 port map( A1 => net42008, A2 => A(3), ZN => net41779);
   U87 : AND3_X1 port map( A1 => net41779, A2 => net41778, A3 => net41780, ZN 
                           => net42103);
   U88 : NAND3_X1 port map( A1 => net41778, A2 => net41780, A3 => net41779, ZN 
                           => net41972);
   U89 : NAND2_X1 port map( A1 => B(3), A2 => A(3), ZN => net41780);
   U90 : XOR2_X1 port map( A => net41945, B => A(3), Z => net41777);
   U91 : NAND2_X1 port map( A1 => carry_2_port, A2 => net42058, ZN => net41982)
                           ;
   U92 : XOR2_X1 port map( A => net42058, B => net42021, Z => n56);
   U93 : NAND2_X1 port map( A1 => carry_2_port, A2 => net42021, ZN => net41983)
                           ;
   U94 : XOR2_X1 port map( A => carry_2_port, B => n56, Z => SUM(2));
   U95 : XNOR2_X1 port map( A => net42242, B => n30, ZN => SUM(7));
   U96 : AND3_X1 port map( A1 => n59, A2 => n57, A3 => n58, ZN => net42242);
   U97 : NAND2_X1 port map( A1 => carry_7_port, A2 => B(7), ZN => net41728);
   U98 : NAND2_X1 port map( A1 => net41837, A2 => A(6), ZN => n59);
   U99 : NAND3_X1 port map( A1 => n59, A2 => n57, A3 => n58, ZN => carry_7_port
                           );
   U100 : NAND3_X1 port map( A1 => n59, A2 => n57, A3 => n58, ZN => net43114);
   U101 : NAND3_X1 port map( A1 => net41783, A2 => net41782, A3 => net41784, ZN
                           => net41837);
   U102 : NAND2_X1 port map( A1 => B(6), A2 => A(6), ZN => n58);
   U103 : XOR2_X1 port map( A => B(6), B => A(6), Z => net41723);
   U104 : AND3_X1 port map( A1 => net41783, A2 => n45, A3 => net41784, ZN => 
                           net42095);
   U105 : NAND3_X1 port map( A1 => net51473, A2 => net41782, A3 => net41784, ZN
                           => net42173);
   U106 : NAND2_X1 port map( A1 => net42173, A2 => B(6), ZN => n57);
   U107 : NAND2_X1 port map( A1 => carry_13_port, A2 => B(13), ZN => n60);
   U108 : NAND2_X1 port map( A1 => n111, A2 => A(10), ZN => n61);
   U109 : XOR2_X1 port map( A => A(26), B => B(26), Z => n62);
   U110 : XOR2_X1 port map( A => n62, B => n5, Z => SUM(26));
   U111 : NAND2_X1 port map( A1 => A(26), A2 => B(26), ZN => n63);
   U112 : NAND2_X1 port map( A1 => A(26), A2 => n15, ZN => n64);
   U113 : NAND2_X1 port map( A1 => B(26), A2 => carry_26_port, ZN => n65);
   U114 : NAND3_X1 port map( A1 => n63, A2 => n64, A3 => n65, ZN => 
                           carry_27_port);
   U115 : XOR2_X1 port map( A => A(27), B => B(27), Z => n66);
   U116 : XOR2_X1 port map( A => n66, B => n23, Z => SUM(27));
   U117 : NAND2_X1 port map( A1 => A(27), A2 => B(27), ZN => n67);
   U118 : NAND2_X1 port map( A1 => A(27), A2 => carry_27_port, ZN => n68);
   U119 : NAND2_X1 port map( A1 => B(27), A2 => carry_27_port, ZN => n69);
   U120 : NAND3_X1 port map( A1 => n67, A2 => n68, A3 => n69, ZN => 
                           carry_28_port);
   U121 : XOR2_X1 port map( A => B(22), B => A(22), Z => n70);
   U122 : XOR2_X1 port map( A => carry_22_port, B => n70, Z => SUM(22));
   U123 : NAND2_X1 port map( A1 => n24, A2 => B(22), ZN => n71);
   U124 : NAND2_X1 port map( A1 => carry_22_port, A2 => A(22), ZN => n72);
   U125 : NAND2_X1 port map( A1 => B(22), A2 => A(22), ZN => n73);
   U126 : NAND3_X1 port map( A1 => n71, A2 => n72, A3 => n73, ZN => 
                           carry_23_port);
   U127 : NAND3_X1 port map( A1 => n115, A2 => n114, A3 => n116, ZN => n74);
   U128 : NAND3_X1 port map( A1 => n135, A2 => n136, A3 => n137, ZN => n75);
   U129 : NAND3_X1 port map( A1 => n91, A2 => n90, A3 => n92, ZN => n76);
   U130 : NAND3_X1 port map( A1 => n90, A2 => n91, A3 => n92, ZN => n77);
   U131 : NAND2_X1 port map( A1 => net42083, A2 => B(4), ZN => n78);
   U132 : AND3_X1 port map( A1 => net43189, A2 => n7, A3 => n79, ZN => net42031
                           );
   U133 : NAND3_X1 port map( A1 => net43189, A2 => n78, A3 => n79, ZN => 
                           carry_5_port);
   U134 : NAND3_X1 port map( A1 => n78, A2 => net41797, A3 => n79, ZN => 
                           net42075);
   U135 : NAND2_X1 port map( A1 => B(4), A2 => net42093, ZN => n79);
   U136 : XOR2_X1 port map( A => A(4), B => B(4), Z => net41795);
   U137 : NAND2_X1 port map( A1 => B(3), A2 => carry_3_port, ZN => net41778);
   U138 : CLKBUF_X1 port map( A => B(3), Z => net41945);
   U139 : NAND3_X1 port map( A1 => n106, A2 => n107, A3 => n108, ZN => n80);
   U140 : NAND2_X1 port map( A1 => n46, A2 => B(20), ZN => n81);
   U141 : NAND2_X1 port map( A1 => carry_20_port, A2 => A(20), ZN => n82);
   U142 : NAND2_X1 port map( A1 => B(20), A2 => A(20), ZN => n83);
   U143 : NAND3_X1 port map( A1 => n81, A2 => n82, A3 => n83, ZN => 
                           carry_21_port);
   U144 : XOR2_X1 port map( A => B(19), B => A(19), Z => n85);
   U145 : XOR2_X1 port map( A => carry_19_port, B => n85, Z => SUM(19));
   U146 : NAND2_X1 port map( A1 => n51, A2 => B(19), ZN => n86);
   U147 : NAND2_X1 port map( A1 => n51, A2 => A(19), ZN => n87);
   U148 : NAND2_X1 port map( A1 => B(19), A2 => A(19), ZN => n88);
   U149 : NAND3_X1 port map( A1 => n86, A2 => n87, A3 => n88, ZN => 
                           carry_20_port);
   U150 : XOR2_X1 port map( A => A(23), B => B(23), Z => n89);
   U151 : XOR2_X1 port map( A => n89, B => n13, Z => SUM(23));
   U152 : NAND2_X1 port map( A1 => A(23), A2 => B(23), ZN => n90);
   U153 : NAND2_X1 port map( A1 => A(23), A2 => n12, ZN => n91);
   U154 : NAND2_X1 port map( A1 => B(23), A2 => carry_23_port, ZN => n92);
   U155 : NAND3_X1 port map( A1 => n90, A2 => n91, A3 => n92, ZN => 
                           carry_24_port);
   U156 : XOR2_X1 port map( A => A(24), B => B(24), Z => n93);
   U157 : XOR2_X1 port map( A => n93, B => n77, Z => SUM(24));
   U158 : NAND2_X1 port map( A1 => A(24), A2 => B(24), ZN => n94);
   U159 : NAND2_X1 port map( A1 => A(24), A2 => n76, ZN => n95);
   U160 : NAND2_X1 port map( A1 => B(24), A2 => carry_24_port, ZN => n96);
   U161 : NAND3_X1 port map( A1 => n94, A2 => n95, A3 => n96, ZN => 
                           carry_25_port);
   U162 : NAND3_X1 port map( A1 => n131, A2 => n130, A3 => n132, ZN => n97);
   U163 : NAND3_X1 port map( A1 => n131, A2 => n130, A3 => n60, ZN => n98);
   U164 : INV_X1 port map( A => B(9), ZN => n99);
   U165 : NAND2_X1 port map( A1 => A(9), A2 => B(9), ZN => net42087);
   U166 : NAND2_X1 port map( A1 => net55590, A2 => B(9), ZN => net42085);
   U167 : NAND2_X1 port map( A1 => net42087, A2 => n100, ZN => net55610);
   U168 : INV_X1 port map( A => A(9), ZN => net55598);
   U169 : XNOR2_X1 port map( A => n113, B => n101, ZN => SUM(12));
   U170 : XNOR2_X1 port map( A => A(12), B => B(12), ZN => n101);
   U171 : XNOR2_X1 port map( A => carry_10_port, B => n102, ZN => SUM(10));
   U172 : XNOR2_X1 port map( A => B(10), B => A(10), ZN => n102);
   U173 : NAND3_X1 port map( A1 => n61, A2 => n123, A3 => n125, ZN => n103);
   U174 : NAND3_X1 port map( A1 => n61, A2 => n123, A3 => n125, ZN => n104);
   U175 : XNOR2_X1 port map( A => n104, B => n105, ZN => SUM(11));
   U176 : XNOR2_X1 port map( A => B(11), B => A(11), ZN => n105);
   U177 : NAND2_X1 port map( A1 => n97, A2 => B(14), ZN => n106);
   U178 : NAND2_X1 port map( A1 => carry_14_port, A2 => A(14), ZN => n107);
   U179 : NAND2_X1 port map( A1 => B(14), A2 => A(14), ZN => n108);
   U180 : NAND3_X1 port map( A1 => n107, A2 => n108, A3 => n106, ZN => 
                           carry_15_port);
   U181 : NAND3_X1 port map( A1 => n115, A2 => n114, A3 => n116, ZN => n109);
   U182 : NAND3_X1 port map( A1 => n114, A2 => n115, A3 => n116, ZN => n110);
   U183 : NAND3_X1 port map( A1 => n6, A2 => n43, A3 => net42087, ZN => n111);
   U184 : NAND3_X1 port map( A1 => net42085, A2 => n84, A3 => net42087, ZN => 
                           n112);
   U185 : NAND3_X1 port map( A1 => n120, A2 => n121, A3 => n122, ZN => n113);
   U186 : NAND2_X1 port map( A1 => carry_15_port, A2 => B(15), ZN => n114);
   U187 : NAND2_X1 port map( A1 => n33, A2 => A(15), ZN => n115);
   U188 : NAND2_X1 port map( A1 => B(15), A2 => A(15), ZN => n116);
   U189 : NAND3_X1 port map( A1 => n128, A2 => n127, A3 => n126, ZN => n117);
   U190 : NAND3_X1 port map( A1 => n128, A2 => n127, A3 => n126, ZN => n118);
   U191 : XNOR2_X1 port map( A => net43087, B => n32, ZN => SUM(8));
   U192 : NAND2_X1 port map( A1 => carry_5_port, A2 => n119, ZN => net51473);
   U193 : CLKBUF_X1 port map( A => A(5), Z => n119);
   U194 : NAND2_X1 port map( A1 => carry_5_port, A2 => n119, ZN => net41783);
   U195 : XOR2_X1 port map( A => B(5), B => A(5), Z => net41781);
   U196 : NAND2_X1 port map( A1 => B(5), A2 => A(5), ZN => net41784);
   U197 : NAND2_X1 port map( A1 => net41972, A2 => net42093, ZN => net43189);
   U198 : NAND2_X1 port map( A1 => net41972, A2 => net42093, ZN => net41797);
   U199 : NAND2_X1 port map( A1 => n103, A2 => B(11), ZN => n120);
   U200 : NAND2_X1 port map( A1 => carry_11_port, A2 => A(11), ZN => n121);
   U201 : NAND2_X1 port map( A1 => B(11), A2 => A(11), ZN => n122);
   U202 : NAND3_X1 port map( A1 => n120, A2 => n121, A3 => n122, ZN => 
                           carry_12_port);
   U203 : NAND2_X1 port map( A1 => n112, A2 => B(10), ZN => n123);
   U204 : NAND2_X1 port map( A1 => n111, A2 => A(10), ZN => n124);
   U205 : NAND2_X1 port map( A1 => B(10), A2 => A(10), ZN => n125);
   U206 : NAND3_X1 port map( A1 => n123, A2 => n124, A3 => n125, ZN => 
                           carry_11_port);
   U207 : XNOR2_X1 port map( A => net42103, B => net41795, ZN => SUM(4));
   U208 : XNOR2_X1 port map( A => net42095, B => net41723, ZN => SUM(6));
   U209 : NAND3_X1 port map( A1 => n6, A2 => n44, A3 => net42087, ZN => 
                           carry_10_port);
   U210 : XNOR2_X1 port map( A => net42031, B => net41781, ZN => SUM(5));
   U211 : CLKBUF_X1 port map( A => B(5), Z => net42000);
   U212 : NAND2_X1 port map( A1 => A(12), A2 => B(12), ZN => n126);
   U213 : NAND2_X1 port map( A1 => A(12), A2 => carry_12_port, ZN => n127);
   U214 : NAND2_X1 port map( A1 => n113, A2 => B(12), ZN => n128);
   U215 : NAND3_X1 port map( A1 => n128, A2 => n127, A3 => n126, ZN => 
                           carry_13_port);
   U216 : XOR2_X1 port map( A => A(13), B => B(13), Z => n129);
   U217 : XOR2_X1 port map( A => n129, B => n118, Z => SUM(13));
   U218 : NAND2_X1 port map( A1 => A(13), A2 => B(13), ZN => n130);
   U219 : NAND2_X1 port map( A1 => n117, A2 => A(13), ZN => n131);
   U220 : NAND2_X1 port map( A1 => carry_13_port, A2 => B(13), ZN => n132);
   U221 : NAND3_X1 port map( A1 => n60, A2 => n131, A3 => n130, ZN => 
                           carry_14_port);
   U222 : NAND3_X1 port map( A1 => n136, A2 => n135, A3 => n137, ZN => n133);
   U223 : XOR2_X1 port map( A => net42248, B => net41777, Z => SUM(3));
   U224 : NAND2_X1 port map( A1 => net42075, A2 => net42000, ZN => net41782);
   U225 : XOR2_X1 port map( A => B(16), B => A(16), Z => n134);
   U226 : XOR2_X1 port map( A => n110, B => n134, Z => SUM(16));
   U227 : NAND2_X1 port map( A1 => n74, A2 => B(16), ZN => n135);
   U228 : NAND2_X1 port map( A1 => n109, A2 => A(16), ZN => n136);
   U229 : NAND2_X1 port map( A1 => B(16), A2 => A(16), ZN => n137);
   U230 : XOR2_X1 port map( A => B(17), B => A(17), Z => n138);
   U231 : NAND2_X1 port map( A1 => n133, A2 => A(17), ZN => n139);
   U232 : NAND2_X1 port map( A1 => B(17), A2 => A(17), ZN => n140);
   U233 : NAND3_X1 port map( A1 => n139, A2 => n17, A3 => n140, ZN => 
                           carry_18_port);
   U234 : XOR2_X1 port map( A => B(33), B => A(33), Z => n141);
   U235 : XOR2_X1 port map( A => carry_33_port, B => n141, Z => SUM(33));
   U236 : NAND2_X1 port map( A1 => carry_33_port, A2 => B(33), ZN => n142);
   U237 : NAND2_X1 port map( A1 => carry_33_port, A2 => A(33), ZN => n143);
   U238 : NAND2_X1 port map( A1 => B(33), A2 => A(33), ZN => n144);
   U239 : NAND3_X1 port map( A1 => n142, A2 => n143, A3 => n144, ZN => 
                           carry_34_port);
   U240 : XOR2_X1 port map( A => B(34), B => A(34), Z => n145);
   U241 : XOR2_X1 port map( A => carry_34_port, B => n145, Z => SUM(34));
   U242 : NAND2_X1 port map( A1 => carry_34_port, A2 => B(34), ZN => n146);
   U243 : NAND2_X1 port map( A1 => carry_34_port, A2 => A(34), ZN => n147);
   U244 : NAND2_X1 port map( A1 => B(34), A2 => A(34), ZN => n148);
   U245 : NAND3_X1 port map( A1 => n146, A2 => n147, A3 => n148, ZN => 
                           carry_35_port);
   U246 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n1);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHMUL_NBIT32_DW01_sub_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end BOOTHMUL_NBIT32_DW01_sub_0;

architecture SYN_rpl of BOOTHMUL_NBIT32_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111, n112, n114, n115, n116, n118, n119, n120, n123, 
      n124, DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, 
      DIFF_2_port, DIFF_1_port, n94, n95, n113, n117, n121, n122, n125, n126, 
      n127, n128, n129 : std_logic;

begin
   DIFF <= ( DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, 
      DIFF_2_port, DIFF_1_port, B(0) );
   
   U42 : XOR2_X1 port map( A => n96, B => B(30), Z => DIFF_30_port);
   U43 : XOR2_X1 port map( A => n98, B => B(27), Z => DIFF_27_port);
   U44 : XOR2_X1 port map( A => n101, B => B(26), Z => DIFF_26_port);
   U45 : XOR2_X1 port map( A => n100, B => B(25), Z => DIFF_25_port);
   U46 : XOR2_X1 port map( A => n102, B => B(23), Z => DIFF_23_port);
   U47 : XOR2_X1 port map( A => n105, B => B(22), Z => DIFF_22_port);
   U48 : XOR2_X1 port map( A => n104, B => B(21), Z => DIFF_21_port);
   U49 : XOR2_X1 port map( A => n106, B => B(19), Z => DIFF_19_port);
   U50 : XOR2_X1 port map( A => n109, B => B(18), Z => DIFF_18_port);
   U51 : XOR2_X1 port map( A => n108, B => B(17), Z => DIFF_17_port);
   U52 : XOR2_X1 port map( A => n110, B => B(15), Z => DIFF_15_port);
   U54 : XOR2_X1 port map( A => n112, B => B(13), Z => DIFF_13_port);
   U55 : XOR2_X1 port map( A => n114, B => B(11), Z => DIFF_11_port);
   U57 : XOR2_X1 port map( A => n116, B => B(9), Z => DIFF_9_port);
   U58 : XOR2_X1 port map( A => n118, B => B(7), Z => DIFF_7_port);
   U60 : XOR2_X1 port map( A => n120, B => B(5), Z => DIFF_5_port);
   U62 : XOR2_X1 port map( A => B(1), B => B(0), Z => DIFF_1_port);
   U1 : AND2_X1 port map( A1 => n117, A2 => n113, ZN => n94);
   U2 : NAND2_X1 port map( A1 => n95, A2 => n94, ZN => n120);
   U3 : OR3_X2 port map( A1 => B(5), A2 => B(6), A3 => n120, ZN => n118);
   U4 : INV_X1 port map( A => n125, ZN => n95);
   U5 : INV_X1 port map( A => B(4), ZN => n113);
   U6 : INV_X1 port map( A => B(3), ZN => n117);
   U7 : XNOR2_X1 port map( A => n121, B => B(6), ZN => DIFF_6_port);
   U8 : NOR2_X1 port map( A1 => n120, A2 => B(5), ZN => n121);
   U9 : NOR3_X1 port map( A1 => B(1), A2 => B(0), A3 => B(2), ZN => n122);
   U10 : XNOR2_X1 port map( A => n122, B => B(3), ZN => DIFF_3_port);
   U11 : OR3_X2 port map( A1 => B(1), A2 => B(2), A3 => B(0), ZN => n125);
   U12 : NAND2_X1 port map( A1 => n97, A2 => n129, ZN => n96);
   U13 : XOR2_X1 port map( A => n97, B => n129, Z => DIFF_29_port);
   U14 : XNOR2_X1 port map( A => n123, B => B(4), ZN => DIFF_4_port);
   U15 : NOR2_X1 port map( A1 => n125, A2 => B(3), ZN => n123);
   U16 : XNOR2_X1 port map( A => B(8), B => n119, ZN => DIFF_8_port);
   U17 : NOR2_X1 port map( A1 => B(7), A2 => n118, ZN => n119);
   U18 : XNOR2_X1 port map( A => n124, B => B(2), ZN => DIFF_2_port);
   U19 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n124);
   U20 : XNOR2_X1 port map( A => n126, B => B(31), ZN => DIFF_31_port);
   U21 : NOR2_X1 port map( A1 => n96, A2 => B(30), ZN => n126);
   U22 : NOR3_X1 port map( A1 => B(27), A2 => B(28), A3 => n98, ZN => n97);
   U23 : OR2_X1 port map( A1 => n100, A2 => B(25), ZN => n101);
   U24 : XNOR2_X1 port map( A => B(20), B => n107, ZN => DIFF_20_port);
   U25 : NOR2_X1 port map( A1 => B(19), A2 => n106, ZN => n107);
   U26 : XNOR2_X1 port map( A => B(24), B => n103, ZN => DIFF_24_port);
   U27 : NOR2_X1 port map( A1 => B(23), A2 => n102, ZN => n103);
   U28 : XNOR2_X1 port map( A => n127, B => B(10), ZN => DIFF_10_port);
   U29 : NOR2_X1 port map( A1 => n116, A2 => B(9), ZN => n127);
   U30 : XNOR2_X1 port map( A => n128, B => B(14), ZN => DIFF_14_port);
   U31 : NOR2_X1 port map( A1 => n112, A2 => B(13), ZN => n128);
   U32 : OR2_X1 port map( A1 => n108, A2 => B(17), ZN => n109);
   U33 : XNOR2_X1 port map( A => B(12), B => n115, ZN => DIFF_12_port);
   U34 : NOR2_X1 port map( A1 => B(11), A2 => n114, ZN => n115);
   U35 : XNOR2_X1 port map( A => B(16), B => n111, ZN => DIFF_16_port);
   U36 : NOR2_X1 port map( A1 => B(15), A2 => n110, ZN => n111);
   U37 : XNOR2_X1 port map( A => B(28), B => n99, ZN => DIFF_28_port);
   U38 : NOR2_X1 port map( A1 => B(27), A2 => n98, ZN => n99);
   U39 : OR3_X1 port map( A1 => B(25), A2 => B(26), A3 => n100, ZN => n98);
   U40 : OR3_X1 port map( A1 => B(17), A2 => B(18), A3 => n108, ZN => n106);
   U41 : OR3_X1 port map( A1 => B(21), A2 => B(22), A3 => n104, ZN => n102);
   U53 : OR3_X1 port map( A1 => B(13), A2 => B(14), A3 => n112, ZN => n110);
   U56 : OR3_X1 port map( A1 => B(10), A2 => B(9), A3 => n116, ZN => n114);
   U59 : OR3_X1 port map( A1 => B(19), A2 => B(20), A3 => n106, ZN => n104);
   U61 : OR3_X1 port map( A1 => B(15), A2 => B(16), A3 => n110, ZN => n108);
   U63 : OR3_X1 port map( A1 => B(23), A2 => B(24), A3 => n102, ZN => n100);
   U64 : OR3_X1 port map( A1 => B(11), A2 => B(12), A3 => n114, ZN => n112);
   U65 : OR3_X1 port map( A1 => B(7), A2 => B(8), A3 => n118, ZN => n116);
   U66 : OR2_X1 port map( A1 => n104, A2 => B(21), ZN => n105);
   U67 : INV_X1 port map( A => B(29), ZN => n129);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT64 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64;

architecture SYN_DIRECT of RCA_NBIT64 is

   component RCA_NBIT64_DW01_add_0
      port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (63 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1065 : std_logic;

begin
   
   Co <= '0';
   n2 <= '0';
   add_95 : RCA_NBIT64_DW01_add_0 port map( A(63) => A(63), A(62) => A(62), 
                           A(61) => A(61), A(60) => A(60), A(59) => A(59), 
                           A(58) => A(58), A(57) => A(57), A(56) => A(56), 
                           A(55) => A(55), A(54) => A(54), A(53) => A(53), 
                           A(52) => A(52), A(51) => A(51), A(50) => A(50), 
                           A(49) => A(49), A(48) => A(48), A(47) => A(47), 
                           A(46) => A(46), A(45) => A(45), A(44) => A(44), 
                           A(43) => A(43), A(42) => A(42), A(41) => A(41), 
                           A(40) => A(40), A(39) => A(39), A(38) => A(38), 
                           A(37) => A(37), A(36) => A(36), A(35) => A(35), 
                           A(34) => A(34), A(33) => A(33), A(32) => A(32), 
                           A(31) => A(31), A(30) => A(30), A(29) => A(29), 
                           A(28) => A(28), A(27) => A(27), A(26) => A(26), 
                           A(25) => A(25), A(24) => A(24), A(23) => A(23), 
                           A(22) => A(22), A(21) => A(21), A(20) => A(20), 
                           A(19) => A(19), A(18) => A(18), A(17) => A(17), 
                           A(16) => A(16), A(15) => A(15), A(14) => A(14), 
                           A(13) => A(13), A(12) => A(12), A(11) => A(11), 
                           A(10) => A(10), A(9) => A(9), A(8) => A(8), A(7) => 
                           A(7), A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3)
                           => A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(63) => B(63), B(62) => B(62), B(61) => B(61), 
                           B(60) => B(60), B(59) => B(59), B(58) => B(58), 
                           B(57) => B(57), B(56) => B(56), B(55) => B(55), 
                           B(54) => B(54), B(53) => B(53), B(52) => B(52), 
                           B(51) => B(51), B(50) => B(50), B(49) => B(49), 
                           B(48) => B(48), B(47) => B(47), B(46) => B(46), 
                           B(45) => B(45), B(44) => B(44), B(43) => B(43), 
                           B(42) => B(42), B(41) => B(41), B(40) => B(40), 
                           B(39) => B(39), B(38) => B(38), B(37) => B(37), 
                           B(36) => B(36), B(35) => B(35), B(34) => B(34), 
                           B(33) => B(33), B(32) => B(32), B(31) => B(31), 
                           B(30) => B(30), B(29) => B(29), B(28) => B(28), 
                           B(27) => B(27), B(26) => B(26), B(25) => B(25), 
                           B(24) => B(24), B(23) => B(23), B(22) => B(22), 
                           B(21) => B(21), B(20) => B(20), B(19) => B(19), 
                           B(18) => B(18), B(17) => B(17), B(16) => B(16), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => B(0), CI => n2, SUM(63) 
                           => S(63), SUM(62) => S(62), SUM(61) => S(61), 
                           SUM(60) => S(60), SUM(59) => S(59), SUM(58) => S(58)
                           , SUM(57) => S(57), SUM(56) => S(56), SUM(55) => 
                           S(55), SUM(54) => S(54), SUM(53) => S(53), SUM(52) 
                           => S(52), SUM(51) => S(51), SUM(50) => S(50), 
                           SUM(49) => S(49), SUM(48) => S(48), SUM(47) => S(47)
                           , SUM(46) => S(46), SUM(45) => S(45), SUM(44) => 
                           S(44), SUM(43) => S(43), SUM(42) => S(42), SUM(41) 
                           => S(41), SUM(40) => S(40), SUM(39) => S(39), 
                           SUM(38) => S(38), SUM(37) => S(37), SUM(36) => S(36)
                           , SUM(35) => S(35), SUM(34) => S(34), SUM(33) => 
                           S(33), SUM(32) => S(32), SUM(31) => S(31), SUM(30) 
                           => S(30), SUM(29) => S(29), SUM(28) => S(28), 
                           SUM(27) => S(27), SUM(26) => S(26), SUM(25) => S(25)
                           , SUM(24) => S(24), SUM(23) => S(23), SUM(22) => 
                           S(22), SUM(21) => S(21), SUM(20) => S(20), SUM(19) 
                           => S(19), SUM(18) => S(18), SUM(17) => S(17), 
                           SUM(16) => S(16), SUM(15) => S(15), SUM(14) => S(14)
                           , SUM(13) => S(13), SUM(12) => S(12), SUM(11) => 
                           S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) => 
                           S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5)
                           , SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1065);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT62 is

   port( A, B : in std_logic_vector (61 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (61 downto 0);  Co : out std_logic);

end RCA_NBIT62;

architecture SYN_DIRECT of RCA_NBIT62 is

   component RCA_NBIT62_DW01_add_0
      port( A, B : in std_logic_vector (61 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (61 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1066 : std_logic;

begin
   
   Co <= '0';
   n2 <= '0';
   add_95 : RCA_NBIT62_DW01_add_0 port map( A(61) => A(61), A(60) => A(60), 
                           A(59) => A(59), A(58) => A(58), A(57) => A(57), 
                           A(56) => A(56), A(55) => A(55), A(54) => A(54), 
                           A(53) => A(53), A(52) => A(52), A(51) => A(51), 
                           A(50) => A(50), A(49) => A(49), A(48) => A(48), 
                           A(47) => A(47), A(46) => A(46), A(45) => A(45), 
                           A(44) => A(44), A(43) => A(43), A(42) => A(42), 
                           A(41) => A(41), A(40) => A(40), A(39) => A(39), 
                           A(38) => A(38), A(37) => A(37), A(36) => A(36), 
                           A(35) => A(35), A(34) => A(34), A(33) => A(33), 
                           A(32) => A(32), A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(61) => B(61), B(60) => B(60), 
                           B(59) => B(59), B(58) => B(58), B(57) => B(57), 
                           B(56) => B(56), B(55) => B(55), B(54) => B(54), 
                           B(53) => B(53), B(52) => B(52), B(51) => B(51), 
                           B(50) => B(50), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => n2, SUM(61) => S(61), 
                           SUM(60) => S(60), SUM(59) => S(59), SUM(58) => S(58)
                           , SUM(57) => S(57), SUM(56) => S(56), SUM(55) => 
                           S(55), SUM(54) => S(54), SUM(53) => S(53), SUM(52) 
                           => S(52), SUM(51) => S(51), SUM(50) => S(50), 
                           SUM(49) => S(49), SUM(48) => S(48), SUM(47) => S(47)
                           , SUM(46) => S(46), SUM(45) => S(45), SUM(44) => 
                           S(44), SUM(43) => S(43), SUM(42) => S(42), SUM(41) 
                           => S(41), SUM(40) => S(40), SUM(39) => S(39), 
                           SUM(38) => S(38), SUM(37) => S(37), SUM(36) => S(36)
                           , SUM(35) => S(35), SUM(34) => S(34), SUM(33) => 
                           S(33), SUM(32) => S(32), SUM(31) => S(31), SUM(30) 
                           => S(30), SUM(29) => S(29), SUM(28) => S(28), 
                           SUM(27) => S(27), SUM(26) => S(26), SUM(25) => S(25)
                           , SUM(24) => S(24), SUM(23) => S(23), SUM(22) => 
                           S(22), SUM(21) => S(21), SUM(20) => S(20), SUM(19) 
                           => S(19), SUM(18) => S(18), SUM(17) => S(17), 
                           SUM(16) => S(16), SUM(15) => S(15), SUM(14) => S(14)
                           , SUM(13) => S(13), SUM(12) => S(12), SUM(11) => 
                           S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) => 
                           S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5)
                           , SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1066);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT60 is

   port( A, B : in std_logic_vector (59 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (59 downto 0);  Co : out std_logic);

end RCA_NBIT60;

architecture SYN_DIRECT of RCA_NBIT60 is

   component RCA_NBIT60_DW01_add_0
      port( A, B : in std_logic_vector (59 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (59 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1067 : std_logic;

begin
   
   Co <= '0';
   n2 <= '0';
   add_95 : RCA_NBIT60_DW01_add_0 port map( A(59) => A(59), A(58) => A(58), 
                           A(57) => A(57), A(56) => A(56), A(55) => A(55), 
                           A(54) => A(54), A(53) => A(53), A(52) => A(52), 
                           A(51) => A(51), A(50) => A(50), A(49) => A(49), 
                           A(48) => A(48), A(47) => A(47), A(46) => A(46), 
                           A(45) => A(45), A(44) => A(44), A(43) => A(43), 
                           A(42) => A(42), A(41) => A(41), A(40) => A(40), 
                           A(39) => A(39), A(38) => A(38), A(37) => A(37), 
                           A(36) => A(36), A(35) => A(35), A(34) => A(34), 
                           A(33) => A(33), A(32) => A(32), A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(59) => B(59), 
                           B(58) => B(58), B(57) => B(57), B(56) => B(56), 
                           B(55) => B(55), B(54) => B(54), B(53) => B(53), 
                           B(52) => B(52), B(51) => B(51), B(50) => B(50), 
                           B(49) => B(49), B(48) => B(48), B(47) => B(47), 
                           B(46) => B(46), B(45) => B(45), B(44) => B(44), 
                           B(43) => B(43), B(42) => B(42), B(41) => B(41), 
                           B(40) => B(40), B(39) => B(39), B(38) => B(38), 
                           B(37) => B(37), B(36) => B(36), B(35) => B(35), 
                           B(34) => B(34), B(33) => B(33), B(32) => B(32), 
                           B(31) => B(31), B(30) => B(30), B(29) => B(29), 
                           B(28) => B(28), B(27) => B(27), B(26) => B(26), 
                           B(25) => B(25), B(24) => B(24), B(23) => B(23), 
                           B(22) => B(22), B(21) => B(21), B(20) => B(20), 
                           B(19) => B(19), B(18) => B(18), B(17) => B(17), 
                           B(16) => B(16), B(15) => B(15), B(14) => B(14), 
                           B(13) => B(13), B(12) => B(12), B(11) => B(11), 
                           B(10) => B(10), B(9) => B(9), B(8) => B(8), B(7) => 
                           B(7), B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3)
                           => B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), 
                           CI => n2, SUM(59) => S(59), SUM(58) => S(58), 
                           SUM(57) => S(57), SUM(56) => S(56), SUM(55) => S(55)
                           , SUM(54) => S(54), SUM(53) => S(53), SUM(52) => 
                           S(52), SUM(51) => S(51), SUM(50) => S(50), SUM(49) 
                           => S(49), SUM(48) => S(48), SUM(47) => S(47), 
                           SUM(46) => S(46), SUM(45) => S(45), SUM(44) => S(44)
                           , SUM(43) => S(43), SUM(42) => S(42), SUM(41) => 
                           S(41), SUM(40) => S(40), SUM(39) => S(39), SUM(38) 
                           => S(38), SUM(37) => S(37), SUM(36) => S(36), 
                           SUM(35) => S(35), SUM(34) => S(34), SUM(33) => S(33)
                           , SUM(32) => S(32), SUM(31) => S(31), SUM(30) => 
                           S(30), SUM(29) => S(29), SUM(28) => S(28), SUM(27) 
                           => S(27), SUM(26) => S(26), SUM(25) => S(25), 
                           SUM(24) => S(24), SUM(23) => S(23), SUM(22) => S(22)
                           , SUM(21) => S(21), SUM(20) => S(20), SUM(19) => 
                           S(19), SUM(18) => S(18), SUM(17) => S(17), SUM(16) 
                           => S(16), SUM(15) => S(15), SUM(14) => S(14), 
                           SUM(13) => S(13), SUM(12) => S(12), SUM(11) => S(11)
                           , SUM(10) => S(10), SUM(9) => S(9), SUM(8) => S(8), 
                           SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5), 
                           SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1067);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT58 is

   port( A, B : in std_logic_vector (57 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (57 downto 0);  Co : out std_logic);

end RCA_NBIT58;

architecture SYN_DIRECT of RCA_NBIT58 is

   component RCA_NBIT58_DW01_add_0
      port( A, B : in std_logic_vector (57 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (57 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1068 : std_logic;

begin
   
   Co <= '0';
   n2 <= '0';
   add_95 : RCA_NBIT58_DW01_add_0 port map( A(57) => A(57), A(56) => A(56), 
                           A(55) => A(55), A(54) => A(54), A(53) => A(53), 
                           A(52) => A(52), A(51) => A(51), A(50) => A(50), 
                           A(49) => A(49), A(48) => A(48), A(47) => A(47), 
                           A(46) => A(46), A(45) => A(45), A(44) => A(44), 
                           A(43) => A(43), A(42) => A(42), A(41) => A(41), 
                           A(40) => A(40), A(39) => A(39), A(38) => A(38), 
                           A(37) => A(37), A(36) => A(36), A(35) => A(35), 
                           A(34) => A(34), A(33) => A(33), A(32) => A(32), 
                           A(31) => A(31), A(30) => A(30), A(29) => A(29), 
                           A(28) => A(28), A(27) => A(27), A(26) => A(26), 
                           A(25) => A(25), A(24) => A(24), A(23) => A(23), 
                           A(22) => A(22), A(21) => A(21), A(20) => A(20), 
                           A(19) => A(19), A(18) => A(18), A(17) => A(17), 
                           A(16) => A(16), A(15) => A(15), A(14) => A(14), 
                           A(13) => A(13), A(12) => A(12), A(11) => A(11), 
                           A(10) => A(10), A(9) => A(9), A(8) => A(8), A(7) => 
                           A(7), A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3)
                           => A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(57) => B(57), B(56) => B(56), B(55) => B(55), 
                           B(54) => B(54), B(53) => B(53), B(52) => B(52), 
                           B(51) => B(51), B(50) => B(50), B(49) => B(49), 
                           B(48) => B(48), B(47) => B(47), B(46) => B(46), 
                           B(45) => B(45), B(44) => B(44), B(43) => B(43), 
                           B(42) => B(42), B(41) => B(41), B(40) => B(40), 
                           B(39) => B(39), B(38) => B(38), B(37) => B(37), 
                           B(36) => B(36), B(35) => B(35), B(34) => B(34), 
                           B(33) => B(33), B(32) => B(32), B(31) => B(31), 
                           B(30) => B(30), B(29) => B(29), B(28) => B(28), 
                           B(27) => B(27), B(26) => B(26), B(25) => B(25), 
                           B(24) => B(24), B(23) => B(23), B(22) => B(22), 
                           B(21) => B(21), B(20) => B(20), B(19) => B(19), 
                           B(18) => B(18), B(17) => B(17), B(16) => B(16), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => B(0), CI => n2, SUM(57) 
                           => S(57), SUM(56) => S(56), SUM(55) => S(55), 
                           SUM(54) => S(54), SUM(53) => S(53), SUM(52) => S(52)
                           , SUM(51) => S(51), SUM(50) => S(50), SUM(49) => 
                           S(49), SUM(48) => S(48), SUM(47) => S(47), SUM(46) 
                           => S(46), SUM(45) => S(45), SUM(44) => S(44), 
                           SUM(43) => S(43), SUM(42) => S(42), SUM(41) => S(41)
                           , SUM(40) => S(40), SUM(39) => S(39), SUM(38) => 
                           S(38), SUM(37) => S(37), SUM(36) => S(36), SUM(35) 
                           => S(35), SUM(34) => S(34), SUM(33) => S(33), 
                           SUM(32) => S(32), SUM(31) => S(31), SUM(30) => S(30)
                           , SUM(29) => S(29), SUM(28) => S(28), SUM(27) => 
                           S(27), SUM(26) => S(26), SUM(25) => S(25), SUM(24) 
                           => S(24), SUM(23) => S(23), SUM(22) => S(22), 
                           SUM(21) => S(21), SUM(20) => S(20), SUM(19) => S(19)
                           , SUM(18) => S(18), SUM(17) => S(17), SUM(16) => 
                           S(16), SUM(15) => S(15), SUM(14) => S(14), SUM(13) 
                           => S(13), SUM(12) => S(12), SUM(11) => S(11), 
                           SUM(10) => S(10), SUM(9) => S(9), SUM(8) => S(8), 
                           SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5), 
                           SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1068);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT56 is

   port( A, B : in std_logic_vector (55 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (55 downto 0);  Co : out std_logic);

end RCA_NBIT56;

architecture SYN_DIRECT of RCA_NBIT56 is

   component RCA_NBIT56_DW01_add_0
      port( A, B : in std_logic_vector (55 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (55 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1069 : std_logic;

begin
   
   Co <= '0';
   n2 <= '0';
   add_95 : RCA_NBIT56_DW01_add_0 port map( A(55) => A(55), A(54) => A(54), 
                           A(53) => A(53), A(52) => A(52), A(51) => A(51), 
                           A(50) => A(50), A(49) => A(49), A(48) => A(48), 
                           A(47) => A(47), A(46) => A(46), A(45) => A(45), 
                           A(44) => A(44), A(43) => A(43), A(42) => A(42), 
                           A(41) => A(41), A(40) => A(40), A(39) => A(39), 
                           A(38) => A(38), A(37) => A(37), A(36) => A(36), 
                           A(35) => A(35), A(34) => A(34), A(33) => A(33), 
                           A(32) => A(32), A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(55) => B(55), B(54) => B(54), 
                           B(53) => B(53), B(52) => B(52), B(51) => B(51), 
                           B(50) => B(50), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => n2, SUM(55) => S(55), 
                           SUM(54) => S(54), SUM(53) => S(53), SUM(52) => S(52)
                           , SUM(51) => S(51), SUM(50) => S(50), SUM(49) => 
                           S(49), SUM(48) => S(48), SUM(47) => S(47), SUM(46) 
                           => S(46), SUM(45) => S(45), SUM(44) => S(44), 
                           SUM(43) => S(43), SUM(42) => S(42), SUM(41) => S(41)
                           , SUM(40) => S(40), SUM(39) => S(39), SUM(38) => 
                           S(38), SUM(37) => S(37), SUM(36) => S(36), SUM(35) 
                           => S(35), SUM(34) => S(34), SUM(33) => S(33), 
                           SUM(32) => S(32), SUM(31) => S(31), SUM(30) => S(30)
                           , SUM(29) => S(29), SUM(28) => S(28), SUM(27) => 
                           S(27), SUM(26) => S(26), SUM(25) => S(25), SUM(24) 
                           => S(24), SUM(23) => S(23), SUM(22) => S(22), 
                           SUM(21) => S(21), SUM(20) => S(20), SUM(19) => S(19)
                           , SUM(18) => S(18), SUM(17) => S(17), SUM(16) => 
                           S(16), SUM(15) => S(15), SUM(14) => S(14), SUM(13) 
                           => S(13), SUM(12) => S(12), SUM(11) => S(11), 
                           SUM(10) => S(10), SUM(9) => S(9), SUM(8) => S(8), 
                           SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5), 
                           SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1069);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT54 is

   port( A, B : in std_logic_vector (53 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (53 downto 0);  Co : out std_logic);

end RCA_NBIT54;

architecture SYN_DIRECT of RCA_NBIT54 is

   component RCA_NBIT54_DW01_add_0
      port( A, B : in std_logic_vector (53 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (53 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1070 : std_logic;

begin
   
   Co <= '0';
   n2 <= '0';
   add_95 : RCA_NBIT54_DW01_add_0 port map( A(53) => A(53), A(52) => A(52), 
                           A(51) => A(51), A(50) => A(50), A(49) => A(49), 
                           A(48) => A(48), A(47) => A(47), A(46) => A(46), 
                           A(45) => A(45), A(44) => A(44), A(43) => A(43), 
                           A(42) => A(42), A(41) => A(41), A(40) => A(40), 
                           A(39) => A(39), A(38) => A(38), A(37) => A(37), 
                           A(36) => A(36), A(35) => A(35), A(34) => A(34), 
                           A(33) => A(33), A(32) => A(32), A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(53) => B(53), 
                           B(52) => B(52), B(51) => B(51), B(50) => B(50), 
                           B(49) => B(49), B(48) => B(48), B(47) => B(47), 
                           B(46) => B(46), B(45) => B(45), B(44) => B(44), 
                           B(43) => B(43), B(42) => B(42), B(41) => B(41), 
                           B(40) => B(40), B(39) => B(39), B(38) => B(38), 
                           B(37) => B(37), B(36) => B(36), B(35) => B(35), 
                           B(34) => B(34), B(33) => B(33), B(32) => B(32), 
                           B(31) => B(31), B(30) => B(30), B(29) => B(29), 
                           B(28) => B(28), B(27) => B(27), B(26) => B(26), 
                           B(25) => B(25), B(24) => B(24), B(23) => B(23), 
                           B(22) => B(22), B(21) => B(21), B(20) => B(20), 
                           B(19) => B(19), B(18) => B(18), B(17) => B(17), 
                           B(16) => B(16), B(15) => B(15), B(14) => B(14), 
                           B(13) => B(13), B(12) => B(12), B(11) => B(11), 
                           B(10) => B(10), B(9) => B(9), B(8) => B(8), B(7) => 
                           B(7), B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3)
                           => B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), 
                           CI => n2, SUM(53) => S(53), SUM(52) => S(52), 
                           SUM(51) => S(51), SUM(50) => S(50), SUM(49) => S(49)
                           , SUM(48) => S(48), SUM(47) => S(47), SUM(46) => 
                           S(46), SUM(45) => S(45), SUM(44) => S(44), SUM(43) 
                           => S(43), SUM(42) => S(42), SUM(41) => S(41), 
                           SUM(40) => S(40), SUM(39) => S(39), SUM(38) => S(38)
                           , SUM(37) => S(37), SUM(36) => S(36), SUM(35) => 
                           S(35), SUM(34) => S(34), SUM(33) => S(33), SUM(32) 
                           => S(32), SUM(31) => S(31), SUM(30) => S(30), 
                           SUM(29) => S(29), SUM(28) => S(28), SUM(27) => S(27)
                           , SUM(26) => S(26), SUM(25) => S(25), SUM(24) => 
                           S(24), SUM(23) => S(23), SUM(22) => S(22), SUM(21) 
                           => S(21), SUM(20) => S(20), SUM(19) => S(19), 
                           SUM(18) => S(18), SUM(17) => S(17), SUM(16) => S(16)
                           , SUM(15) => S(15), SUM(14) => S(14), SUM(13) => 
                           S(13), SUM(12) => S(12), SUM(11) => S(11), SUM(10) 
                           => S(10), SUM(9) => S(9), SUM(8) => S(8), SUM(7) => 
                           S(7), SUM(6) => S(6), SUM(5) => S(5), SUM(4) => S(4)
                           , SUM(3) => S(3), SUM(2) => S(2), SUM(1) => S(1), 
                           SUM(0) => S(0), CO => n_1070);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT52 is

   port( A, B : in std_logic_vector (51 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (51 downto 0);  Co : out std_logic);

end RCA_NBIT52;

architecture SYN_DIRECT of RCA_NBIT52 is

   component RCA_NBIT52_DW01_add_0
      port( A, B : in std_logic_vector (51 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (51 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1071 : std_logic;

begin
   
   Co <= '0';
   n2 <= '0';
   add_95 : RCA_NBIT52_DW01_add_0 port map( A(51) => A(51), A(50) => A(50), 
                           A(49) => A(49), A(48) => A(48), A(47) => A(47), 
                           A(46) => A(46), A(45) => A(45), A(44) => A(44), 
                           A(43) => A(43), A(42) => A(42), A(41) => A(41), 
                           A(40) => A(40), A(39) => A(39), A(38) => A(38), 
                           A(37) => A(37), A(36) => A(36), A(35) => A(35), 
                           A(34) => A(34), A(33) => A(33), A(32) => A(32), 
                           A(31) => A(31), A(30) => A(30), A(29) => A(29), 
                           A(28) => A(28), A(27) => A(27), A(26) => A(26), 
                           A(25) => A(25), A(24) => A(24), A(23) => A(23), 
                           A(22) => A(22), A(21) => A(21), A(20) => A(20), 
                           A(19) => A(19), A(18) => A(18), A(17) => A(17), 
                           A(16) => A(16), A(15) => A(15), A(14) => A(14), 
                           A(13) => A(13), A(12) => A(12), A(11) => A(11), 
                           A(10) => A(10), A(9) => A(9), A(8) => A(8), A(7) => 
                           A(7), A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3)
                           => A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(51) => B(51), B(50) => B(50), B(49) => B(49), 
                           B(48) => B(48), B(47) => B(47), B(46) => B(46), 
                           B(45) => B(45), B(44) => B(44), B(43) => B(43), 
                           B(42) => B(42), B(41) => B(41), B(40) => B(40), 
                           B(39) => B(39), B(38) => B(38), B(37) => B(37), 
                           B(36) => B(36), B(35) => B(35), B(34) => B(34), 
                           B(33) => B(33), B(32) => B(32), B(31) => B(31), 
                           B(30) => B(30), B(29) => B(29), B(28) => B(28), 
                           B(27) => B(27), B(26) => B(26), B(25) => B(25), 
                           B(24) => B(24), B(23) => B(23), B(22) => B(22), 
                           B(21) => B(21), B(20) => B(20), B(19) => B(19), 
                           B(18) => B(18), B(17) => B(17), B(16) => B(16), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => B(0), CI => n2, SUM(51) 
                           => S(51), SUM(50) => S(50), SUM(49) => S(49), 
                           SUM(48) => S(48), SUM(47) => S(47), SUM(46) => S(46)
                           , SUM(45) => S(45), SUM(44) => S(44), SUM(43) => 
                           S(43), SUM(42) => S(42), SUM(41) => S(41), SUM(40) 
                           => S(40), SUM(39) => S(39), SUM(38) => S(38), 
                           SUM(37) => S(37), SUM(36) => S(36), SUM(35) => S(35)
                           , SUM(34) => S(34), SUM(33) => S(33), SUM(32) => 
                           S(32), SUM(31) => S(31), SUM(30) => S(30), SUM(29) 
                           => S(29), SUM(28) => S(28), SUM(27) => S(27), 
                           SUM(26) => S(26), SUM(25) => S(25), SUM(24) => S(24)
                           , SUM(23) => S(23), SUM(22) => S(22), SUM(21) => 
                           S(21), SUM(20) => S(20), SUM(19) => S(19), SUM(18) 
                           => S(18), SUM(17) => S(17), SUM(16) => S(16), 
                           SUM(15) => S(15), SUM(14) => S(14), SUM(13) => S(13)
                           , SUM(12) => S(12), SUM(11) => S(11), SUM(10) => 
                           S(10), SUM(9) => S(9), SUM(8) => S(8), SUM(7) => 
                           S(7), SUM(6) => S(6), SUM(5) => S(5), SUM(4) => S(4)
                           , SUM(3) => S(3), SUM(2) => S(2), SUM(1) => S(1), 
                           SUM(0) => S(0), CO => n_1071);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT50 is

   port( A, B : in std_logic_vector (49 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (49 downto 0);  Co : out std_logic);

end RCA_NBIT50;

architecture SYN_DIRECT of RCA_NBIT50 is

   component RCA_NBIT50_DW01_add_0
      port( A, B : in std_logic_vector (49 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (49 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1072 : std_logic;

begin
   
   Co <= '0';
   n2 <= '0';
   add_95 : RCA_NBIT50_DW01_add_0 port map( A(49) => A(49), A(48) => A(48), 
                           A(47) => A(47), A(46) => A(46), A(45) => A(45), 
                           A(44) => A(44), A(43) => A(43), A(42) => A(42), 
                           A(41) => A(41), A(40) => A(40), A(39) => A(39), 
                           A(38) => A(38), A(37) => A(37), A(36) => A(36), 
                           A(35) => A(35), A(34) => A(34), A(33) => A(33), 
                           A(32) => A(32), A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => n2, SUM(49) => S(49), 
                           SUM(48) => S(48), SUM(47) => S(47), SUM(46) => S(46)
                           , SUM(45) => S(45), SUM(44) => S(44), SUM(43) => 
                           S(43), SUM(42) => S(42), SUM(41) => S(41), SUM(40) 
                           => S(40), SUM(39) => S(39), SUM(38) => S(38), 
                           SUM(37) => S(37), SUM(36) => S(36), SUM(35) => S(35)
                           , SUM(34) => S(34), SUM(33) => S(33), SUM(32) => 
                           S(32), SUM(31) => S(31), SUM(30) => S(30), SUM(29) 
                           => S(29), SUM(28) => S(28), SUM(27) => S(27), 
                           SUM(26) => S(26), SUM(25) => S(25), SUM(24) => S(24)
                           , SUM(23) => S(23), SUM(22) => S(22), SUM(21) => 
                           S(21), SUM(20) => S(20), SUM(19) => S(19), SUM(18) 
                           => S(18), SUM(17) => S(17), SUM(16) => S(16), 
                           SUM(15) => S(15), SUM(14) => S(14), SUM(13) => S(13)
                           , SUM(12) => S(12), SUM(11) => S(11), SUM(10) => 
                           S(10), SUM(9) => S(9), SUM(8) => S(8), SUM(7) => 
                           S(7), SUM(6) => S(6), SUM(5) => S(5), SUM(4) => S(4)
                           , SUM(3) => S(3), SUM(2) => S(2), SUM(1) => S(1), 
                           SUM(0) => S(0), CO => n_1072);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT48 is

   port( A, B : in std_logic_vector (47 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (47 downto 0);  Co : out std_logic);

end RCA_NBIT48;

architecture SYN_DIRECT of RCA_NBIT48 is

   component RCA_NBIT48_DW01_add_0
      port( A, B : in std_logic_vector (47 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (47 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1073 : std_logic;

begin
   
   Co <= '0';
   n2 <= '0';
   add_95 : RCA_NBIT48_DW01_add_0 port map( A(47) => A(47), A(46) => A(46), 
                           A(45) => A(45), A(44) => A(44), A(43) => A(43), 
                           A(42) => A(42), A(41) => A(41), A(40) => A(40), 
                           A(39) => A(39), A(38) => A(38), A(37) => A(37), 
                           A(36) => A(36), A(35) => A(35), A(34) => A(34), 
                           A(33) => A(33), A(32) => A(32), A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(47) => B(47), 
                           B(46) => B(46), B(45) => B(45), B(44) => B(44), 
                           B(43) => B(43), B(42) => B(42), B(41) => B(41), 
                           B(40) => B(40), B(39) => B(39), B(38) => B(38), 
                           B(37) => B(37), B(36) => B(36), B(35) => B(35), 
                           B(34) => B(34), B(33) => B(33), B(32) => B(32), 
                           B(31) => B(31), B(30) => B(30), B(29) => B(29), 
                           B(28) => B(28), B(27) => B(27), B(26) => B(26), 
                           B(25) => B(25), B(24) => B(24), B(23) => B(23), 
                           B(22) => B(22), B(21) => B(21), B(20) => B(20), 
                           B(19) => B(19), B(18) => B(18), B(17) => B(17), 
                           B(16) => B(16), B(15) => B(15), B(14) => B(14), 
                           B(13) => B(13), B(12) => B(12), B(11) => B(11), 
                           B(10) => B(10), B(9) => B(9), B(8) => B(8), B(7) => 
                           B(7), B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3)
                           => B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), 
                           CI => n2, SUM(47) => S(47), SUM(46) => S(46), 
                           SUM(45) => S(45), SUM(44) => S(44), SUM(43) => S(43)
                           , SUM(42) => S(42), SUM(41) => S(41), SUM(40) => 
                           S(40), SUM(39) => S(39), SUM(38) => S(38), SUM(37) 
                           => S(37), SUM(36) => S(36), SUM(35) => S(35), 
                           SUM(34) => S(34), SUM(33) => S(33), SUM(32) => S(32)
                           , SUM(31) => S(31), SUM(30) => S(30), SUM(29) => 
                           S(29), SUM(28) => S(28), SUM(27) => S(27), SUM(26) 
                           => S(26), SUM(25) => S(25), SUM(24) => S(24), 
                           SUM(23) => S(23), SUM(22) => S(22), SUM(21) => S(21)
                           , SUM(20) => S(20), SUM(19) => S(19), SUM(18) => 
                           S(18), SUM(17) => S(17), SUM(16) => S(16), SUM(15) 
                           => S(15), SUM(14) => S(14), SUM(13) => S(13), 
                           SUM(12) => S(12), SUM(11) => S(11), SUM(10) => S(10)
                           , SUM(9) => S(9), SUM(8) => S(8), SUM(7) => S(7), 
                           SUM(6) => S(6), SUM(5) => S(5), SUM(4) => S(4), 
                           SUM(3) => S(3), SUM(2) => S(2), SUM(1) => S(1), 
                           SUM(0) => S(0), CO => n_1073);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT46 is

   port( A, B : in std_logic_vector (45 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (45 downto 0);  Co : out std_logic);

end RCA_NBIT46;

architecture SYN_DIRECT of RCA_NBIT46 is

   component RCA_NBIT46_DW01_add_0
      port( A, B : in std_logic_vector (45 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (45 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1074 : std_logic;

begin
   
   Co <= '0';
   n2 <= '0';
   add_95 : RCA_NBIT46_DW01_add_0 port map( A(45) => A(45), A(44) => A(44), 
                           A(43) => A(43), A(42) => A(42), A(41) => A(41), 
                           A(40) => A(40), A(39) => A(39), A(38) => A(38), 
                           A(37) => A(37), A(36) => A(36), A(35) => A(35), 
                           A(34) => A(34), A(33) => A(33), A(32) => A(32), 
                           A(31) => A(31), A(30) => A(30), A(29) => A(29), 
                           A(28) => A(28), A(27) => A(27), A(26) => A(26), 
                           A(25) => A(25), A(24) => A(24), A(23) => A(23), 
                           A(22) => A(22), A(21) => A(21), A(20) => A(20), 
                           A(19) => A(19), A(18) => A(18), A(17) => A(17), 
                           A(16) => A(16), A(15) => A(15), A(14) => A(14), 
                           A(13) => A(13), A(12) => A(12), A(11) => A(11), 
                           A(10) => A(10), A(9) => A(9), A(8) => A(8), A(7) => 
                           A(7), A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3)
                           => A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(45) => B(45), B(44) => B(44), B(43) => B(43), 
                           B(42) => B(42), B(41) => B(41), B(40) => B(40), 
                           B(39) => B(39), B(38) => B(38), B(37) => B(37), 
                           B(36) => B(36), B(35) => B(35), B(34) => B(34), 
                           B(33) => B(33), B(32) => B(32), B(31) => B(31), 
                           B(30) => B(30), B(29) => B(29), B(28) => B(28), 
                           B(27) => B(27), B(26) => B(26), B(25) => B(25), 
                           B(24) => B(24), B(23) => B(23), B(22) => B(22), 
                           B(21) => B(21), B(20) => B(20), B(19) => B(19), 
                           B(18) => B(18), B(17) => B(17), B(16) => B(16), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => B(0), CI => n2, SUM(45) 
                           => S(45), SUM(44) => S(44), SUM(43) => S(43), 
                           SUM(42) => S(42), SUM(41) => S(41), SUM(40) => S(40)
                           , SUM(39) => S(39), SUM(38) => S(38), SUM(37) => 
                           S(37), SUM(36) => S(36), SUM(35) => S(35), SUM(34) 
                           => S(34), SUM(33) => S(33), SUM(32) => S(32), 
                           SUM(31) => S(31), SUM(30) => S(30), SUM(29) => S(29)
                           , SUM(28) => S(28), SUM(27) => S(27), SUM(26) => 
                           S(26), SUM(25) => S(25), SUM(24) => S(24), SUM(23) 
                           => S(23), SUM(22) => S(22), SUM(21) => S(21), 
                           SUM(20) => S(20), SUM(19) => S(19), SUM(18) => S(18)
                           , SUM(17) => S(17), SUM(16) => S(16), SUM(15) => 
                           S(15), SUM(14) => S(14), SUM(13) => S(13), SUM(12) 
                           => S(12), SUM(11) => S(11), SUM(10) => S(10), SUM(9)
                           => S(9), SUM(8) => S(8), SUM(7) => S(7), SUM(6) => 
                           S(6), SUM(5) => S(5), SUM(4) => S(4), SUM(3) => S(3)
                           , SUM(2) => S(2), SUM(1) => S(1), SUM(0) => S(0), CO
                           => n_1074);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT44 is

   port( A, B : in std_logic_vector (43 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (43 downto 0);  Co : out std_logic);

end RCA_NBIT44;

architecture SYN_DIRECT of RCA_NBIT44 is

   component RCA_NBIT44_DW01_add_0
      port( A, B : in std_logic_vector (43 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (43 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1075 : std_logic;

begin
   
   Co <= '0';
   n2 <= '0';
   add_95 : RCA_NBIT44_DW01_add_0 port map( A(43) => A(43), A(42) => A(42), 
                           A(41) => A(41), A(40) => A(40), A(39) => A(39), 
                           A(38) => A(38), A(37) => A(37), A(36) => A(36), 
                           A(35) => A(35), A(34) => A(34), A(33) => A(33), 
                           A(32) => A(32), A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => n2, SUM(43) => S(43), 
                           SUM(42) => S(42), SUM(41) => S(41), SUM(40) => S(40)
                           , SUM(39) => S(39), SUM(38) => S(38), SUM(37) => 
                           S(37), SUM(36) => S(36), SUM(35) => S(35), SUM(34) 
                           => S(34), SUM(33) => S(33), SUM(32) => S(32), 
                           SUM(31) => S(31), SUM(30) => S(30), SUM(29) => S(29)
                           , SUM(28) => S(28), SUM(27) => S(27), SUM(26) => 
                           S(26), SUM(25) => S(25), SUM(24) => S(24), SUM(23) 
                           => S(23), SUM(22) => S(22), SUM(21) => S(21), 
                           SUM(20) => S(20), SUM(19) => S(19), SUM(18) => S(18)
                           , SUM(17) => S(17), SUM(16) => S(16), SUM(15) => 
                           S(15), SUM(14) => S(14), SUM(13) => S(13), SUM(12) 
                           => S(12), SUM(11) => S(11), SUM(10) => S(10), SUM(9)
                           => S(9), SUM(8) => S(8), SUM(7) => S(7), SUM(6) => 
                           S(6), SUM(5) => S(5), SUM(4) => S(4), SUM(3) => S(3)
                           , SUM(2) => S(2), SUM(1) => S(1), SUM(0) => S(0), CO
                           => n_1075);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT42 is

   port( A, B : in std_logic_vector (41 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (41 downto 0);  Co : out std_logic);

end RCA_NBIT42;

architecture SYN_DIRECT of RCA_NBIT42 is

   component RCA_NBIT42_DW01_add_0
      port( A, B : in std_logic_vector (41 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (41 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1076 : std_logic;

begin
   
   Co <= '0';
   n2 <= '0';
   add_95 : RCA_NBIT42_DW01_add_0 port map( A(41) => A(41), A(40) => A(40), 
                           A(39) => A(39), A(38) => A(38), A(37) => A(37), 
                           A(36) => A(36), A(35) => A(35), A(34) => A(34), 
                           A(33) => A(33), A(32) => A(32), A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(41) => B(41), 
                           B(40) => B(40), B(39) => B(39), B(38) => B(38), 
                           B(37) => B(37), B(36) => B(36), B(35) => B(35), 
                           B(34) => B(34), B(33) => B(33), B(32) => B(32), 
                           B(31) => B(31), B(30) => B(30), B(29) => B(29), 
                           B(28) => B(28), B(27) => B(27), B(26) => B(26), 
                           B(25) => B(25), B(24) => B(24), B(23) => B(23), 
                           B(22) => B(22), B(21) => B(21), B(20) => B(20), 
                           B(19) => B(19), B(18) => B(18), B(17) => B(17), 
                           B(16) => B(16), B(15) => B(15), B(14) => B(14), 
                           B(13) => B(13), B(12) => B(12), B(11) => B(11), 
                           B(10) => B(10), B(9) => B(9), B(8) => B(8), B(7) => 
                           B(7), B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3)
                           => B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), 
                           CI => n2, SUM(41) => S(41), SUM(40) => S(40), 
                           SUM(39) => S(39), SUM(38) => S(38), SUM(37) => S(37)
                           , SUM(36) => S(36), SUM(35) => S(35), SUM(34) => 
                           S(34), SUM(33) => S(33), SUM(32) => S(32), SUM(31) 
                           => S(31), SUM(30) => S(30), SUM(29) => S(29), 
                           SUM(28) => S(28), SUM(27) => S(27), SUM(26) => S(26)
                           , SUM(25) => S(25), SUM(24) => S(24), SUM(23) => 
                           S(23), SUM(22) => S(22), SUM(21) => S(21), SUM(20) 
                           => S(20), SUM(19) => S(19), SUM(18) => S(18), 
                           SUM(17) => S(17), SUM(16) => S(16), SUM(15) => S(15)
                           , SUM(14) => S(14), SUM(13) => S(13), SUM(12) => 
                           S(12), SUM(11) => S(11), SUM(10) => S(10), SUM(9) =>
                           S(9), SUM(8) => S(8), SUM(7) => S(7), SUM(6) => S(6)
                           , SUM(5) => S(5), SUM(4) => S(4), SUM(3) => S(3), 
                           SUM(2) => S(2), SUM(1) => S(1), SUM(0) => S(0), CO 
                           => n_1076);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT40 is

   port( A, B : in std_logic_vector (39 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (39 downto 0);  Co : out std_logic);

end RCA_NBIT40;

architecture SYN_DIRECT of RCA_NBIT40 is

   component RCA_NBIT40_DW01_add_0
      port( A, B : in std_logic_vector (39 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (39 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1077 : std_logic;

begin
   
   Co <= '0';
   n2 <= '0';
   add_95 : RCA_NBIT40_DW01_add_0 port map( A(39) => A(39), A(38) => A(38), 
                           A(37) => A(37), A(36) => A(36), A(35) => A(35), 
                           A(34) => A(34), A(33) => A(33), A(32) => A(32), 
                           A(31) => A(31), A(30) => A(30), A(29) => A(29), 
                           A(28) => A(28), A(27) => A(27), A(26) => A(26), 
                           A(25) => A(25), A(24) => A(24), A(23) => A(23), 
                           A(22) => A(22), A(21) => A(21), A(20) => A(20), 
                           A(19) => A(19), A(18) => A(18), A(17) => A(17), 
                           A(16) => A(16), A(15) => A(15), A(14) => A(14), 
                           A(13) => A(13), A(12) => A(12), A(11) => A(11), 
                           A(10) => A(10), A(9) => A(9), A(8) => A(8), A(7) => 
                           A(7), A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3)
                           => A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(39) => B(39), B(38) => B(38), B(37) => B(37), 
                           B(36) => B(36), B(35) => B(35), B(34) => B(34), 
                           B(33) => B(33), B(32) => B(32), B(31) => B(31), 
                           B(30) => B(30), B(29) => B(29), B(28) => B(28), 
                           B(27) => B(27), B(26) => B(26), B(25) => B(25), 
                           B(24) => B(24), B(23) => B(23), B(22) => B(22), 
                           B(21) => B(21), B(20) => B(20), B(19) => B(19), 
                           B(18) => B(18), B(17) => B(17), B(16) => B(16), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => B(0), CI => n2, SUM(39) 
                           => S(39), SUM(38) => S(38), SUM(37) => S(37), 
                           SUM(36) => S(36), SUM(35) => S(35), SUM(34) => S(34)
                           , SUM(33) => S(33), SUM(32) => S(32), SUM(31) => 
                           S(31), SUM(30) => S(30), SUM(29) => S(29), SUM(28) 
                           => S(28), SUM(27) => S(27), SUM(26) => S(26), 
                           SUM(25) => S(25), SUM(24) => S(24), SUM(23) => S(23)
                           , SUM(22) => S(22), SUM(21) => S(21), SUM(20) => 
                           S(20), SUM(19) => S(19), SUM(18) => S(18), SUM(17) 
                           => S(17), SUM(16) => S(16), SUM(15) => S(15), 
                           SUM(14) => S(14), SUM(13) => S(13), SUM(12) => S(12)
                           , SUM(11) => S(11), SUM(10) => S(10), SUM(9) => S(9)
                           , SUM(8) => S(8), SUM(7) => S(7), SUM(6) => S(6), 
                           SUM(5) => S(5), SUM(4) => S(4), SUM(3) => S(3), 
                           SUM(2) => S(2), SUM(1) => S(1), SUM(0) => S(0), CO 
                           => n_1077);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT38 is

   port( A, B : in std_logic_vector (37 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (37 downto 0);  Co : out std_logic);

end RCA_NBIT38;

architecture SYN_DIRECT of RCA_NBIT38 is

   component RCA_NBIT38_DW01_add_0
      port( A, B : in std_logic_vector (37 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (37 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1078 : std_logic;

begin
   
   Co <= '0';
   n2 <= '0';
   add_95 : RCA_NBIT38_DW01_add_0 port map( A(37) => A(37), A(36) => A(36), 
                           A(35) => A(35), A(34) => A(34), A(33) => A(33), 
                           A(32) => A(32), A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => n2, SUM(37) => S(37), 
                           SUM(36) => S(36), SUM(35) => S(35), SUM(34) => S(34)
                           , SUM(33) => S(33), SUM(32) => S(32), SUM(31) => 
                           S(31), SUM(30) => S(30), SUM(29) => S(29), SUM(28) 
                           => S(28), SUM(27) => S(27), SUM(26) => S(26), 
                           SUM(25) => S(25), SUM(24) => S(24), SUM(23) => S(23)
                           , SUM(22) => S(22), SUM(21) => S(21), SUM(20) => 
                           S(20), SUM(19) => S(19), SUM(18) => S(18), SUM(17) 
                           => S(17), SUM(16) => S(16), SUM(15) => S(15), 
                           SUM(14) => S(14), SUM(13) => S(13), SUM(12) => S(12)
                           , SUM(11) => S(11), SUM(10) => S(10), SUM(9) => S(9)
                           , SUM(8) => S(8), SUM(7) => S(7), SUM(6) => S(6), 
                           SUM(5) => S(5), SUM(4) => S(4), SUM(3) => S(3), 
                           SUM(2) => S(2), SUM(1) => S(1), SUM(0) => S(0), CO 
                           => n_1078);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT36 is

   port( A, B : in std_logic_vector (35 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (35 downto 0);  Co : out std_logic);

end RCA_NBIT36;

architecture SYN_DIRECT of RCA_NBIT36 is

   component RCA_NBIT36_DW01_add_0
      port( A, B : in std_logic_vector (35 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (35 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1079 : std_logic;

begin
   
   Co <= '0';
   n2 <= '0';
   add_95 : RCA_NBIT36_DW01_add_0 port map( A(35) => A(35), A(34) => A(34), 
                           A(33) => A(33), A(32) => A(32), A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(35) => B(35), 
                           B(34) => B(34), B(33) => B(33), B(32) => B(32), 
                           B(31) => B(31), B(30) => B(30), B(29) => B(29), 
                           B(28) => B(28), B(27) => B(27), B(26) => B(26), 
                           B(25) => B(25), B(24) => B(24), B(23) => B(23), 
                           B(22) => B(22), B(21) => B(21), B(20) => B(20), 
                           B(19) => B(19), B(18) => B(18), B(17) => B(17), 
                           B(16) => B(16), B(15) => B(15), B(14) => B(14), 
                           B(13) => B(13), B(12) => B(12), B(11) => B(11), 
                           B(10) => B(10), B(9) => B(9), B(8) => B(8), B(7) => 
                           B(7), B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3)
                           => B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), 
                           CI => n2, SUM(35) => S(35), SUM(34) => S(34), 
                           SUM(33) => S(33), SUM(32) => S(32), SUM(31) => S(31)
                           , SUM(30) => S(30), SUM(29) => S(29), SUM(28) => 
                           S(28), SUM(27) => S(27), SUM(26) => S(26), SUM(25) 
                           => S(25), SUM(24) => S(24), SUM(23) => S(23), 
                           SUM(22) => S(22), SUM(21) => S(21), SUM(20) => S(20)
                           , SUM(19) => S(19), SUM(18) => S(18), SUM(17) => 
                           S(17), SUM(16) => S(16), SUM(15) => S(15), SUM(14) 
                           => S(14), SUM(13) => S(13), SUM(12) => S(12), 
                           SUM(11) => S(11), SUM(10) => S(10), SUM(9) => S(9), 
                           SUM(8) => S(8), SUM(7) => S(7), SUM(6) => S(6), 
                           SUM(5) => S(5), SUM(4) => S(4), SUM(3) => S(3), 
                           SUM(2) => S(2), SUM(1) => S(1), SUM(0) => S(0), CO 
                           => n_1079);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT64_i30 is

   port( A_s, A_ns, B : in std_logic_vector (63 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (63 downto 0));

end BOOTHENC_NBIT64_i30;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT64_i30 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, O_63_port, O_62_port, O_61_port, O_60_port, O_59_port,
      O_58_port, O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, 
      O_52_port, O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, 
      O_46_port, O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, 
      O_40_port, O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, 
      O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, 
      O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, 
      O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, 
      O_16_port, O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, 
      O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, 
      O_3_port, O_2_port, O_1_port, n128, n129, n130, n131, n132, n133, n134, 
      n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, 
      n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, 
      n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, 
      n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, 
      n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, 
      n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, 
      n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, 
      n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, 
      n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, 
      n340, n341, n342, n343, n344, n345, n346, n347 : std_logic;

begin
   O <= ( O_63_port, O_62_port, O_61_port, O_60_port, O_59_port, O_58_port, 
      O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, O_52_port, 
      O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, O_46_port, 
      O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, O_40_port, 
      O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, 
      O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, 
      O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, 
      O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, O_16_port, 
      O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, O_10_port, 
      O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, O_3_port, 
      O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(61), A_s(60), A_s(59), A_s(58), A_s(57), A_s(56), A_s(55), 
      A_s(54), A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), 
      A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), 
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   A_nso <= ( A_ns(61), A_ns(60), A_ns(59), A_ns(58), A_ns(57), A_ns(56), 
      A_ns(55), A_ns(54), A_ns(53), A_ns(52), A_ns(51), A_ns(50), A_ns(49), 
      A_ns(48), A_ns(47), A_ns(46), A_ns(45), A_ns(44), A_ns(43), A_ns(42), 
      A_ns(41), A_ns(40), A_ns(39), A_ns(38), A_ns(37), A_ns(36), A_ns(35), 
      A_ns(34), A_ns(33), A_ns(32), A_ns(31), A_ns(30), A_ns(29), A_ns(28), 
      A_ns(27), A_ns(26), A_ns(25), A_ns(24), A_ns(23), A_ns(22), A_ns(21), 
      A_ns(20), A_ns(19), A_ns(18), A_ns(17), A_ns(16), A_ns(15), A_ns(14), 
      A_ns(13), A_ns(12), A_ns(11), A_ns(10), A_ns(9), A_ns(8), A_ns(7), 
      A_ns(6), A_ns(5), A_ns(4), A_ns(3), A_ns(2), A_ns(1), A_ns(0), 
      X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U257 : XOR2_X1 port map( A => B(29), B => B(30), Z => n194);
   U258 : NAND3_X1 port map( A1 => B(30), A2 => n347, A3 => B(29), ZN => n128);
   U2 : OAI221_X1 port map( B1 => n215, B2 => n281, C1 => n211, C2 => n247, A 
                           => n140, ZN => O_58_port);
   U3 : OAI221_X1 port map( B1 => n215, B2 => n282, C1 => n212, C2 => n248, A 
                           => n139, ZN => O_59_port);
   U4 : OAI221_X1 port map( B1 => n215, B2 => n285, C1 => n212, C2 => n251, A 
                           => n135, ZN => O_62_port);
   U5 : OAI221_X1 port map( B1 => n216, B2 => n279, C1 => n211, C2 => n245, A 
                           => n142, ZN => O_56_port);
   U6 : AOI22_X1 port map( A1 => A_ns(29), A2 => n203, B1 => A_s(29), B2 => 
                           n197, ZN => n170);
   U7 : AOI22_X1 port map( A1 => A_ns(30), A2 => n203, B1 => A_s(30), B2 => 
                           n197, ZN => n169);
   U8 : AOI22_X1 port map( A1 => A_ns(31), A2 => n203, B1 => A_s(31), B2 => 
                           n197, ZN => n168);
   U9 : AOI22_X1 port map( A1 => A_ns(32), A2 => n204, B1 => A_s(32), B2 => 
                           n198, ZN => n167);
   U10 : AOI22_X1 port map( A1 => A_ns(33), A2 => n204, B1 => A_s(33), B2 => 
                           n198, ZN => n166);
   U11 : AOI22_X1 port map( A1 => A_ns(34), A2 => n204, B1 => A_s(34), B2 => 
                           n198, ZN => n165);
   U12 : AOI22_X1 port map( A1 => A_ns(43), A2 => n205, B1 => A_s(43), B2 => 
                           n199, ZN => n155);
   U13 : AOI22_X1 port map( A1 => A_ns(44), A2 => n205, B1 => A_s(44), B2 => 
                           n199, ZN => n154);
   U14 : AOI22_X1 port map( A1 => A_ns(45), A2 => n205, B1 => A_s(45), B2 => 
                           n199, ZN => n153);
   U15 : AOI22_X1 port map( A1 => A_ns(46), A2 => n205, B1 => A_s(46), B2 => 
                           n199, ZN => n152);
   U16 : AOI22_X1 port map( A1 => A_ns(47), A2 => n205, B1 => A_s(47), B2 => 
                           n199, ZN => n151);
   U17 : AOI22_X1 port map( A1 => A_ns(48), A2 => n205, B1 => A_s(48), B2 => 
                           n199, ZN => n150);
   U18 : AOI22_X1 port map( A1 => A_ns(49), A2 => n205, B1 => A_s(49), B2 => 
                           n199, ZN => n148);
   U19 : AOI22_X1 port map( A1 => A_ns(50), A2 => n205, B1 => A_s(50), B2 => 
                           n199, ZN => n147);
   U20 : AOI22_X1 port map( A1 => A_ns(51), A2 => n205, B1 => A_s(51), B2 => 
                           n199, ZN => n146);
   U21 : AOI22_X1 port map( A1 => A_ns(52), A2 => n205, B1 => A_s(52), B2 => 
                           n199, ZN => n145);
   U22 : AOI22_X1 port map( A1 => A_ns(53), A2 => n205, B1 => A_s(53), B2 => 
                           n199, ZN => n144);
   U23 : AOI22_X1 port map( A1 => A_ns(54), A2 => n206, B1 => A_s(54), B2 => 
                           n200, ZN => n143);
   U24 : AOI22_X1 port map( A1 => A_ns(55), A2 => n206, B1 => A_s(55), B2 => 
                           n200, ZN => n142);
   U25 : AOI22_X1 port map( A1 => A_ns(56), A2 => n206, B1 => A_s(56), B2 => 
                           n200, ZN => n141);
   U26 : AOI22_X1 port map( A1 => A_ns(57), A2 => n206, B1 => A_s(57), B2 => 
                           n200, ZN => n140);
   U27 : AOI22_X1 port map( A1 => A_ns(58), A2 => n206, B1 => A_s(58), B2 => 
                           n200, ZN => n139);
   U28 : AOI22_X1 port map( A1 => A_ns(59), A2 => n206, B1 => A_s(59), B2 => 
                           n200, ZN => n137);
   U29 : AOI22_X1 port map( A1 => A_ns(60), A2 => n206, B1 => A_s(60), B2 => 
                           n200, ZN => n136);
   U30 : AOI22_X1 port map( A1 => A_ns(61), A2 => n206, B1 => A_s(61), B2 => 
                           n200, ZN => n135);
   U31 : AOI22_X1 port map( A1 => A_ns(35), A2 => n204, B1 => A_s(35), B2 => 
                           n198, ZN => n164);
   U32 : AOI22_X1 port map( A1 => A_ns(36), A2 => n204, B1 => A_s(36), B2 => 
                           n198, ZN => n163);
   U33 : AOI22_X1 port map( A1 => A_ns(37), A2 => n204, B1 => A_s(37), B2 => 
                           n198, ZN => n162);
   U34 : AOI22_X1 port map( A1 => A_ns(38), A2 => n204, B1 => A_s(38), B2 => 
                           n198, ZN => n161);
   U35 : AOI22_X1 port map( A1 => A_ns(39), A2 => n204, B1 => A_s(39), B2 => 
                           n198, ZN => n159);
   U36 : AOI22_X1 port map( A1 => A_ns(40), A2 => n204, B1 => A_s(40), B2 => 
                           n198, ZN => n158);
   U37 : AOI22_X1 port map( A1 => A_ns(41), A2 => n204, B1 => A_s(41), B2 => 
                           n198, ZN => n157);
   U38 : AOI22_X1 port map( A1 => A_ns(42), A2 => n204, B1 => A_s(42), B2 => 
                           n198, ZN => n156);
   U39 : AOI22_X1 port map( A1 => A_ns(62), A2 => n206, B1 => A_s(62), B2 => 
                           n200, ZN => n134);
   U40 : BUF_X1 port map( A => n346, Z => n203);
   U41 : BUF_X1 port map( A => n346, Z => n204);
   U42 : BUF_X1 port map( A => n345, Z => n197);
   U43 : BUF_X1 port map( A => n345, Z => n198);
   U44 : BUF_X1 port map( A => n345, Z => n199);
   U45 : BUF_X1 port map( A => n346, Z => n205);
   U46 : BUF_X1 port map( A => n345, Z => n200);
   U47 : BUF_X1 port map( A => n346, Z => n206);
   U48 : BUF_X1 port map( A => n346, Z => n202);
   U49 : BUF_X1 port map( A => n345, Z => n196);
   U50 : OAI221_X1 port map( B1 => n215, B2 => n284, C1 => n212, C2 => n250, A 
                           => n136, ZN => O_61_port);
   U51 : OAI221_X1 port map( B1 => n215, B2 => n283, C1 => n212, C2 => n249, A 
                           => n137, ZN => O_60_port);
   U52 : OAI221_X1 port map( B1 => n215, B2 => n280, C1 => n211, C2 => n246, A 
                           => n141, ZN => O_57_port);
   U53 : OAI221_X1 port map( B1 => n216, B2 => n278, C1 => n211, C2 => n244, A 
                           => n143, ZN => O_55_port);
   U54 : OAI221_X1 port map( B1 => n216, B2 => n277, C1 => n211, C2 => n243, A 
                           => n144, ZN => O_54_port);
   U55 : OAI221_X1 port map( B1 => n216, B2 => n276, C1 => n211, C2 => n242, A 
                           => n145, ZN => O_53_port);
   U56 : OAI221_X1 port map( B1 => n216, B2 => n272, C1 => n211, C2 => n238, A 
                           => n150, ZN => O_49_port);
   U57 : OAI221_X1 port map( B1 => n216, B2 => n271, C1 => n211, C2 => n237, A 
                           => n151, ZN => O_48_port);
   U58 : OAI221_X1 port map( B1 => n216, B2 => n275, C1 => n211, C2 => n241, A 
                           => n146, ZN => O_52_port);
   U59 : OAI221_X1 port map( B1 => n216, B2 => n274, C1 => n211, C2 => n240, A 
                           => n147, ZN => O_51_port);
   U60 : OAI221_X1 port map( B1 => n216, B2 => n273, C1 => n211, C2 => n239, A 
                           => n148, ZN => O_50_port);
   U61 : OAI221_X1 port map( B1 => n216, B2 => n270, C1 => n211, C2 => n236, A 
                           => n152, ZN => O_47_port);
   U62 : OAI221_X1 port map( B1 => n216, B2 => n269, C1 => n210, C2 => n235, A 
                           => n153, ZN => O_46_port);
   U63 : OAI221_X1 port map( B1 => n217, B2 => n268, C1 => n210, C2 => n234, A 
                           => n154, ZN => O_45_port);
   U64 : OAI221_X1 port map( B1 => n217, B2 => n267, C1 => n210, C2 => n233, A 
                           => n155, ZN => O_44_port);
   U65 : OAI221_X1 port map( B1 => n217, B2 => n266, C1 => n210, C2 => n232, A 
                           => n156, ZN => O_43_port);
   U66 : OAI221_X1 port map( B1 => n217, B2 => n265, C1 => n210, C2 => n231, A 
                           => n157, ZN => O_42_port);
   U67 : OAI221_X1 port map( B1 => n217, B2 => n264, C1 => n210, C2 => n230, A 
                           => n158, ZN => O_41_port);
   U68 : OAI221_X1 port map( B1 => n217, B2 => n263, C1 => n210, C2 => n229, A 
                           => n159, ZN => O_40_port);
   U69 : OAI221_X1 port map( B1 => n217, B2 => n262, C1 => n210, C2 => n228, A 
                           => n161, ZN => O_39_port);
   U70 : OAI221_X1 port map( B1 => n218, B2 => n255, C1 => n209, C2 => n221, A 
                           => n168, ZN => O_32_port);
   U71 : OAI221_X1 port map( B1 => n218, B2 => n256, C1 => n209, C2 => n222, A 
                           => n167, ZN => O_33_port);
   U72 : OAI221_X1 port map( B1 => n218, B2 => n257, C1 => n209, C2 => n223, A 
                           => n166, ZN => O_34_port);
   U73 : OAI221_X1 port map( B1 => n217, B2 => n258, C1 => n210, C2 => n224, A 
                           => n165, ZN => O_35_port);
   U74 : OAI221_X1 port map( B1 => n217, B2 => n259, C1 => n210, C2 => n225, A 
                           => n164, ZN => O_36_port);
   U75 : OAI221_X1 port map( B1 => n217, B2 => n260, C1 => n210, C2 => n226, A 
                           => n163, ZN => O_37_port);
   U76 : OAI221_X1 port map( B1 => n217, B2 => n261, C1 => n210, C2 => n227, A 
                           => n162, ZN => O_38_port);
   U77 : OAI221_X1 port map( B1 => n215, B2 => n286, C1 => n212, C2 => n252, A 
                           => n134, ZN => O_63_port);
   U78 : BUF_X1 port map( A => n214, Z => n209);
   U79 : BUF_X1 port map( A => n213, Z => n210);
   U80 : INV_X1 port map( A => n183, ZN => n346);
   U81 : INV_X1 port map( A => n182, ZN => n345);
   U82 : BUF_X1 port map( A => n213, Z => n211);
   U83 : BUF_X1 port map( A => n213, Z => n212);
   U84 : BUF_X1 port map( A => n214, Z => n208);
   U85 : OAI221_X1 port map( B1 => n218, B2 => n254, C1 => n209, C2 => n253, A 
                           => n169, ZN => O_31_port);
   U86 : BUF_X1 port map( A => n128, Z => n217);
   U87 : BUF_X1 port map( A => n128, Z => n218);
   U88 : NAND2_X1 port map( A1 => n194, A2 => n347, ZN => n182);
   U89 : NAND2_X1 port map( A1 => n194, A2 => n182, ZN => n183);
   U90 : BUF_X1 port map( A => n129, Z => n213);
   U91 : BUF_X1 port map( A => n129, Z => n214);
   U92 : BUF_X1 port map( A => n128, Z => n216);
   U93 : BUF_X1 port map( A => n128, Z => n215);
   U94 : BUF_X1 port map( A => n128, Z => n219);
   U95 : OAI221_X1 port map( B1 => n218, B2 => n344, C1 => n209, C2 => n343, A 
                           => n170, ZN => O_30_port);
   U96 : INV_X1 port map( A => A_s(28), ZN => n344);
   U97 : INV_X1 port map( A => A_ns(28), ZN => n343);
   U98 : OAI221_X1 port map( B1 => n218, B2 => n342, C1 => n209, C2 => n340, A 
                           => n172, ZN => O_29_port);
   U99 : INV_X1 port map( A => A_s(27), ZN => n342);
   U100 : INV_X1 port map( A => A_ns(27), ZN => n340);
   U101 : OAI221_X1 port map( B1 => n219, B2 => n322, C1 => n208, C2 => n320, A
                           => n184, ZN => O_19_port);
   U102 : INV_X1 port map( A => A_s(17), ZN => n322);
   U103 : INV_X1 port map( A => A_ns(17), ZN => n320);
   U104 : OAI221_X1 port map( B1 => n219, B2 => n325, C1 => n208, C2 => n323, A
                           => n181, ZN => O_20_port);
   U105 : INV_X1 port map( A => A_s(18), ZN => n325);
   U106 : INV_X1 port map( A => A_ns(18), ZN => n323);
   U107 : OAI221_X1 port map( B1 => n219, B2 => n326, C1 => n208, C2 => n324, A
                           => n180, ZN => O_21_port);
   U108 : INV_X1 port map( A => A_s(19), ZN => n326);
   U109 : INV_X1 port map( A => A_ns(19), ZN => n324);
   U110 : OAI221_X1 port map( B1 => n219, B2 => n329, C1 => n208, C2 => n327, A
                           => n179, ZN => O_22_port);
   U111 : INV_X1 port map( A => A_s(20), ZN => n329);
   U112 : INV_X1 port map( A => A_ns(20), ZN => n327);
   U113 : OAI221_X1 port map( B1 => n219, B2 => n330, C1 => n209, C2 => n328, A
                           => n178, ZN => O_23_port);
   U114 : INV_X1 port map( A => A_s(21), ZN => n330);
   U115 : INV_X1 port map( A => A_ns(21), ZN => n328);
   U116 : OAI221_X1 port map( B1 => n218, B2 => n333, C1 => n209, C2 => n331, A
                           => n177, ZN => O_24_port);
   U117 : INV_X1 port map( A => A_s(22), ZN => n333);
   U118 : INV_X1 port map( A => A_ns(22), ZN => n331);
   U119 : OAI221_X1 port map( B1 => n218, B2 => n334, C1 => n209, C2 => n332, A
                           => n176, ZN => O_25_port);
   U120 : INV_X1 port map( A => A_s(23), ZN => n334);
   U121 : INV_X1 port map( A => A_ns(23), ZN => n332);
   U122 : OAI221_X1 port map( B1 => n218, B2 => n337, C1 => n209, C2 => n335, A
                           => n175, ZN => O_26_port);
   U123 : INV_X1 port map( A => A_s(24), ZN => n337);
   U124 : INV_X1 port map( A => A_ns(24), ZN => n335);
   U125 : OAI221_X1 port map( B1 => n218, B2 => n338, C1 => n209, C2 => n336, A
                           => n174, ZN => O_27_port);
   U126 : INV_X1 port map( A => A_s(25), ZN => n338);
   U127 : INV_X1 port map( A => A_ns(25), ZN => n336);
   U128 : OAI221_X1 port map( B1 => n218, B2 => n341, C1 => n209, C2 => n339, A
                           => n173, ZN => O_28_port);
   U129 : INV_X1 port map( A => A_s(26), ZN => n341);
   U130 : INV_X1 port map( A => A_ns(26), ZN => n339);
   U131 : INV_X1 port map( A => B(31), ZN => n347);
   U132 : OAI221_X1 port map( B1 => n215, B2 => n301, C1 => n212, C2 => n299, A
                           => n131, ZN => O_8_port);
   U133 : INV_X1 port map( A => A_s(6), ZN => n301);
   U134 : INV_X1 port map( A => A_ns(6), ZN => n299);
   U135 : OAI221_X1 port map( B1 => n215, B2 => n302, C1 => n212, C2 => n300, A
                           => n130, ZN => O_9_port);
   U136 : INV_X1 port map( A => A_s(7), ZN => n302);
   U137 : INV_X1 port map( A => A_ns(7), ZN => n300);
   U138 : OAI221_X1 port map( B1 => n305, B2 => n220, C1 => n303, C2 => n208, A
                           => n193, ZN => O_10_port);
   U139 : INV_X1 port map( A => A_ns(8), ZN => n303);
   U140 : INV_X1 port map( A => A_s(8), ZN => n305);
   U141 : OAI221_X1 port map( B1 => n220, B2 => n306, C1 => n208, C2 => n304, A
                           => n192, ZN => O_11_port);
   U142 : INV_X1 port map( A => A_s(9), ZN => n306);
   U143 : INV_X1 port map( A => A_ns(9), ZN => n304);
   U144 : OAI221_X1 port map( B1 => n219, B2 => n309, C1 => n208, C2 => n307, A
                           => n191, ZN => O_12_port);
   U145 : INV_X1 port map( A => A_s(10), ZN => n309);
   U146 : INV_X1 port map( A => A_ns(10), ZN => n307);
   U147 : OAI221_X1 port map( B1 => n219, B2 => n310, C1 => n208, C2 => n308, A
                           => n190, ZN => O_13_port);
   U148 : INV_X1 port map( A => A_s(11), ZN => n310);
   U149 : INV_X1 port map( A => A_ns(11), ZN => n308);
   U150 : OAI221_X1 port map( B1 => n219, B2 => n313, C1 => n208, C2 => n311, A
                           => n189, ZN => O_14_port);
   U151 : INV_X1 port map( A => A_s(12), ZN => n313);
   U152 : INV_X1 port map( A => A_ns(12), ZN => n311);
   U153 : OAI221_X1 port map( B1 => n219, B2 => n314, C1 => n208, C2 => n312, A
                           => n188, ZN => O_15_port);
   U154 : INV_X1 port map( A => A_s(13), ZN => n314);
   U155 : INV_X1 port map( A => A_ns(13), ZN => n312);
   U156 : OAI221_X1 port map( B1 => n219, B2 => n317, C1 => n208, C2 => n315, A
                           => n187, ZN => O_16_port);
   U157 : INV_X1 port map( A => A_s(14), ZN => n317);
   U158 : INV_X1 port map( A => A_ns(14), ZN => n315);
   U159 : OAI221_X1 port map( B1 => n219, B2 => n318, C1 => n208, C2 => n316, A
                           => n186, ZN => O_17_port);
   U160 : INV_X1 port map( A => A_s(15), ZN => n318);
   U161 : INV_X1 port map( A => A_ns(15), ZN => n316);
   U162 : OAI221_X1 port map( B1 => n219, B2 => n321, C1 => n208, C2 => n319, A
                           => n185, ZN => O_18_port);
   U163 : INV_X1 port map( A => A_s(16), ZN => n321);
   U164 : INV_X1 port map( A => A_ns(16), ZN => n319);
   U165 : OR3_X1 port map( A1 => B(29), A2 => B(30), A3 => n347, ZN => n129);
   U166 : OAI22_X1 port map( A1 => n182, A2 => n289, B1 => n183, B2 => n287, ZN
                           => O_1_port);
   U167 : OAI221_X1 port map( B1 => n218, B2 => n289, C1 => n209, C2 => n287, A
                           => n171, ZN => O_2_port);
   U168 : AOI22_X1 port map( A1 => A_ns(1), A2 => n203, B1 => A_s(1), B2 => 
                           n197, ZN => n171);
   U169 : OAI221_X1 port map( B1 => n217, B2 => n290, C1 => n210, C2 => n288, A
                           => n160, ZN => O_3_port);
   U170 : INV_X1 port map( A => A_s(1), ZN => n290);
   U171 : INV_X1 port map( A => A_ns(1), ZN => n288);
   U172 : OAI221_X1 port map( B1 => n216, B2 => n293, C1 => n211, C2 => n291, A
                           => n149, ZN => O_4_port);
   U173 : INV_X1 port map( A => A_s(2), ZN => n293);
   U174 : INV_X1 port map( A => A_ns(2), ZN => n291);
   U175 : OAI221_X1 port map( B1 => n215, B2 => n294, C1 => n212, C2 => n292, A
                           => n138, ZN => O_5_port);
   U176 : INV_X1 port map( A => A_s(3), ZN => n294);
   U177 : INV_X1 port map( A => A_ns(3), ZN => n292);
   U178 : OAI221_X1 port map( B1 => n215, B2 => n297, C1 => n212, C2 => n295, A
                           => n133, ZN => O_6_port);
   U179 : INV_X1 port map( A => A_s(4), ZN => n297);
   U180 : INV_X1 port map( A => A_ns(4), ZN => n295);
   U181 : OAI221_X1 port map( B1 => n215, B2 => n298, C1 => n212, C2 => n296, A
                           => n132, ZN => O_7_port);
   U182 : INV_X1 port map( A => A_s(5), ZN => n298);
   U183 : INV_X1 port map( A => A_ns(5), ZN => n296);
   U184 : INV_X1 port map( A => A_ns(0), ZN => n287);
   U185 : INV_X1 port map( A => A_s(0), ZN => n289);
   U186 : AOI22_X1 port map( A1 => A_ns(2), A2 => n204, B1 => A_s(2), B2 => 
                           n198, ZN => n160);
   U187 : AOI22_X1 port map( A1 => A_ns(3), A2 => n205, B1 => A_s(3), B2 => 
                           n199, ZN => n149);
   U188 : AOI22_X1 port map( A1 => A_ns(4), A2 => n206, B1 => A_s(4), B2 => 
                           n200, ZN => n138);
   U189 : AOI22_X1 port map( A1 => A_ns(5), A2 => n206, B1 => A_s(5), B2 => 
                           n200, ZN => n133);
   U190 : AOI22_X1 port map( A1 => A_ns(6), A2 => n206, B1 => A_s(6), B2 => 
                           n200, ZN => n132);
   U191 : AOI22_X1 port map( A1 => A_ns(7), A2 => n207, B1 => A_s(7), B2 => 
                           n201, ZN => n131);
   U192 : AOI22_X1 port map( A1 => A_ns(8), A2 => n207, B1 => A_s(8), B2 => 
                           n201, ZN => n130);
   U193 : AOI22_X1 port map( A1 => A_ns(9), A2 => n202, B1 => A_s(9), B2 => 
                           n196, ZN => n193);
   U194 : AOI22_X1 port map( A1 => A_ns(10), A2 => n202, B1 => A_s(10), B2 => 
                           n196, ZN => n192);
   U195 : AOI22_X1 port map( A1 => A_ns(11), A2 => n202, B1 => A_s(11), B2 => 
                           n196, ZN => n191);
   U196 : AOI22_X1 port map( A1 => A_ns(12), A2 => n202, B1 => A_s(12), B2 => 
                           n196, ZN => n190);
   U197 : AOI22_X1 port map( A1 => A_ns(13), A2 => n202, B1 => A_s(13), B2 => 
                           n196, ZN => n189);
   U198 : AOI22_X1 port map( A1 => A_ns(14), A2 => n202, B1 => A_s(14), B2 => 
                           n196, ZN => n188);
   U199 : AOI22_X1 port map( A1 => A_ns(15), A2 => n202, B1 => A_s(15), B2 => 
                           n196, ZN => n187);
   U200 : AOI22_X1 port map( A1 => A_ns(16), A2 => n202, B1 => A_s(16), B2 => 
                           n196, ZN => n186);
   U201 : AOI22_X1 port map( A1 => A_ns(17), A2 => n202, B1 => A_s(17), B2 => 
                           n196, ZN => n185);
   U202 : AOI22_X1 port map( A1 => A_ns(18), A2 => n202, B1 => A_s(18), B2 => 
                           n196, ZN => n184);
   U203 : AOI22_X1 port map( A1 => A_ns(19), A2 => n202, B1 => A_s(19), B2 => 
                           n196, ZN => n181);
   U204 : AOI22_X1 port map( A1 => A_ns(20), A2 => n202, B1 => A_s(20), B2 => 
                           n196, ZN => n180);
   U205 : AOI22_X1 port map( A1 => A_ns(21), A2 => n203, B1 => A_s(21), B2 => 
                           n197, ZN => n179);
   U206 : AOI22_X1 port map( A1 => A_ns(22), A2 => n203, B1 => A_s(22), B2 => 
                           n197, ZN => n178);
   U207 : AOI22_X1 port map( A1 => A_ns(23), A2 => n203, B1 => A_s(23), B2 => 
                           n197, ZN => n177);
   U208 : AOI22_X1 port map( A1 => A_ns(24), A2 => n203, B1 => A_s(24), B2 => 
                           n197, ZN => n176);
   U209 : AOI22_X1 port map( A1 => A_ns(25), A2 => n203, B1 => A_s(25), B2 => 
                           n197, ZN => n175);
   U210 : AOI22_X1 port map( A1 => A_ns(26), A2 => n203, B1 => A_s(26), B2 => 
                           n197, ZN => n174);
   U211 : AOI22_X1 port map( A1 => A_ns(27), A2 => n203, B1 => A_s(27), B2 => 
                           n197, ZN => n173);
   U212 : AOI22_X1 port map( A1 => A_ns(28), A2 => n203, B1 => A_s(28), B2 => 
                           n197, ZN => n172);
   U213 : CLKBUF_X1 port map( A => n345, Z => n201);
   U214 : CLKBUF_X1 port map( A => n346, Z => n207);
   U215 : CLKBUF_X1 port map( A => n128, Z => n220);
   U216 : INV_X1 port map( A => A_ns(30), ZN => n221);
   U217 : INV_X1 port map( A => A_ns(31), ZN => n222);
   U218 : INV_X1 port map( A => A_ns(32), ZN => n223);
   U219 : INV_X1 port map( A => A_ns(33), ZN => n224);
   U220 : INV_X1 port map( A => A_ns(34), ZN => n225);
   U221 : INV_X1 port map( A => A_ns(35), ZN => n226);
   U222 : INV_X1 port map( A => A_ns(36), ZN => n227);
   U223 : INV_X1 port map( A => A_ns(37), ZN => n228);
   U224 : INV_X1 port map( A => A_ns(38), ZN => n229);
   U225 : INV_X1 port map( A => A_ns(39), ZN => n230);
   U226 : INV_X1 port map( A => A_ns(40), ZN => n231);
   U227 : INV_X1 port map( A => A_ns(41), ZN => n232);
   U228 : INV_X1 port map( A => A_ns(42), ZN => n233);
   U229 : INV_X1 port map( A => A_ns(43), ZN => n234);
   U230 : INV_X1 port map( A => A_ns(44), ZN => n235);
   U231 : INV_X1 port map( A => A_ns(45), ZN => n236);
   U232 : INV_X1 port map( A => A_ns(46), ZN => n237);
   U233 : INV_X1 port map( A => A_ns(47), ZN => n238);
   U234 : INV_X1 port map( A => A_ns(48), ZN => n239);
   U235 : INV_X1 port map( A => A_ns(49), ZN => n240);
   U236 : INV_X1 port map( A => A_ns(50), ZN => n241);
   U237 : INV_X1 port map( A => A_ns(51), ZN => n242);
   U238 : INV_X1 port map( A => A_ns(52), ZN => n243);
   U239 : INV_X1 port map( A => A_ns(53), ZN => n244);
   U240 : INV_X1 port map( A => A_ns(54), ZN => n245);
   U241 : INV_X1 port map( A => A_ns(55), ZN => n246);
   U242 : INV_X1 port map( A => A_ns(56), ZN => n247);
   U243 : INV_X1 port map( A => A_ns(57), ZN => n248);
   U244 : INV_X1 port map( A => A_ns(58), ZN => n249);
   U245 : INV_X1 port map( A => A_ns(59), ZN => n250);
   U246 : INV_X1 port map( A => A_ns(60), ZN => n251);
   U247 : INV_X1 port map( A => A_ns(61), ZN => n252);
   U248 : INV_X1 port map( A => A_ns(29), ZN => n253);
   U249 : INV_X1 port map( A => A_s(29), ZN => n254);
   U250 : INV_X1 port map( A => A_s(30), ZN => n255);
   U251 : INV_X1 port map( A => A_s(31), ZN => n256);
   U252 : INV_X1 port map( A => A_s(32), ZN => n257);
   U253 : INV_X1 port map( A => A_s(33), ZN => n258);
   U254 : INV_X1 port map( A => A_s(34), ZN => n259);
   U255 : INV_X1 port map( A => A_s(35), ZN => n260);
   U256 : INV_X1 port map( A => A_s(36), ZN => n261);
   U259 : INV_X1 port map( A => A_s(37), ZN => n262);
   U260 : INV_X1 port map( A => A_s(38), ZN => n263);
   U261 : INV_X1 port map( A => A_s(39), ZN => n264);
   U262 : INV_X1 port map( A => A_s(40), ZN => n265);
   U263 : INV_X1 port map( A => A_s(41), ZN => n266);
   U264 : INV_X1 port map( A => A_s(42), ZN => n267);
   U265 : INV_X1 port map( A => A_s(43), ZN => n268);
   U266 : INV_X1 port map( A => A_s(44), ZN => n269);
   U267 : INV_X1 port map( A => A_s(45), ZN => n270);
   U268 : INV_X1 port map( A => A_s(46), ZN => n271);
   U269 : INV_X1 port map( A => A_s(47), ZN => n272);
   U270 : INV_X1 port map( A => A_s(48), ZN => n273);
   U271 : INV_X1 port map( A => A_s(49), ZN => n274);
   U272 : INV_X1 port map( A => A_s(50), ZN => n275);
   U273 : INV_X1 port map( A => A_s(51), ZN => n276);
   U274 : INV_X1 port map( A => A_s(52), ZN => n277);
   U275 : INV_X1 port map( A => A_s(53), ZN => n278);
   U276 : INV_X1 port map( A => A_s(54), ZN => n279);
   U277 : INV_X1 port map( A => A_s(55), ZN => n280);
   U278 : INV_X1 port map( A => A_s(56), ZN => n281);
   U279 : INV_X1 port map( A => A_s(57), ZN => n282);
   U280 : INV_X1 port map( A => A_s(58), ZN => n283);
   U281 : INV_X1 port map( A => A_s(59), ZN => n284);
   U282 : INV_X1 port map( A => A_s(60), ZN => n285);
   U283 : INV_X1 port map( A => A_s(61), ZN => n286);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT62_i28 is

   port( A_s, A_ns, B : in std_logic_vector (61 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (61 downto 0));

end BOOTHENC_NBIT62_i28;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT62_i28 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, O_61_port, O_60_port, O_59_port, O_58_port, O_57_port,
      O_56_port, O_55_port, O_54_port, O_53_port, O_52_port, O_51_port, 
      O_50_port, O_49_port, O_48_port, O_47_port, O_46_port, O_45_port, 
      O_44_port, O_43_port, O_42_port, O_41_port, O_40_port, O_39_port, 
      O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, O_33_port, 
      O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, O_27_port, 
      O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, O_21_port, 
      O_20_port, O_19_port, O_18_port, O_17_port, O_16_port, O_15_port, 
      O_14_port, O_13_port, O_12_port, O_11_port, O_10_port, O_9_port, O_8_port
      , O_7_port, O_6_port, O_5_port, O_4_port, O_3_port, O_2_port, O_1_port, 
      n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, 
      n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, 
      n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, 
      n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, 
      n184, n185, n186, n187, n188, n190, n191, n192, n193, n194, n195, n196, 
      n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, 
      n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, 
      n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, 
      n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, 
      n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, 
      n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, 
      n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, 
      n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, 
      n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, 
      n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, 
      n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, 
      n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340 : 
      std_logic;

begin
   O <= ( O_61_port, O_60_port, O_59_port, O_58_port, O_57_port, O_56_port, 
      O_55_port, O_54_port, O_53_port, O_52_port, O_51_port, O_50_port, 
      O_49_port, O_48_port, O_47_port, O_46_port, O_45_port, O_44_port, 
      O_43_port, O_42_port, O_41_port, O_40_port, O_39_port, O_38_port, 
      O_37_port, O_36_port, O_35_port, O_34_port, O_33_port, O_32_port, 
      O_31_port, O_30_port, O_29_port, O_28_port, O_27_port, O_26_port, 
      O_25_port, O_24_port, O_23_port, O_22_port, O_21_port, O_20_port, 
      O_19_port, O_18_port, O_17_port, O_16_port, O_15_port, O_14_port, 
      O_13_port, O_12_port, O_11_port, O_10_port, O_9_port, O_8_port, O_7_port,
      O_6_port, O_5_port, O_4_port, O_3_port, O_2_port, O_1_port, X_Logic0_port
      );
   A_so <= ( A_s(59), A_s(58), A_s(57), A_s(56), A_s(55), A_s(54), A_s(53), 
      A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), A_s(46), A_s(45), 
      A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), A_s(38), A_s(37), 
      A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), A_s(30), A_s(29), 
      A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), A_s(22), A_s(21), 
      A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), A_s(14), A_s(13), 
      A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), A_s(6), A_s(5), A_s(4)
      , A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, X_Logic0_port );
   A_nso <= ( A_ns(59), A_ns(58), A_ns(57), A_ns(56), A_ns(55), A_ns(54), 
      A_ns(53), A_ns(52), A_ns(51), A_ns(50), A_ns(49), A_ns(48), A_ns(47), 
      A_ns(46), A_ns(45), A_ns(44), A_ns(43), A_ns(42), A_ns(41), A_ns(40), 
      A_ns(39), A_ns(38), A_ns(37), A_ns(36), A_ns(35), A_ns(34), A_ns(33), 
      A_ns(32), A_ns(31), A_ns(30), A_ns(29), A_ns(28), A_ns(27), A_ns(26), 
      A_ns(25), A_ns(24), A_ns(23), A_ns(22), A_ns(21), A_ns(20), A_ns(19), 
      A_ns(18), A_ns(17), A_ns(16), A_ns(15), A_ns(14), A_ns(13), A_ns(12), 
      A_ns(11), A_ns(10), A_ns(9), A_ns(8), A_ns(7), A_ns(6), A_ns(5), A_ns(4),
      A_ns(3), A_ns(2), A_ns(1), A_ns(0), X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U249 : XOR2_X1 port map( A => B(27), B => B(28), Z => n188);
   U250 : NAND3_X1 port map( A1 => B(28), A2 => n340, A3 => B(27), ZN => n124);
   U2 : OAI221_X1 port map( B1 => n213, B2 => n278, C1 => n207, C2 => n244, A 
                           => n136, ZN => O_56_port);
   U3 : OAI221_X1 port map( B1 => n213, B2 => n282, C1 => n208, C2 => n248, A 
                           => n131, ZN => O_60_port);
   U4 : OAI221_X1 port map( B1 => n213, B2 => n281, C1 => n208, C2 => n247, A 
                           => n133, ZN => O_59_port);
   U5 : AOI22_X1 port map( A1 => A_ns(27), A2 => n200, B1 => A_s(27), B2 => 
                           n193, ZN => n167);
   U6 : BUF_X1 port map( A => n197, Z => n200);
   U7 : BUF_X1 port map( A => n190, Z => n193);
   U8 : BUF_X1 port map( A => n197, Z => n201);
   U9 : BUF_X1 port map( A => n190, Z => n194);
   U10 : BUF_X1 port map( A => n198, Z => n202);
   U11 : BUF_X1 port map( A => n191, Z => n195);
   U12 : BUF_X1 port map( A => n198, Z => n203);
   U13 : BUF_X1 port map( A => n191, Z => n196);
   U14 : BUF_X1 port map( A => n197, Z => n199);
   U15 : BUF_X1 port map( A => n190, Z => n192);
   U16 : OAI221_X1 port map( B1 => n213, B2 => n283, C1 => n208, C2 => n249, A 
                           => n130, ZN => O_61_port);
   U17 : AOI22_X1 port map( A1 => A_ns(60), A2 => n203, B1 => A_s(60), B2 => 
                           n196, ZN => n130);
   U18 : AOI22_X1 port map( A1 => A_ns(58), A2 => n203, B1 => A_s(58), B2 => 
                           n196, ZN => n133);
   U19 : OAI221_X1 port map( B1 => n213, B2 => n279, C1 => n207, C2 => n245, A 
                           => n135, ZN => O_57_port);
   U20 : AOI22_X1 port map( A1 => A_ns(56), A2 => n203, B1 => A_s(56), B2 => 
                           n196, ZN => n135);
   U21 : OAI221_X1 port map( B1 => n213, B2 => n280, C1 => n207, C2 => n246, A 
                           => n134, ZN => O_58_port);
   U22 : AOI22_X1 port map( A1 => A_ns(57), A2 => n203, B1 => A_s(57), B2 => 
                           n196, ZN => n134);
   U23 : AOI22_X1 port map( A1 => A_ns(55), A2 => n203, B1 => A_s(55), B2 => 
                           n196, ZN => n136);
   U24 : OAI221_X1 port map( B1 => n214, B2 => n276, C1 => n207, C2 => n242, A 
                           => n138, ZN => O_54_port);
   U25 : AOI22_X1 port map( A1 => A_ns(53), A2 => n202, B1 => A_s(53), B2 => 
                           n195, ZN => n138);
   U26 : OAI221_X1 port map( B1 => n214, B2 => n275, C1 => n207, C2 => n241, A 
                           => n139, ZN => O_53_port);
   U27 : AOI22_X1 port map( A1 => A_ns(52), A2 => n202, B1 => A_s(52), B2 => 
                           n195, ZN => n139);
   U28 : OAI221_X1 port map( B1 => n215, B2 => n260, C1 => n206, C2 => n226, A 
                           => n156, ZN => O_38_port);
   U29 : AOI22_X1 port map( A1 => A_ns(37), A2 => n201, B1 => A_s(37), B2 => 
                           n194, ZN => n156);
   U30 : OAI221_X1 port map( B1 => n215, B2 => n259, C1 => n206, C2 => n225, A 
                           => n157, ZN => O_37_port);
   U31 : AOI22_X1 port map( A1 => A_ns(36), A2 => n201, B1 => A_s(36), B2 => 
                           n194, ZN => n157);
   U32 : OAI221_X1 port map( B1 => n215, B2 => n258, C1 => n206, C2 => n224, A 
                           => n158, ZN => O_36_port);
   U33 : AOI22_X1 port map( A1 => A_ns(35), A2 => n201, B1 => A_s(35), B2 => 
                           n194, ZN => n158);
   U34 : OAI221_X1 port map( B1 => n215, B2 => n257, C1 => n206, C2 => n223, A 
                           => n159, ZN => O_35_port);
   U35 : AOI22_X1 port map( A1 => A_ns(34), A2 => n201, B1 => A_s(34), B2 => 
                           n194, ZN => n159);
   U36 : OAI221_X1 port map( B1 => n215, B2 => n256, C1 => n205, C2 => n222, A 
                           => n160, ZN => O_34_port);
   U37 : AOI22_X1 port map( A1 => A_ns(33), A2 => n201, B1 => A_s(33), B2 => 
                           n194, ZN => n160);
   U38 : OAI221_X1 port map( B1 => n215, B2 => n255, C1 => n205, C2 => n221, A 
                           => n161, ZN => O_33_port);
   U39 : AOI22_X1 port map( A1 => A_ns(32), A2 => n201, B1 => A_s(32), B2 => 
                           n194, ZN => n161);
   U40 : OAI221_X1 port map( B1 => n216, B2 => n254, C1 => n205, C2 => n220, A 
                           => n162, ZN => O_32_port);
   U41 : AOI22_X1 port map( A1 => A_ns(31), A2 => n200, B1 => A_s(31), B2 => 
                           n193, ZN => n162);
   U42 : OAI221_X1 port map( B1 => n216, B2 => n253, C1 => n205, C2 => n219, A 
                           => n163, ZN => O_31_port);
   U43 : AOI22_X1 port map( A1 => A_ns(30), A2 => n200, B1 => A_s(30), B2 => 
                           n193, ZN => n163);
   U44 : AOI22_X1 port map( A1 => A_ns(59), A2 => n203, B1 => A_s(59), B2 => 
                           n196, ZN => n131);
   U45 : OAI221_X1 port map( B1 => n213, B2 => n277, C1 => n207, C2 => n243, A 
                           => n137, ZN => O_55_port);
   U46 : AOI22_X1 port map( A1 => A_ns(54), A2 => n203, B1 => A_s(54), B2 => 
                           n196, ZN => n137);
   U47 : OAI221_X1 port map( B1 => n214, B2 => n274, C1 => n207, C2 => n240, A 
                           => n140, ZN => O_52_port);
   U48 : AOI22_X1 port map( A1 => A_ns(51), A2 => n202, B1 => A_s(51), B2 => 
                           n195, ZN => n140);
   U49 : OAI221_X1 port map( B1 => n214, B2 => n273, C1 => n207, C2 => n239, A 
                           => n141, ZN => O_51_port);
   U50 : AOI22_X1 port map( A1 => A_ns(50), A2 => n202, B1 => A_s(50), B2 => 
                           n195, ZN => n141);
   U51 : OAI221_X1 port map( B1 => n214, B2 => n272, C1 => n207, C2 => n238, A 
                           => n142, ZN => O_50_port);
   U52 : AOI22_X1 port map( A1 => A_ns(49), A2 => n202, B1 => A_s(49), B2 => 
                           n195, ZN => n142);
   U53 : OAI221_X1 port map( B1 => n214, B2 => n271, C1 => n207, C2 => n237, A 
                           => n144, ZN => O_49_port);
   U54 : AOI22_X1 port map( A1 => A_ns(48), A2 => n202, B1 => A_s(48), B2 => 
                           n195, ZN => n144);
   U55 : OAI221_X1 port map( B1 => n214, B2 => n270, C1 => n207, C2 => n236, A 
                           => n145, ZN => O_48_port);
   U56 : AOI22_X1 port map( A1 => A_ns(47), A2 => n202, B1 => A_s(47), B2 => 
                           n195, ZN => n145);
   U57 : OAI221_X1 port map( B1 => n214, B2 => n269, C1 => n207, C2 => n235, A 
                           => n146, ZN => O_47_port);
   U58 : AOI22_X1 port map( A1 => A_ns(46), A2 => n202, B1 => A_s(46), B2 => 
                           n195, ZN => n146);
   U59 : OAI221_X1 port map( B1 => n214, B2 => n268, C1 => n206, C2 => n234, A 
                           => n147, ZN => O_46_port);
   U60 : AOI22_X1 port map( A1 => A_ns(45), A2 => n202, B1 => A_s(45), B2 => 
                           n195, ZN => n147);
   U61 : OAI221_X1 port map( B1 => n214, B2 => n267, C1 => n206, C2 => n233, A 
                           => n148, ZN => O_45_port);
   U62 : AOI22_X1 port map( A1 => A_ns(44), A2 => n202, B1 => A_s(44), B2 => 
                           n195, ZN => n148);
   U63 : OAI221_X1 port map( B1 => n214, B2 => n266, C1 => n206, C2 => n232, A 
                           => n149, ZN => O_44_port);
   U64 : AOI22_X1 port map( A1 => A_ns(43), A2 => n202, B1 => A_s(43), B2 => 
                           n195, ZN => n149);
   U65 : OAI221_X1 port map( B1 => n215, B2 => n265, C1 => n206, C2 => n231, A 
                           => n150, ZN => O_43_port);
   U66 : AOI22_X1 port map( A1 => A_ns(42), A2 => n201, B1 => A_s(42), B2 => 
                           n194, ZN => n150);
   U67 : OAI221_X1 port map( B1 => n215, B2 => n264, C1 => n206, C2 => n230, A 
                           => n151, ZN => O_42_port);
   U68 : AOI22_X1 port map( A1 => A_ns(41), A2 => n201, B1 => A_s(41), B2 => 
                           n194, ZN => n151);
   U69 : OAI221_X1 port map( B1 => n215, B2 => n263, C1 => n206, C2 => n229, A 
                           => n152, ZN => O_41_port);
   U70 : AOI22_X1 port map( A1 => A_ns(40), A2 => n201, B1 => A_s(40), B2 => 
                           n194, ZN => n152);
   U71 : OAI221_X1 port map( B1 => n215, B2 => n262, C1 => n206, C2 => n228, A 
                           => n153, ZN => O_40_port);
   U72 : AOI22_X1 port map( A1 => A_ns(39), A2 => n201, B1 => A_s(39), B2 => 
                           n194, ZN => n153);
   U73 : OAI221_X1 port map( B1 => n215, B2 => n261, C1 => n206, C2 => n227, A 
                           => n155, ZN => O_39_port);
   U74 : AOI22_X1 port map( A1 => A_ns(38), A2 => n201, B1 => A_s(38), B2 => 
                           n194, ZN => n155);
   U75 : BUF_X1 port map( A => n338, Z => n190);
   U76 : BUF_X1 port map( A => n339, Z => n197);
   U77 : BUF_X1 port map( A => n338, Z => n191);
   U78 : BUF_X1 port map( A => n339, Z => n198);
   U79 : OAI221_X1 port map( B1 => n216, B2 => n252, C1 => n205, C2 => n218, A 
                           => n164, ZN => O_30_port);
   U80 : AOI22_X1 port map( A1 => A_ns(29), A2 => n200, B1 => A_s(29), B2 => 
                           n193, ZN => n164);
   U81 : INV_X1 port map( A => n176, ZN => n338);
   U82 : INV_X1 port map( A => n177, ZN => n339);
   U83 : BUF_X1 port map( A => n212, Z => n216);
   U84 : BUF_X1 port map( A => n211, Z => n215);
   U85 : BUF_X1 port map( A => n210, Z => n205);
   U86 : BUF_X1 port map( A => n209, Z => n206);
   U87 : BUF_X1 port map( A => n211, Z => n214);
   U88 : BUF_X1 port map( A => n209, Z => n207);
   U89 : BUF_X1 port map( A => n211, Z => n213);
   U90 : BUF_X1 port map( A => n209, Z => n208);
   U91 : BUF_X1 port map( A => n212, Z => n217);
   U92 : BUF_X1 port map( A => n210, Z => n204);
   U93 : OAI221_X1 port map( B1 => n216, B2 => n251, C1 => n205, C2 => n250, A 
                           => n166, ZN => O_29_port);
   U94 : AOI22_X1 port map( A1 => A_ns(28), A2 => n200, B1 => A_s(28), B2 => 
                           n193, ZN => n166);
   U95 : NAND2_X1 port map( A1 => n188, A2 => n340, ZN => n176);
   U96 : NAND2_X1 port map( A1 => n188, A2 => n176, ZN => n177);
   U97 : BUF_X1 port map( A => n124, Z => n211);
   U98 : BUF_X1 port map( A => n125, Z => n209);
   U99 : BUF_X1 port map( A => n124, Z => n212);
   U100 : BUF_X1 port map( A => n125, Z => n210);
   U101 : OAI221_X1 port map( B1 => n216, B2 => n337, C1 => n205, C2 => n336, A
                           => n167, ZN => O_28_port);
   U102 : INV_X1 port map( A => A_s(26), ZN => n337);
   U103 : INV_X1 port map( A => A_ns(26), ZN => n336);
   U104 : OAI221_X1 port map( B1 => n217, B2 => n319, C1 => n204, C2 => n317, A
                           => n178, ZN => O_19_port);
   U105 : INV_X1 port map( A => A_s(17), ZN => n319);
   U106 : INV_X1 port map( A => A_ns(17), ZN => n317);
   U107 : OAI221_X1 port map( B1 => n217, B2 => n322, C1 => n204, C2 => n320, A
                           => n175, ZN => O_20_port);
   U108 : INV_X1 port map( A => A_s(18), ZN => n322);
   U109 : INV_X1 port map( A => A_ns(18), ZN => n320);
   U110 : OAI221_X1 port map( B1 => n217, B2 => n323, C1 => n204, C2 => n321, A
                           => n174, ZN => O_21_port);
   U111 : INV_X1 port map( A => A_s(19), ZN => n323);
   U112 : INV_X1 port map( A => A_ns(19), ZN => n321);
   U113 : OAI221_X1 port map( B1 => n216, B2 => n326, C1 => n204, C2 => n324, A
                           => n173, ZN => O_22_port);
   U114 : INV_X1 port map( A => A_s(20), ZN => n326);
   U115 : INV_X1 port map( A => A_ns(20), ZN => n324);
   U116 : OAI221_X1 port map( B1 => n216, B2 => n327, C1 => n205, C2 => n325, A
                           => n172, ZN => O_23_port);
   U117 : INV_X1 port map( A => A_s(21), ZN => n327);
   U118 : INV_X1 port map( A => A_ns(21), ZN => n325);
   U119 : OAI221_X1 port map( B1 => n216, B2 => n330, C1 => n205, C2 => n328, A
                           => n171, ZN => O_24_port);
   U120 : INV_X1 port map( A => A_s(22), ZN => n330);
   U121 : INV_X1 port map( A => A_ns(22), ZN => n328);
   U122 : OAI221_X1 port map( B1 => n216, B2 => n331, C1 => n205, C2 => n329, A
                           => n170, ZN => O_25_port);
   U123 : INV_X1 port map( A => A_s(23), ZN => n331);
   U124 : INV_X1 port map( A => A_ns(23), ZN => n329);
   U125 : OAI221_X1 port map( B1 => n216, B2 => n334, C1 => n205, C2 => n332, A
                           => n169, ZN => O_26_port);
   U126 : INV_X1 port map( A => A_s(24), ZN => n334);
   U127 : INV_X1 port map( A => A_ns(24), ZN => n332);
   U128 : OAI221_X1 port map( B1 => n216, B2 => n335, C1 => n205, C2 => n333, A
                           => n168, ZN => O_27_port);
   U129 : INV_X1 port map( A => A_s(25), ZN => n335);
   U130 : INV_X1 port map( A => A_ns(25), ZN => n333);
   U131 : INV_X1 port map( A => B(29), ZN => n340);
   U132 : OAI221_X1 port map( B1 => n213, B2 => n298, C1 => n208, C2 => n296, A
                           => n127, ZN => O_8_port);
   U133 : INV_X1 port map( A => A_s(6), ZN => n298);
   U134 : INV_X1 port map( A => A_ns(6), ZN => n296);
   U135 : OAI221_X1 port map( B1 => n213, B2 => n299, C1 => n208, C2 => n297, A
                           => n126, ZN => O_9_port);
   U136 : INV_X1 port map( A => A_s(7), ZN => n299);
   U137 : INV_X1 port map( A => A_ns(7), ZN => n297);
   U138 : OAI221_X1 port map( B1 => n302, B2 => n217, C1 => n300, C2 => n204, A
                           => n187, ZN => O_10_port);
   U139 : INV_X1 port map( A => A_ns(8), ZN => n300);
   U140 : INV_X1 port map( A => A_s(8), ZN => n302);
   U141 : OAI221_X1 port map( B1 => n217, B2 => n303, C1 => n204, C2 => n301, A
                           => n186, ZN => O_11_port);
   U142 : INV_X1 port map( A => A_s(9), ZN => n303);
   U143 : INV_X1 port map( A => A_ns(9), ZN => n301);
   U144 : OAI221_X1 port map( B1 => n217, B2 => n306, C1 => n204, C2 => n304, A
                           => n185, ZN => O_12_port);
   U145 : INV_X1 port map( A => A_s(10), ZN => n306);
   U146 : INV_X1 port map( A => A_ns(10), ZN => n304);
   U147 : OAI221_X1 port map( B1 => n217, B2 => n307, C1 => n204, C2 => n305, A
                           => n184, ZN => O_13_port);
   U148 : INV_X1 port map( A => A_s(11), ZN => n307);
   U149 : INV_X1 port map( A => A_ns(11), ZN => n305);
   U150 : OAI221_X1 port map( B1 => n217, B2 => n310, C1 => n204, C2 => n308, A
                           => n183, ZN => O_14_port);
   U151 : INV_X1 port map( A => A_s(12), ZN => n310);
   U152 : INV_X1 port map( A => A_ns(12), ZN => n308);
   U153 : OAI221_X1 port map( B1 => n217, B2 => n311, C1 => n204, C2 => n309, A
                           => n182, ZN => O_15_port);
   U154 : INV_X1 port map( A => A_s(13), ZN => n311);
   U155 : INV_X1 port map( A => A_ns(13), ZN => n309);
   U156 : OAI221_X1 port map( B1 => n217, B2 => n314, C1 => n204, C2 => n312, A
                           => n181, ZN => O_16_port);
   U157 : INV_X1 port map( A => A_s(14), ZN => n314);
   U158 : INV_X1 port map( A => A_ns(14), ZN => n312);
   U159 : OAI221_X1 port map( B1 => n217, B2 => n315, C1 => n204, C2 => n313, A
                           => n180, ZN => O_17_port);
   U160 : INV_X1 port map( A => A_s(15), ZN => n315);
   U161 : INV_X1 port map( A => A_ns(15), ZN => n313);
   U162 : OAI221_X1 port map( B1 => n217, B2 => n318, C1 => n204, C2 => n316, A
                           => n179, ZN => O_18_port);
   U163 : INV_X1 port map( A => A_s(16), ZN => n318);
   U164 : INV_X1 port map( A => A_ns(16), ZN => n316);
   U165 : OR3_X1 port map( A1 => B(27), A2 => B(28), A3 => n340, ZN => n125);
   U166 : OAI22_X1 port map( A1 => n176, A2 => n286, B1 => n177, B2 => n284, ZN
                           => O_1_port);
   U167 : OAI221_X1 port map( B1 => n216, B2 => n286, C1 => n205, C2 => n284, A
                           => n165, ZN => O_2_port);
   U168 : AOI22_X1 port map( A1 => A_ns(1), A2 => n200, B1 => A_s(1), B2 => 
                           n193, ZN => n165);
   U169 : OAI221_X1 port map( B1 => n215, B2 => n287, C1 => n206, C2 => n285, A
                           => n154, ZN => O_3_port);
   U170 : INV_X1 port map( A => A_s(1), ZN => n287);
   U171 : INV_X1 port map( A => A_ns(1), ZN => n285);
   U172 : OAI221_X1 port map( B1 => n214, B2 => n290, C1 => n207, C2 => n288, A
                           => n143, ZN => O_4_port);
   U173 : INV_X1 port map( A => A_s(2), ZN => n290);
   U174 : INV_X1 port map( A => A_ns(2), ZN => n288);
   U175 : OAI221_X1 port map( B1 => n213, B2 => n291, C1 => n208, C2 => n289, A
                           => n132, ZN => O_5_port);
   U176 : INV_X1 port map( A => A_s(3), ZN => n291);
   U177 : INV_X1 port map( A => A_ns(3), ZN => n289);
   U178 : OAI221_X1 port map( B1 => n213, B2 => n294, C1 => n208, C2 => n292, A
                           => n129, ZN => O_6_port);
   U179 : INV_X1 port map( A => A_s(4), ZN => n294);
   U180 : INV_X1 port map( A => A_ns(4), ZN => n292);
   U181 : OAI221_X1 port map( B1 => n213, B2 => n295, C1 => n208, C2 => n293, A
                           => n128, ZN => O_7_port);
   U182 : INV_X1 port map( A => A_s(5), ZN => n295);
   U183 : INV_X1 port map( A => A_ns(5), ZN => n293);
   U184 : INV_X1 port map( A => A_ns(0), ZN => n284);
   U185 : INV_X1 port map( A => A_s(0), ZN => n286);
   U186 : AOI22_X1 port map( A1 => A_ns(2), A2 => n201, B1 => A_s(2), B2 => 
                           n194, ZN => n154);
   U187 : AOI22_X1 port map( A1 => A_ns(3), A2 => n202, B1 => A_s(3), B2 => 
                           n195, ZN => n143);
   U188 : AOI22_X1 port map( A1 => A_ns(4), A2 => n203, B1 => A_s(4), B2 => 
                           n196, ZN => n132);
   U189 : AOI22_X1 port map( A1 => A_ns(5), A2 => n203, B1 => A_s(5), B2 => 
                           n196, ZN => n129);
   U190 : AOI22_X1 port map( A1 => A_ns(6), A2 => n203, B1 => A_s(6), B2 => 
                           n196, ZN => n128);
   U191 : AOI22_X1 port map( A1 => A_ns(7), A2 => n203, B1 => A_s(7), B2 => 
                           n196, ZN => n127);
   U192 : AOI22_X1 port map( A1 => A_ns(8), A2 => n203, B1 => A_s(8), B2 => 
                           n196, ZN => n126);
   U193 : AOI22_X1 port map( A1 => A_ns(9), A2 => n199, B1 => A_s(9), B2 => 
                           n192, ZN => n187);
   U194 : AOI22_X1 port map( A1 => A_ns(10), A2 => n199, B1 => A_s(10), B2 => 
                           n192, ZN => n186);
   U195 : AOI22_X1 port map( A1 => A_ns(11), A2 => n199, B1 => A_s(11), B2 => 
                           n192, ZN => n185);
   U196 : AOI22_X1 port map( A1 => A_ns(12), A2 => n199, B1 => A_s(12), B2 => 
                           n192, ZN => n184);
   U197 : AOI22_X1 port map( A1 => A_ns(13), A2 => n199, B1 => A_s(13), B2 => 
                           n192, ZN => n183);
   U198 : AOI22_X1 port map( A1 => A_ns(14), A2 => n199, B1 => A_s(14), B2 => 
                           n192, ZN => n182);
   U199 : AOI22_X1 port map( A1 => A_ns(15), A2 => n199, B1 => A_s(15), B2 => 
                           n192, ZN => n181);
   U200 : AOI22_X1 port map( A1 => A_ns(16), A2 => n199, B1 => A_s(16), B2 => 
                           n192, ZN => n180);
   U201 : AOI22_X1 port map( A1 => A_ns(17), A2 => n199, B1 => A_s(17), B2 => 
                           n192, ZN => n179);
   U202 : AOI22_X1 port map( A1 => A_ns(18), A2 => n199, B1 => A_s(18), B2 => 
                           n192, ZN => n178);
   U203 : AOI22_X1 port map( A1 => A_ns(19), A2 => n199, B1 => A_s(19), B2 => 
                           n192, ZN => n175);
   U204 : AOI22_X1 port map( A1 => A_ns(20), A2 => n199, B1 => A_s(20), B2 => 
                           n192, ZN => n174);
   U205 : AOI22_X1 port map( A1 => A_ns(21), A2 => n200, B1 => A_s(21), B2 => 
                           n193, ZN => n173);
   U206 : AOI22_X1 port map( A1 => A_ns(22), A2 => n200, B1 => A_s(22), B2 => 
                           n193, ZN => n172);
   U207 : AOI22_X1 port map( A1 => A_ns(23), A2 => n200, B1 => A_s(23), B2 => 
                           n193, ZN => n171);
   U208 : AOI22_X1 port map( A1 => A_ns(24), A2 => n200, B1 => A_s(24), B2 => 
                           n193, ZN => n170);
   U209 : AOI22_X1 port map( A1 => A_ns(25), A2 => n200, B1 => A_s(25), B2 => 
                           n193, ZN => n169);
   U210 : AOI22_X1 port map( A1 => A_ns(26), A2 => n200, B1 => A_s(26), B2 => 
                           n193, ZN => n168);
   U211 : INV_X1 port map( A => A_ns(28), ZN => n218);
   U212 : INV_X1 port map( A => A_ns(29), ZN => n219);
   U213 : INV_X1 port map( A => A_ns(30), ZN => n220);
   U214 : INV_X1 port map( A => A_ns(31), ZN => n221);
   U215 : INV_X1 port map( A => A_ns(32), ZN => n222);
   U216 : INV_X1 port map( A => A_ns(33), ZN => n223);
   U217 : INV_X1 port map( A => A_ns(34), ZN => n224);
   U218 : INV_X1 port map( A => A_ns(35), ZN => n225);
   U219 : INV_X1 port map( A => A_ns(36), ZN => n226);
   U220 : INV_X1 port map( A => A_ns(37), ZN => n227);
   U221 : INV_X1 port map( A => A_ns(38), ZN => n228);
   U222 : INV_X1 port map( A => A_ns(39), ZN => n229);
   U223 : INV_X1 port map( A => A_ns(40), ZN => n230);
   U224 : INV_X1 port map( A => A_ns(41), ZN => n231);
   U225 : INV_X1 port map( A => A_ns(42), ZN => n232);
   U226 : INV_X1 port map( A => A_ns(43), ZN => n233);
   U227 : INV_X1 port map( A => A_ns(44), ZN => n234);
   U228 : INV_X1 port map( A => A_ns(45), ZN => n235);
   U229 : INV_X1 port map( A => A_ns(46), ZN => n236);
   U230 : INV_X1 port map( A => A_ns(47), ZN => n237);
   U231 : INV_X1 port map( A => A_ns(48), ZN => n238);
   U232 : INV_X1 port map( A => A_ns(49), ZN => n239);
   U233 : INV_X1 port map( A => A_ns(50), ZN => n240);
   U234 : INV_X1 port map( A => A_ns(51), ZN => n241);
   U235 : INV_X1 port map( A => A_ns(52), ZN => n242);
   U236 : INV_X1 port map( A => A_ns(53), ZN => n243);
   U237 : INV_X1 port map( A => A_ns(54), ZN => n244);
   U238 : INV_X1 port map( A => A_ns(55), ZN => n245);
   U239 : INV_X1 port map( A => A_ns(56), ZN => n246);
   U240 : INV_X1 port map( A => A_ns(57), ZN => n247);
   U241 : INV_X1 port map( A => A_ns(58), ZN => n248);
   U242 : INV_X1 port map( A => A_ns(59), ZN => n249);
   U243 : INV_X1 port map( A => A_ns(27), ZN => n250);
   U244 : INV_X1 port map( A => A_s(27), ZN => n251);
   U245 : INV_X1 port map( A => A_s(28), ZN => n252);
   U246 : INV_X1 port map( A => A_s(29), ZN => n253);
   U247 : INV_X1 port map( A => A_s(30), ZN => n254);
   U248 : INV_X1 port map( A => A_s(31), ZN => n255);
   U251 : INV_X1 port map( A => A_s(32), ZN => n256);
   U252 : INV_X1 port map( A => A_s(33), ZN => n257);
   U253 : INV_X1 port map( A => A_s(34), ZN => n258);
   U254 : INV_X1 port map( A => A_s(35), ZN => n259);
   U255 : INV_X1 port map( A => A_s(36), ZN => n260);
   U256 : INV_X1 port map( A => A_s(37), ZN => n261);
   U257 : INV_X1 port map( A => A_s(38), ZN => n262);
   U258 : INV_X1 port map( A => A_s(39), ZN => n263);
   U259 : INV_X1 port map( A => A_s(40), ZN => n264);
   U260 : INV_X1 port map( A => A_s(41), ZN => n265);
   U261 : INV_X1 port map( A => A_s(42), ZN => n266);
   U262 : INV_X1 port map( A => A_s(43), ZN => n267);
   U263 : INV_X1 port map( A => A_s(44), ZN => n268);
   U264 : INV_X1 port map( A => A_s(45), ZN => n269);
   U265 : INV_X1 port map( A => A_s(46), ZN => n270);
   U266 : INV_X1 port map( A => A_s(47), ZN => n271);
   U267 : INV_X1 port map( A => A_s(48), ZN => n272);
   U268 : INV_X1 port map( A => A_s(49), ZN => n273);
   U269 : INV_X1 port map( A => A_s(50), ZN => n274);
   U270 : INV_X1 port map( A => A_s(51), ZN => n275);
   U271 : INV_X1 port map( A => A_s(52), ZN => n276);
   U272 : INV_X1 port map( A => A_s(53), ZN => n277);
   U273 : INV_X1 port map( A => A_s(54), ZN => n278);
   U274 : INV_X1 port map( A => A_s(55), ZN => n279);
   U275 : INV_X1 port map( A => A_s(56), ZN => n280);
   U276 : INV_X1 port map( A => A_s(57), ZN => n281);
   U277 : INV_X1 port map( A => A_s(58), ZN => n282);
   U278 : INV_X1 port map( A => A_s(59), ZN => n283);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT60_i26 is

   port( A_s, A_ns, B : in std_logic_vector (59 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (59 downto 0));

end BOOTHENC_NBIT60_i26;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT60_i26 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, O_59_port, O_58_port, O_57_port, O_56_port, O_55_port,
      O_54_port, O_53_port, O_52_port, O_51_port, O_50_port, O_49_port, 
      O_48_port, O_47_port, O_46_port, O_45_port, O_44_port, O_43_port, 
      O_42_port, O_41_port, O_40_port, O_39_port, O_38_port, O_37_port, 
      O_36_port, O_35_port, O_34_port, O_33_port, O_32_port, O_31_port, 
      O_30_port, O_29_port, O_28_port, O_27_port, O_26_port, O_25_port, 
      O_24_port, O_23_port, O_22_port, O_21_port, O_20_port, O_19_port, 
      O_18_port, O_17_port, O_16_port, O_15_port, O_14_port, O_13_port, 
      O_12_port, O_11_port, O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, 
      O_5_port, O_4_port, O_3_port, O_2_port, O_1_port, n120, n121, n122, n123,
      n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, 
      n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, 
      n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, 
      n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n184, 
      n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, 
      n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, 
      n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, 
      n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, 
      n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, 
      n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, 
      n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, 
      n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, 
      n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, 
      n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, 
      n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, 
      n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, 
      n329, n330 : std_logic;

begin
   O <= ( O_59_port, O_58_port, O_57_port, O_56_port, O_55_port, O_54_port, 
      O_53_port, O_52_port, O_51_port, O_50_port, O_49_port, O_48_port, 
      O_47_port, O_46_port, O_45_port, O_44_port, O_43_port, O_42_port, 
      O_41_port, O_40_port, O_39_port, O_38_port, O_37_port, O_36_port, 
      O_35_port, O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, 
      O_29_port, O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, 
      O_23_port, O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, 
      O_17_port, O_16_port, O_15_port, O_14_port, O_13_port, O_12_port, 
      O_11_port, O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, 
      O_4_port, O_3_port, O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(57), A_s(56), A_s(55), A_s(54), A_s(53), A_s(52), A_s(51), 
      A_s(50), A_s(49), A_s(48), A_s(47), A_s(46), A_s(45), A_s(44), A_s(43), 
      A_s(42), A_s(41), A_s(40), A_s(39), A_s(38), A_s(37), A_s(36), A_s(35), 
      A_s(34), A_s(33), A_s(32), A_s(31), A_s(30), A_s(29), A_s(28), A_s(27), 
      A_s(26), A_s(25), A_s(24), A_s(23), A_s(22), A_s(21), A_s(20), A_s(19), 
      A_s(18), A_s(17), A_s(16), A_s(15), A_s(14), A_s(13), A_s(12), A_s(11), 
      A_s(10), A_s(9), A_s(8), A_s(7), A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), 
      A_s(1), A_s(0), X_Logic0_port, X_Logic0_port );
   A_nso <= ( A_ns(57), A_ns(56), A_ns(55), A_ns(54), A_ns(53), A_ns(52), 
      A_ns(51), A_ns(50), A_ns(49), A_ns(48), A_ns(47), A_ns(46), A_ns(45), 
      A_ns(44), A_ns(43), A_ns(42), A_ns(41), A_ns(40), A_ns(39), A_ns(38), 
      A_ns(37), A_ns(36), A_ns(35), A_ns(34), A_ns(33), A_ns(32), A_ns(31), 
      A_ns(30), A_ns(29), A_ns(28), A_ns(27), A_ns(26), A_ns(25), A_ns(24), 
      A_ns(23), A_ns(22), A_ns(21), A_ns(20), A_ns(19), A_ns(18), A_ns(17), 
      A_ns(16), A_ns(15), A_ns(14), A_ns(13), A_ns(12), A_ns(11), A_ns(10), 
      A_ns(9), A_ns(8), A_ns(7), A_ns(6), A_ns(5), A_ns(4), A_ns(3), A_ns(2), 
      A_ns(1), A_ns(0), X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U241 : XOR2_X1 port map( A => B(25), B => B(26), Z => n182);
   U242 : NAND3_X1 port map( A1 => B(26), A2 => n330, A3 => B(25), ZN => n120);
   U2 : OAI221_X1 port map( B1 => n210, B2 => n327, C1 => n199, C2 => n326, A 
                           => n163, ZN => O_26_port);
   U3 : AOI22_X1 port map( A1 => A_ns(25), A2 => n194, B1 => A_s(25), B2 => 
                           n187, ZN => n163);
   U4 : BUF_X1 port map( A => n191, Z => n194);
   U5 : BUF_X1 port map( A => n184, Z => n187);
   U6 : BUF_X1 port map( A => n191, Z => n195);
   U7 : BUF_X1 port map( A => n184, Z => n188);
   U8 : BUF_X1 port map( A => n192, Z => n196);
   U9 : BUF_X1 port map( A => n185, Z => n189);
   U10 : BUF_X1 port map( A => n192, Z => n197);
   U11 : BUF_X1 port map( A => n185, Z => n190);
   U12 : BUF_X1 port map( A => n191, Z => n193);
   U13 : BUF_X1 port map( A => n184, Z => n186);
   U14 : OAI221_X1 port map( B1 => n207, B2 => n277, C1 => n202, C2 => n243, A 
                           => n127, ZN => O_59_port);
   U15 : AOI22_X1 port map( A1 => A_ns(58), A2 => n197, B1 => A_s(58), B2 => 
                           n190, ZN => n127);
   U16 : OAI221_X1 port map( B1 => n207, B2 => n276, C1 => n201, C2 => n242, A 
                           => n128, ZN => O_58_port);
   U17 : AOI22_X1 port map( A1 => A_ns(57), A2 => n197, B1 => A_s(57), B2 => 
                           n190, ZN => n128);
   U18 : OAI221_X1 port map( B1 => n207, B2 => n275, C1 => n201, C2 => n241, A 
                           => n129, ZN => O_57_port);
   U19 : AOI22_X1 port map( A1 => A_ns(56), A2 => n197, B1 => A_s(56), B2 => 
                           n190, ZN => n129);
   U20 : OAI221_X1 port map( B1 => n207, B2 => n274, C1 => n201, C2 => n240, A 
                           => n130, ZN => O_56_port);
   U21 : AOI22_X1 port map( A1 => A_ns(55), A2 => n197, B1 => A_s(55), B2 => 
                           n190, ZN => n130);
   U22 : OAI221_X1 port map( B1 => n207, B2 => n273, C1 => n201, C2 => n239, A 
                           => n131, ZN => O_55_port);
   U23 : AOI22_X1 port map( A1 => A_ns(54), A2 => n197, B1 => A_s(54), B2 => 
                           n190, ZN => n131);
   U24 : OAI221_X1 port map( B1 => n207, B2 => n272, C1 => n201, C2 => n238, A 
                           => n132, ZN => O_54_port);
   U25 : AOI22_X1 port map( A1 => A_ns(53), A2 => n196, B1 => A_s(53), B2 => 
                           n189, ZN => n132);
   U26 : OAI221_X1 port map( B1 => n207, B2 => n271, C1 => n201, C2 => n237, A 
                           => n133, ZN => O_53_port);
   U27 : AOI22_X1 port map( A1 => A_ns(52), A2 => n196, B1 => A_s(52), B2 => 
                           n189, ZN => n133);
   U28 : OAI221_X1 port map( B1 => n208, B2 => n270, C1 => n201, C2 => n236, A 
                           => n134, ZN => O_52_port);
   U29 : AOI22_X1 port map( A1 => A_ns(51), A2 => n196, B1 => A_s(51), B2 => 
                           n189, ZN => n134);
   U30 : OAI221_X1 port map( B1 => n208, B2 => n269, C1 => n201, C2 => n235, A 
                           => n135, ZN => O_51_port);
   U31 : AOI22_X1 port map( A1 => A_ns(50), A2 => n196, B1 => A_s(50), B2 => 
                           n189, ZN => n135);
   U32 : OAI221_X1 port map( B1 => n208, B2 => n268, C1 => n201, C2 => n234, A 
                           => n136, ZN => O_50_port);
   U33 : AOI22_X1 port map( A1 => A_ns(49), A2 => n196, B1 => A_s(49), B2 => 
                           n189, ZN => n136);
   U34 : OAI221_X1 port map( B1 => n208, B2 => n267, C1 => n201, C2 => n233, A 
                           => n138, ZN => O_49_port);
   U35 : AOI22_X1 port map( A1 => A_ns(48), A2 => n196, B1 => A_s(48), B2 => 
                           n189, ZN => n138);
   U36 : OAI221_X1 port map( B1 => n208, B2 => n266, C1 => n201, C2 => n232, A 
                           => n139, ZN => O_48_port);
   U37 : AOI22_X1 port map( A1 => A_ns(47), A2 => n196, B1 => A_s(47), B2 => 
                           n189, ZN => n139);
   U38 : OAI221_X1 port map( B1 => n208, B2 => n265, C1 => n201, C2 => n231, A 
                           => n140, ZN => O_47_port);
   U39 : AOI22_X1 port map( A1 => A_ns(46), A2 => n196, B1 => A_s(46), B2 => 
                           n189, ZN => n140);
   U40 : OAI221_X1 port map( B1 => n208, B2 => n264, C1 => n200, C2 => n230, A 
                           => n141, ZN => O_46_port);
   U41 : AOI22_X1 port map( A1 => A_ns(45), A2 => n196, B1 => A_s(45), B2 => 
                           n189, ZN => n141);
   U42 : OAI221_X1 port map( B1 => n208, B2 => n263, C1 => n200, C2 => n229, A 
                           => n142, ZN => O_45_port);
   U43 : AOI22_X1 port map( A1 => A_ns(44), A2 => n196, B1 => A_s(44), B2 => 
                           n189, ZN => n142);
   U44 : OAI221_X1 port map( B1 => n208, B2 => n262, C1 => n200, C2 => n228, A 
                           => n143, ZN => O_44_port);
   U45 : AOI22_X1 port map( A1 => A_ns(43), A2 => n196, B1 => A_s(43), B2 => 
                           n189, ZN => n143);
   U46 : OAI221_X1 port map( B1 => n208, B2 => n261, C1 => n200, C2 => n227, A 
                           => n144, ZN => O_43_port);
   U47 : AOI22_X1 port map( A1 => A_ns(42), A2 => n195, B1 => A_s(42), B2 => 
                           n188, ZN => n144);
   U48 : OAI221_X1 port map( B1 => n208, B2 => n260, C1 => n200, C2 => n226, A 
                           => n145, ZN => O_42_port);
   U49 : AOI22_X1 port map( A1 => A_ns(41), A2 => n195, B1 => A_s(41), B2 => 
                           n188, ZN => n145);
   U50 : OAI221_X1 port map( B1 => n209, B2 => n259, C1 => n200, C2 => n225, A 
                           => n146, ZN => O_41_port);
   U51 : AOI22_X1 port map( A1 => A_ns(40), A2 => n195, B1 => A_s(40), B2 => 
                           n188, ZN => n146);
   U52 : OAI221_X1 port map( B1 => n209, B2 => n257, C1 => n200, C2 => n223, A 
                           => n149, ZN => O_39_port);
   U53 : AOI22_X1 port map( A1 => A_ns(38), A2 => n195, B1 => A_s(38), B2 => 
                           n188, ZN => n149);
   U54 : OAI221_X1 port map( B1 => n209, B2 => n258, C1 => n200, C2 => n224, A 
                           => n147, ZN => O_40_port);
   U55 : AOI22_X1 port map( A1 => A_ns(39), A2 => n195, B1 => A_s(39), B2 => 
                           n188, ZN => n147);
   U56 : OAI221_X1 port map( B1 => n209, B2 => n256, C1 => n200, C2 => n222, A 
                           => n150, ZN => O_38_port);
   U57 : AOI22_X1 port map( A1 => A_ns(37), A2 => n195, B1 => A_s(37), B2 => 
                           n188, ZN => n150);
   U58 : OAI221_X1 port map( B1 => n209, B2 => n255, C1 => n200, C2 => n221, A 
                           => n151, ZN => O_37_port);
   U59 : AOI22_X1 port map( A1 => A_ns(36), A2 => n195, B1 => A_s(36), B2 => 
                           n188, ZN => n151);
   U60 : OAI221_X1 port map( B1 => n209, B2 => n254, C1 => n200, C2 => n220, A 
                           => n152, ZN => O_36_port);
   U61 : AOI22_X1 port map( A1 => A_ns(35), A2 => n195, B1 => A_s(35), B2 => 
                           n188, ZN => n152);
   U62 : OAI221_X1 port map( B1 => n209, B2 => n253, C1 => n200, C2 => n219, A 
                           => n153, ZN => O_35_port);
   U63 : AOI22_X1 port map( A1 => A_ns(34), A2 => n195, B1 => A_s(34), B2 => 
                           n188, ZN => n153);
   U64 : OAI221_X1 port map( B1 => n209, B2 => n252, C1 => n199, C2 => n218, A 
                           => n154, ZN => O_34_port);
   U65 : AOI22_X1 port map( A1 => A_ns(33), A2 => n195, B1 => A_s(33), B2 => 
                           n188, ZN => n154);
   U66 : OAI221_X1 port map( B1 => n209, B2 => n251, C1 => n199, C2 => n217, A 
                           => n155, ZN => O_33_port);
   U67 : AOI22_X1 port map( A1 => A_ns(32), A2 => n195, B1 => A_s(32), B2 => 
                           n188, ZN => n155);
   U68 : OAI221_X1 port map( B1 => n209, B2 => n250, C1 => n199, C2 => n216, A 
                           => n156, ZN => O_32_port);
   U69 : AOI22_X1 port map( A1 => A_ns(31), A2 => n194, B1 => A_s(31), B2 => 
                           n187, ZN => n156);
   U70 : OAI221_X1 port map( B1 => n209, B2 => n249, C1 => n199, C2 => n215, A 
                           => n157, ZN => O_31_port);
   U71 : AOI22_X1 port map( A1 => A_ns(30), A2 => n194, B1 => A_s(30), B2 => 
                           n187, ZN => n157);
   U72 : OAI221_X1 port map( B1 => n210, B2 => n247, C1 => n199, C2 => n213, A 
                           => n160, ZN => O_29_port);
   U73 : AOI22_X1 port map( A1 => A_ns(28), A2 => n194, B1 => A_s(28), B2 => 
                           n187, ZN => n160);
   U74 : OAI221_X1 port map( B1 => n210, B2 => n248, C1 => n199, C2 => n214, A 
                           => n158, ZN => O_30_port);
   U75 : AOI22_X1 port map( A1 => A_ns(29), A2 => n194, B1 => A_s(29), B2 => 
                           n187, ZN => n158);
   U76 : BUF_X1 port map( A => n328, Z => n184);
   U77 : BUF_X1 port map( A => n329, Z => n191);
   U78 : BUF_X1 port map( A => n328, Z => n185);
   U79 : BUF_X1 port map( A => n329, Z => n192);
   U80 : OAI221_X1 port map( B1 => n210, B2 => n246, C1 => n199, C2 => n212, A 
                           => n161, ZN => O_28_port);
   U81 : AOI22_X1 port map( A1 => A_ns(27), A2 => n194, B1 => A_s(27), B2 => 
                           n187, ZN => n161);
   U82 : BUF_X1 port map( A => n206, Z => n210);
   U83 : BUF_X1 port map( A => n204, Z => n199);
   U84 : INV_X1 port map( A => n170, ZN => n328);
   U85 : INV_X1 port map( A => n171, ZN => n329);
   U86 : BUF_X1 port map( A => n205, Z => n209);
   U87 : BUF_X1 port map( A => n203, Z => n200);
   U88 : BUF_X1 port map( A => n205, Z => n208);
   U89 : BUF_X1 port map( A => n203, Z => n201);
   U90 : BUF_X1 port map( A => n205, Z => n207);
   U91 : BUF_X1 port map( A => n203, Z => n202);
   U92 : BUF_X1 port map( A => n204, Z => n198);
   U93 : BUF_X1 port map( A => n206, Z => n211);
   U94 : OAI221_X1 port map( B1 => n210, B2 => n245, C1 => n199, C2 => n244, A 
                           => n162, ZN => O_27_port);
   U95 : AOI22_X1 port map( A1 => A_ns(26), A2 => n194, B1 => A_s(26), B2 => 
                           n187, ZN => n162);
   U96 : NAND2_X1 port map( A1 => n182, A2 => n330, ZN => n170);
   U97 : NAND2_X1 port map( A1 => n182, A2 => n170, ZN => n171);
   U98 : BUF_X1 port map( A => n120, Z => n206);
   U99 : BUF_X1 port map( A => n121, Z => n204);
   U100 : BUF_X1 port map( A => n120, Z => n205);
   U101 : BUF_X1 port map( A => n121, Z => n203);
   U102 : INV_X1 port map( A => A_s(24), ZN => n327);
   U103 : INV_X1 port map( A => A_ns(24), ZN => n326);
   U104 : OAI221_X1 port map( B1 => n211, B2 => n313, C1 => n198, C2 => n311, A
                           => n172, ZN => O_19_port);
   U105 : INV_X1 port map( A => A_s(17), ZN => n313);
   U106 : INV_X1 port map( A => A_ns(17), ZN => n311);
   U107 : OAI221_X1 port map( B1 => n210, B2 => n316, C1 => n198, C2 => n314, A
                           => n169, ZN => O_20_port);
   U108 : INV_X1 port map( A => A_s(18), ZN => n316);
   U109 : INV_X1 port map( A => A_ns(18), ZN => n314);
   U110 : OAI221_X1 port map( B1 => n210, B2 => n317, C1 => n198, C2 => n315, A
                           => n168, ZN => O_21_port);
   U111 : INV_X1 port map( A => A_s(19), ZN => n317);
   U112 : INV_X1 port map( A => A_ns(19), ZN => n315);
   U113 : OAI221_X1 port map( B1 => n210, B2 => n320, C1 => n198, C2 => n318, A
                           => n167, ZN => O_22_port);
   U114 : INV_X1 port map( A => A_s(20), ZN => n320);
   U115 : INV_X1 port map( A => A_ns(20), ZN => n318);
   U116 : OAI221_X1 port map( B1 => n210, B2 => n321, C1 => n199, C2 => n319, A
                           => n166, ZN => O_23_port);
   U117 : INV_X1 port map( A => A_s(21), ZN => n321);
   U118 : INV_X1 port map( A => A_ns(21), ZN => n319);
   U119 : OAI221_X1 port map( B1 => n210, B2 => n324, C1 => n199, C2 => n322, A
                           => n165, ZN => O_24_port);
   U120 : INV_X1 port map( A => A_s(22), ZN => n324);
   U121 : INV_X1 port map( A => A_ns(22), ZN => n322);
   U122 : OAI221_X1 port map( B1 => n210, B2 => n325, C1 => n199, C2 => n323, A
                           => n164, ZN => O_25_port);
   U123 : INV_X1 port map( A => A_s(23), ZN => n325);
   U124 : INV_X1 port map( A => A_ns(23), ZN => n323);
   U125 : INV_X1 port map( A => B(27), ZN => n330);
   U126 : OR3_X1 port map( A1 => B(25), A2 => B(26), A3 => n330, ZN => n121);
   U127 : OAI221_X1 port map( B1 => n207, B2 => n292, C1 => n202, C2 => n290, A
                           => n123, ZN => O_8_port);
   U128 : INV_X1 port map( A => A_s(6), ZN => n292);
   U129 : INV_X1 port map( A => A_ns(6), ZN => n290);
   U130 : OAI221_X1 port map( B1 => n207, B2 => n293, C1 => n202, C2 => n291, A
                           => n122, ZN => O_9_port);
   U131 : INV_X1 port map( A => A_s(7), ZN => n293);
   U132 : INV_X1 port map( A => A_ns(7), ZN => n291);
   U133 : OAI221_X1 port map( B1 => n296, B2 => n211, C1 => n294, C2 => n198, A
                           => n181, ZN => O_10_port);
   U134 : INV_X1 port map( A => A_ns(8), ZN => n294);
   U135 : INV_X1 port map( A => A_s(8), ZN => n296);
   U136 : OAI221_X1 port map( B1 => n211, B2 => n297, C1 => n198, C2 => n295, A
                           => n180, ZN => O_11_port);
   U137 : INV_X1 port map( A => A_s(9), ZN => n297);
   U138 : INV_X1 port map( A => A_ns(9), ZN => n295);
   U139 : OAI221_X1 port map( B1 => n211, B2 => n300, C1 => n198, C2 => n298, A
                           => n179, ZN => O_12_port);
   U140 : INV_X1 port map( A => A_s(10), ZN => n300);
   U141 : INV_X1 port map( A => A_ns(10), ZN => n298);
   U142 : OAI221_X1 port map( B1 => n211, B2 => n301, C1 => n198, C2 => n299, A
                           => n178, ZN => O_13_port);
   U143 : INV_X1 port map( A => A_s(11), ZN => n301);
   U144 : INV_X1 port map( A => A_ns(11), ZN => n299);
   U145 : OAI221_X1 port map( B1 => n211, B2 => n304, C1 => n198, C2 => n302, A
                           => n177, ZN => O_14_port);
   U146 : INV_X1 port map( A => A_s(12), ZN => n304);
   U147 : INV_X1 port map( A => A_ns(12), ZN => n302);
   U148 : OAI221_X1 port map( B1 => n211, B2 => n305, C1 => n198, C2 => n303, A
                           => n176, ZN => O_15_port);
   U149 : INV_X1 port map( A => A_s(13), ZN => n305);
   U150 : INV_X1 port map( A => A_ns(13), ZN => n303);
   U151 : OAI221_X1 port map( B1 => n211, B2 => n308, C1 => n198, C2 => n306, A
                           => n175, ZN => O_16_port);
   U152 : INV_X1 port map( A => A_s(14), ZN => n308);
   U153 : INV_X1 port map( A => A_ns(14), ZN => n306);
   U154 : OAI221_X1 port map( B1 => n211, B2 => n309, C1 => n198, C2 => n307, A
                           => n174, ZN => O_17_port);
   U155 : INV_X1 port map( A => A_s(15), ZN => n309);
   U156 : INV_X1 port map( A => A_ns(15), ZN => n307);
   U157 : OAI221_X1 port map( B1 => n211, B2 => n312, C1 => n198, C2 => n310, A
                           => n173, ZN => O_18_port);
   U158 : INV_X1 port map( A => A_s(16), ZN => n312);
   U159 : INV_X1 port map( A => A_ns(16), ZN => n310);
   U160 : OAI22_X1 port map( A1 => n170, A2 => n280, B1 => n171, B2 => n278, ZN
                           => O_1_port);
   U161 : OAI221_X1 port map( B1 => n210, B2 => n280, C1 => n199, C2 => n278, A
                           => n159, ZN => O_2_port);
   U162 : AOI22_X1 port map( A1 => A_ns(1), A2 => n194, B1 => A_s(1), B2 => 
                           n187, ZN => n159);
   U163 : OAI221_X1 port map( B1 => n209, B2 => n281, C1 => n200, C2 => n279, A
                           => n148, ZN => O_3_port);
   U164 : INV_X1 port map( A => A_s(1), ZN => n281);
   U165 : INV_X1 port map( A => A_ns(1), ZN => n279);
   U166 : OAI221_X1 port map( B1 => n208, B2 => n284, C1 => n201, C2 => n282, A
                           => n137, ZN => O_4_port);
   U167 : INV_X1 port map( A => A_s(2), ZN => n284);
   U168 : INV_X1 port map( A => A_ns(2), ZN => n282);
   U169 : OAI221_X1 port map( B1 => n207, B2 => n285, C1 => n202, C2 => n283, A
                           => n126, ZN => O_5_port);
   U170 : INV_X1 port map( A => A_s(3), ZN => n285);
   U171 : INV_X1 port map( A => A_ns(3), ZN => n283);
   U172 : OAI221_X1 port map( B1 => n207, B2 => n288, C1 => n202, C2 => n286, A
                           => n125, ZN => O_6_port);
   U173 : INV_X1 port map( A => A_s(4), ZN => n288);
   U174 : INV_X1 port map( A => A_ns(4), ZN => n286);
   U175 : OAI221_X1 port map( B1 => n207, B2 => n289, C1 => n202, C2 => n287, A
                           => n124, ZN => O_7_port);
   U176 : INV_X1 port map( A => A_s(5), ZN => n289);
   U177 : INV_X1 port map( A => A_ns(5), ZN => n287);
   U178 : INV_X1 port map( A => A_ns(0), ZN => n278);
   U179 : INV_X1 port map( A => A_s(0), ZN => n280);
   U180 : AOI22_X1 port map( A1 => A_ns(2), A2 => n195, B1 => A_s(2), B2 => 
                           n188, ZN => n148);
   U181 : AOI22_X1 port map( A1 => A_ns(3), A2 => n196, B1 => A_s(3), B2 => 
                           n189, ZN => n137);
   U182 : AOI22_X1 port map( A1 => A_ns(4), A2 => n197, B1 => A_s(4), B2 => 
                           n190, ZN => n126);
   U183 : AOI22_X1 port map( A1 => A_ns(5), A2 => n197, B1 => A_s(5), B2 => 
                           n190, ZN => n125);
   U184 : AOI22_X1 port map( A1 => A_ns(6), A2 => n197, B1 => A_s(6), B2 => 
                           n190, ZN => n124);
   U185 : AOI22_X1 port map( A1 => A_ns(7), A2 => n197, B1 => A_s(7), B2 => 
                           n190, ZN => n123);
   U186 : AOI22_X1 port map( A1 => A_ns(8), A2 => n197, B1 => A_s(8), B2 => 
                           n190, ZN => n122);
   U187 : AOI22_X1 port map( A1 => A_ns(9), A2 => n193, B1 => A_s(9), B2 => 
                           n186, ZN => n181);
   U188 : AOI22_X1 port map( A1 => A_ns(10), A2 => n193, B1 => A_s(10), B2 => 
                           n186, ZN => n180);
   U189 : AOI22_X1 port map( A1 => A_ns(11), A2 => n193, B1 => A_s(11), B2 => 
                           n186, ZN => n179);
   U190 : AOI22_X1 port map( A1 => A_ns(12), A2 => n193, B1 => A_s(12), B2 => 
                           n186, ZN => n178);
   U191 : AOI22_X1 port map( A1 => A_ns(13), A2 => n193, B1 => A_s(13), B2 => 
                           n186, ZN => n177);
   U192 : AOI22_X1 port map( A1 => A_ns(14), A2 => n193, B1 => A_s(14), B2 => 
                           n186, ZN => n176);
   U193 : AOI22_X1 port map( A1 => A_ns(15), A2 => n193, B1 => A_s(15), B2 => 
                           n186, ZN => n175);
   U194 : AOI22_X1 port map( A1 => A_ns(16), A2 => n193, B1 => A_s(16), B2 => 
                           n186, ZN => n174);
   U195 : AOI22_X1 port map( A1 => A_ns(17), A2 => n193, B1 => A_s(17), B2 => 
                           n186, ZN => n173);
   U196 : AOI22_X1 port map( A1 => A_ns(18), A2 => n193, B1 => A_s(18), B2 => 
                           n186, ZN => n172);
   U197 : AOI22_X1 port map( A1 => A_ns(19), A2 => n193, B1 => A_s(19), B2 => 
                           n186, ZN => n169);
   U198 : AOI22_X1 port map( A1 => A_ns(20), A2 => n193, B1 => A_s(20), B2 => 
                           n186, ZN => n168);
   U199 : AOI22_X1 port map( A1 => A_ns(21), A2 => n194, B1 => A_s(21), B2 => 
                           n187, ZN => n167);
   U200 : AOI22_X1 port map( A1 => A_ns(22), A2 => n194, B1 => A_s(22), B2 => 
                           n187, ZN => n166);
   U201 : AOI22_X1 port map( A1 => A_ns(23), A2 => n194, B1 => A_s(23), B2 => 
                           n187, ZN => n165);
   U202 : AOI22_X1 port map( A1 => A_ns(24), A2 => n194, B1 => A_s(24), B2 => 
                           n187, ZN => n164);
   U203 : INV_X1 port map( A => A_ns(26), ZN => n212);
   U204 : INV_X1 port map( A => A_ns(27), ZN => n213);
   U205 : INV_X1 port map( A => A_ns(28), ZN => n214);
   U206 : INV_X1 port map( A => A_ns(29), ZN => n215);
   U207 : INV_X1 port map( A => A_ns(30), ZN => n216);
   U208 : INV_X1 port map( A => A_ns(31), ZN => n217);
   U209 : INV_X1 port map( A => A_ns(32), ZN => n218);
   U210 : INV_X1 port map( A => A_ns(33), ZN => n219);
   U211 : INV_X1 port map( A => A_ns(34), ZN => n220);
   U212 : INV_X1 port map( A => A_ns(35), ZN => n221);
   U213 : INV_X1 port map( A => A_ns(36), ZN => n222);
   U214 : INV_X1 port map( A => A_ns(37), ZN => n223);
   U215 : INV_X1 port map( A => A_ns(38), ZN => n224);
   U216 : INV_X1 port map( A => A_ns(39), ZN => n225);
   U217 : INV_X1 port map( A => A_ns(40), ZN => n226);
   U218 : INV_X1 port map( A => A_ns(41), ZN => n227);
   U219 : INV_X1 port map( A => A_ns(42), ZN => n228);
   U220 : INV_X1 port map( A => A_ns(43), ZN => n229);
   U221 : INV_X1 port map( A => A_ns(44), ZN => n230);
   U222 : INV_X1 port map( A => A_ns(45), ZN => n231);
   U223 : INV_X1 port map( A => A_ns(46), ZN => n232);
   U224 : INV_X1 port map( A => A_ns(47), ZN => n233);
   U225 : INV_X1 port map( A => A_ns(48), ZN => n234);
   U226 : INV_X1 port map( A => A_ns(49), ZN => n235);
   U227 : INV_X1 port map( A => A_ns(50), ZN => n236);
   U228 : INV_X1 port map( A => A_ns(51), ZN => n237);
   U229 : INV_X1 port map( A => A_ns(52), ZN => n238);
   U230 : INV_X1 port map( A => A_ns(53), ZN => n239);
   U231 : INV_X1 port map( A => A_ns(54), ZN => n240);
   U232 : INV_X1 port map( A => A_ns(55), ZN => n241);
   U233 : INV_X1 port map( A => A_ns(56), ZN => n242);
   U234 : INV_X1 port map( A => A_ns(57), ZN => n243);
   U235 : INV_X1 port map( A => A_ns(25), ZN => n244);
   U236 : INV_X1 port map( A => A_s(25), ZN => n245);
   U237 : INV_X1 port map( A => A_s(26), ZN => n246);
   U238 : INV_X1 port map( A => A_s(27), ZN => n247);
   U239 : INV_X1 port map( A => A_s(28), ZN => n248);
   U240 : INV_X1 port map( A => A_s(29), ZN => n249);
   U243 : INV_X1 port map( A => A_s(30), ZN => n250);
   U244 : INV_X1 port map( A => A_s(31), ZN => n251);
   U245 : INV_X1 port map( A => A_s(32), ZN => n252);
   U246 : INV_X1 port map( A => A_s(33), ZN => n253);
   U247 : INV_X1 port map( A => A_s(34), ZN => n254);
   U248 : INV_X1 port map( A => A_s(35), ZN => n255);
   U249 : INV_X1 port map( A => A_s(36), ZN => n256);
   U250 : INV_X1 port map( A => A_s(37), ZN => n257);
   U251 : INV_X1 port map( A => A_s(38), ZN => n258);
   U252 : INV_X1 port map( A => A_s(39), ZN => n259);
   U253 : INV_X1 port map( A => A_s(40), ZN => n260);
   U254 : INV_X1 port map( A => A_s(41), ZN => n261);
   U255 : INV_X1 port map( A => A_s(42), ZN => n262);
   U256 : INV_X1 port map( A => A_s(43), ZN => n263);
   U257 : INV_X1 port map( A => A_s(44), ZN => n264);
   U258 : INV_X1 port map( A => A_s(45), ZN => n265);
   U259 : INV_X1 port map( A => A_s(46), ZN => n266);
   U260 : INV_X1 port map( A => A_s(47), ZN => n267);
   U261 : INV_X1 port map( A => A_s(48), ZN => n268);
   U262 : INV_X1 port map( A => A_s(49), ZN => n269);
   U263 : INV_X1 port map( A => A_s(50), ZN => n270);
   U264 : INV_X1 port map( A => A_s(51), ZN => n271);
   U265 : INV_X1 port map( A => A_s(52), ZN => n272);
   U266 : INV_X1 port map( A => A_s(53), ZN => n273);
   U267 : INV_X1 port map( A => A_s(54), ZN => n274);
   U268 : INV_X1 port map( A => A_s(55), ZN => n275);
   U269 : INV_X1 port map( A => A_s(56), ZN => n276);
   U270 : INV_X1 port map( A => A_s(57), ZN => n277);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT58_i24 is

   port( A_s, A_ns, B : in std_logic_vector (57 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (57 downto 0));

end BOOTHENC_NBIT58_i24;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT58_i24 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, O_57_port, O_56_port, O_55_port, O_54_port, O_53_port,
      O_52_port, O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, 
      O_46_port, O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, 
      O_40_port, O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, 
      O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, 
      O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, 
      O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, 
      O_16_port, O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, 
      O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, 
      O_3_port, O_2_port, O_1_port, n116, n117, n118, n119, n120, n121, n122, 
      n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, 
      n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n178, n179, n180, n181, n182, n183, 
      n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, A_nso_48_port, n229, 
      A_nso_49_port, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240
      , n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
      n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, 
      n265, n266, n267, n268, n269, n270, n271, n272, A_so_57_port, n274, n275,
      n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, 
      n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, 
      n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, 
      n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323 : 
      std_logic;

begin
   O <= ( O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, O_52_port, 
      O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, O_46_port, 
      O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, O_40_port, 
      O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, 
      O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, 
      O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, 
      O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, O_16_port, 
      O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, O_10_port, 
      O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, O_3_port, 
      O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_so_57_port, A_s(54), A_s(53), A_s(52), A_s(51), A_s(50), A_s(49)
      , A_s(48), A_s(47), A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41),
      A_s(40), A_s(39), A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), 
      A_s(32), A_s(31), A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), 
      A_s(24), A_s(23), A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), 
      A_s(16), A_s(15), A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), 
      A_s(8), A_s(7), A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), 
      X_Logic0_port, X_Logic0_port );
   A_nso <= ( A_ns(55), A_ns(54), A_ns(53), A_ns(52), A_ns(51), A_ns(50), 
      A_ns(49), A_ns(48), A_nso_49_port, A_nso_48_port, A_ns(45), A_ns(44), 
      A_ns(43), A_ns(42), A_ns(41), A_ns(40), A_ns(39), A_ns(38), A_ns(37), 
      A_ns(36), A_ns(35), A_ns(34), A_ns(33), A_ns(32), A_ns(31), A_ns(30), 
      A_ns(29), A_ns(28), A_ns(27), A_ns(26), A_ns(25), A_ns(24), A_ns(23), 
      A_ns(22), A_ns(21), A_ns(20), A_ns(19), A_ns(18), A_ns(17), A_ns(16), 
      A_ns(15), A_ns(14), A_ns(13), A_ns(12), A_ns(11), A_ns(10), A_ns(9), 
      A_ns(8), A_ns(7), A_ns(6), A_ns(5), A_ns(4), A_ns(3), A_ns(2), A_ns(1), 
      A_ns(0), X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U233 : XOR2_X1 port map( A => B(23), B => B(24), Z => n176);
   U234 : NAND3_X1 port map( A1 => B(24), A2 => n323, A3 => B(23), ZN => n116);
   U2 : OAI221_X1 port map( B1 => n201, B2 => n269, C1 => n195, C2 => n235, A 
                           => n127, ZN => O_53_port);
   U3 : OAI221_X1 port map( B1 => n201, B2 => n270, C1 => n195, C2 => n236, A 
                           => n126, ZN => O_54_port);
   U4 : OAI221_X1 port map( B1 => n201, B2 => n271, C1 => n195, C2 => n237, A 
                           => n125, ZN => O_55_port);
   U5 : AOI22_X1 port map( A1 => A_ns(23), A2 => n188, B1 => A_s(23), B2 => 
                           n181, ZN => n159);
   U6 : BUF_X1 port map( A => n185, Z => n188);
   U7 : BUF_X1 port map( A => n185, Z => n189);
   U8 : BUF_X1 port map( A => n178, Z => n181);
   U9 : BUF_X1 port map( A => n186, Z => n190);
   U10 : BUF_X1 port map( A => n178, Z => n182);
   U11 : BUF_X1 port map( A => n179, Z => n183);
   U12 : BUF_X1 port map( A => n186, Z => n191);
   U13 : BUF_X1 port map( A => n179, Z => n184);
   U14 : BUF_X1 port map( A => n185, Z => n187);
   U15 : BUF_X1 port map( A => n178, Z => n180);
   U16 : OAI221_X1 port map( B1 => n201, B2 => n274, C1 => n195, C2 => n239, A 
                           => n123, ZN => O_57_port);
   U17 : AOI22_X1 port map( A1 => A_ns(56), A2 => n191, B1 => A_s(56), B2 => 
                           n184, ZN => n123);
   U18 : AOI22_X1 port map( A1 => A_ns(53), A2 => n190, B1 => A_s(53), B2 => 
                           n183, ZN => n126);
   U19 : AOI22_X1 port map( A1 => A_ns(52), A2 => n190, B1 => A_s(52), B2 => 
                           n183, ZN => n127);
   U20 : OAI221_X1 port map( B1 => n201, B2 => n268, C1 => n195, C2 => n234, A 
                           => n128, ZN => O_52_port);
   U21 : AOI22_X1 port map( A1 => A_ns(51), A2 => n190, B1 => A_s(51), B2 => 
                           n183, ZN => n128);
   U22 : OAI221_X1 port map( B1 => n202, B2 => n262, C1 => n194, C2 => n226, A 
                           => n135, ZN => O_46_port);
   U23 : AOI22_X1 port map( A1 => A_ns(45), A2 => n190, B1 => A_s(45), B2 => 
                           n183, ZN => n135);
   U24 : OAI221_X1 port map( B1 => n203, B2 => n253, C1 => n194, C2 => n217, A 
                           => n145, ZN => O_37_port);
   U25 : AOI22_X1 port map( A1 => A_ns(36), A2 => n189, B1 => A_s(36), B2 => 
                           n182, ZN => n145);
   U26 : OAI221_X1 port map( B1 => n203, B2 => n252, C1 => n194, C2 => n216, A 
                           => n146, ZN => O_36_port);
   U27 : AOI22_X1 port map( A1 => A_ns(35), A2 => n189, B1 => A_s(35), B2 => 
                           n182, ZN => n146);
   U28 : OAI221_X1 port map( B1 => n203, B2 => n251, C1 => n194, C2 => n215, A 
                           => n147, ZN => O_35_port);
   U29 : AOI22_X1 port map( A1 => A_ns(34), A2 => n189, B1 => A_s(34), B2 => 
                           n182, ZN => n147);
   U30 : OAI221_X1 port map( B1 => n203, B2 => n250, C1 => n193, C2 => n214, A 
                           => n148, ZN => O_34_port);
   U31 : AOI22_X1 port map( A1 => A_ns(33), A2 => n189, B1 => A_s(33), B2 => 
                           n182, ZN => n148);
   U32 : OAI221_X1 port map( B1 => n203, B2 => n249, C1 => n193, C2 => n213, A 
                           => n149, ZN => O_33_port);
   U33 : AOI22_X1 port map( A1 => A_ns(32), A2 => n189, B1 => A_s(32), B2 => 
                           n182, ZN => n149);
   U34 : OAI221_X1 port map( B1 => n203, B2 => n248, C1 => n193, C2 => n212, A 
                           => n150, ZN => O_32_port);
   U35 : AOI22_X1 port map( A1 => A_ns(31), A2 => n188, B1 => A_s(31), B2 => 
                           n181, ZN => n150);
   U36 : OAI221_X1 port map( B1 => n203, B2 => n247, C1 => n193, C2 => n211, A 
                           => n151, ZN => O_31_port);
   U37 : AOI22_X1 port map( A1 => A_ns(30), A2 => n188, B1 => A_s(30), B2 => 
                           n181, ZN => n151);
   U38 : OAI221_X1 port map( B1 => n203, B2 => n246, C1 => n193, C2 => n210, A 
                           => n152, ZN => O_30_port);
   U39 : AOI22_X1 port map( A1 => A_ns(29), A2 => n188, B1 => A_s(29), B2 => 
                           n181, ZN => n152);
   U40 : OAI221_X1 port map( B1 => n204, B2 => n245, C1 => n193, C2 => n209, A 
                           => n154, ZN => O_29_port);
   U41 : AOI22_X1 port map( A1 => A_ns(28), A2 => n188, B1 => A_s(28), B2 => 
                           n181, ZN => n154);
   U42 : OAI221_X1 port map( B1 => n204, B2 => n244, C1 => n193, C2 => n208, A 
                           => n155, ZN => O_28_port);
   U43 : AOI22_X1 port map( A1 => A_ns(27), A2 => n188, B1 => A_s(27), B2 => 
                           n181, ZN => n155);
   U44 : OAI221_X1 port map( B1 => n204, B2 => n243, C1 => n193, C2 => n207, A 
                           => n156, ZN => O_27_port);
   U45 : AOI22_X1 port map( A1 => A_ns(26), A2 => n188, B1 => A_s(26), B2 => 
                           n181, ZN => n156);
   U46 : OAI221_X1 port map( B1 => n201, B2 => n272, C1 => n195, C2 => n238, A 
                           => n124, ZN => O_56_port);
   U47 : AOI22_X1 port map( A1 => A_ns(55), A2 => n191, B1 => A_so_57_port, B2 
                           => n184, ZN => n124);
   U48 : OAI221_X1 port map( B1 => n201, B2 => n267, C1 => n195, C2 => n233, A 
                           => n129, ZN => O_51_port);
   U49 : AOI22_X1 port map( A1 => A_ns(50), A2 => n190, B1 => A_s(50), B2 => 
                           n183, ZN => n129);
   U50 : OAI221_X1 port map( B1 => n202, B2 => n266, C1 => n195, C2 => n232, A 
                           => n130, ZN => O_50_port);
   U51 : AOI22_X1 port map( A1 => A_ns(49), A2 => n190, B1 => A_s(49), B2 => 
                           n183, ZN => n130);
   U52 : OAI221_X1 port map( B1 => n202, B2 => n265, C1 => n195, C2 => n231, A 
                           => n132, ZN => O_49_port);
   U53 : AOI22_X1 port map( A1 => A_ns(48), A2 => n190, B1 => A_s(48), B2 => 
                           n183, ZN => n132);
   U54 : OAI221_X1 port map( B1 => n202, B2 => n264, C1 => n195, C2 => n229, A 
                           => n133, ZN => O_48_port);
   U55 : AOI22_X1 port map( A1 => A_nso_49_port, A2 => n190, B1 => A_s(47), B2 
                           => n183, ZN => n133);
   U56 : OAI221_X1 port map( B1 => n202, B2 => n263, C1 => n195, C2 => n227, A 
                           => n134, ZN => O_47_port);
   U57 : AOI22_X1 port map( A1 => A_nso_48_port, A2 => n190, B1 => A_s(46), B2 
                           => n183, ZN => n134);
   U58 : OAI221_X1 port map( B1 => n202, B2 => n261, C1 => n194, C2 => n225, A 
                           => n136, ZN => O_45_port);
   U59 : AOI22_X1 port map( A1 => A_ns(44), A2 => n190, B1 => A_s(44), B2 => 
                           n183, ZN => n136);
   U60 : OAI221_X1 port map( B1 => n202, B2 => n260, C1 => n194, C2 => n224, A 
                           => n137, ZN => O_44_port);
   U61 : AOI22_X1 port map( A1 => A_ns(43), A2 => n190, B1 => A_s(43), B2 => 
                           n183, ZN => n137);
   U62 : OAI221_X1 port map( B1 => n202, B2 => n259, C1 => n194, C2 => n223, A 
                           => n138, ZN => O_43_port);
   U63 : AOI22_X1 port map( A1 => A_ns(42), A2 => n189, B1 => A_s(42), B2 => 
                           n182, ZN => n138);
   U64 : OAI221_X1 port map( B1 => n202, B2 => n258, C1 => n194, C2 => n222, A 
                           => n139, ZN => O_42_port);
   U65 : AOI22_X1 port map( A1 => A_ns(41), A2 => n189, B1 => A_s(41), B2 => 
                           n182, ZN => n139);
   U66 : OAI221_X1 port map( B1 => n202, B2 => n257, C1 => n194, C2 => n221, A 
                           => n140, ZN => O_41_port);
   U67 : AOI22_X1 port map( A1 => A_ns(40), A2 => n189, B1 => A_s(40), B2 => 
                           n182, ZN => n140);
   U68 : OAI221_X1 port map( B1 => n203, B2 => n255, C1 => n194, C2 => n219, A 
                           => n143, ZN => O_39_port);
   U69 : AOI22_X1 port map( A1 => A_ns(38), A2 => n189, B1 => A_s(38), B2 => 
                           n182, ZN => n143);
   U70 : OAI221_X1 port map( B1 => n202, B2 => n256, C1 => n194, C2 => n220, A 
                           => n141, ZN => O_40_port);
   U71 : AOI22_X1 port map( A1 => A_ns(39), A2 => n189, B1 => A_s(39), B2 => 
                           n182, ZN => n141);
   U72 : OAI221_X1 port map( B1 => n203, B2 => n254, C1 => n194, C2 => n218, A 
                           => n144, ZN => O_38_port);
   U73 : AOI22_X1 port map( A1 => A_ns(37), A2 => n189, B1 => A_s(37), B2 => 
                           n182, ZN => n144);
   U74 : BUF_X1 port map( A => n321, Z => n178);
   U75 : BUF_X1 port map( A => n322, Z => n185);
   U76 : BUF_X1 port map( A => n322, Z => n186);
   U77 : BUF_X1 port map( A => n321, Z => n179);
   U78 : AOI22_X1 port map( A1 => A_ns(54), A2 => n191, B1 => A_s(54), B2 => 
                           n184, ZN => n125);
   U79 : OAI221_X1 port map( B1 => n204, B2 => n242, C1 => n193, C2 => n206, A 
                           => n157, ZN => O_26_port);
   U80 : AOI22_X1 port map( A1 => A_ns(25), A2 => n188, B1 => A_s(25), B2 => 
                           n181, ZN => n157);
   U81 : BUF_X1 port map( A => n199, Z => n203);
   U82 : BUF_X1 port map( A => n200, Z => n204);
   U83 : BUF_X1 port map( A => n198, Z => n193);
   U84 : INV_X1 port map( A => n164, ZN => n321);
   U85 : INV_X1 port map( A => n165, ZN => n322);
   U86 : BUF_X1 port map( A => n199, Z => n202);
   U87 : BUF_X1 port map( A => n197, Z => n194);
   U88 : BUF_X1 port map( A => n199, Z => n201);
   U89 : BUF_X1 port map( A => n197, Z => n195);
   U90 : BUF_X1 port map( A => n198, Z => n192);
   U91 : BUF_X1 port map( A => n200, Z => n205);
   U92 : BUF_X1 port map( A => n197, Z => n196);
   U93 : OAI221_X1 port map( B1 => n204, B2 => n241, C1 => n193, C2 => n240, A 
                           => n158, ZN => O_25_port);
   U94 : AOI22_X1 port map( A1 => A_ns(24), A2 => n188, B1 => A_s(24), B2 => 
                           n181, ZN => n158);
   U95 : NAND2_X1 port map( A1 => n176, A2 => n323, ZN => n164);
   U96 : NAND2_X1 port map( A1 => n176, A2 => n164, ZN => n165);
   U97 : BUF_X1 port map( A => n116, Z => n199);
   U98 : BUF_X1 port map( A => n117, Z => n198);
   U99 : BUF_X1 port map( A => n116, Z => n200);
   U100 : BUF_X1 port map( A => n117, Z => n197);
   U101 : OAI221_X1 port map( B1 => n204, B2 => n320, C1 => n193, C2 => n319, A
                           => n159, ZN => O_24_port);
   U102 : INV_X1 port map( A => A_s(22), ZN => n320);
   U103 : INV_X1 port map( A => A_ns(22), ZN => n319);
   U104 : OAI221_X1 port map( B1 => n204, B2 => n310, C1 => n192, C2 => n308, A
                           => n166, ZN => O_19_port);
   U105 : INV_X1 port map( A => A_s(17), ZN => n310);
   U106 : INV_X1 port map( A => A_ns(17), ZN => n308);
   U107 : OAI221_X1 port map( B1 => n204, B2 => n313, C1 => n192, C2 => n311, A
                           => n163, ZN => O_20_port);
   U108 : INV_X1 port map( A => A_s(18), ZN => n313);
   U109 : INV_X1 port map( A => A_ns(18), ZN => n311);
   U110 : OAI221_X1 port map( B1 => n204, B2 => n314, C1 => n192, C2 => n312, A
                           => n162, ZN => O_21_port);
   U111 : INV_X1 port map( A => A_s(19), ZN => n314);
   U112 : INV_X1 port map( A => A_ns(19), ZN => n312);
   U113 : OAI221_X1 port map( B1 => n204, B2 => n317, C1 => n192, C2 => n315, A
                           => n161, ZN => O_22_port);
   U114 : INV_X1 port map( A => A_s(20), ZN => n317);
   U115 : INV_X1 port map( A => A_ns(20), ZN => n315);
   U116 : OAI221_X1 port map( B1 => n204, B2 => n318, C1 => n193, C2 => n316, A
                           => n160, ZN => O_23_port);
   U117 : INV_X1 port map( A => A_s(21), ZN => n318);
   U118 : INV_X1 port map( A => A_ns(21), ZN => n316);
   U119 : INV_X1 port map( A => B(25), ZN => n323);
   U120 : OR3_X1 port map( A1 => B(23), A2 => B(24), A3 => n323, ZN => n117);
   U121 : OAI221_X1 port map( B1 => n201, B2 => n289, C1 => n196, C2 => n287, A
                           => n119, ZN => O_8_port);
   U122 : INV_X1 port map( A => A_s(6), ZN => n289);
   U123 : INV_X1 port map( A => A_ns(6), ZN => n287);
   U124 : OAI221_X1 port map( B1 => n201, B2 => n290, C1 => n196, C2 => n288, A
                           => n118, ZN => O_9_port);
   U125 : INV_X1 port map( A => A_s(7), ZN => n290);
   U126 : INV_X1 port map( A => A_ns(7), ZN => n288);
   U127 : OAI221_X1 port map( B1 => n293, B2 => n205, C1 => n291, C2 => n192, A
                           => n175, ZN => O_10_port);
   U128 : INV_X1 port map( A => A_ns(8), ZN => n291);
   U129 : INV_X1 port map( A => A_s(8), ZN => n293);
   U130 : OAI221_X1 port map( B1 => n205, B2 => n294, C1 => n192, C2 => n292, A
                           => n174, ZN => O_11_port);
   U131 : INV_X1 port map( A => A_s(9), ZN => n294);
   U132 : INV_X1 port map( A => A_ns(9), ZN => n292);
   U133 : OAI221_X1 port map( B1 => n205, B2 => n297, C1 => n192, C2 => n295, A
                           => n173, ZN => O_12_port);
   U134 : INV_X1 port map( A => A_s(10), ZN => n297);
   U135 : INV_X1 port map( A => A_ns(10), ZN => n295);
   U136 : OAI221_X1 port map( B1 => n205, B2 => n298, C1 => n192, C2 => n296, A
                           => n172, ZN => O_13_port);
   U137 : INV_X1 port map( A => A_s(11), ZN => n298);
   U138 : INV_X1 port map( A => A_ns(11), ZN => n296);
   U139 : OAI221_X1 port map( B1 => n205, B2 => n301, C1 => n192, C2 => n299, A
                           => n171, ZN => O_14_port);
   U140 : INV_X1 port map( A => A_s(12), ZN => n301);
   U141 : INV_X1 port map( A => A_ns(12), ZN => n299);
   U142 : OAI221_X1 port map( B1 => n205, B2 => n302, C1 => n192, C2 => n300, A
                           => n170, ZN => O_15_port);
   U143 : INV_X1 port map( A => A_s(13), ZN => n302);
   U144 : INV_X1 port map( A => A_ns(13), ZN => n300);
   U145 : OAI221_X1 port map( B1 => n205, B2 => n305, C1 => n192, C2 => n303, A
                           => n169, ZN => O_16_port);
   U146 : INV_X1 port map( A => A_s(14), ZN => n305);
   U147 : INV_X1 port map( A => A_ns(14), ZN => n303);
   U148 : OAI221_X1 port map( B1 => n205, B2 => n306, C1 => n192, C2 => n304, A
                           => n168, ZN => O_17_port);
   U149 : INV_X1 port map( A => A_s(15), ZN => n306);
   U150 : INV_X1 port map( A => A_ns(15), ZN => n304);
   U151 : OAI221_X1 port map( B1 => n204, B2 => n309, C1 => n192, C2 => n307, A
                           => n167, ZN => O_18_port);
   U152 : INV_X1 port map( A => A_s(16), ZN => n309);
   U153 : INV_X1 port map( A => A_ns(16), ZN => n307);
   U154 : OAI22_X1 port map( A1 => n164, A2 => n277, B1 => n165, B2 => n275, ZN
                           => O_1_port);
   U155 : OAI221_X1 port map( B1 => n203, B2 => n277, C1 => n193, C2 => n275, A
                           => n153, ZN => O_2_port);
   U156 : AOI22_X1 port map( A1 => A_ns(1), A2 => n188, B1 => A_s(1), B2 => 
                           n181, ZN => n153);
   U157 : OAI221_X1 port map( B1 => n203, B2 => n278, C1 => n194, C2 => n276, A
                           => n142, ZN => O_3_port);
   U158 : INV_X1 port map( A => A_s(1), ZN => n278);
   U159 : INV_X1 port map( A => A_ns(1), ZN => n276);
   U160 : OAI221_X1 port map( B1 => n202, B2 => n281, C1 => n195, C2 => n279, A
                           => n131, ZN => O_4_port);
   U161 : INV_X1 port map( A => A_s(2), ZN => n281);
   U162 : INV_X1 port map( A => A_ns(2), ZN => n279);
   U163 : OAI221_X1 port map( B1 => n201, B2 => n282, C1 => n195, C2 => n280, A
                           => n122, ZN => O_5_port);
   U164 : INV_X1 port map( A => A_s(3), ZN => n282);
   U165 : INV_X1 port map( A => A_ns(3), ZN => n280);
   U166 : OAI221_X1 port map( B1 => n201, B2 => n285, C1 => n196, C2 => n283, A
                           => n121, ZN => O_6_port);
   U167 : INV_X1 port map( A => A_s(4), ZN => n285);
   U168 : INV_X1 port map( A => A_ns(4), ZN => n283);
   U169 : OAI221_X1 port map( B1 => n201, B2 => n286, C1 => n196, C2 => n284, A
                           => n120, ZN => O_7_port);
   U170 : INV_X1 port map( A => A_s(5), ZN => n286);
   U171 : INV_X1 port map( A => A_ns(5), ZN => n284);
   U172 : INV_X1 port map( A => A_ns(0), ZN => n275);
   U173 : INV_X1 port map( A => A_s(0), ZN => n277);
   U174 : AOI22_X1 port map( A1 => A_ns(2), A2 => n189, B1 => A_s(2), B2 => 
                           n182, ZN => n142);
   U175 : AOI22_X1 port map( A1 => A_ns(3), A2 => n190, B1 => A_s(3), B2 => 
                           n183, ZN => n131);
   U176 : AOI22_X1 port map( A1 => A_ns(4), A2 => n191, B1 => A_s(4), B2 => 
                           n184, ZN => n122);
   U177 : AOI22_X1 port map( A1 => A_ns(5), A2 => n191, B1 => A_s(5), B2 => 
                           n184, ZN => n121);
   U178 : AOI22_X1 port map( A1 => A_ns(6), A2 => n191, B1 => A_s(6), B2 => 
                           n184, ZN => n120);
   U179 : AOI22_X1 port map( A1 => A_ns(7), A2 => n191, B1 => A_s(7), B2 => 
                           n184, ZN => n119);
   U180 : AOI22_X1 port map( A1 => A_ns(8), A2 => n191, B1 => A_s(8), B2 => 
                           n184, ZN => n118);
   U181 : AOI22_X1 port map( A1 => A_ns(9), A2 => n187, B1 => A_s(9), B2 => 
                           n180, ZN => n175);
   U182 : AOI22_X1 port map( A1 => A_ns(10), A2 => n187, B1 => A_s(10), B2 => 
                           n180, ZN => n174);
   U183 : AOI22_X1 port map( A1 => A_ns(11), A2 => n187, B1 => A_s(11), B2 => 
                           n180, ZN => n173);
   U184 : AOI22_X1 port map( A1 => A_ns(12), A2 => n187, B1 => A_s(12), B2 => 
                           n180, ZN => n172);
   U185 : AOI22_X1 port map( A1 => A_ns(13), A2 => n187, B1 => A_s(13), B2 => 
                           n180, ZN => n171);
   U186 : AOI22_X1 port map( A1 => A_ns(14), A2 => n187, B1 => A_s(14), B2 => 
                           n180, ZN => n170);
   U187 : AOI22_X1 port map( A1 => A_ns(15), A2 => n187, B1 => A_s(15), B2 => 
                           n180, ZN => n169);
   U188 : AOI22_X1 port map( A1 => A_ns(16), A2 => n187, B1 => A_s(16), B2 => 
                           n180, ZN => n168);
   U189 : AOI22_X1 port map( A1 => A_ns(17), A2 => n187, B1 => A_s(17), B2 => 
                           n180, ZN => n167);
   U190 : AOI22_X1 port map( A1 => A_ns(18), A2 => n187, B1 => A_s(18), B2 => 
                           n180, ZN => n166);
   U191 : AOI22_X1 port map( A1 => A_ns(19), A2 => n187, B1 => A_s(19), B2 => 
                           n180, ZN => n163);
   U192 : AOI22_X1 port map( A1 => A_ns(20), A2 => n187, B1 => A_s(20), B2 => 
                           n180, ZN => n162);
   U193 : AOI22_X1 port map( A1 => A_ns(21), A2 => n188, B1 => A_s(21), B2 => 
                           n181, ZN => n161);
   U194 : AOI22_X1 port map( A1 => A_ns(22), A2 => n188, B1 => A_s(22), B2 => 
                           n181, ZN => n160);
   U195 : INV_X1 port map( A => A_ns(24), ZN => n206);
   U196 : INV_X1 port map( A => A_ns(25), ZN => n207);
   U197 : INV_X1 port map( A => A_ns(26), ZN => n208);
   U198 : INV_X1 port map( A => A_ns(27), ZN => n209);
   U199 : INV_X1 port map( A => A_ns(28), ZN => n210);
   U200 : INV_X1 port map( A => A_ns(29), ZN => n211);
   U201 : INV_X1 port map( A => A_ns(30), ZN => n212);
   U202 : INV_X1 port map( A => A_ns(31), ZN => n213);
   U203 : INV_X1 port map( A => A_ns(32), ZN => n214);
   U204 : INV_X1 port map( A => A_ns(33), ZN => n215);
   U205 : INV_X1 port map( A => A_ns(34), ZN => n216);
   U206 : INV_X1 port map( A => A_ns(35), ZN => n217);
   U207 : INV_X1 port map( A => A_ns(36), ZN => n218);
   U208 : INV_X1 port map( A => A_ns(37), ZN => n219);
   U209 : INV_X1 port map( A => A_ns(38), ZN => n220);
   U210 : INV_X1 port map( A => A_ns(39), ZN => n221);
   U211 : INV_X1 port map( A => A_ns(40), ZN => n222);
   U212 : INV_X1 port map( A => A_ns(41), ZN => n223);
   U213 : INV_X1 port map( A => A_ns(42), ZN => n224);
   U214 : INV_X1 port map( A => A_ns(43), ZN => n225);
   U215 : INV_X1 port map( A => A_ns(44), ZN => n226);
   U216 : INV_X1 port map( A => A_ns(45), ZN => n227);
   U217 : INV_X1 port map( A => n229, ZN => A_nso_48_port);
   U218 : INV_X1 port map( A => A_ns(46), ZN => n229);
   U219 : INV_X1 port map( A => n231, ZN => A_nso_49_port);
   U220 : INV_X1 port map( A => A_ns(47), ZN => n231);
   U221 : INV_X1 port map( A => A_ns(48), ZN => n232);
   U222 : INV_X1 port map( A => A_ns(49), ZN => n233);
   U223 : INV_X1 port map( A => A_ns(50), ZN => n234);
   U224 : INV_X1 port map( A => A_ns(51), ZN => n235);
   U225 : INV_X1 port map( A => A_ns(52), ZN => n236);
   U226 : INV_X1 port map( A => A_ns(53), ZN => n237);
   U227 : INV_X1 port map( A => A_ns(54), ZN => n238);
   U228 : INV_X1 port map( A => A_ns(55), ZN => n239);
   U229 : INV_X1 port map( A => A_ns(23), ZN => n240);
   U230 : INV_X1 port map( A => A_s(23), ZN => n241);
   U231 : INV_X1 port map( A => A_s(24), ZN => n242);
   U232 : INV_X1 port map( A => A_s(25), ZN => n243);
   U235 : INV_X1 port map( A => A_s(26), ZN => n244);
   U236 : INV_X1 port map( A => A_s(27), ZN => n245);
   U237 : INV_X1 port map( A => A_s(28), ZN => n246);
   U238 : INV_X1 port map( A => A_s(29), ZN => n247);
   U239 : INV_X1 port map( A => A_s(30), ZN => n248);
   U240 : INV_X1 port map( A => A_s(31), ZN => n249);
   U241 : INV_X1 port map( A => A_s(32), ZN => n250);
   U242 : INV_X1 port map( A => A_s(33), ZN => n251);
   U243 : INV_X1 port map( A => A_s(34), ZN => n252);
   U244 : INV_X1 port map( A => A_s(35), ZN => n253);
   U245 : INV_X1 port map( A => A_s(36), ZN => n254);
   U246 : INV_X1 port map( A => A_s(37), ZN => n255);
   U247 : INV_X1 port map( A => A_s(38), ZN => n256);
   U248 : INV_X1 port map( A => A_s(39), ZN => n257);
   U249 : INV_X1 port map( A => A_s(40), ZN => n258);
   U250 : INV_X1 port map( A => A_s(41), ZN => n259);
   U251 : INV_X1 port map( A => A_s(42), ZN => n260);
   U252 : INV_X1 port map( A => A_s(43), ZN => n261);
   U253 : INV_X1 port map( A => A_s(44), ZN => n262);
   U254 : INV_X1 port map( A => A_s(45), ZN => n263);
   U255 : INV_X1 port map( A => A_s(46), ZN => n264);
   U256 : INV_X1 port map( A => A_s(47), ZN => n265);
   U257 : INV_X1 port map( A => A_s(48), ZN => n266);
   U258 : INV_X1 port map( A => A_s(49), ZN => n267);
   U259 : INV_X1 port map( A => A_s(50), ZN => n268);
   U260 : INV_X1 port map( A => A_s(51), ZN => n269);
   U261 : INV_X1 port map( A => A_s(52), ZN => n270);
   U262 : INV_X1 port map( A => A_s(53), ZN => n271);
   U263 : INV_X1 port map( A => A_s(54), ZN => n272);
   U264 : INV_X1 port map( A => n274, ZN => A_so_57_port);
   U265 : INV_X1 port map( A => A_s(55), ZN => n274);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT56_i22 is

   port( A_s, A_ns, B : in std_logic_vector (55 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (55 downto 0));

end BOOTHENC_NBIT56_i22;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT56_i22 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, O_55_port, O_54_port, O_53_port, O_52_port, O_51_port,
      O_50_port, O_49_port, O_48_port, O_47_port, O_46_port, O_45_port, 
      O_44_port, O_43_port, O_42_port, O_41_port, O_40_port, O_39_port, 
      O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, O_33_port, 
      O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, O_27_port, 
      O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, O_21_port, 
      O_20_port, O_19_port, O_18_port, O_17_port, O_16_port, O_15_port, 
      O_14_port, O_13_port, O_12_port, O_11_port, O_9_port, O_8_port, O_7_port,
      O_6_port, O_5_port, O_4_port, O_3_port, O_2_port, O_10_port, n111, n112, 
      n113, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n167, n168, n169, n170, n174, n175, n176, 
      n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, 
      n189, n190, A_nso_25_port, n192, n193, n194, n195, n196, n197, n198, n199
      , n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, O_1_port, n258, 
      n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, 
      n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, 
      n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, 
      n295, n296, n297 : std_logic;

begin
   O <= ( O_55_port, O_54_port, O_53_port, O_52_port, O_51_port, O_50_port, 
      O_49_port, O_48_port, O_47_port, O_46_port, O_45_port, O_44_port, 
      O_43_port, O_42_port, O_41_port, O_40_port, O_39_port, O_38_port, 
      O_37_port, O_36_port, O_35_port, O_34_port, O_33_port, O_32_port, 
      O_31_port, O_30_port, O_29_port, O_28_port, O_27_port, O_26_port, 
      O_25_port, O_24_port, O_23_port, O_22_port, O_21_port, O_20_port, 
      O_19_port, O_18_port, O_17_port, O_16_port, O_15_port, O_14_port, 
      O_13_port, O_12_port, O_11_port, O_10_port, O_9_port, O_8_port, O_7_port,
      O_6_port, O_5_port, O_4_port, O_3_port, O_2_port, O_1_port, X_Logic0_port
      );
   A_so <= ( A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), 
      A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), 
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   A_nso <= ( A_ns(53), A_ns(52), A_ns(51), A_ns(50), A_ns(49), A_ns(48), 
      A_ns(47), A_ns(46), A_ns(45), A_ns(44), A_ns(43), A_ns(42), A_ns(41), 
      A_ns(40), A_ns(39), A_ns(38), A_ns(37), A_ns(36), A_ns(35), A_ns(34), 
      A_ns(33), A_ns(32), A_ns(31), A_ns(30), A_ns(29), A_ns(28), A_ns(27), 
      A_ns(26), A_ns(25), A_ns(24), A_nso_25_port, A_ns(22), A_ns(21), A_ns(20)
      , A_ns(19), A_ns(18), A_ns(17), A_ns(16), A_ns(15), A_ns(14), A_ns(13), 
      A_ns(12), A_ns(11), A_ns(10), A_ns(9), A_ns(8), A_ns(7), A_ns(6), A_ns(5)
      , A_ns(4), A_ns(3), A_ns(2), A_ns(1), A_ns(0), X_Logic0_port, 
      X_Logic0_port );
   
   X_Logic0_port <= '0';
   U224 : XOR2_X1 port map( A => B(21), B => B(22), Z => n170);
   U225 : NAND3_X1 port map( A1 => B(22), A2 => n297, A3 => B(21), ZN => n119);
   U2 : OAI221_X1 port map( B1 => n111, B2 => n220, C1 => n112, C2 => n254, A 
                           => n123, ZN => O_52_port);
   U3 : OAI221_X1 port map( B1 => n111, B2 => n221, C1 => n112, C2 => n255, A 
                           => n122, ZN => O_53_port);
   U4 : OAI221_X1 port map( B1 => n111, B2 => n222, C1 => n112, C2 => n256, A 
                           => n121, ZN => O_54_port);
   U5 : OAI221_X1 port map( B1 => n187, B2 => n223, C1 => n184, C2 => n224, A 
                           => n156, ZN => O_22_port);
   U6 : INV_X1 port map( A => n189, ZN => n187);
   U7 : INV_X1 port map( A => n189, ZN => n188);
   U8 : INV_X1 port map( A => n186, ZN => n184);
   U9 : BUF_X1 port map( A => n175, Z => n178);
   U10 : INV_X1 port map( A => n186, ZN => n185);
   U11 : BUF_X1 port map( A => n175, Z => n179);
   U12 : BUF_X1 port map( A => n176, Z => n180);
   U13 : BUF_X1 port map( A => n175, Z => n177);
   U14 : BUF_X1 port map( A => n176, Z => n181);
   U15 : AOI22_X1 port map( A1 => A_s(52), A2 => n180, B1 => A_ns(52), B2 => 
                           n183, ZN => n121);
   U16 : AOI22_X1 port map( A1 => A_s(51), A2 => n180, B1 => A_ns(51), B2 => 
                           n183, ZN => n122);
   U17 : AOI22_X1 port map( A1 => A_s(50), A2 => n180, B1 => A_ns(50), B2 => 
                           n183, ZN => n123);
   U18 : OAI221_X1 port map( B1 => n111, B2 => n219, C1 => n112, C2 => n253, A 
                           => n124, ZN => O_51_port);
   U19 : AOI22_X1 port map( A1 => A_s(49), A2 => n180, B1 => A_ns(49), B2 => 
                           n183, ZN => n124);
   U20 : OAI221_X1 port map( B1 => n111, B2 => n218, C1 => n112, C2 => n252, A 
                           => n125, ZN => O_50_port);
   U21 : AOI22_X1 port map( A1 => A_s(48), A2 => n180, B1 => A_ns(48), B2 => 
                           n183, ZN => n125);
   U22 : OAI221_X1 port map( B1 => n111, B2 => n217, C1 => n112, C2 => n251, A 
                           => n127, ZN => O_49_port);
   U23 : AOI22_X1 port map( A1 => A_s(47), A2 => n180, B1 => A_ns(47), B2 => 
                           n183, ZN => n127);
   U24 : OAI221_X1 port map( B1 => n111, B2 => n216, C1 => n112, C2 => n250, A 
                           => n128, ZN => O_48_port);
   U25 : AOI22_X1 port map( A1 => A_s(46), A2 => n180, B1 => A_ns(46), B2 => 
                           n183, ZN => n128);
   U26 : OAI221_X1 port map( B1 => n111, B2 => n215, C1 => n184, C2 => n249, A 
                           => n129, ZN => O_47_port);
   U27 : AOI22_X1 port map( A1 => A_s(45), A2 => n180, B1 => A_ns(45), B2 => 
                           n183, ZN => n129);
   U28 : OAI221_X1 port map( B1 => n111, B2 => n214, C1 => n185, C2 => n248, A 
                           => n130, ZN => O_46_port);
   U29 : AOI22_X1 port map( A1 => A_s(44), A2 => n180, B1 => A_ns(44), B2 => 
                           n183, ZN => n130);
   U30 : OAI221_X1 port map( B1 => n188, B2 => n213, C1 => n185, C2 => n247, A 
                           => n131, ZN => O_45_port);
   U31 : AOI22_X1 port map( A1 => A_s(43), A2 => n180, B1 => A_ns(43), B2 => 
                           n183, ZN => n131);
   U32 : OAI221_X1 port map( B1 => n188, B2 => n212, C1 => n185, C2 => n246, A 
                           => n132, ZN => O_44_port);
   U33 : AOI22_X1 port map( A1 => A_s(42), A2 => n179, B1 => A_ns(42), B2 => 
                           n182, ZN => n132);
   U34 : OAI221_X1 port map( B1 => n188, B2 => n211, C1 => n185, C2 => n245, A 
                           => n133, ZN => O_43_port);
   U35 : AOI22_X1 port map( A1 => A_s(41), A2 => n179, B1 => A_ns(41), B2 => 
                           n182, ZN => n133);
   U36 : OAI221_X1 port map( B1 => n188, B2 => n210, C1 => n185, C2 => n244, A 
                           => n134, ZN => O_42_port);
   U37 : AOI22_X1 port map( A1 => A_s(40), A2 => n179, B1 => A_ns(40), B2 => 
                           n182, ZN => n134);
   U38 : OAI221_X1 port map( B1 => n188, B2 => n209, C1 => n185, C2 => n243, A 
                           => n135, ZN => O_41_port);
   U39 : AOI22_X1 port map( A1 => A_s(39), A2 => n179, B1 => A_ns(39), B2 => 
                           n182, ZN => n135);
   U40 : OAI221_X1 port map( B1 => n188, B2 => n208, C1 => n185, C2 => n242, A 
                           => n136, ZN => O_40_port);
   U41 : AOI22_X1 port map( A1 => A_s(38), A2 => n179, B1 => A_ns(38), B2 => 
                           n182, ZN => n136);
   U42 : OAI221_X1 port map( B1 => n188, B2 => n207, C1 => n185, C2 => n241, A 
                           => n138, ZN => O_39_port);
   U43 : AOI22_X1 port map( A1 => A_s(37), A2 => n179, B1 => A_ns(37), B2 => 
                           n182, ZN => n138);
   U44 : OAI221_X1 port map( B1 => n188, B2 => n206, C1 => n185, C2 => n240, A 
                           => n139, ZN => O_38_port);
   U45 : AOI22_X1 port map( A1 => A_s(36), A2 => n179, B1 => A_ns(36), B2 => 
                           n182, ZN => n139);
   U46 : OAI221_X1 port map( B1 => n188, B2 => n205, C1 => n185, C2 => n239, A 
                           => n140, ZN => O_37_port);
   U47 : AOI22_X1 port map( A1 => A_s(35), A2 => n179, B1 => A_ns(35), B2 => 
                           n182, ZN => n140);
   U48 : OAI221_X1 port map( B1 => n188, B2 => n204, C1 => n185, C2 => n238, A 
                           => n141, ZN => O_36_port);
   U49 : AOI22_X1 port map( A1 => A_s(34), A2 => n179, B1 => A_ns(34), B2 => 
                           n182, ZN => n141);
   U50 : OAI221_X1 port map( B1 => n188, B2 => n203, C1 => n185, C2 => n237, A 
                           => n142, ZN => O_35_port);
   U51 : AOI22_X1 port map( A1 => A_s(33), A2 => n179, B1 => A_ns(33), B2 => 
                           n182, ZN => n142);
   U52 : OAI221_X1 port map( B1 => n188, B2 => n202, C1 => n185, C2 => n236, A 
                           => n143, ZN => O_34_port);
   U53 : AOI22_X1 port map( A1 => A_s(32), A2 => n179, B1 => A_ns(32), B2 => 
                           n182, ZN => n143);
   U54 : OAI221_X1 port map( B1 => n188, B2 => n201, C1 => n185, C2 => n235, A 
                           => n144, ZN => O_33_port);
   U55 : AOI22_X1 port map( A1 => A_s(31), A2 => n178, B1 => A_ns(31), B2 => 
                           n182, ZN => n144);
   U56 : OAI221_X1 port map( B1 => n188, B2 => n200, C1 => n185, C2 => n234, A 
                           => n145, ZN => O_32_port);
   U57 : AOI22_X1 port map( A1 => A_s(30), A2 => n178, B1 => A_ns(30), B2 => 
                           n182, ZN => n145);
   U58 : OAI221_X1 port map( B1 => n188, B2 => n199, C1 => n185, C2 => n233, A 
                           => n146, ZN => O_31_port);
   U59 : AOI22_X1 port map( A1 => A_s(29), A2 => n178, B1 => A_ns(29), B2 => 
                           n182, ZN => n146);
   U60 : OAI221_X1 port map( B1 => n188, B2 => n198, C1 => n185, C2 => n232, A 
                           => n147, ZN => O_30_port);
   U61 : AOI22_X1 port map( A1 => A_s(28), A2 => n178, B1 => A_ns(28), B2 => 
                           n182, ZN => n147);
   U62 : OAI221_X1 port map( B1 => n188, B2 => n197, C1 => n185, C2 => n231, A 
                           => n149, ZN => O_29_port);
   U63 : AOI22_X1 port map( A1 => A_s(27), A2 => n178, B1 => A_ns(27), B2 => 
                           n182, ZN => n149);
   U64 : OAI221_X1 port map( B1 => n188, B2 => n196, C1 => n185, C2 => n230, A 
                           => n150, ZN => O_28_port);
   U65 : AOI22_X1 port map( A1 => A_s(26), A2 => n178, B1 => A_ns(26), B2 => 
                           n182, ZN => n150);
   U66 : OAI221_X1 port map( B1 => n188, B2 => n195, C1 => n185, C2 => n229, A 
                           => n151, ZN => O_27_port);
   U67 : AOI22_X1 port map( A1 => A_s(25), A2 => n178, B1 => A_ns(25), B2 => 
                           n182, ZN => n151);
   U68 : OAI221_X1 port map( B1 => n188, B2 => n193, C1 => n185, C2 => n227, A 
                           => n153, ZN => O_25_port);
   U69 : AOI22_X1 port map( A1 => A_s(23), A2 => n178, B1 => A_nso_25_port, B2 
                           => n182, ZN => n153);
   U70 : OAI221_X1 port map( B1 => n188, B2 => n194, C1 => n185, C2 => n228, A 
                           => n152, ZN => O_26_port);
   U71 : AOI22_X1 port map( A1 => A_s(24), A2 => n178, B1 => A_ns(24), B2 => 
                           n182, ZN => n152);
   U72 : OAI221_X1 port map( B1 => n188, B2 => n192, C1 => n185, C2 => n226, A 
                           => n154, ZN => O_24_port);
   U73 : AOI22_X1 port map( A1 => A_s(22), A2 => n178, B1 => A_ns(22), B2 => 
                           n182, ZN => n154);
   U74 : BUF_X1 port map( A => n296, Z => n175);
   U75 : BUF_X1 port map( A => n296, Z => n176);
   U76 : OAI221_X1 port map( B1 => n119, B2 => n256, C1 => n174, C2 => n222, A 
                           => n120, ZN => O_55_port);
   U77 : AOI22_X1 port map( A1 => A_ns(54), A2 => n189, B1 => A_s(54), B2 => 
                           n186, ZN => n120);
   U78 : OAI221_X1 port map( B1 => n188, B2 => n190, C1 => n185, C2 => n225, A 
                           => n155, ZN => O_23_port);
   U79 : AOI22_X1 port map( A1 => A_s(21), A2 => n178, B1 => A_ns(21), B2 => 
                           n182, ZN => n155);
   U80 : NAND2_X1 port map( A1 => n170, A2 => n184, ZN => n111);
   U81 : NAND2_X1 port map( A1 => n170, A2 => n297, ZN => n112);
   U82 : INV_X1 port map( A => n119, ZN => n296);
   U83 : INV_X1 port map( A => n174, ZN => n182);
   U84 : INV_X1 port map( A => n174, ZN => n183);
   U85 : AOI22_X1 port map( A1 => A_s(20), A2 => n177, B1 => A_ns(20), B2 => 
                           n183, ZN => n156);
   U86 : INV_X1 port map( A => B(23), ZN => n297);
   U87 : OAI221_X1 port map( B1 => n187, B2 => n290, C1 => n184, C2 => n292, A 
                           => n160, ZN => O_19_port);
   U88 : INV_X1 port map( A => A_ns(18), ZN => n290);
   U89 : INV_X1 port map( A => A_s(18), ZN => n292);
   U90 : OAI221_X1 port map( B1 => n187, B2 => n291, C1 => n184, C2 => n293, A 
                           => n158, ZN => O_20_port);
   U91 : INV_X1 port map( A => A_ns(19), ZN => n291);
   U92 : INV_X1 port map( A => A_s(19), ZN => n293);
   U93 : OAI221_X1 port map( B1 => n187, B2 => n294, C1 => n184, C2 => n295, A 
                           => n157, ZN => O_21_port);
   U94 : INV_X1 port map( A => A_ns(20), ZN => n294);
   U95 : INV_X1 port map( A => A_s(20), ZN => n295);
   U96 : OR3_X1 port map( A1 => B(21), A2 => B(22), A3 => n297, ZN => n174);
   U97 : OAI221_X1 port map( B1 => n111, B2 => n269, C1 => n112, C2 => n271, A 
                           => n115, ZN => O_8_port);
   U98 : INV_X1 port map( A => A_ns(7), ZN => n269);
   U99 : INV_X1 port map( A => A_s(7), ZN => n271);
   U100 : OAI221_X1 port map( B1 => n111, B2 => n272, C1 => n112, C2 => n273, A
                           => n113, ZN => O_9_port);
   U101 : AOI22_X1 port map( A1 => A_s(7), A2 => n181, B1 => A_ns(7), B2 => 
                           n183, ZN => n113);
   U102 : OAI221_X1 port map( B1 => n273, B2 => n119, C1 => n272, C2 => n174, A
                           => n169, ZN => O_10_port);
   U103 : AOI22_X1 port map( A1 => A_ns(9), A2 => n189, B1 => A_s(9), B2 => 
                           n186, ZN => n169);
   U104 : OAI221_X1 port map( B1 => n187, B2 => n274, C1 => n184, C2 => n276, A
                           => n168, ZN => O_11_port);
   U105 : INV_X1 port map( A => A_ns(10), ZN => n274);
   U106 : INV_X1 port map( A => A_s(10), ZN => n276);
   U107 : OAI221_X1 port map( B1 => n187, B2 => n275, C1 => n184, C2 => n277, A
                           => n167, ZN => O_12_port);
   U108 : INV_X1 port map( A => A_ns(11), ZN => n275);
   U109 : INV_X1 port map( A => A_s(11), ZN => n277);
   U110 : OAI221_X1 port map( B1 => n187, B2 => n278, C1 => n184, C2 => n280, A
                           => n166, ZN => O_13_port);
   U111 : INV_X1 port map( A => A_ns(12), ZN => n278);
   U112 : INV_X1 port map( A => A_s(12), ZN => n280);
   U113 : OAI221_X1 port map( B1 => n187, B2 => n279, C1 => n184, C2 => n281, A
                           => n165, ZN => O_14_port);
   U114 : INV_X1 port map( A => A_ns(13), ZN => n279);
   U115 : INV_X1 port map( A => A_s(13), ZN => n281);
   U116 : OAI221_X1 port map( B1 => n187, B2 => n282, C1 => n184, C2 => n284, A
                           => n164, ZN => O_15_port);
   U117 : INV_X1 port map( A => A_ns(14), ZN => n282);
   U118 : INV_X1 port map( A => A_s(14), ZN => n284);
   U119 : OAI221_X1 port map( B1 => n187, B2 => n283, C1 => n184, C2 => n285, A
                           => n163, ZN => O_16_port);
   U120 : INV_X1 port map( A => A_ns(15), ZN => n283);
   U121 : INV_X1 port map( A => A_s(15), ZN => n285);
   U122 : OAI221_X1 port map( B1 => n187, B2 => n286, C1 => n184, C2 => n288, A
                           => n162, ZN => O_17_port);
   U123 : INV_X1 port map( A => A_ns(16), ZN => n286);
   U124 : INV_X1 port map( A => A_s(16), ZN => n288);
   U125 : OAI221_X1 port map( B1 => n187, B2 => n287, C1 => n184, C2 => n289, A
                           => n161, ZN => O_18_port);
   U126 : INV_X1 port map( A => A_ns(17), ZN => n287);
   U127 : INV_X1 port map( A => A_s(17), ZN => n289);
   U128 : INV_X1 port map( A => n159, ZN => O_1_port);
   U129 : AOI22_X1 port map( A1 => n186, A2 => A_s(0), B1 => n189, B2 => 
                           A_ns(0), ZN => n159);
   U130 : OAI221_X1 port map( B1 => n188, B2 => n258, C1 => n185, C2 => n259, A
                           => n148, ZN => O_2_port);
   U131 : INV_X1 port map( A => A_ns(1), ZN => n258);
   U132 : INV_X1 port map( A => A_s(1), ZN => n259);
   U133 : OAI221_X1 port map( B1 => n188, B2 => n260, C1 => n112, C2 => n262, A
                           => n137, ZN => O_3_port);
   U134 : INV_X1 port map( A => A_ns(2), ZN => n260);
   U135 : INV_X1 port map( A => A_s(2), ZN => n262);
   U136 : OAI221_X1 port map( B1 => n111, B2 => n261, C1 => n112, C2 => n263, A
                           => n126, ZN => O_4_port);
   U137 : INV_X1 port map( A => A_ns(3), ZN => n261);
   U138 : INV_X1 port map( A => A_s(3), ZN => n263);
   U139 : OAI221_X1 port map( B1 => n111, B2 => n264, C1 => n112, C2 => n266, A
                           => n118, ZN => O_5_port);
   U140 : INV_X1 port map( A => A_ns(4), ZN => n264);
   U141 : INV_X1 port map( A => A_s(4), ZN => n266);
   U142 : OAI221_X1 port map( B1 => n111, B2 => n265, C1 => n112, C2 => n267, A
                           => n117, ZN => O_6_port);
   U143 : INV_X1 port map( A => A_ns(5), ZN => n265);
   U144 : INV_X1 port map( A => A_s(5), ZN => n267);
   U145 : OAI221_X1 port map( B1 => n111, B2 => n268, C1 => n185, C2 => n270, A
                           => n116, ZN => O_7_port);
   U146 : INV_X1 port map( A => A_ns(6), ZN => n268);
   U147 : INV_X1 port map( A => A_s(6), ZN => n270);
   U148 : INV_X1 port map( A => A_s(8), ZN => n273);
   U149 : INV_X1 port map( A => A_ns(8), ZN => n272);
   U150 : AOI22_X1 port map( A1 => A_s(0), A2 => n178, B1 => A_ns(0), B2 => 
                           n182, ZN => n148);
   U151 : AOI22_X1 port map( A1 => A_s(1), A2 => n179, B1 => A_ns(1), B2 => 
                           n182, ZN => n137);
   U152 : AOI22_X1 port map( A1 => A_s(2), A2 => n180, B1 => A_ns(2), B2 => 
                           n183, ZN => n126);
   U153 : AOI22_X1 port map( A1 => A_s(3), A2 => n180, B1 => A_ns(3), B2 => 
                           n183, ZN => n118);
   U154 : AOI22_X1 port map( A1 => A_s(4), A2 => n181, B1 => A_ns(4), B2 => 
                           n183, ZN => n117);
   U155 : AOI22_X1 port map( A1 => A_s(5), A2 => n181, B1 => A_ns(5), B2 => 
                           n183, ZN => n116);
   U156 : AOI22_X1 port map( A1 => A_s(6), A2 => n181, B1 => A_ns(6), B2 => 
                           n183, ZN => n115);
   U157 : AOI22_X1 port map( A1 => A_s(9), A2 => n177, B1 => A_ns(9), B2 => 
                           n183, ZN => n168);
   U158 : AOI22_X1 port map( A1 => A_s(10), A2 => n177, B1 => A_ns(10), B2 => 
                           n183, ZN => n167);
   U159 : AOI22_X1 port map( A1 => A_s(11), A2 => n177, B1 => A_ns(11), B2 => 
                           n183, ZN => n166);
   U160 : AOI22_X1 port map( A1 => A_s(12), A2 => n177, B1 => A_ns(12), B2 => 
                           n183, ZN => n165);
   U161 : AOI22_X1 port map( A1 => A_s(13), A2 => n177, B1 => A_ns(13), B2 => 
                           n183, ZN => n164);
   U162 : AOI22_X1 port map( A1 => A_s(14), A2 => n177, B1 => A_ns(14), B2 => 
                           n183, ZN => n163);
   U163 : AOI22_X1 port map( A1 => A_s(15), A2 => n177, B1 => A_ns(15), B2 => 
                           n183, ZN => n162);
   U164 : AOI22_X1 port map( A1 => A_s(16), A2 => n177, B1 => A_ns(16), B2 => 
                           n183, ZN => n161);
   U165 : AOI22_X1 port map( A1 => A_s(17), A2 => n177, B1 => A_ns(17), B2 => 
                           n183, ZN => n160);
   U166 : AOI22_X1 port map( A1 => A_s(18), A2 => n177, B1 => A_ns(18), B2 => 
                           n182, ZN => n158);
   U167 : AOI22_X1 port map( A1 => A_s(19), A2 => n177, B1 => A_ns(19), B2 => 
                           n182, ZN => n157);
   U168 : INV_X1 port map( A => n112, ZN => n186);
   U169 : INV_X1 port map( A => n111, ZN => n189);
   U170 : INV_X1 port map( A => A_ns(22), ZN => n190);
   U171 : INV_X1 port map( A => n192, ZN => A_nso_25_port);
   U172 : INV_X1 port map( A => A_ns(23), ZN => n192);
   U173 : INV_X1 port map( A => A_ns(24), ZN => n193);
   U174 : INV_X1 port map( A => A_ns(25), ZN => n194);
   U175 : INV_X1 port map( A => A_ns(26), ZN => n195);
   U176 : INV_X1 port map( A => A_ns(27), ZN => n196);
   U177 : INV_X1 port map( A => A_ns(28), ZN => n197);
   U178 : INV_X1 port map( A => A_ns(29), ZN => n198);
   U179 : INV_X1 port map( A => A_ns(30), ZN => n199);
   U180 : INV_X1 port map( A => A_ns(31), ZN => n200);
   U181 : INV_X1 port map( A => A_ns(32), ZN => n201);
   U182 : INV_X1 port map( A => A_ns(33), ZN => n202);
   U183 : INV_X1 port map( A => A_ns(34), ZN => n203);
   U184 : INV_X1 port map( A => A_ns(35), ZN => n204);
   U185 : INV_X1 port map( A => A_ns(36), ZN => n205);
   U186 : INV_X1 port map( A => A_ns(37), ZN => n206);
   U187 : INV_X1 port map( A => A_ns(38), ZN => n207);
   U188 : INV_X1 port map( A => A_ns(39), ZN => n208);
   U189 : INV_X1 port map( A => A_ns(40), ZN => n209);
   U190 : INV_X1 port map( A => A_ns(41), ZN => n210);
   U191 : INV_X1 port map( A => A_ns(42), ZN => n211);
   U192 : INV_X1 port map( A => A_ns(43), ZN => n212);
   U193 : INV_X1 port map( A => A_ns(44), ZN => n213);
   U194 : INV_X1 port map( A => A_ns(45), ZN => n214);
   U195 : INV_X1 port map( A => A_ns(46), ZN => n215);
   U196 : INV_X1 port map( A => A_ns(47), ZN => n216);
   U197 : INV_X1 port map( A => A_ns(48), ZN => n217);
   U198 : INV_X1 port map( A => A_ns(49), ZN => n218);
   U199 : INV_X1 port map( A => A_ns(50), ZN => n219);
   U200 : INV_X1 port map( A => A_ns(51), ZN => n220);
   U201 : INV_X1 port map( A => A_ns(52), ZN => n221);
   U202 : INV_X1 port map( A => A_ns(53), ZN => n222);
   U203 : INV_X1 port map( A => A_ns(21), ZN => n223);
   U204 : INV_X1 port map( A => A_s(21), ZN => n224);
   U205 : INV_X1 port map( A => A_s(22), ZN => n225);
   U206 : INV_X1 port map( A => A_s(23), ZN => n226);
   U207 : INV_X1 port map( A => A_s(24), ZN => n227);
   U208 : INV_X1 port map( A => A_s(25), ZN => n228);
   U209 : INV_X1 port map( A => A_s(26), ZN => n229);
   U210 : INV_X1 port map( A => A_s(27), ZN => n230);
   U211 : INV_X1 port map( A => A_s(28), ZN => n231);
   U212 : INV_X1 port map( A => A_s(29), ZN => n232);
   U213 : INV_X1 port map( A => A_s(30), ZN => n233);
   U214 : INV_X1 port map( A => A_s(31), ZN => n234);
   U215 : INV_X1 port map( A => A_s(32), ZN => n235);
   U216 : INV_X1 port map( A => A_s(33), ZN => n236);
   U217 : INV_X1 port map( A => A_s(34), ZN => n237);
   U218 : INV_X1 port map( A => A_s(35), ZN => n238);
   U219 : INV_X1 port map( A => A_s(36), ZN => n239);
   U220 : INV_X1 port map( A => A_s(37), ZN => n240);
   U221 : INV_X1 port map( A => A_s(38), ZN => n241);
   U222 : INV_X1 port map( A => A_s(39), ZN => n242);
   U223 : INV_X1 port map( A => A_s(40), ZN => n243);
   U226 : INV_X1 port map( A => A_s(41), ZN => n244);
   U227 : INV_X1 port map( A => A_s(42), ZN => n245);
   U228 : INV_X1 port map( A => A_s(43), ZN => n246);
   U229 : INV_X1 port map( A => A_s(44), ZN => n247);
   U230 : INV_X1 port map( A => A_s(45), ZN => n248);
   U231 : INV_X1 port map( A => A_s(46), ZN => n249);
   U232 : INV_X1 port map( A => A_s(47), ZN => n250);
   U233 : INV_X1 port map( A => A_s(48), ZN => n251);
   U234 : INV_X1 port map( A => A_s(49), ZN => n252);
   U235 : INV_X1 port map( A => A_s(50), ZN => n253);
   U236 : INV_X1 port map( A => A_s(51), ZN => n254);
   U237 : INV_X1 port map( A => A_s(52), ZN => n255);
   U238 : INV_X1 port map( A => A_s(53), ZN => n256);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT54_i20 is

   port( A_s, A_ns, B : in std_logic_vector (53 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (53 downto 0));

end BOOTHENC_NBIT54_i20;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT54_i20 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, O_53_port, O_52_port, O_51_port, O_50_port, O_49_port,
      O_48_port, O_47_port, O_46_port, O_45_port, O_44_port, O_43_port, 
      O_42_port, O_41_port, O_40_port, O_39_port, O_38_port, O_37_port, 
      O_36_port, O_35_port, O_34_port, O_33_port, O_32_port, O_31_port, 
      O_30_port, O_29_port, O_28_port, O_27_port, O_26_port, O_25_port, 
      O_24_port, O_23_port, O_22_port, O_21_port, O_20_port, O_19_port, 
      O_18_port, O_17_port, O_16_port, O_15_port, O_14_port, O_13_port, 
      O_12_port, O_11_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, 
      O_4_port, O_3_port, O_2_port, O_10_port, n107, n109, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n169, n170, n171, n172, n173, n174, n175, n176, n177, 
      n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, 
      n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, 
      n202, n203, n204, A_nso_42_port, n206, A_nso_43_port, n208, n209, n210, 
      n211, A_nso_47_port, n213, A_nso_48_port, n215, A_nso_49_port, n217, n218
      , n219, n220, A_nso_53_port, n222, n223, n224, n225, n226, n227, n228, 
      n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, 
      n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, 
      n253, n254, n255, n256, O_1_port, n258, n259, n260, n261, n262, n263, 
      n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, 
      n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, 
      n288, n289, n290, n291, n292, n293 : std_logic;

begin
   O <= ( O_53_port, O_52_port, O_51_port, O_50_port, O_49_port, O_48_port, 
      O_47_port, O_46_port, O_45_port, O_44_port, O_43_port, O_42_port, 
      O_41_port, O_40_port, O_39_port, O_38_port, O_37_port, O_36_port, 
      O_35_port, O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, 
      O_29_port, O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, 
      O_23_port, O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, 
      O_17_port, O_16_port, O_15_port, O_14_port, O_13_port, O_12_port, 
      O_11_port, O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, 
      O_4_port, O_3_port, O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), A_s(46), A_s(45), 
      A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), A_s(38), A_s(37), 
      A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), A_s(30), A_s(29), 
      A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), A_s(22), A_s(21), 
      A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), A_s(14), A_s(13), 
      A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), A_s(6), A_s(5), A_s(4)
      , A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, X_Logic0_port );
   A_nso <= ( A_nso_53_port, A_ns(50), A_ns(49), A_ns(48), A_nso_49_port, 
      A_nso_48_port, A_nso_47_port, A_ns(44), A_ns(43), A_ns(42), A_nso_43_port
      , A_nso_42_port, A_ns(39), A_ns(38), A_ns(37), A_ns(36), A_ns(35), 
      A_ns(34), A_ns(33), A_ns(32), A_ns(31), A_ns(30), A_ns(29), A_ns(28), 
      A_ns(27), A_ns(26), A_ns(25), A_ns(24), A_ns(23), A_ns(22), A_ns(21), 
      A_ns(20), A_ns(19), A_ns(18), A_ns(17), A_ns(16), A_ns(15), A_ns(14), 
      A_ns(13), A_ns(12), A_ns(11), A_ns(10), A_ns(9), A_ns(8), A_ns(7), 
      A_ns(6), A_ns(5), A_ns(4), A_ns(3), A_ns(2), A_ns(1), A_ns(0), 
      X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U216 : XOR2_X1 port map( A => B(19), B => B(20), Z => n164);
   U217 : NAND3_X1 port map( A1 => B(20), A2 => n293, A3 => B(19), ZN => n115);
   U2 : OAI221_X1 port map( B1 => n107, B2 => n220, C1 => n180, C2 => n255, A 
                           => n118, ZN => O_51_port);
   U3 : OAI221_X1 port map( B1 => n107, B2 => n218, C1 => n180, C2 => n253, A 
                           => n121, ZN => O_49_port);
   U4 : INV_X1 port map( A => A_ns(51), ZN => n222);
   U5 : INV_X1 port map( A => A_s(51), ZN => n256);
   U6 : INV_X1 port map( A => n184, ZN => n182);
   U7 : INV_X1 port map( A => n184, ZN => n183);
   U8 : BUF_X1 port map( A => n171, Z => n173);
   U9 : BUF_X1 port map( A => n171, Z => n174);
   U10 : BUF_X1 port map( A => n171, Z => n175);
   U11 : BUF_X1 port map( A => n172, Z => n176);
   U12 : BUF_X1 port map( A => n172, Z => n177);
   U13 : AOI22_X1 port map( A1 => A_s(49), A2 => n176, B1 => A_ns(49), B2 => 
                           n179, ZN => n118);
   U14 : OAI221_X1 port map( B1 => n107, B2 => n222, C1 => n180, C2 => n256, A 
                           => n117, ZN => O_52_port);
   U15 : AOI22_X1 port map( A1 => A_s(50), A2 => n176, B1 => A_ns(50), B2 => 
                           n179, ZN => n117);
   U16 : AOI22_X1 port map( A1 => A_s(47), A2 => n176, B1 => A_nso_49_port, B2 
                           => n179, ZN => n121);
   U17 : OAI221_X1 port map( B1 => n107, B2 => n219, C1 => n180, C2 => n254, A 
                           => n119, ZN => O_50_port);
   U18 : AOI22_X1 port map( A1 => A_s(48), A2 => n176, B1 => A_ns(48), B2 => 
                           n179, ZN => n119);
   U19 : OAI221_X1 port map( B1 => n107, B2 => n217, C1 => n180, C2 => n252, A 
                           => n122, ZN => O_48_port);
   U20 : AOI22_X1 port map( A1 => A_s(46), A2 => n176, B1 => A_nso_48_port, B2 
                           => n179, ZN => n122);
   U21 : OAI221_X1 port map( B1 => n107, B2 => n215, C1 => n181, C2 => n251, A 
                           => n123, ZN => O_47_port);
   U22 : AOI22_X1 port map( A1 => A_s(45), A2 => n176, B1 => A_nso_47_port, B2 
                           => n179, ZN => n123);
   U23 : OAI221_X1 port map( B1 => n182, B2 => n213, C1 => n181, C2 => n250, A 
                           => n124, ZN => O_46_port);
   U24 : AOI22_X1 port map( A1 => A_s(44), A2 => n176, B1 => A_ns(44), B2 => 
                           n179, ZN => n124);
   U25 : OAI221_X1 port map( B1 => n183, B2 => n211, C1 => n181, C2 => n249, A 
                           => n125, ZN => O_45_port);
   U26 : AOI22_X1 port map( A1 => A_s(43), A2 => n176, B1 => A_ns(43), B2 => 
                           n179, ZN => n125);
   U27 : OAI221_X1 port map( B1 => n183, B2 => n210, C1 => n181, C2 => n248, A 
                           => n126, ZN => O_44_port);
   U28 : AOI22_X1 port map( A1 => A_s(42), A2 => n175, B1 => A_ns(42), B2 => 
                           n179, ZN => n126);
   U29 : OAI221_X1 port map( B1 => n183, B2 => n209, C1 => n181, C2 => n247, A 
                           => n127, ZN => O_43_port);
   U30 : AOI22_X1 port map( A1 => A_s(41), A2 => n175, B1 => A_nso_43_port, B2 
                           => n179, ZN => n127);
   U31 : OAI221_X1 port map( B1 => n183, B2 => n208, C1 => n181, C2 => n246, A 
                           => n128, ZN => O_42_port);
   U32 : AOI22_X1 port map( A1 => A_s(40), A2 => n175, B1 => A_nso_42_port, B2 
                           => n179, ZN => n128);
   U33 : OAI221_X1 port map( B1 => n183, B2 => n206, C1 => n181, C2 => n245, A 
                           => n129, ZN => O_41_port);
   U34 : AOI22_X1 port map( A1 => A_s(39), A2 => n175, B1 => A_ns(39), B2 => 
                           n179, ZN => n129);
   U35 : OAI221_X1 port map( B1 => n183, B2 => n204, C1 => n181, C2 => n244, A 
                           => n130, ZN => O_40_port);
   U36 : AOI22_X1 port map( A1 => A_s(38), A2 => n175, B1 => A_ns(38), B2 => 
                           n179, ZN => n130);
   U37 : OAI221_X1 port map( B1 => n183, B2 => n203, C1 => n181, C2 => n243, A 
                           => n132, ZN => O_39_port);
   U38 : AOI22_X1 port map( A1 => A_s(37), A2 => n175, B1 => A_ns(37), B2 => 
                           n179, ZN => n132);
   U39 : OAI221_X1 port map( B1 => n183, B2 => n202, C1 => n181, C2 => n242, A 
                           => n133, ZN => O_38_port);
   U40 : AOI22_X1 port map( A1 => A_s(36), A2 => n175, B1 => A_ns(36), B2 => 
                           n179, ZN => n133);
   U41 : OAI221_X1 port map( B1 => n183, B2 => n201, C1 => n181, C2 => n241, A 
                           => n134, ZN => O_37_port);
   U42 : AOI22_X1 port map( A1 => A_s(35), A2 => n175, B1 => A_ns(35), B2 => 
                           n179, ZN => n134);
   U43 : OAI221_X1 port map( B1 => n183, B2 => n200, C1 => n181, C2 => n240, A 
                           => n135, ZN => O_36_port);
   U44 : AOI22_X1 port map( A1 => A_s(34), A2 => n175, B1 => A_ns(34), B2 => 
                           n179, ZN => n135);
   U45 : OAI221_X1 port map( B1 => n183, B2 => n199, C1 => n181, C2 => n239, A 
                           => n136, ZN => O_35_port);
   U46 : AOI22_X1 port map( A1 => A_s(33), A2 => n175, B1 => A_ns(33), B2 => 
                           n179, ZN => n136);
   U47 : OAI221_X1 port map( B1 => n183, B2 => n198, C1 => n181, C2 => n238, A 
                           => n137, ZN => O_34_port);
   U48 : AOI22_X1 port map( A1 => A_s(32), A2 => n175, B1 => A_ns(32), B2 => 
                           n179, ZN => n137);
   U49 : OAI221_X1 port map( B1 => n183, B2 => n197, C1 => n181, C2 => n237, A 
                           => n138, ZN => O_33_port);
   U50 : AOI22_X1 port map( A1 => A_s(31), A2 => n174, B1 => A_ns(31), B2 => 
                           n178, ZN => n138);
   U51 : OAI221_X1 port map( B1 => n183, B2 => n196, C1 => n181, C2 => n236, A 
                           => n139, ZN => O_32_port);
   U52 : AOI22_X1 port map( A1 => A_s(30), A2 => n174, B1 => A_ns(30), B2 => 
                           n178, ZN => n139);
   U53 : OAI221_X1 port map( B1 => n183, B2 => n187, C1 => n181, C2 => n227, A 
                           => n149, ZN => O_23_port);
   U54 : AOI22_X1 port map( A1 => A_s(21), A2 => n174, B1 => A_ns(21), B2 => 
                           n178, ZN => n149);
   U55 : OAI221_X1 port map( B1 => n183, B2 => n188, C1 => n181, C2 => n228, A 
                           => n148, ZN => O_24_port);
   U56 : AOI22_X1 port map( A1 => A_s(22), A2 => n174, B1 => A_ns(22), B2 => 
                           n178, ZN => n148);
   U57 : OAI221_X1 port map( B1 => n183, B2 => n189, C1 => n181, C2 => n229, A 
                           => n147, ZN => O_25_port);
   U58 : AOI22_X1 port map( A1 => A_s(23), A2 => n174, B1 => A_ns(23), B2 => 
                           n178, ZN => n147);
   U59 : OAI221_X1 port map( B1 => n183, B2 => n190, C1 => n181, C2 => n230, A 
                           => n146, ZN => O_26_port);
   U60 : AOI22_X1 port map( A1 => A_s(24), A2 => n174, B1 => A_ns(24), B2 => 
                           n178, ZN => n146);
   U61 : OAI221_X1 port map( B1 => n183, B2 => n191, C1 => n181, C2 => n231, A 
                           => n145, ZN => O_27_port);
   U62 : AOI22_X1 port map( A1 => A_s(25), A2 => n174, B1 => A_ns(25), B2 => 
                           n178, ZN => n145);
   U63 : OAI221_X1 port map( B1 => n183, B2 => n192, C1 => n181, C2 => n232, A 
                           => n144, ZN => O_28_port);
   U64 : AOI22_X1 port map( A1 => A_s(26), A2 => n174, B1 => A_ns(26), B2 => 
                           n178, ZN => n144);
   U65 : OAI221_X1 port map( B1 => n183, B2 => n193, C1 => n181, C2 => n233, A 
                           => n143, ZN => O_29_port);
   U66 : AOI22_X1 port map( A1 => A_s(27), A2 => n174, B1 => A_ns(27), B2 => 
                           n178, ZN => n143);
   U67 : OAI221_X1 port map( B1 => n183, B2 => n194, C1 => n181, C2 => n234, A 
                           => n141, ZN => O_30_port);
   U68 : AOI22_X1 port map( A1 => A_s(28), A2 => n174, B1 => A_ns(28), B2 => 
                           n178, ZN => n141);
   U69 : OAI221_X1 port map( B1 => n183, B2 => n195, C1 => n181, C2 => n235, A 
                           => n140, ZN => O_31_port);
   U70 : AOI22_X1 port map( A1 => A_s(29), A2 => n174, B1 => A_ns(29), B2 => 
                           n178, ZN => n140);
   U71 : OAI221_X1 port map( B1 => n182, B2 => n186, C1 => n180, C2 => n226, A 
                           => n150, ZN => O_22_port);
   U72 : AOI22_X1 port map( A1 => A_s(20), A2 => n173, B1 => A_ns(20), B2 => 
                           n179, ZN => n150);
   U73 : BUF_X1 port map( A => n292, Z => n171);
   U74 : BUF_X1 port map( A => n292, Z => n172);
   U75 : OAI221_X1 port map( B1 => n115, B2 => n256, C1 => n170, C2 => n222, A 
                           => n116, ZN => O_53_port);
   U76 : AOI22_X1 port map( A1 => A_ns(52), A2 => n184, B1 => A_s(52), B2 => 
                           n169, ZN => n116);
   U77 : OAI221_X1 port map( B1 => n182, B2 => n185, C1 => n180, C2 => n225, A 
                           => n151, ZN => O_21_port);
   U78 : AOI22_X1 port map( A1 => A_s(19), A2 => n173, B1 => A_ns(19), B2 => 
                           n178, ZN => n151);
   U79 : INV_X1 port map( A => n170, ZN => n178);
   U80 : NAND2_X1 port map( A1 => n164, A2 => n180, ZN => n107);
   U81 : AND2_X1 port map( A1 => n164, A2 => n293, ZN => n169);
   U82 : INV_X1 port map( A => n115, ZN => n292);
   U83 : INV_X1 port map( A => n170, ZN => n179);
   U84 : OAI221_X1 port map( B1 => n182, B2 => n223, C1 => n180, C2 => n224, A 
                           => n152, ZN => O_20_port);
   U85 : AOI22_X1 port map( A1 => A_s(18), A2 => n173, B1 => A_ns(18), B2 => 
                           n179, ZN => n152);
   U86 : OR3_X1 port map( A1 => B(19), A2 => B(20), A3 => n293, ZN => n170);
   U87 : INV_X1 port map( A => B(21), ZN => n293);
   U88 : OAI221_X1 port map( B1 => n182, B2 => n290, C1 => n180, C2 => n291, A 
                           => n154, ZN => O_19_port);
   U89 : INV_X1 port map( A => A_ns(18), ZN => n290);
   U90 : INV_X1 port map( A => A_s(18), ZN => n291);
   U91 : OAI221_X1 port map( B1 => n107, B2 => n269, C1 => n180, C2 => n271, A 
                           => n111, ZN => O_8_port);
   U92 : INV_X1 port map( A => A_ns(7), ZN => n269);
   U93 : INV_X1 port map( A => A_s(7), ZN => n271);
   U94 : OAI221_X1 port map( B1 => n107, B2 => n272, C1 => n180, C2 => n273, A 
                           => n109, ZN => O_9_port);
   U95 : AOI22_X1 port map( A1 => A_s(7), A2 => n177, B1 => A_ns(7), B2 => n178
                           , ZN => n109);
   U96 : OAI221_X1 port map( B1 => n273, B2 => n115, C1 => n272, C2 => n170, A 
                           => n163, ZN => O_10_port);
   U97 : AOI22_X1 port map( A1 => A_ns(9), A2 => n184, B1 => A_s(9), B2 => n169
                           , ZN => n163);
   U98 : OAI221_X1 port map( B1 => n182, B2 => n274, C1 => n180, C2 => n276, A 
                           => n162, ZN => O_11_port);
   U99 : INV_X1 port map( A => A_ns(10), ZN => n274);
   U100 : INV_X1 port map( A => A_s(10), ZN => n276);
   U101 : OAI221_X1 port map( B1 => n182, B2 => n275, C1 => n180, C2 => n277, A
                           => n161, ZN => O_12_port);
   U102 : INV_X1 port map( A => A_ns(11), ZN => n275);
   U103 : INV_X1 port map( A => A_s(11), ZN => n277);
   U104 : OAI221_X1 port map( B1 => n182, B2 => n278, C1 => n180, C2 => n280, A
                           => n160, ZN => O_13_port);
   U105 : INV_X1 port map( A => A_ns(12), ZN => n278);
   U106 : INV_X1 port map( A => A_s(12), ZN => n280);
   U107 : OAI221_X1 port map( B1 => n182, B2 => n279, C1 => n180, C2 => n281, A
                           => n159, ZN => O_14_port);
   U108 : INV_X1 port map( A => A_ns(13), ZN => n279);
   U109 : INV_X1 port map( A => A_s(13), ZN => n281);
   U110 : OAI221_X1 port map( B1 => n182, B2 => n282, C1 => n180, C2 => n284, A
                           => n158, ZN => O_15_port);
   U111 : INV_X1 port map( A => A_ns(14), ZN => n282);
   U112 : INV_X1 port map( A => A_s(14), ZN => n284);
   U113 : OAI221_X1 port map( B1 => n182, B2 => n283, C1 => n180, C2 => n285, A
                           => n157, ZN => O_16_port);
   U114 : INV_X1 port map( A => A_ns(15), ZN => n283);
   U115 : INV_X1 port map( A => A_s(15), ZN => n285);
   U116 : OAI221_X1 port map( B1 => n182, B2 => n286, C1 => n180, C2 => n288, A
                           => n156, ZN => O_17_port);
   U117 : INV_X1 port map( A => A_ns(16), ZN => n286);
   U118 : INV_X1 port map( A => A_s(16), ZN => n288);
   U119 : OAI221_X1 port map( B1 => n182, B2 => n287, C1 => n180, C2 => n289, A
                           => n155, ZN => O_18_port);
   U120 : INV_X1 port map( A => A_ns(17), ZN => n287);
   U121 : INV_X1 port map( A => A_s(17), ZN => n289);
   U122 : INV_X1 port map( A => n153, ZN => O_1_port);
   U123 : AOI22_X1 port map( A1 => n169, A2 => A_s(0), B1 => n184, B2 => 
                           A_ns(0), ZN => n153);
   U124 : OAI221_X1 port map( B1 => n183, B2 => n258, C1 => n181, C2 => n259, A
                           => n142, ZN => O_2_port);
   U125 : INV_X1 port map( A => A_ns(1), ZN => n258);
   U126 : INV_X1 port map( A => A_s(1), ZN => n259);
   U127 : OAI221_X1 port map( B1 => n107, B2 => n260, C1 => n180, C2 => n262, A
                           => n131, ZN => O_3_port);
   U128 : INV_X1 port map( A => A_ns(2), ZN => n260);
   U129 : INV_X1 port map( A => A_s(2), ZN => n262);
   U130 : OAI221_X1 port map( B1 => n107, B2 => n261, C1 => n180, C2 => n263, A
                           => n120, ZN => O_4_port);
   U131 : INV_X1 port map( A => A_ns(3), ZN => n261);
   U132 : INV_X1 port map( A => A_s(3), ZN => n263);
   U133 : OAI221_X1 port map( B1 => n107, B2 => n264, C1 => n180, C2 => n266, A
                           => n114, ZN => O_5_port);
   U134 : INV_X1 port map( A => A_ns(4), ZN => n264);
   U135 : INV_X1 port map( A => A_s(4), ZN => n266);
   U136 : OAI221_X1 port map( B1 => n107, B2 => n265, C1 => n180, C2 => n267, A
                           => n113, ZN => O_6_port);
   U137 : INV_X1 port map( A => A_ns(5), ZN => n265);
   U138 : INV_X1 port map( A => A_s(5), ZN => n267);
   U139 : OAI221_X1 port map( B1 => n183, B2 => n268, C1 => n180, C2 => n270, A
                           => n112, ZN => O_7_port);
   U140 : INV_X1 port map( A => A_ns(6), ZN => n268);
   U141 : INV_X1 port map( A => A_s(6), ZN => n270);
   U142 : INV_X1 port map( A => A_s(8), ZN => n273);
   U143 : INV_X1 port map( A => A_ns(8), ZN => n272);
   U144 : AOI22_X1 port map( A1 => A_s(0), A2 => n174, B1 => A_ns(0), B2 => 
                           n178, ZN => n142);
   U145 : AOI22_X1 port map( A1 => A_s(1), A2 => n175, B1 => A_ns(1), B2 => 
                           n179, ZN => n131);
   U146 : AOI22_X1 port map( A1 => A_s(2), A2 => n176, B1 => A_ns(2), B2 => 
                           n178, ZN => n120);
   U147 : AOI22_X1 port map( A1 => A_s(3), A2 => n176, B1 => A_ns(3), B2 => 
                           n178, ZN => n114);
   U148 : AOI22_X1 port map( A1 => A_s(4), A2 => n176, B1 => A_ns(4), B2 => 
                           n178, ZN => n113);
   U149 : AOI22_X1 port map( A1 => A_s(5), A2 => n176, B1 => A_ns(5), B2 => 
                           n178, ZN => n112);
   U150 : AOI22_X1 port map( A1 => A_s(6), A2 => n177, B1 => A_ns(6), B2 => 
                           n178, ZN => n111);
   U151 : AOI22_X1 port map( A1 => A_s(9), A2 => n173, B1 => A_ns(9), B2 => 
                           n179, ZN => n162);
   U152 : AOI22_X1 port map( A1 => A_s(10), A2 => n173, B1 => A_ns(10), B2 => 
                           n179, ZN => n161);
   U153 : AOI22_X1 port map( A1 => A_s(11), A2 => n173, B1 => A_ns(11), B2 => 
                           n179, ZN => n160);
   U154 : AOI22_X1 port map( A1 => A_s(12), A2 => n173, B1 => A_ns(12), B2 => 
                           n179, ZN => n159);
   U155 : AOI22_X1 port map( A1 => A_s(13), A2 => n173, B1 => A_ns(13), B2 => 
                           n178, ZN => n158);
   U156 : AOI22_X1 port map( A1 => A_s(14), A2 => n173, B1 => A_ns(14), B2 => 
                           n178, ZN => n157);
   U157 : AOI22_X1 port map( A1 => A_s(15), A2 => n173, B1 => A_ns(15), B2 => 
                           n178, ZN => n156);
   U158 : AOI22_X1 port map( A1 => A_s(16), A2 => n173, B1 => A_ns(16), B2 => 
                           n178, ZN => n155);
   U159 : AOI22_X1 port map( A1 => A_s(17), A2 => n173, B1 => A_ns(17), B2 => 
                           n178, ZN => n154);
   U160 : INV_X1 port map( A => n169, ZN => n180);
   U161 : INV_X1 port map( A => n169, ZN => n181);
   U162 : INV_X1 port map( A => n107, ZN => n184);
   U163 : INV_X1 port map( A => A_ns(20), ZN => n185);
   U164 : INV_X1 port map( A => A_ns(21), ZN => n186);
   U165 : INV_X1 port map( A => A_ns(22), ZN => n187);
   U166 : INV_X1 port map( A => A_ns(23), ZN => n188);
   U167 : INV_X1 port map( A => A_ns(24), ZN => n189);
   U168 : INV_X1 port map( A => A_ns(25), ZN => n190);
   U169 : INV_X1 port map( A => A_ns(26), ZN => n191);
   U170 : INV_X1 port map( A => A_ns(27), ZN => n192);
   U171 : INV_X1 port map( A => A_ns(28), ZN => n193);
   U172 : INV_X1 port map( A => A_ns(29), ZN => n194);
   U173 : INV_X1 port map( A => A_ns(30), ZN => n195);
   U174 : INV_X1 port map( A => A_ns(31), ZN => n196);
   U175 : INV_X1 port map( A => A_ns(32), ZN => n197);
   U176 : INV_X1 port map( A => A_ns(33), ZN => n198);
   U177 : INV_X1 port map( A => A_ns(34), ZN => n199);
   U178 : INV_X1 port map( A => A_ns(35), ZN => n200);
   U179 : INV_X1 port map( A => A_ns(36), ZN => n201);
   U180 : INV_X1 port map( A => A_ns(37), ZN => n202);
   U181 : INV_X1 port map( A => A_ns(38), ZN => n203);
   U182 : INV_X1 port map( A => A_ns(39), ZN => n204);
   U183 : INV_X1 port map( A => n206, ZN => A_nso_42_port);
   U184 : INV_X1 port map( A => A_ns(40), ZN => n206);
   U185 : INV_X1 port map( A => n208, ZN => A_nso_43_port);
   U186 : INV_X1 port map( A => A_ns(41), ZN => n208);
   U187 : INV_X1 port map( A => A_ns(42), ZN => n209);
   U188 : INV_X1 port map( A => A_ns(43), ZN => n210);
   U189 : INV_X1 port map( A => A_ns(44), ZN => n211);
   U190 : INV_X1 port map( A => n213, ZN => A_nso_47_port);
   U191 : INV_X1 port map( A => A_ns(45), ZN => n213);
   U192 : INV_X1 port map( A => n215, ZN => A_nso_48_port);
   U193 : INV_X1 port map( A => A_ns(46), ZN => n215);
   U194 : INV_X1 port map( A => n217, ZN => A_nso_49_port);
   U195 : INV_X1 port map( A => A_ns(47), ZN => n217);
   U196 : INV_X1 port map( A => A_ns(48), ZN => n218);
   U197 : INV_X1 port map( A => A_ns(49), ZN => n219);
   U198 : INV_X1 port map( A => A_ns(50), ZN => n220);
   U199 : INV_X1 port map( A => n222, ZN => A_nso_53_port);
   U200 : INV_X1 port map( A => A_ns(19), ZN => n223);
   U201 : INV_X1 port map( A => A_s(19), ZN => n224);
   U202 : INV_X1 port map( A => A_s(20), ZN => n225);
   U203 : INV_X1 port map( A => A_s(21), ZN => n226);
   U204 : INV_X1 port map( A => A_s(22), ZN => n227);
   U205 : INV_X1 port map( A => A_s(23), ZN => n228);
   U206 : INV_X1 port map( A => A_s(24), ZN => n229);
   U207 : INV_X1 port map( A => A_s(25), ZN => n230);
   U208 : INV_X1 port map( A => A_s(26), ZN => n231);
   U209 : INV_X1 port map( A => A_s(27), ZN => n232);
   U210 : INV_X1 port map( A => A_s(28), ZN => n233);
   U211 : INV_X1 port map( A => A_s(29), ZN => n234);
   U212 : INV_X1 port map( A => A_s(30), ZN => n235);
   U213 : INV_X1 port map( A => A_s(31), ZN => n236);
   U214 : INV_X1 port map( A => A_s(32), ZN => n237);
   U215 : INV_X1 port map( A => A_s(33), ZN => n238);
   U218 : INV_X1 port map( A => A_s(34), ZN => n239);
   U219 : INV_X1 port map( A => A_s(35), ZN => n240);
   U220 : INV_X1 port map( A => A_s(36), ZN => n241);
   U221 : INV_X1 port map( A => A_s(37), ZN => n242);
   U222 : INV_X1 port map( A => A_s(38), ZN => n243);
   U223 : INV_X1 port map( A => A_s(39), ZN => n244);
   U224 : INV_X1 port map( A => A_s(40), ZN => n245);
   U225 : INV_X1 port map( A => A_s(41), ZN => n246);
   U226 : INV_X1 port map( A => A_s(42), ZN => n247);
   U227 : INV_X1 port map( A => A_s(43), ZN => n248);
   U228 : INV_X1 port map( A => A_s(44), ZN => n249);
   U229 : INV_X1 port map( A => A_s(45), ZN => n250);
   U230 : INV_X1 port map( A => A_s(46), ZN => n251);
   U231 : INV_X1 port map( A => A_s(47), ZN => n252);
   U232 : INV_X1 port map( A => A_s(48), ZN => n253);
   U233 : INV_X1 port map( A => A_s(49), ZN => n254);
   U234 : INV_X1 port map( A => A_s(50), ZN => n255);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT52_i18 is

   port( A_s, A_ns, B : in std_logic_vector (51 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (51 downto 0));

end BOOTHENC_NBIT52_i18;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT52_i18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, O_49_port, O_50_port, O_51_port, O_48_port, O_47_port,
      O_46_port, O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, 
      O_40_port, O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, 
      O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, 
      O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, 
      O_22_port, O_21_port, O_20_port, O_19_port, O_2_port, O_3_port, O_4_port,
      O_5_port, O_6_port, O_7_port, O_8_port, O_9_port, O_10_port, O_11_port, 
      O_12_port, O_13_port, O_14_port, O_15_port, O_16_port, O_17_port, 
      O_18_port, n105, n107, n108, n109, n110, n111, n112, n113, n114, n115, 
      n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, 
      n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, 
      n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n211, n212, n213, n214, n215, 
      n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, A_nso_20_port
      , n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
      n239, n240, n241, n242, n243, A_nso_37_port, n245, A_nso_38_port, n247, 
      A_nso_39_port, n249, n250, n251, n252, n253, A_nso_44_port, n255, n256, 
      n257, n258, A_nso_48_port, n260, A_nso_49_port, n262, A_nso_50_port, n264
      , n265, A_nso_19_port, n267, n268, n269, n270, n271, n272, n273, n274, 
      n275, A_so_27_port, n277, n278, n279, n280, n281, n282, n283, 
      A_so_34_port, n285, A_so_35_port, n287, A_so_36_port, n289, n290, n291, 
      A_so_39_port, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
      n303, n304, n305, O_1_port, n307, n308, n309, n310, n311, n312, n313, 
      n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, 
      n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, 
      n338 : std_logic;

begin
   O <= ( O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, O_46_port, 
      O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, O_40_port, 
      O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, 
      O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, 
      O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, 
      O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, O_16_port, 
      O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, O_10_port, 
      O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, O_3_port, 
      O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(49), A_s(48), A_s(47), A_s(46), A_s(45), A_s(44), A_s(43), 
      A_s(42), A_s(41), A_s(40), A_s(39), A_s(38), A_so_39_port, A_s(36), 
      A_s(35), A_so_36_port, A_so_35_port, A_so_34_port, A_s(31), A_s(30), 
      A_s(29), A_s(28), A_s(27), A_s(26), A_so_27_port, A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   A_nso <= ( A_ns(49), A_nso_50_port, A_nso_49_port, A_nso_48_port, A_ns(45), 
      A_ns(44), A_ns(43), A_nso_44_port, A_ns(41), A_ns(40), A_ns(39), A_ns(38)
      , A_nso_39_port, A_nso_38_port, A_nso_37_port, A_ns(34), A_ns(33), 
      A_ns(32), A_ns(31), A_ns(30), A_ns(29), A_ns(28), A_ns(27), A_ns(26), 
      A_ns(25), A_ns(24), A_ns(23), A_ns(22), A_ns(21), A_ns(20), A_ns(19), 
      A_nso_20_port, A_nso_19_port, A_ns(16), A_ns(15), A_ns(14), A_ns(13), 
      A_ns(12), A_ns(11), A_ns(10), A_ns(9), A_ns(8), A_ns(7), A_ns(6), A_ns(5)
      , A_ns(4), A_ns(3), A_ns(2), A_ns(1), A_ns(0), X_Logic0_port, 
      X_Logic0_port );
   
   X_Logic0_port <= '0';
   U208 : XOR2_X1 port map( A => B(17), B => B(18), Z => n158);
   U209 : NAND3_X1 port map( A1 => B(18), A2 => n338, A3 => B(17), ZN => n111);
   U2 : OAI221_X1 port map( B1 => n225, B2 => n264, C1 => n222, C2 => n304, A 
                           => n115, ZN => O_49_port);
   U3 : OAI221_X1 port map( B1 => n224, B2 => n267, C1 => n222, C2 => n268, A 
                           => n149, ZN => O_18_port);
   U4 : INV_X1 port map( A => A_ns(49), ZN => n265);
   U5 : BUF_X1 port map( A => n214, Z => n216);
   U6 : BUF_X1 port map( A => n214, Z => n217);
   U7 : BUF_X1 port map( A => n215, Z => n218);
   U8 : BUF_X1 port map( A => n215, Z => n219);
   U9 : INV_X1 port map( A => A_s(49), ZN => n305);
   U10 : OAI221_X1 port map( B1 => n225, B2 => n265, C1 => n222, C2 => n305, A 
                           => n113, ZN => O_50_port);
   U11 : AOI22_X1 port map( A1 => A_s(48), A2 => n219, B1 => A_nso_50_port, B2 
                           => n221, ZN => n113);
   U12 : AOI22_X1 port map( A1 => A_s(47), A2 => n219, B1 => A_nso_49_port, B2 
                           => n221, ZN => n115);
   U13 : OAI221_X1 port map( B1 => n225, B2 => n260, C1 => n223, C2 => n302, A 
                           => n117, ZN => O_47_port);
   U14 : AOI22_X1 port map( A1 => A_s(45), A2 => n219, B1 => A_ns(45), B2 => 
                           n221, ZN => n117);
   U15 : OAI221_X1 port map( B1 => n225, B2 => n258, C1 => n223, C2 => n301, A 
                           => n118, ZN => O_46_port);
   U16 : AOI22_X1 port map( A1 => A_s(44), A2 => n219, B1 => A_ns(44), B2 => 
                           n221, ZN => n118);
   U17 : OAI221_X1 port map( B1 => n225, B2 => n262, C1 => n222, C2 => n303, A 
                           => n116, ZN => O_48_port);
   U18 : AOI22_X1 port map( A1 => A_s(46), A2 => n219, B1 => A_nso_48_port, B2 
                           => n221, ZN => n116);
   U19 : OAI221_X1 port map( B1 => n225, B2 => n257, C1 => n223, C2 => n300, A 
                           => n119, ZN => O_45_port);
   U20 : AOI22_X1 port map( A1 => A_s(43), A2 => n219, B1 => A_ns(43), B2 => 
                           n221, ZN => n119);
   U21 : OAI221_X1 port map( B1 => n225, B2 => n256, C1 => n223, C2 => n299, A 
                           => n120, ZN => O_44_port);
   U22 : AOI22_X1 port map( A1 => A_s(42), A2 => n218, B1 => A_nso_44_port, B2 
                           => n221, ZN => n120);
   U23 : OAI221_X1 port map( B1 => n225, B2 => n255, C1 => n223, C2 => n298, A 
                           => n121, ZN => O_43_port);
   U24 : AOI22_X1 port map( A1 => A_s(41), A2 => n218, B1 => A_ns(41), B2 => 
                           n221, ZN => n121);
   U25 : OAI221_X1 port map( B1 => n225, B2 => n253, C1 => n223, C2 => n297, A 
                           => n122, ZN => O_42_port);
   U26 : AOI22_X1 port map( A1 => A_s(40), A2 => n218, B1 => A_ns(40), B2 => 
                           n221, ZN => n122);
   U27 : OAI221_X1 port map( B1 => n225, B2 => n252, C1 => n223, C2 => n296, A 
                           => n123, ZN => O_41_port);
   U28 : AOI22_X1 port map( A1 => A_s(39), A2 => n218, B1 => A_ns(39), B2 => 
                           n221, ZN => n123);
   U29 : OAI221_X1 port map( B1 => n225, B2 => n251, C1 => n223, C2 => n295, A 
                           => n124, ZN => O_40_port);
   U30 : AOI22_X1 port map( A1 => A_s(38), A2 => n218, B1 => A_ns(38), B2 => 
                           n221, ZN => n124);
   U31 : OAI221_X1 port map( B1 => n225, B2 => n250, C1 => n223, C2 => n294, A 
                           => n126, ZN => O_39_port);
   U32 : AOI22_X1 port map( A1 => A_so_39_port, A2 => n218, B1 => A_nso_39_port
                           , B2 => n221, ZN => n126);
   U33 : OAI221_X1 port map( B1 => n225, B2 => n249, C1 => n223, C2 => n293, A 
                           => n127, ZN => O_38_port);
   U34 : AOI22_X1 port map( A1 => A_s(36), A2 => n218, B1 => A_nso_38_port, B2 
                           => n221, ZN => n127);
   U35 : OAI221_X1 port map( B1 => n225, B2 => n247, C1 => n223, C2 => n291, A 
                           => n128, ZN => O_37_port);
   U36 : AOI22_X1 port map( A1 => A_s(35), A2 => n218, B1 => A_nso_37_port, B2 
                           => n221, ZN => n128);
   U37 : OAI221_X1 port map( B1 => n225, B2 => n245, C1 => n223, C2 => n290, A 
                           => n129, ZN => O_36_port);
   U38 : AOI22_X1 port map( A1 => A_so_36_port, A2 => n218, B1 => A_ns(34), B2 
                           => n221, ZN => n129);
   U39 : OAI221_X1 port map( B1 => n225, B2 => n243, C1 => n223, C2 => n289, A 
                           => n130, ZN => O_35_port);
   U40 : AOI22_X1 port map( A1 => A_so_35_port, A2 => n218, B1 => A_ns(33), B2 
                           => n221, ZN => n130);
   U41 : OAI221_X1 port map( B1 => n225, B2 => n242, C1 => n223, C2 => n287, A 
                           => n131, ZN => O_34_port);
   U42 : AOI22_X1 port map( A1 => A_so_34_port, A2 => n218, B1 => A_ns(32), B2 
                           => n221, ZN => n131);
   U43 : OAI221_X1 port map( B1 => n224, B2 => n241, C1 => n223, C2 => n285, A 
                           => n132, ZN => O_33_port);
   U44 : AOI22_X1 port map( A1 => A_s(31), A2 => n217, B1 => A_ns(31), B2 => 
                           n220, ZN => n132);
   U45 : OAI221_X1 port map( B1 => n224, B2 => n229, C1 => n222, C2 => n271, A 
                           => n145, ZN => O_21_port);
   U46 : AOI22_X1 port map( A1 => A_s(19), A2 => n216, B1 => A_ns(19), B2 => 
                           n220, ZN => n145);
   U47 : OAI221_X1 port map( B1 => n224, B2 => n230, C1 => n222, C2 => n272, A 
                           => n144, ZN => O_22_port);
   U48 : AOI22_X1 port map( A1 => A_s(20), A2 => n216, B1 => A_ns(20), B2 => 
                           n221, ZN => n144);
   U49 : OAI221_X1 port map( B1 => n225, B2 => n231, C1 => n223, C2 => n273, A 
                           => n143, ZN => O_23_port);
   U50 : AOI22_X1 port map( A1 => A_s(21), A2 => n217, B1 => A_ns(21), B2 => 
                           n220, ZN => n143);
   U51 : OAI221_X1 port map( B1 => n224, B2 => n232, C1 => n223, C2 => n274, A 
                           => n142, ZN => O_24_port);
   U52 : AOI22_X1 port map( A1 => A_s(22), A2 => n217, B1 => A_ns(22), B2 => 
                           n220, ZN => n142);
   U53 : OAI221_X1 port map( B1 => n224, B2 => n233, C1 => n223, C2 => n275, A 
                           => n141, ZN => O_25_port);
   U54 : AOI22_X1 port map( A1 => A_s(23), A2 => n217, B1 => A_ns(23), B2 => 
                           n220, ZN => n141);
   U55 : OAI221_X1 port map( B1 => n224, B2 => n234, C1 => n223, C2 => n277, A 
                           => n140, ZN => O_26_port);
   U56 : AOI22_X1 port map( A1 => A_s(24), A2 => n217, B1 => A_ns(24), B2 => 
                           n220, ZN => n140);
   U57 : OAI221_X1 port map( B1 => n224, B2 => n235, C1 => n223, C2 => n278, A 
                           => n139, ZN => O_27_port);
   U58 : AOI22_X1 port map( A1 => A_so_27_port, A2 => n217, B1 => A_ns(25), B2 
                           => n220, ZN => n139);
   U59 : OAI221_X1 port map( B1 => n224, B2 => n236, C1 => n223, C2 => n279, A 
                           => n138, ZN => O_28_port);
   U60 : AOI22_X1 port map( A1 => A_s(26), A2 => n217, B1 => A_ns(26), B2 => 
                           n220, ZN => n138);
   U61 : OAI221_X1 port map( B1 => n224, B2 => n237, C1 => n223, C2 => n280, A 
                           => n137, ZN => O_29_port);
   U62 : AOI22_X1 port map( A1 => A_s(27), A2 => n217, B1 => A_ns(27), B2 => 
                           n220, ZN => n137);
   U63 : OAI221_X1 port map( B1 => n224, B2 => n238, C1 => n223, C2 => n281, A 
                           => n135, ZN => O_30_port);
   U64 : AOI22_X1 port map( A1 => A_s(28), A2 => n217, B1 => A_ns(28), B2 => 
                           n220, ZN => n135);
   U65 : OAI221_X1 port map( B1 => n224, B2 => n239, C1 => n223, C2 => n282, A 
                           => n134, ZN => O_31_port);
   U66 : AOI22_X1 port map( A1 => A_s(29), A2 => n217, B1 => A_ns(29), B2 => 
                           n220, ZN => n134);
   U67 : OAI221_X1 port map( B1 => n224, B2 => n240, C1 => n223, C2 => n283, A 
                           => n133, ZN => O_32_port);
   U68 : AOI22_X1 port map( A1 => A_s(30), A2 => n217, B1 => A_ns(30), B2 => 
                           n220, ZN => n133);
   U69 : OAI221_X1 port map( B1 => n224, B2 => n228, C1 => n222, C2 => n270, A 
                           => n146, ZN => O_20_port);
   U70 : AOI22_X1 port map( A1 => A_s(18), A2 => n216, B1 => A_nso_20_port, B2 
                           => n221, ZN => n146);
   U71 : INV_X1 port map( A => n212, ZN => n223);
   U72 : BUF_X1 port map( A => n337, Z => n214);
   U73 : BUF_X1 port map( A => n337, Z => n215);
   U74 : INV_X1 port map( A => n211, ZN => n225);
   U75 : OAI221_X1 port map( B1 => n111, B2 => n305, C1 => n213, C2 => n265, A 
                           => n112, ZN => O_51_port);
   U76 : AOI22_X1 port map( A1 => A_ns(50), A2 => n211, B1 => A_s(50), B2 => 
                           n212, ZN => n112);
   U77 : OAI221_X1 port map( B1 => n224, B2 => n227, C1 => n222, C2 => n269, A 
                           => n148, ZN => O_19_port);
   U78 : AOI22_X1 port map( A1 => A_s(17), A2 => n216, B1 => A_nso_19_port, B2 
                           => n220, ZN => n148);
   U79 : AND2_X1 port map( A1 => n158, A2 => n222, ZN => n211);
   U80 : AND2_X1 port map( A1 => n158, A2 => n338, ZN => n212);
   U81 : INV_X1 port map( A => n111, ZN => n337);
   U82 : INV_X1 port map( A => n213, ZN => n221);
   U83 : AOI22_X1 port map( A1 => A_s(16), A2 => n216, B1 => A_ns(16), B2 => 
                           n220, ZN => n149);
   U84 : OR3_X1 port map( A1 => B(17), A2 => B(18), A3 => n338, ZN => n213);
   U85 : INV_X1 port map( A => B(19), ZN => n338);
   U86 : OAI221_X1 port map( B1 => n225, B2 => n318, C1 => n222, C2 => n320, A 
                           => n107, ZN => O_8_port);
   U87 : INV_X1 port map( A => A_ns(7), ZN => n318);
   U88 : INV_X1 port map( A => A_s(7), ZN => n320);
   U89 : OAI221_X1 port map( B1 => n225, B2 => n321, C1 => n222, C2 => n322, A 
                           => n105, ZN => O_9_port);
   U90 : AOI22_X1 port map( A1 => A_s(7), A2 => n219, B1 => A_ns(7), B2 => n221
                           , ZN => n105);
   U91 : OAI221_X1 port map( B1 => n322, B2 => n111, C1 => n321, C2 => n213, A 
                           => n157, ZN => O_10_port);
   U92 : AOI22_X1 port map( A1 => A_ns(9), A2 => n211, B1 => A_s(9), B2 => n212
                           , ZN => n157);
   U93 : OAI221_X1 port map( B1 => n224, B2 => n323, C1 => n222, C2 => n325, A 
                           => n156, ZN => O_11_port);
   U94 : INV_X1 port map( A => A_ns(10), ZN => n323);
   U95 : INV_X1 port map( A => A_s(10), ZN => n325);
   U96 : OAI221_X1 port map( B1 => n224, B2 => n324, C1 => n222, C2 => n326, A 
                           => n155, ZN => O_12_port);
   U97 : INV_X1 port map( A => A_ns(11), ZN => n324);
   U98 : INV_X1 port map( A => A_s(11), ZN => n326);
   U99 : OAI221_X1 port map( B1 => n224, B2 => n327, C1 => n222, C2 => n329, A 
                           => n154, ZN => O_13_port);
   U100 : INV_X1 port map( A => A_ns(12), ZN => n327);
   U101 : INV_X1 port map( A => A_s(12), ZN => n329);
   U102 : OAI221_X1 port map( B1 => n224, B2 => n328, C1 => n222, C2 => n330, A
                           => n153, ZN => O_14_port);
   U103 : INV_X1 port map( A => A_ns(13), ZN => n328);
   U104 : INV_X1 port map( A => A_s(13), ZN => n330);
   U105 : OAI221_X1 port map( B1 => n224, B2 => n331, C1 => n222, C2 => n333, A
                           => n152, ZN => O_15_port);
   U106 : INV_X1 port map( A => A_ns(14), ZN => n331);
   U107 : INV_X1 port map( A => A_s(14), ZN => n333);
   U108 : OAI221_X1 port map( B1 => n224, B2 => n332, C1 => n222, C2 => n334, A
                           => n151, ZN => O_16_port);
   U109 : INV_X1 port map( A => A_ns(15), ZN => n332);
   U110 : INV_X1 port map( A => A_s(15), ZN => n334);
   U111 : OAI221_X1 port map( B1 => n224, B2 => n335, C1 => n222, C2 => n336, A
                           => n150, ZN => O_17_port);
   U112 : INV_X1 port map( A => A_ns(16), ZN => n335);
   U113 : INV_X1 port map( A => A_s(16), ZN => n336);
   U114 : INV_X1 port map( A => n147, ZN => O_1_port);
   U115 : AOI22_X1 port map( A1 => n212, A2 => A_s(0), B1 => n211, B2 => 
                           A_ns(0), ZN => n147);
   U116 : OAI221_X1 port map( B1 => n224, B2 => n307, C1 => n223, C2 => n308, A
                           => n136, ZN => O_2_port);
   U117 : INV_X1 port map( A => A_ns(1), ZN => n307);
   U118 : INV_X1 port map( A => A_s(1), ZN => n308);
   U119 : OAI221_X1 port map( B1 => n225, B2 => n309, C1 => n222, C2 => n311, A
                           => n125, ZN => O_3_port);
   U120 : INV_X1 port map( A => A_ns(2), ZN => n309);
   U121 : INV_X1 port map( A => A_s(2), ZN => n311);
   U122 : OAI221_X1 port map( B1 => n225, B2 => n310, C1 => n222, C2 => n312, A
                           => n114, ZN => O_4_port);
   U123 : INV_X1 port map( A => A_ns(3), ZN => n310);
   U124 : INV_X1 port map( A => A_s(3), ZN => n312);
   U125 : OAI221_X1 port map( B1 => n225, B2 => n313, C1 => n222, C2 => n315, A
                           => n110, ZN => O_5_port);
   U126 : INV_X1 port map( A => A_ns(4), ZN => n313);
   U127 : INV_X1 port map( A => A_s(4), ZN => n315);
   U128 : OAI221_X1 port map( B1 => n225, B2 => n314, C1 => n222, C2 => n316, A
                           => n109, ZN => O_6_port);
   U129 : INV_X1 port map( A => A_ns(5), ZN => n314);
   U130 : INV_X1 port map( A => A_s(5), ZN => n316);
   U131 : OAI221_X1 port map( B1 => n225, B2 => n317, C1 => n222, C2 => n319, A
                           => n108, ZN => O_7_port);
   U132 : INV_X1 port map( A => A_ns(6), ZN => n317);
   U133 : INV_X1 port map( A => A_s(6), ZN => n319);
   U134 : INV_X1 port map( A => A_s(8), ZN => n322);
   U135 : INV_X1 port map( A => A_ns(8), ZN => n321);
   U136 : AOI22_X1 port map( A1 => A_s(0), A2 => n217, B1 => A_ns(0), B2 => 
                           n220, ZN => n136);
   U137 : AOI22_X1 port map( A1 => A_s(1), A2 => n218, B1 => A_ns(1), B2 => 
                           n221, ZN => n125);
   U138 : AOI22_X1 port map( A1 => A_s(2), A2 => n219, B1 => A_ns(2), B2 => 
                           n221, ZN => n114);
   U139 : AOI22_X1 port map( A1 => A_s(3), A2 => n219, B1 => A_ns(3), B2 => 
                           n221, ZN => n110);
   U140 : AOI22_X1 port map( A1 => A_s(4), A2 => n219, B1 => A_ns(4), B2 => 
                           n221, ZN => n109);
   U141 : AOI22_X1 port map( A1 => A_s(5), A2 => n219, B1 => A_ns(5), B2 => 
                           n221, ZN => n108);
   U142 : AOI22_X1 port map( A1 => A_s(6), A2 => n219, B1 => A_ns(6), B2 => 
                           n221, ZN => n107);
   U143 : AOI22_X1 port map( A1 => A_s(9), A2 => n216, B1 => A_ns(9), B2 => 
                           n220, ZN => n156);
   U144 : AOI22_X1 port map( A1 => A_s(10), A2 => n216, B1 => A_ns(10), B2 => 
                           n220, ZN => n155);
   U145 : AOI22_X1 port map( A1 => A_s(11), A2 => n216, B1 => A_ns(11), B2 => 
                           n220, ZN => n154);
   U146 : AOI22_X1 port map( A1 => A_s(12), A2 => n216, B1 => A_ns(12), B2 => 
                           n220, ZN => n153);
   U147 : AOI22_X1 port map( A1 => A_s(13), A2 => n216, B1 => A_ns(13), B2 => 
                           n220, ZN => n152);
   U148 : AOI22_X1 port map( A1 => A_s(14), A2 => n216, B1 => A_ns(14), B2 => 
                           n220, ZN => n151);
   U149 : AOI22_X1 port map( A1 => A_s(15), A2 => n216, B1 => A_ns(15), B2 => 
                           n220, ZN => n150);
   U150 : INV_X1 port map( A => n213, ZN => n220);
   U151 : INV_X1 port map( A => n212, ZN => n222);
   U152 : INV_X1 port map( A => n211, ZN => n224);
   U153 : INV_X1 port map( A => n227, ZN => A_nso_20_port);
   U154 : INV_X1 port map( A => A_ns(18), ZN => n227);
   U155 : INV_X1 port map( A => A_ns(19), ZN => n228);
   U156 : INV_X1 port map( A => A_ns(20), ZN => n229);
   U157 : INV_X1 port map( A => A_ns(21), ZN => n230);
   U158 : INV_X1 port map( A => A_ns(22), ZN => n231);
   U159 : INV_X1 port map( A => A_ns(23), ZN => n232);
   U160 : INV_X1 port map( A => A_ns(24), ZN => n233);
   U161 : INV_X1 port map( A => A_ns(25), ZN => n234);
   U162 : INV_X1 port map( A => A_ns(26), ZN => n235);
   U163 : INV_X1 port map( A => A_ns(27), ZN => n236);
   U164 : INV_X1 port map( A => A_ns(28), ZN => n237);
   U165 : INV_X1 port map( A => A_ns(29), ZN => n238);
   U166 : INV_X1 port map( A => A_ns(30), ZN => n239);
   U167 : INV_X1 port map( A => A_ns(31), ZN => n240);
   U168 : INV_X1 port map( A => A_ns(32), ZN => n241);
   U169 : INV_X1 port map( A => A_ns(33), ZN => n242);
   U170 : INV_X1 port map( A => A_ns(34), ZN => n243);
   U171 : INV_X1 port map( A => n245, ZN => A_nso_37_port);
   U172 : INV_X1 port map( A => A_ns(35), ZN => n245);
   U173 : INV_X1 port map( A => n247, ZN => A_nso_38_port);
   U174 : INV_X1 port map( A => A_ns(36), ZN => n247);
   U175 : INV_X1 port map( A => n249, ZN => A_nso_39_port);
   U176 : INV_X1 port map( A => A_ns(37), ZN => n249);
   U177 : INV_X1 port map( A => A_ns(38), ZN => n250);
   U178 : INV_X1 port map( A => A_ns(39), ZN => n251);
   U179 : INV_X1 port map( A => A_ns(40), ZN => n252);
   U180 : INV_X1 port map( A => A_ns(41), ZN => n253);
   U181 : INV_X1 port map( A => n255, ZN => A_nso_44_port);
   U182 : INV_X1 port map( A => A_ns(42), ZN => n255);
   U183 : INV_X1 port map( A => A_ns(43), ZN => n256);
   U184 : INV_X1 port map( A => A_ns(44), ZN => n257);
   U185 : INV_X1 port map( A => A_ns(45), ZN => n258);
   U186 : INV_X1 port map( A => n260, ZN => A_nso_48_port);
   U187 : INV_X1 port map( A => A_ns(46), ZN => n260);
   U188 : INV_X1 port map( A => n262, ZN => A_nso_49_port);
   U189 : INV_X1 port map( A => A_ns(47), ZN => n262);
   U190 : INV_X1 port map( A => n264, ZN => A_nso_50_port);
   U191 : INV_X1 port map( A => A_ns(48), ZN => n264);
   U192 : INV_X1 port map( A => n267, ZN => A_nso_19_port);
   U193 : INV_X1 port map( A => A_ns(17), ZN => n267);
   U194 : INV_X1 port map( A => A_s(17), ZN => n268);
   U195 : INV_X1 port map( A => A_s(18), ZN => n269);
   U196 : INV_X1 port map( A => A_s(19), ZN => n270);
   U197 : INV_X1 port map( A => A_s(20), ZN => n271);
   U198 : INV_X1 port map( A => A_s(21), ZN => n272);
   U199 : INV_X1 port map( A => A_s(22), ZN => n273);
   U200 : INV_X1 port map( A => A_s(23), ZN => n274);
   U201 : INV_X1 port map( A => A_s(24), ZN => n275);
   U202 : INV_X1 port map( A => n277, ZN => A_so_27_port);
   U203 : INV_X1 port map( A => A_s(25), ZN => n277);
   U204 : INV_X1 port map( A => A_s(26), ZN => n278);
   U205 : INV_X1 port map( A => A_s(27), ZN => n279);
   U206 : INV_X1 port map( A => A_s(28), ZN => n280);
   U207 : INV_X1 port map( A => A_s(29), ZN => n281);
   U210 : INV_X1 port map( A => A_s(30), ZN => n282);
   U211 : INV_X1 port map( A => A_s(31), ZN => n283);
   U212 : INV_X1 port map( A => n285, ZN => A_so_34_port);
   U213 : INV_X1 port map( A => A_s(32), ZN => n285);
   U214 : INV_X1 port map( A => n287, ZN => A_so_35_port);
   U215 : INV_X1 port map( A => A_s(33), ZN => n287);
   U216 : INV_X1 port map( A => n289, ZN => A_so_36_port);
   U217 : INV_X1 port map( A => A_s(34), ZN => n289);
   U218 : INV_X1 port map( A => A_s(35), ZN => n290);
   U219 : INV_X1 port map( A => A_s(36), ZN => n291);
   U220 : INV_X1 port map( A => n293, ZN => A_so_39_port);
   U221 : INV_X1 port map( A => A_s(37), ZN => n293);
   U222 : INV_X1 port map( A => A_s(38), ZN => n294);
   U223 : INV_X1 port map( A => A_s(39), ZN => n295);
   U224 : INV_X1 port map( A => A_s(40), ZN => n296);
   U225 : INV_X1 port map( A => A_s(41), ZN => n297);
   U226 : INV_X1 port map( A => A_s(42), ZN => n298);
   U227 : INV_X1 port map( A => A_s(43), ZN => n299);
   U228 : INV_X1 port map( A => A_s(44), ZN => n300);
   U229 : INV_X1 port map( A => A_s(45), ZN => n301);
   U230 : INV_X1 port map( A => A_s(46), ZN => n302);
   U231 : INV_X1 port map( A => A_s(47), ZN => n303);
   U232 : INV_X1 port map( A => A_s(48), ZN => n304);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT50_i16 is

   port( A_s, A_ns, B : in std_logic_vector (49 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (49 downto 0));

end BOOTHENC_NBIT50_i16;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT50_i16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI221_X4
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, O_47_port, O_48_port, O_49_port, O_46_port, O_45_port,
      O_44_port, O_43_port, O_42_port, O_41_port, O_40_port, O_39_port, 
      O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, O_33_port, 
      O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, O_27_port, 
      O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, O_21_port, 
      O_20_port, O_19_port, O_18_port, O_17_port, O_2_port, O_3_port, O_4_port,
      O_5_port, O_6_port, O_7_port, O_8_port, O_9_port, O_10_port, O_11_port, 
      O_12_port, O_13_port, O_14_port, O_15_port, O_16_port, n101, n103, n104, 
      n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, 
      n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, 
      n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, 
      n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, 
      n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, 
      n214, n215, n216, A_nso_18_port, n218, n219, A_nso_20_port, n221, n222, 
      n223, A_nso_23_port, n225, A_nso_24_port, n227, A_nso_25_port, n229, 
      A_nso_26_port, n231, A_nso_27_port, n233, A_nso_28_port, n235, 
      A_nso_29_port, n237, A_nso_30_port, n239, A_nso_31_port, n241, 
      A_nso_32_port, n243, A_nso_33_port, n245, A_nso_34_port, n247, n248, n249
      , n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
      n262, A_nso_17_port, n264, A_so_17_port, n266, A_so_18_port, n268, 
      A_so_19_port, n270, A_so_20_port, n272, A_so_21_port, n274, A_so_22_port,
      n276, A_so_23_port, n278, n279, n280, n281, n282, n283, n284, 
      A_so_30_port, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
      n296, A_so_41_port, n298, A_so_42_port, n300, n301, n302, n303, n304, 
      n305, n306, n307, O_1_port, n309, n310, n311, n312, n313, n314, n315, 
      n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, 
      n328, n329, n330, n331, n332, n333, n334, n335, n336 : std_logic;

begin
   O <= ( O_49_port, O_48_port, O_47_port, O_46_port, O_45_port, O_44_port, 
      O_43_port, O_42_port, O_41_port, O_40_port, O_39_port, O_38_port, 
      O_37_port, O_36_port, O_35_port, O_34_port, O_33_port, O_32_port, 
      O_31_port, O_30_port, O_29_port, O_28_port, O_27_port, O_26_port, 
      O_25_port, O_24_port, O_23_port, O_22_port, O_21_port, O_20_port, 
      O_19_port, O_18_port, O_17_port, O_16_port, O_15_port, O_14_port, 
      O_13_port, O_12_port, O_11_port, O_10_port, O_9_port, O_8_port, O_7_port,
      O_6_port, O_5_port, O_4_port, O_3_port, O_2_port, O_1_port, X_Logic0_port
      );
   A_so <= ( A_s(47), A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), 
      A_so_42_port, A_so_41_port, A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), 
      A_s(33), A_s(32), A_s(31), A_s(30), A_s(29), A_so_30_port, A_s(27), 
      A_s(26), A_s(25), A_s(24), A_s(23), A_s(22), A_so_23_port, A_so_22_port, 
      A_so_21_port, A_so_20_port, A_so_19_port, A_so_18_port, A_so_17_port, 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   A_nso <= ( A_ns(47), A_ns(46), A_ns(45), A_ns(44), A_ns(43), A_ns(42), 
      A_ns(41), A_ns(40), A_ns(39), A_ns(38), A_ns(37), A_ns(36), A_ns(35), 
      A_ns(34), A_ns(33), A_nso_34_port, A_nso_33_port, A_nso_32_port, 
      A_nso_31_port, A_nso_30_port, A_nso_29_port, A_nso_28_port, A_nso_27_port
      , A_nso_26_port, A_nso_25_port, A_nso_24_port, A_nso_23_port, A_ns(20), 
      A_ns(19), A_nso_20_port, A_ns(17), A_nso_18_port, A_nso_17_port, A_ns(14)
      , A_ns(13), A_ns(12), A_ns(11), A_ns(10), A_ns(9), A_ns(8), A_ns(7), 
      A_ns(6), A_ns(5), A_ns(4), A_ns(3), A_ns(2), A_ns(1), A_ns(0), 
      X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U200 : XOR2_X1 port map( A => B(15), B => B(16), Z => n152);
   U201 : NAND3_X1 port map( A1 => B(16), A2 => n336, A3 => B(15), ZN => n108);
   U2 : OAI221_X4 port map( B1 => n216, B2 => n262, C1 => n213, C2 => n307, A 
                           => n110, ZN => O_48_port);
   U3 : OAI221_X1 port map( B1 => n215, B2 => n254, C1 => n214, C2 => n298, A 
                           => n118, ZN => O_40_port);
   U4 : OAI221_X1 port map( B1 => n216, B2 => n259, C1 => n214, C2 => n304, A 
                           => n113, ZN => O_45_port);
   U5 : OAI221_X1 port map( B1 => n216, B2 => n261, C1 => n214, C2 => n306, A 
                           => n111, ZN => O_47_port);
   U6 : OAI221_X1 port map( B1 => n215, B2 => n218, C1 => n213, C2 => n268, A 
                           => n144, ZN => O_17_port);
   U7 : OAI221_X1 port map( B1 => n216, B2 => n264, C1 => n213, C2 => n266, A 
                           => n145, ZN => O_16_port);
   U8 : OAI221_X1 port map( B1 => n216, B2 => n260, C1 => n214, C2 => n305, A 
                           => n112, ZN => O_46_port);
   U9 : INV_X1 port map( A => A_ns(47), ZN => n262);
   U10 : BUF_X1 port map( A => n205, Z => n207);
   U11 : BUF_X1 port map( A => n205, Z => n208);
   U12 : BUF_X1 port map( A => n206, Z => n209);
   U13 : BUF_X1 port map( A => n206, Z => n210);
   U14 : AOI22_X1 port map( A1 => A_s(46), A2 => n210, B1 => A_ns(46), B2 => 
                           n211, ZN => n110);
   U15 : BUF_X1 port map( A => n335, Z => n205);
   U16 : INV_X1 port map( A => n203, ZN => n214);
   U17 : INV_X1 port map( A => n202, ZN => n215);
   U18 : BUF_X1 port map( A => n335, Z => n206);
   U19 : INV_X1 port map( A => n202, ZN => n216);
   U20 : OAI221_X1 port map( B1 => n108, B2 => n307, C1 => n204, C2 => n262, A 
                           => n109, ZN => O_49_port);
   U21 : AOI22_X1 port map( A1 => A_ns(48), A2 => n202, B1 => A_s(48), B2 => 
                           n203, ZN => n109);
   U22 : AOI22_X1 port map( A1 => A_s(45), A2 => n210, B1 => A_ns(45), B2 => 
                           n212, ZN => n111);
   U23 : AOI22_X1 port map( A1 => A_s(43), A2 => n210, B1 => A_ns(43), B2 => 
                           n212, ZN => n113);
   U24 : OAI221_X1 port map( B1 => n215, B2 => n258, C1 => n214, C2 => n303, A 
                           => n114, ZN => O_44_port);
   U25 : AOI22_X1 port map( A1 => A_s(42), A2 => n209, B1 => A_ns(42), B2 => 
                           n212, ZN => n114);
   U26 : AOI22_X1 port map( A1 => A_s(44), A2 => n210, B1 => A_ns(44), B2 => 
                           n212, ZN => n112);
   U27 : OAI221_X1 port map( B1 => n215, B2 => n257, C1 => n214, C2 => n302, A 
                           => n115, ZN => O_43_port);
   U28 : AOI22_X1 port map( A1 => A_s(41), A2 => n209, B1 => A_ns(41), B2 => 
                           n212, ZN => n115);
   U29 : OAI221_X1 port map( B1 => n215, B2 => n256, C1 => n214, C2 => n301, A 
                           => n116, ZN => O_42_port);
   U30 : AOI22_X1 port map( A1 => A_so_42_port, A2 => n209, B1 => A_ns(40), B2 
                           => n212, ZN => n116);
   U31 : OAI221_X1 port map( B1 => n215, B2 => n255, C1 => n214, C2 => n300, A 
                           => n117, ZN => O_41_port);
   U32 : AOI22_X1 port map( A1 => A_so_41_port, A2 => n209, B1 => A_ns(39), B2 
                           => n212, ZN => n117);
   U33 : AOI22_X1 port map( A1 => A_s(38), A2 => n209, B1 => A_ns(38), B2 => 
                           n212, ZN => n118);
   U34 : OAI221_X1 port map( B1 => n215, B2 => n253, C1 => n214, C2 => n296, A 
                           => n120, ZN => O_39_port);
   U35 : AOI22_X1 port map( A1 => A_s(37), A2 => n209, B1 => A_ns(37), B2 => 
                           n212, ZN => n120);
   U36 : OAI221_X1 port map( B1 => n215, B2 => n252, C1 => n214, C2 => n295, A 
                           => n121, ZN => O_38_port);
   U37 : AOI22_X1 port map( A1 => A_s(36), A2 => n209, B1 => A_ns(36), B2 => 
                           n212, ZN => n121);
   U38 : OAI221_X1 port map( B1 => n215, B2 => n251, C1 => n214, C2 => n294, A 
                           => n122, ZN => O_37_port);
   U39 : AOI22_X1 port map( A1 => A_s(35), A2 => n209, B1 => A_ns(35), B2 => 
                           n212, ZN => n122);
   U40 : OAI221_X1 port map( B1 => n215, B2 => n250, C1 => n214, C2 => n293, A 
                           => n123, ZN => O_36_port);
   U41 : AOI22_X1 port map( A1 => A_s(34), A2 => n209, B1 => A_ns(34), B2 => 
                           n212, ZN => n123);
   U42 : OAI221_X1 port map( B1 => n215, B2 => n249, C1 => n214, C2 => n292, A 
                           => n124, ZN => O_35_port);
   U43 : AOI22_X1 port map( A1 => A_s(33), A2 => n209, B1 => A_ns(33), B2 => 
                           n212, ZN => n124);
   U44 : OAI221_X1 port map( B1 => n215, B2 => n248, C1 => n214, C2 => n291, A 
                           => n125, ZN => O_34_port);
   U45 : AOI22_X1 port map( A1 => A_s(32), A2 => n209, B1 => A_nso_34_port, B2 
                           => n212, ZN => n125);
   U46 : OAI221_X1 port map( B1 => n215, B2 => n221, C1 => n213, C2 => n272, A 
                           => n142, ZN => O_19_port);
   U47 : AOI22_X1 port map( A1 => A_so_19_port, A2 => n207, B1 => A_ns(17), B2 
                           => n211, ZN => n142);
   U48 : OAI221_X1 port map( B1 => n216, B2 => n222, C1 => n213, C2 => n274, A 
                           => n140, ZN => O_20_port);
   U49 : AOI22_X1 port map( A1 => A_so_20_port, A2 => n207, B1 => A_nso_20_port
                           , B2 => n211, ZN => n140);
   U50 : OAI221_X1 port map( B1 => n216, B2 => n223, C1 => n213, C2 => n276, A 
                           => n139, ZN => O_21_port);
   U51 : AOI22_X1 port map( A1 => A_so_21_port, A2 => n207, B1 => A_ns(19), B2 
                           => n211, ZN => n139);
   U52 : OAI221_X1 port map( B1 => n216, B2 => n225, C1 => n213, C2 => n278, A 
                           => n138, ZN => O_22_port);
   U53 : AOI22_X1 port map( A1 => A_so_22_port, A2 => n207, B1 => A_ns(20), B2 
                           => n211, ZN => n138);
   U54 : OAI221_X1 port map( B1 => n216, B2 => n227, C1 => n214, C2 => n279, A 
                           => n137, ZN => O_23_port);
   U55 : AOI22_X1 port map( A1 => A_so_23_port, A2 => n208, B1 => A_nso_23_port
                           , B2 => n212, ZN => n137);
   U56 : OAI221_X1 port map( B1 => n215, B2 => n229, C1 => n214, C2 => n280, A 
                           => n136, ZN => O_24_port);
   U57 : AOI22_X1 port map( A1 => A_s(22), A2 => n208, B1 => A_nso_24_port, B2 
                           => n212, ZN => n136);
   U58 : OAI221_X1 port map( B1 => n215, B2 => n231, C1 => n214, C2 => n281, A 
                           => n135, ZN => O_25_port);
   U59 : AOI22_X1 port map( A1 => A_s(23), A2 => n208, B1 => A_nso_25_port, B2 
                           => n212, ZN => n135);
   U60 : OAI221_X1 port map( B1 => n215, B2 => n233, C1 => n214, C2 => n282, A 
                           => n134, ZN => O_26_port);
   U61 : AOI22_X1 port map( A1 => A_s(24), A2 => n208, B1 => A_nso_26_port, B2 
                           => n212, ZN => n134);
   U62 : OAI221_X1 port map( B1 => n215, B2 => n235, C1 => n214, C2 => n283, A 
                           => n133, ZN => O_27_port);
   U63 : AOI22_X1 port map( A1 => A_s(25), A2 => n208, B1 => A_nso_27_port, B2 
                           => n212, ZN => n133);
   U64 : OAI221_X1 port map( B1 => n215, B2 => n237, C1 => n214, C2 => n284, A 
                           => n132, ZN => O_28_port);
   U65 : AOI22_X1 port map( A1 => A_s(26), A2 => n208, B1 => A_nso_28_port, B2 
                           => n212, ZN => n132);
   U66 : OAI221_X1 port map( B1 => n215, B2 => n239, C1 => n214, C2 => n286, A 
                           => n131, ZN => O_29_port);
   U67 : AOI22_X1 port map( A1 => A_s(27), A2 => n208, B1 => A_nso_29_port, B2 
                           => n212, ZN => n131);
   U68 : OAI221_X1 port map( B1 => n215, B2 => n241, C1 => n214, C2 => n287, A 
                           => n129, ZN => O_30_port);
   U69 : AOI22_X1 port map( A1 => A_so_30_port, A2 => n208, B1 => A_nso_30_port
                           , B2 => n212, ZN => n129);
   U70 : OAI221_X1 port map( B1 => n215, B2 => n243, C1 => n214, C2 => n288, A 
                           => n128, ZN => O_31_port);
   U71 : AOI22_X1 port map( A1 => A_s(29), A2 => n208, B1 => A_nso_31_port, B2 
                           => n212, ZN => n128);
   U72 : OAI221_X1 port map( B1 => n215, B2 => n245, C1 => n214, C2 => n289, A 
                           => n127, ZN => O_32_port);
   U73 : AOI22_X1 port map( A1 => A_s(30), A2 => n208, B1 => A_nso_32_port, B2 
                           => n212, ZN => n127);
   U74 : OAI221_X1 port map( B1 => n215, B2 => n247, C1 => n214, C2 => n290, A 
                           => n126, ZN => O_33_port);
   U75 : AOI22_X1 port map( A1 => A_s(31), A2 => n208, B1 => A_nso_33_port, B2 
                           => n212, ZN => n126);
   U76 : OAI221_X1 port map( B1 => n215, B2 => n219, C1 => n213, C2 => n270, A 
                           => n143, ZN => O_18_port);
   U77 : AOI22_X1 port map( A1 => A_so_18_port, A2 => n207, B1 => A_nso_18_port
                           , B2 => n211, ZN => n143);
   U78 : AOI22_X1 port map( A1 => A_so_17_port, A2 => n207, B1 => A_nso_17_port
                           , B2 => n211, ZN => n144);
   U79 : AND2_X1 port map( A1 => n152, A2 => n213, ZN => n202);
   U80 : AND2_X1 port map( A1 => n152, A2 => n336, ZN => n203);
   U81 : INV_X1 port map( A => n108, ZN => n335);
   U82 : INV_X1 port map( A => n204, ZN => n212);
   U83 : INV_X1 port map( A => A_s(47), ZN => n307);
   U84 : AOI22_X1 port map( A1 => A_s(14), A2 => n207, B1 => A_ns(14), B2 => 
                           n211, ZN => n145);
   U85 : OR3_X1 port map( A1 => B(15), A2 => B(16), A3 => n336, ZN => n204);
   U86 : INV_X1 port map( A => B(17), ZN => n336);
   U87 : OAI221_X1 port map( B1 => n216, B2 => n320, C1 => n213, C2 => n322, A 
                           => n103, ZN => O_8_port);
   U88 : INV_X1 port map( A => A_ns(7), ZN => n320);
   U89 : INV_X1 port map( A => A_s(7), ZN => n322);
   U90 : OAI221_X1 port map( B1 => n216, B2 => n323, C1 => n213, C2 => n324, A 
                           => n101, ZN => O_9_port);
   U91 : AOI22_X1 port map( A1 => A_s(7), A2 => n210, B1 => A_ns(7), B2 => n211
                           , ZN => n101);
   U92 : OAI221_X1 port map( B1 => n324, B2 => n108, C1 => n323, C2 => n204, A 
                           => n151, ZN => O_10_port);
   U93 : AOI22_X1 port map( A1 => A_ns(9), A2 => n202, B1 => A_s(9), B2 => n203
                           , ZN => n151);
   U94 : OAI221_X1 port map( B1 => n216, B2 => n325, C1 => n213, C2 => n327, A 
                           => n150, ZN => O_11_port);
   U95 : INV_X1 port map( A => A_ns(10), ZN => n325);
   U96 : INV_X1 port map( A => A_s(10), ZN => n327);
   U97 : OAI221_X1 port map( B1 => n216, B2 => n326, C1 => n213, C2 => n328, A 
                           => n149, ZN => O_12_port);
   U98 : INV_X1 port map( A => A_ns(11), ZN => n326);
   U99 : INV_X1 port map( A => A_s(11), ZN => n328);
   U100 : OAI221_X1 port map( B1 => n216, B2 => n329, C1 => n213, C2 => n331, A
                           => n148, ZN => O_13_port);
   U101 : INV_X1 port map( A => A_ns(12), ZN => n329);
   U102 : INV_X1 port map( A => A_s(12), ZN => n331);
   U103 : OAI221_X1 port map( B1 => n216, B2 => n330, C1 => n213, C2 => n332, A
                           => n147, ZN => O_14_port);
   U104 : INV_X1 port map( A => A_ns(13), ZN => n330);
   U105 : INV_X1 port map( A => A_s(13), ZN => n332);
   U106 : OAI221_X1 port map( B1 => n216, B2 => n333, C1 => n213, C2 => n334, A
                           => n146, ZN => O_15_port);
   U107 : INV_X1 port map( A => A_ns(14), ZN => n333);
   U108 : INV_X1 port map( A => A_s(14), ZN => n334);
   U109 : INV_X1 port map( A => n141, ZN => O_1_port);
   U110 : AOI22_X1 port map( A1 => n203, A2 => A_s(0), B1 => n202, B2 => 
                           A_ns(0), ZN => n141);
   U111 : OAI221_X1 port map( B1 => n216, B2 => n309, C1 => n214, C2 => n310, A
                           => n130, ZN => O_2_port);
   U112 : INV_X1 port map( A => A_ns(1), ZN => n309);
   U113 : INV_X1 port map( A => A_s(1), ZN => n310);
   U114 : OAI221_X1 port map( B1 => n215, B2 => n311, C1 => n213, C2 => n313, A
                           => n119, ZN => O_3_port);
   U115 : INV_X1 port map( A => A_ns(2), ZN => n311);
   U116 : INV_X1 port map( A => A_s(2), ZN => n313);
   U117 : OAI221_X1 port map( B1 => n216, B2 => n312, C1 => n213, C2 => n314, A
                           => n107, ZN => O_4_port);
   U118 : INV_X1 port map( A => A_ns(3), ZN => n312);
   U119 : INV_X1 port map( A => A_s(3), ZN => n314);
   U120 : OAI221_X1 port map( B1 => n216, B2 => n315, C1 => n213, C2 => n317, A
                           => n106, ZN => O_5_port);
   U121 : INV_X1 port map( A => A_ns(4), ZN => n315);
   U122 : INV_X1 port map( A => A_s(4), ZN => n317);
   U123 : OAI221_X1 port map( B1 => n216, B2 => n316, C1 => n213, C2 => n318, A
                           => n105, ZN => O_6_port);
   U124 : INV_X1 port map( A => A_ns(5), ZN => n316);
   U125 : INV_X1 port map( A => A_s(5), ZN => n318);
   U126 : OAI221_X1 port map( B1 => n216, B2 => n319, C1 => n213, C2 => n321, A
                           => n104, ZN => O_7_port);
   U127 : INV_X1 port map( A => A_ns(6), ZN => n319);
   U128 : INV_X1 port map( A => A_s(6), ZN => n321);
   U129 : INV_X1 port map( A => A_s(8), ZN => n324);
   U130 : INV_X1 port map( A => A_ns(8), ZN => n323);
   U131 : AOI22_X1 port map( A1 => A_s(0), A2 => n208, B1 => A_ns(0), B2 => 
                           n212, ZN => n130);
   U132 : AOI22_X1 port map( A1 => A_s(1), A2 => n209, B1 => A_ns(1), B2 => 
                           n211, ZN => n119);
   U133 : AOI22_X1 port map( A1 => A_s(2), A2 => n210, B1 => A_ns(2), B2 => 
                           n211, ZN => n107);
   U134 : AOI22_X1 port map( A1 => A_s(3), A2 => n210, B1 => A_ns(3), B2 => 
                           n211, ZN => n106);
   U135 : AOI22_X1 port map( A1 => A_s(4), A2 => n210, B1 => A_ns(4), B2 => 
                           n211, ZN => n105);
   U136 : AOI22_X1 port map( A1 => A_s(5), A2 => n210, B1 => A_ns(5), B2 => 
                           n211, ZN => n104);
   U137 : AOI22_X1 port map( A1 => A_s(6), A2 => n210, B1 => A_ns(6), B2 => 
                           n211, ZN => n103);
   U138 : AOI22_X1 port map( A1 => A_s(9), A2 => n207, B1 => A_ns(9), B2 => 
                           n211, ZN => n150);
   U139 : AOI22_X1 port map( A1 => A_s(10), A2 => n207, B1 => A_ns(10), B2 => 
                           n211, ZN => n149);
   U140 : AOI22_X1 port map( A1 => A_s(11), A2 => n207, B1 => A_ns(11), B2 => 
                           n211, ZN => n148);
   U141 : AOI22_X1 port map( A1 => A_s(12), A2 => n207, B1 => A_ns(12), B2 => 
                           n211, ZN => n147);
   U142 : AOI22_X1 port map( A1 => A_s(13), A2 => n207, B1 => A_ns(13), B2 => 
                           n211, ZN => n146);
   U143 : INV_X1 port map( A => n204, ZN => n211);
   U144 : INV_X1 port map( A => n203, ZN => n213);
   U145 : INV_X1 port map( A => n218, ZN => A_nso_18_port);
   U146 : INV_X1 port map( A => A_ns(16), ZN => n218);
   U147 : INV_X1 port map( A => A_ns(17), ZN => n219);
   U148 : INV_X1 port map( A => n221, ZN => A_nso_20_port);
   U149 : INV_X1 port map( A => A_ns(18), ZN => n221);
   U150 : INV_X1 port map( A => A_ns(19), ZN => n222);
   U151 : INV_X1 port map( A => A_ns(20), ZN => n223);
   U152 : INV_X1 port map( A => n225, ZN => A_nso_23_port);
   U153 : INV_X1 port map( A => A_ns(21), ZN => n225);
   U154 : INV_X1 port map( A => n227, ZN => A_nso_24_port);
   U155 : INV_X1 port map( A => A_ns(22), ZN => n227);
   U156 : INV_X1 port map( A => n229, ZN => A_nso_25_port);
   U157 : INV_X1 port map( A => A_ns(23), ZN => n229);
   U158 : INV_X1 port map( A => n231, ZN => A_nso_26_port);
   U159 : INV_X1 port map( A => A_ns(24), ZN => n231);
   U160 : INV_X1 port map( A => n233, ZN => A_nso_27_port);
   U161 : INV_X1 port map( A => A_ns(25), ZN => n233);
   U162 : INV_X1 port map( A => n235, ZN => A_nso_28_port);
   U163 : INV_X1 port map( A => A_ns(26), ZN => n235);
   U164 : INV_X1 port map( A => n237, ZN => A_nso_29_port);
   U165 : INV_X1 port map( A => A_ns(27), ZN => n237);
   U166 : INV_X1 port map( A => n239, ZN => A_nso_30_port);
   U167 : INV_X1 port map( A => A_ns(28), ZN => n239);
   U168 : INV_X1 port map( A => n241, ZN => A_nso_31_port);
   U169 : INV_X1 port map( A => A_ns(29), ZN => n241);
   U170 : INV_X1 port map( A => n243, ZN => A_nso_32_port);
   U171 : INV_X1 port map( A => A_ns(30), ZN => n243);
   U172 : INV_X1 port map( A => n245, ZN => A_nso_33_port);
   U173 : INV_X1 port map( A => A_ns(31), ZN => n245);
   U174 : INV_X1 port map( A => n247, ZN => A_nso_34_port);
   U175 : INV_X1 port map( A => A_ns(32), ZN => n247);
   U176 : INV_X1 port map( A => A_ns(33), ZN => n248);
   U177 : INV_X1 port map( A => A_ns(34), ZN => n249);
   U178 : INV_X1 port map( A => A_ns(35), ZN => n250);
   U179 : INV_X1 port map( A => A_ns(36), ZN => n251);
   U180 : INV_X1 port map( A => A_ns(37), ZN => n252);
   U181 : INV_X1 port map( A => A_ns(38), ZN => n253);
   U182 : INV_X1 port map( A => A_ns(39), ZN => n254);
   U183 : INV_X1 port map( A => A_ns(40), ZN => n255);
   U184 : INV_X1 port map( A => A_ns(41), ZN => n256);
   U185 : INV_X1 port map( A => A_ns(42), ZN => n257);
   U186 : INV_X1 port map( A => A_ns(43), ZN => n258);
   U187 : INV_X1 port map( A => A_ns(44), ZN => n259);
   U188 : INV_X1 port map( A => A_ns(45), ZN => n260);
   U189 : INV_X1 port map( A => A_ns(46), ZN => n261);
   U190 : INV_X1 port map( A => n264, ZN => A_nso_17_port);
   U191 : INV_X1 port map( A => A_ns(15), ZN => n264);
   U192 : INV_X1 port map( A => n266, ZN => A_so_17_port);
   U193 : INV_X1 port map( A => A_s(15), ZN => n266);
   U194 : INV_X1 port map( A => n268, ZN => A_so_18_port);
   U195 : INV_X1 port map( A => A_s(16), ZN => n268);
   U196 : INV_X1 port map( A => n270, ZN => A_so_19_port);
   U197 : INV_X1 port map( A => A_s(17), ZN => n270);
   U198 : INV_X1 port map( A => n272, ZN => A_so_20_port);
   U199 : INV_X1 port map( A => A_s(18), ZN => n272);
   U202 : INV_X1 port map( A => n274, ZN => A_so_21_port);
   U203 : INV_X1 port map( A => A_s(19), ZN => n274);
   U204 : INV_X1 port map( A => n276, ZN => A_so_22_port);
   U205 : INV_X1 port map( A => A_s(20), ZN => n276);
   U206 : INV_X1 port map( A => n278, ZN => A_so_23_port);
   U207 : INV_X1 port map( A => A_s(21), ZN => n278);
   U208 : INV_X1 port map( A => A_s(22), ZN => n279);
   U209 : INV_X1 port map( A => A_s(23), ZN => n280);
   U210 : INV_X1 port map( A => A_s(24), ZN => n281);
   U211 : INV_X1 port map( A => A_s(25), ZN => n282);
   U212 : INV_X1 port map( A => A_s(26), ZN => n283);
   U213 : INV_X1 port map( A => A_s(27), ZN => n284);
   U214 : INV_X1 port map( A => n286, ZN => A_so_30_port);
   U215 : INV_X1 port map( A => A_s(28), ZN => n286);
   U216 : INV_X1 port map( A => A_s(29), ZN => n287);
   U217 : INV_X1 port map( A => A_s(30), ZN => n288);
   U218 : INV_X1 port map( A => A_s(31), ZN => n289);
   U219 : INV_X1 port map( A => A_s(32), ZN => n290);
   U220 : INV_X1 port map( A => A_s(33), ZN => n291);
   U221 : INV_X1 port map( A => A_s(34), ZN => n292);
   U222 : INV_X1 port map( A => A_s(35), ZN => n293);
   U223 : INV_X1 port map( A => A_s(36), ZN => n294);
   U224 : INV_X1 port map( A => A_s(37), ZN => n295);
   U225 : INV_X1 port map( A => A_s(38), ZN => n296);
   U226 : INV_X1 port map( A => n298, ZN => A_so_41_port);
   U227 : INV_X1 port map( A => A_s(39), ZN => n298);
   U228 : INV_X1 port map( A => n300, ZN => A_so_42_port);
   U229 : INV_X1 port map( A => A_s(40), ZN => n300);
   U230 : INV_X1 port map( A => A_s(41), ZN => n301);
   U231 : INV_X1 port map( A => A_s(42), ZN => n302);
   U232 : INV_X1 port map( A => A_s(43), ZN => n303);
   U233 : INV_X1 port map( A => A_s(44), ZN => n304);
   U234 : INV_X1 port map( A => A_s(45), ZN => n305);
   U235 : INV_X1 port map( A => A_s(46), ZN => n306);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT48_i14 is

   port( A_s, A_ns, B : in std_logic_vector (47 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (47 downto 0));

end BOOTHENC_NBIT48_i14;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT48_i14 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105
      , n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
      n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, 
      n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, 
      n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
      n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, 
      n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, 
      n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, 
      n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, 
      n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, 
      n214, n215, n216, n217, O_2_port, n219, O_1_port, O_3_port, n222, 
      O_4_port, n224, O_5_port, n226, O_6_port, n228, O_7_port, n230, O_8_port,
      n232, O_9_port, n234, O_10_port, n236, O_11_port, n238, O_12_port, n240, 
      O_13_port, n242, O_14_port, n244, O_45_port, O_46_port, n247, O_47_port, 
      n249, O_44_port, n251, O_43_port, n253, O_42_port, n255, O_41_port, n257,
      O_40_port, n259, O_39_port, n261, O_38_port, n263, O_37_port, n265, 
      O_36_port, n267, O_35_port, n269, O_34_port, n271, O_33_port, n273, 
      O_32_port, n275, O_31_port, n277, O_30_port, n279, O_29_port, n281, 
      O_28_port, n283, O_27_port, n285, O_26_port, n287, O_25_port, n289, 
      O_24_port, n291, O_23_port, n293, O_22_port, n295, O_21_port, n297, 
      O_20_port, n299, O_19_port, n301, O_18_port, n303, O_17_port, n305, 
      O_16_port, n307, O_15_port, n309, n310, n311, n312 : std_logic;

begin
   O <= ( O_47_port, O_46_port, O_45_port, O_44_port, O_43_port, O_42_port, 
      O_41_port, O_40_port, O_39_port, O_38_port, O_37_port, O_36_port, 
      O_35_port, O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, 
      O_29_port, O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, 
      O_23_port, O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, 
      O_17_port, O_16_port, O_15_port, O_14_port, O_13_port, O_12_port, 
      O_11_port, O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, 
      O_4_port, O_3_port, O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), 
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   A_nso <= ( A_ns(45), A_ns(44), A_ns(43), A_ns(42), A_ns(41), A_ns(40), 
      A_ns(39), A_ns(38), A_ns(37), A_ns(36), A_ns(35), A_ns(34), A_ns(33), 
      A_ns(32), A_ns(31), A_ns(30), A_ns(29), A_ns(28), A_ns(27), A_ns(26), 
      A_ns(25), A_ns(24), A_ns(23), A_ns(22), A_ns(21), A_ns(20), A_ns(19), 
      A_ns(18), A_ns(17), A_ns(16), A_ns(15), A_ns(14), A_ns(13), A_ns(12), 
      A_ns(11), A_ns(10), A_ns(9), A_ns(8), A_ns(7), A_ns(6), A_ns(5), A_ns(4),
      A_ns(3), A_ns(2), A_ns(1), A_ns(0), X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U194 : XOR2_X1 port map( A => B(13), B => B(14), Z => n193);
   U2 : BUF_X1 port map( A => n195, Z => n199);
   U3 : BUF_X1 port map( A => n195, Z => n198);
   U4 : BUF_X1 port map( A => n194, Z => n197);
   U5 : BUF_X1 port map( A => n194, Z => n196);
   U6 : BUF_X1 port map( A => n213, Z => n217);
   U7 : BUF_X1 port map( A => n311, Z => n195);
   U8 : BUF_X1 port map( A => n213, Z => n216);
   U9 : BUF_X1 port map( A => n212, Z => n215);
   U10 : BUF_X1 port map( A => n311, Z => n194);
   U11 : BUF_X1 port map( A => n212, Z => n214);
   U12 : BUF_X1 port map( A => n207, Z => n211);
   U13 : BUF_X1 port map( A => n201, Z => n205);
   U14 : BUF_X1 port map( A => n97, Z => n213);
   U15 : INV_X1 port map( A => n192, ZN => n311);
   U16 : BUF_X1 port map( A => n207, Z => n210);
   U17 : BUF_X1 port map( A => n201, Z => n204);
   U18 : BUF_X1 port map( A => n206, Z => n209);
   U19 : BUF_X1 port map( A => n200, Z => n203);
   U20 : BUF_X1 port map( A => n97, Z => n212);
   U21 : BUF_X1 port map( A => n206, Z => n208);
   U22 : BUF_X1 port map( A => n200, Z => n202);
   U23 : INV_X1 port map( A => n118, ZN => O_47_port);
   U24 : AOI221_X1 port map( B1 => n211, B2 => A_s(45), C1 => n205, C2 => 
                           A_ns(45), A => n249, ZN => n118);
   U25 : INV_X1 port map( A => n119, ZN => n249);
   U26 : INV_X1 port map( A => n120, ZN => O_46_port);
   U27 : AOI221_X1 port map( B1 => n214, B2 => A_ns(45), C1 => n196, C2 => 
                           A_s(45), A => n247, ZN => n120);
   U28 : INV_X1 port map( A => n121, ZN => n247);
   U29 : NAND2_X1 port map( A1 => n193, A2 => n312, ZN => n192);
   U30 : BUF_X1 port map( A => n100, Z => n201);
   U31 : BUF_X1 port map( A => n99, Z => n207);
   U32 : AND2_X1 port map( A1 => n193, A2 => n192, ZN => n97);
   U33 : AOI22_X1 port map( A1 => A_ns(46), A2 => n214, B1 => A_s(46), B2 => 
                           n196, ZN => n119);
   U34 : BUF_X1 port map( A => n100, Z => n200);
   U35 : BUF_X1 port map( A => n99, Z => n206);
   U36 : INV_X1 port map( A => n122, ZN => O_45_port);
   U37 : AOI221_X1 port map( B1 => n214, B2 => A_ns(44), C1 => n197, C2 => 
                           A_s(44), A => n251, ZN => n122);
   U38 : INV_X1 port map( A => n123, ZN => n251);
   U39 : INV_X1 port map( A => n124, ZN => O_44_port);
   U40 : AOI221_X1 port map( B1 => n214, B2 => A_ns(43), C1 => n197, C2 => 
                           A_s(43), A => n253, ZN => n124);
   U41 : INV_X1 port map( A => n125, ZN => n253);
   U42 : INV_X1 port map( A => n126, ZN => O_43_port);
   U43 : AOI221_X1 port map( B1 => n215, B2 => A_ns(42), C1 => n197, C2 => 
                           A_s(42), A => n255, ZN => n126);
   U44 : INV_X1 port map( A => n127, ZN => n255);
   U45 : INV_X1 port map( A => n128, ZN => O_42_port);
   U46 : AOI221_X1 port map( B1 => n215, B2 => A_ns(41), C1 => n197, C2 => 
                           A_s(41), A => n257, ZN => n128);
   U47 : INV_X1 port map( A => n129, ZN => n257);
   U48 : INV_X1 port map( A => n130, ZN => O_41_port);
   U49 : AOI221_X1 port map( B1 => n215, B2 => A_ns(40), C1 => n197, C2 => 
                           A_s(40), A => n259, ZN => n130);
   U50 : INV_X1 port map( A => n131, ZN => n259);
   U51 : INV_X1 port map( A => n132, ZN => O_40_port);
   U52 : AOI221_X1 port map( B1 => n215, B2 => A_ns(39), C1 => n197, C2 => 
                           A_s(39), A => n261, ZN => n132);
   U53 : INV_X1 port map( A => n133, ZN => n261);
   U54 : INV_X1 port map( A => n134, ZN => O_39_port);
   U55 : AOI221_X1 port map( B1 => n215, B2 => A_ns(38), C1 => n197, C2 => 
                           A_s(38), A => n263, ZN => n134);
   U56 : INV_X1 port map( A => n135, ZN => n263);
   U57 : INV_X1 port map( A => n136, ZN => O_38_port);
   U58 : AOI221_X1 port map( B1 => n215, B2 => A_ns(37), C1 => n197, C2 => 
                           A_s(37), A => n265, ZN => n136);
   U59 : INV_X1 port map( A => n137, ZN => n265);
   U60 : INV_X1 port map( A => n138, ZN => O_37_port);
   U61 : AOI221_X1 port map( B1 => n215, B2 => A_ns(36), C1 => n197, C2 => 
                           A_s(36), A => n267, ZN => n138);
   U62 : INV_X1 port map( A => n139, ZN => n267);
   U63 : INV_X1 port map( A => n140, ZN => O_36_port);
   U64 : AOI221_X1 port map( B1 => n215, B2 => A_ns(35), C1 => n197, C2 => 
                           A_s(35), A => n269, ZN => n140);
   U65 : INV_X1 port map( A => n141, ZN => n269);
   U66 : INV_X1 port map( A => n142, ZN => O_35_port);
   U67 : AOI221_X1 port map( B1 => n215, B2 => A_ns(34), C1 => n197, C2 => 
                           A_s(34), A => n271, ZN => n142);
   U68 : INV_X1 port map( A => n143, ZN => n271);
   U69 : INV_X1 port map( A => n180, ZN => O_17_port);
   U70 : AOI221_X1 port map( B1 => n217, B2 => A_ns(16), C1 => n199, C2 => 
                           A_s(16), A => n307, ZN => n180);
   U71 : INV_X1 port map( A => n181, ZN => n307);
   U72 : INV_X1 port map( A => n178, ZN => O_18_port);
   U73 : AOI221_X1 port map( B1 => n217, B2 => A_ns(17), C1 => n199, C2 => 
                           A_s(17), A => n305, ZN => n178);
   U74 : INV_X1 port map( A => n179, ZN => n305);
   U75 : INV_X1 port map( A => n176, ZN => O_19_port);
   U76 : AOI221_X1 port map( B1 => n217, B2 => A_ns(18), C1 => n199, C2 => 
                           A_s(18), A => n303, ZN => n176);
   U77 : INV_X1 port map( A => n177, ZN => n303);
   U78 : INV_X1 port map( A => n174, ZN => O_20_port);
   U79 : AOI221_X1 port map( B1 => n216, B2 => A_ns(19), C1 => n199, C2 => 
                           A_s(19), A => n301, ZN => n174);
   U80 : INV_X1 port map( A => n175, ZN => n301);
   U81 : INV_X1 port map( A => n172, ZN => O_21_port);
   U82 : AOI221_X1 port map( B1 => n216, B2 => A_ns(20), C1 => n199, C2 => 
                           A_s(20), A => n299, ZN => n172);
   U83 : INV_X1 port map( A => n173, ZN => n299);
   U84 : INV_X1 port map( A => n170, ZN => O_22_port);
   U85 : AOI221_X1 port map( B1 => n216, B2 => A_ns(21), C1 => n198, C2 => 
                           A_s(21), A => n297, ZN => n170);
   U86 : INV_X1 port map( A => n171, ZN => n297);
   U87 : INV_X1 port map( A => n168, ZN => O_23_port);
   U88 : AOI221_X1 port map( B1 => n216, B2 => A_ns(22), C1 => n198, C2 => 
                           A_s(22), A => n295, ZN => n168);
   U89 : INV_X1 port map( A => n169, ZN => n295);
   U90 : INV_X1 port map( A => n166, ZN => O_24_port);
   U91 : AOI221_X1 port map( B1 => n216, B2 => A_ns(23), C1 => n198, C2 => 
                           A_s(23), A => n293, ZN => n166);
   U92 : INV_X1 port map( A => n167, ZN => n293);
   U93 : INV_X1 port map( A => n164, ZN => O_25_port);
   U94 : AOI221_X1 port map( B1 => n216, B2 => A_ns(24), C1 => n198, C2 => 
                           A_s(24), A => n291, ZN => n164);
   U95 : INV_X1 port map( A => n165, ZN => n291);
   U96 : INV_X1 port map( A => n162, ZN => O_26_port);
   U97 : AOI221_X1 port map( B1 => n216, B2 => A_ns(25), C1 => n198, C2 => 
                           A_s(25), A => n289, ZN => n162);
   U98 : INV_X1 port map( A => n163, ZN => n289);
   U99 : INV_X1 port map( A => n160, ZN => O_27_port);
   U100 : AOI221_X1 port map( B1 => n216, B2 => A_ns(26), C1 => n198, C2 => 
                           A_s(26), A => n287, ZN => n160);
   U101 : INV_X1 port map( A => n161, ZN => n287);
   U102 : INV_X1 port map( A => n158, ZN => O_28_port);
   U103 : AOI221_X1 port map( B1 => n216, B2 => A_ns(27), C1 => n198, C2 => 
                           A_s(27), A => n285, ZN => n158);
   U104 : INV_X1 port map( A => n159, ZN => n285);
   U105 : INV_X1 port map( A => n156, ZN => O_29_port);
   U106 : AOI221_X1 port map( B1 => n216, B2 => A_ns(28), C1 => n198, C2 => 
                           A_s(28), A => n283, ZN => n156);
   U107 : INV_X1 port map( A => n157, ZN => n283);
   U108 : INV_X1 port map( A => n152, ZN => O_30_port);
   U109 : AOI221_X1 port map( B1 => n216, B2 => A_ns(29), C1 => n198, C2 => 
                           A_s(29), A => n281, ZN => n152);
   U110 : INV_X1 port map( A => n153, ZN => n281);
   U111 : INV_X1 port map( A => n150, ZN => O_31_port);
   U112 : AOI221_X1 port map( B1 => n216, B2 => A_ns(30), C1 => n198, C2 => 
                           A_s(30), A => n279, ZN => n150);
   U113 : INV_X1 port map( A => n151, ZN => n279);
   U114 : INV_X1 port map( A => n148, ZN => O_32_port);
   U115 : AOI221_X1 port map( B1 => n215, B2 => A_ns(31), C1 => n198, C2 => 
                           A_s(31), A => n277, ZN => n148);
   U116 : INV_X1 port map( A => n149, ZN => n277);
   U117 : INV_X1 port map( A => n146, ZN => O_33_port);
   U118 : AOI221_X1 port map( B1 => n215, B2 => A_ns(32), C1 => n198, C2 => 
                           A_s(32), A => n275, ZN => n146);
   U119 : INV_X1 port map( A => n147, ZN => n275);
   U120 : INV_X1 port map( A => n144, ZN => O_34_port);
   U121 : AOI221_X1 port map( B1 => n215, B2 => A_ns(33), C1 => n197, C2 => 
                           A_s(33), A => n273, ZN => n144);
   U122 : INV_X1 port map( A => n145, ZN => n273);
   U123 : INV_X1 port map( A => n182, ZN => O_16_port);
   U124 : AOI221_X1 port map( B1 => n217, B2 => A_ns(15), C1 => n199, C2 => 
                           A_s(15), A => n309, ZN => n182);
   U125 : INV_X1 port map( A => n183, ZN => n309);
   U126 : INV_X1 port map( A => n184, ZN => O_15_port);
   U127 : INV_X1 port map( A => n185, ZN => n310);
   U128 : INV_X1 port map( A => n186, ZN => O_14_port);
   U129 : INV_X1 port map( A => n187, ZN => n244);
   U130 : AOI22_X1 port map( A1 => A_s(19), A2 => n211, B1 => A_ns(19), B2 => 
                           n205, ZN => n173);
   U131 : AOI22_X1 port map( A1 => A_s(21), A2 => n210, B1 => A_ns(21), B2 => 
                           n204, ZN => n169);
   U132 : AOI22_X1 port map( A1 => A_s(22), A2 => n210, B1 => A_ns(22), B2 => 
                           n204, ZN => n167);
   U133 : AOI22_X1 port map( A1 => A_s(23), A2 => n210, B1 => A_ns(23), B2 => 
                           n204, ZN => n165);
   U134 : AOI22_X1 port map( A1 => A_s(15), A2 => n211, B1 => A_ns(15), B2 => 
                           n205, ZN => n181);
   U135 : AOI22_X1 port map( A1 => A_s(16), A2 => n211, B1 => A_ns(16), B2 => 
                           n205, ZN => n179);
   U136 : AOI22_X1 port map( A1 => A_s(18), A2 => n211, B1 => A_ns(18), B2 => 
                           n205, ZN => n175);
   U137 : AOI22_X1 port map( A1 => A_s(20), A2 => n210, B1 => A_ns(20), B2 => 
                           n204, ZN => n171);
   U138 : AOI22_X1 port map( A1 => A_s(17), A2 => n211, B1 => A_ns(17), B2 => 
                           n205, ZN => n177);
   U139 : NOR3_X1 port map( A1 => B(13), A2 => B(14), A3 => n312, ZN => n100);
   U140 : INV_X1 port map( A => B(15), ZN => n312);
   U141 : AND3_X1 port map( A1 => B(13), A2 => n312, A3 => B(14), ZN => n99);
   U142 : AOI22_X1 port map( A1 => A_s(24), A2 => n210, B1 => A_ns(24), B2 => 
                           n204, ZN => n163);
   U143 : AOI22_X1 port map( A1 => A_s(25), A2 => n210, B1 => A_ns(25), B2 => 
                           n204, ZN => n161);
   U144 : AOI22_X1 port map( A1 => A_s(26), A2 => n210, B1 => A_ns(26), B2 => 
                           n204, ZN => n159);
   U145 : AOI22_X1 port map( A1 => A_s(27), A2 => n210, B1 => A_ns(27), B2 => 
                           n204, ZN => n157);
   U146 : AOI22_X1 port map( A1 => A_s(28), A2 => n210, B1 => A_ns(28), B2 => 
                           n204, ZN => n153);
   U147 : AOI22_X1 port map( A1 => A_s(29), A2 => n210, B1 => A_ns(29), B2 => 
                           n204, ZN => n151);
   U148 : AOI22_X1 port map( A1 => A_s(41), A2 => n209, B1 => A_ns(41), B2 => 
                           n203, ZN => n127);
   U149 : AOI22_X1 port map( A1 => A_s(42), A2 => n208, B1 => A_ns(42), B2 => 
                           n202, ZN => n125);
   U150 : AOI22_X1 port map( A1 => A_s(43), A2 => n208, B1 => A_ns(43), B2 => 
                           n202, ZN => n123);
   U151 : AOI22_X1 port map( A1 => A_s(44), A2 => n208, B1 => A_ns(44), B2 => 
                           n202, ZN => n121);
   U152 : AOI22_X1 port map( A1 => A_s(32), A2 => n209, B1 => A_ns(32), B2 => 
                           n203, ZN => n145);
   U153 : AOI22_X1 port map( A1 => A_s(30), A2 => n210, B1 => A_ns(30), B2 => 
                           n204, ZN => n149);
   U154 : AOI22_X1 port map( A1 => A_s(31), A2 => n209, B1 => A_ns(31), B2 => 
                           n203, ZN => n147);
   U155 : AOI22_X1 port map( A1 => A_s(33), A2 => n209, B1 => A_ns(33), B2 => 
                           n203, ZN => n143);
   U156 : AOI22_X1 port map( A1 => A_s(34), A2 => n209, B1 => A_ns(34), B2 => 
                           n203, ZN => n141);
   U157 : AOI22_X1 port map( A1 => A_s(35), A2 => n209, B1 => A_ns(35), B2 => 
                           n203, ZN => n139);
   U158 : AOI22_X1 port map( A1 => A_s(36), A2 => n209, B1 => A_ns(36), B2 => 
                           n203, ZN => n137);
   U159 : AOI22_X1 port map( A1 => A_s(37), A2 => n209, B1 => A_ns(37), B2 => 
                           n203, ZN => n135);
   U160 : AOI22_X1 port map( A1 => A_s(38), A2 => n209, B1 => A_ns(38), B2 => 
                           n203, ZN => n133);
   U161 : AOI22_X1 port map( A1 => A_s(39), A2 => n209, B1 => A_ns(39), B2 => 
                           n203, ZN => n131);
   U162 : AOI22_X1 port map( A1 => A_s(40), A2 => n209, B1 => A_ns(40), B2 => 
                           n203, ZN => n129);
   U163 : INV_X1 port map( A => n112, ZN => O_8_port);
   U164 : AOI221_X1 port map( B1 => n214, B2 => A_ns(7), C1 => n196, C2 => 
                           A_s(7), A => n232, ZN => n112);
   U165 : INV_X1 port map( A => n113, ZN => n232);
   U166 : INV_X1 port map( A => n103, ZN => O_9_port);
   U167 : AOI221_X1 port map( B1 => n214, B2 => A_ns(8), C1 => n196, C2 => 
                           A_s(8), A => n234, ZN => n103);
   U168 : INV_X1 port map( A => n104, ZN => n234);
   U169 : INV_X1 port map( A => n190, ZN => O_10_port);
   U170 : AOI221_X1 port map( B1 => n214, B2 => A_ns(9), C1 => n196, C2 => 
                           A_s(9), A => n236, ZN => n190);
   U171 : INV_X1 port map( A => n191, ZN => n236);
   U172 : INV_X1 port map( A => n101, ZN => O_11_port);
   U173 : AOI221_X1 port map( B1 => n214, B2 => A_ns(10), C1 => n196, C2 => 
                           A_s(10), A => n238, ZN => n101);
   U174 : INV_X1 port map( A => n102, ZN => n238);
   U175 : INV_X1 port map( A => n188, ZN => O_12_port);
   U176 : AOI221_X1 port map( B1 => A_ns(11), B2 => n217, C1 => A_s(11), C2 => 
                           n196, A => n240, ZN => n188);
   U177 : INV_X1 port map( A => n189, ZN => n240);
   U178 : INV_X1 port map( A => n96, ZN => O_13_port);
   U179 : AOI221_X1 port map( B1 => n215, B2 => A_ns(12), C1 => n197, C2 => 
                           A_s(12), A => n242, ZN => n96);
   U180 : INV_X1 port map( A => n98, ZN => n242);
   U181 : INV_X1 port map( A => n111, ZN => O_1_port);
   U182 : AOI22_X1 port map( A1 => n196, A2 => A_s(0), B1 => n217, B2 => 
                           A_ns(0), ZN => n111);
   U183 : INV_X1 port map( A => n154, ZN => O_2_port);
   U184 : AOI221_X1 port map( B1 => n216, B2 => A_ns(1), C1 => n198, C2 => 
                           A_s(1), A => n219, ZN => n154);
   U185 : INV_X1 port map( A => n155, ZN => n219);
   U186 : INV_X1 port map( A => n109, ZN => O_3_port);
   U187 : AOI221_X1 port map( B1 => n214, B2 => A_ns(2), C1 => n196, C2 => 
                           A_s(2), A => n222, ZN => n109);
   U188 : INV_X1 port map( A => n110, ZN => n222);
   U189 : INV_X1 port map( A => n116, ZN => O_4_port);
   U190 : AOI221_X1 port map( B1 => n214, B2 => A_ns(3), C1 => n196, C2 => 
                           A_s(3), A => n224, ZN => n116);
   U191 : INV_X1 port map( A => n117, ZN => n224);
   U192 : INV_X1 port map( A => n107, ZN => O_5_port);
   U193 : AOI221_X1 port map( B1 => n214, B2 => A_ns(4), C1 => n196, C2 => 
                           A_s(4), A => n226, ZN => n107);
   U195 : INV_X1 port map( A => n108, ZN => n226);
   U196 : INV_X1 port map( A => n114, ZN => O_6_port);
   U197 : AOI221_X1 port map( B1 => n214, B2 => A_ns(5), C1 => n196, C2 => 
                           A_s(5), A => n228, ZN => n114);
   U198 : INV_X1 port map( A => n115, ZN => n228);
   U199 : INV_X1 port map( A => n105, ZN => O_7_port);
   U200 : AOI221_X1 port map( B1 => n214, B2 => A_ns(6), C1 => n196, C2 => 
                           A_s(6), A => n230, ZN => n105);
   U201 : INV_X1 port map( A => n106, ZN => n230);
   U202 : AOI22_X1 port map( A1 => A_s(0), A2 => n210, B1 => A_ns(0), B2 => 
                           n204, ZN => n155);
   U203 : AOI22_X1 port map( A1 => A_s(1), A2 => n208, B1 => A_ns(1), B2 => 
                           n202, ZN => n110);
   U204 : AOI22_X1 port map( A1 => A_s(2), A2 => n208, B1 => A_ns(2), B2 => 
                           n202, ZN => n117);
   U205 : AOI22_X1 port map( A1 => A_s(3), A2 => n208, B1 => A_ns(3), B2 => 
                           n202, ZN => n108);
   U206 : AOI22_X1 port map( A1 => A_s(4), A2 => n208, B1 => A_ns(4), B2 => 
                           n202, ZN => n115);
   U207 : AOI22_X1 port map( A1 => A_s(5), A2 => n208, B1 => A_ns(5), B2 => 
                           n202, ZN => n106);
   U208 : AOI22_X1 port map( A1 => A_s(6), A2 => n208, B1 => A_ns(6), B2 => 
                           n202, ZN => n113);
   U209 : AOI22_X1 port map( A1 => A_s(7), A2 => n208, B1 => A_ns(7), B2 => 
                           n202, ZN => n104);
   U210 : AOI22_X1 port map( A1 => A_s(8), A2 => n208, B1 => A_ns(8), B2 => 
                           n202, ZN => n191);
   U211 : AOI22_X1 port map( A1 => A_s(9), A2 => n208, B1 => A_ns(9), B2 => 
                           n202, ZN => n102);
   U212 : AOI22_X1 port map( A1 => A_s(10), A2 => n211, B1 => A_ns(10), B2 => 
                           n205, ZN => n189);
   U213 : AOI22_X1 port map( A1 => A_s(11), A2 => n209, B1 => A_ns(11), B2 => 
                           n203, ZN => n98);
   U214 : AOI22_X1 port map( A1 => A_s(12), A2 => n211, B1 => A_ns(12), B2 => 
                           n205, ZN => n187);
   U215 : AOI221_X1 port map( B1 => n217, B2 => A_ns(14), C1 => n199, C2 => 
                           A_s(14), A => n310, ZN => n184);
   U216 : AOI22_X1 port map( A1 => A_s(14), A2 => n211, B1 => A_ns(14), B2 => 
                           n205, ZN => n183);
   U217 : AOI221_X1 port map( B1 => n217, B2 => A_ns(13), C1 => n199, C2 => 
                           A_s(13), A => n244, ZN => n186);
   U218 : AOI22_X1 port map( A1 => A_s(13), A2 => n211, B1 => A_ns(13), B2 => 
                           n205, ZN => n185);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT46_i12 is

   port( A_s, A_ns, B : in std_logic_vector (45 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (45 downto 0));

end BOOTHENC_NBIT46_i12;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT46_i12 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, 
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, 
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, 
      n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, 
      O_2_port, n211, O_1_port, O_3_port, n214, O_4_port, n216, O_5_port, n218,
      O_6_port, n220, O_7_port, n222, O_8_port, n224, O_9_port, n226, O_10_port
      , n228, O_11_port, n230, O_12_port, n232, O_43_port, O_44_port, n235, 
      O_45_port, n237, O_42_port, n239, O_41_port, n241, O_40_port, n243, 
      O_39_port, n245, O_38_port, n247, O_37_port, n249, O_36_port, n251, 
      O_35_port, n253, O_34_port, n255, O_33_port, n257, O_32_port, n259, 
      O_31_port, n261, O_30_port, n263, O_29_port, n265, O_28_port, n267, 
      O_27_port, n269, O_26_port, n271, O_25_port, n273, O_24_port, n275, 
      O_23_port, n277, O_22_port, n279, O_21_port, n281, O_20_port, n283, 
      O_19_port, n285, O_18_port, n287, O_17_port, n289, O_16_port, n291, 
      O_15_port, n293, O_14_port, n295, O_13_port, n297, n298, n299, n300 : 
      std_logic;

begin
   O <= ( O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, O_40_port, 
      O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, 
      O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, 
      O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, 
      O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, O_16_port, 
      O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, O_10_port, 
      O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, O_3_port, 
      O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), A_s(38), A_s(37), 
      A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), A_s(30), A_s(29), 
      A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), A_s(22), A_s(21), 
      A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), A_s(14), A_s(13), 
      A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), A_s(6), A_s(5), A_s(4)
      , A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, X_Logic0_port );
   A_nso <= ( A_ns(43), A_ns(42), A_ns(41), A_ns(40), A_ns(39), A_ns(38), 
      A_ns(37), A_ns(36), A_ns(35), A_ns(34), A_ns(33), A_ns(32), A_ns(31), 
      A_ns(30), A_ns(29), A_ns(28), A_ns(27), A_ns(26), A_ns(25), A_ns(24), 
      A_ns(23), A_ns(22), A_ns(21), A_ns(20), A_ns(19), A_ns(18), A_ns(17), 
      A_ns(16), A_ns(15), A_ns(14), A_ns(13), A_ns(12), A_ns(11), A_ns(10), 
      A_ns(9), A_ns(8), A_ns(7), A_ns(6), A_ns(5), A_ns(4), A_ns(3), A_ns(2), 
      A_ns(1), A_ns(0), X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U186 : XOR2_X1 port map( A => B(11), B => B(12), Z => n185);
   U2 : BUF_X1 port map( A => n187, Z => n190);
   U3 : BUF_X1 port map( A => n186, Z => n188);
   U4 : BUF_X1 port map( A => n187, Z => n191);
   U5 : BUF_X1 port map( A => n186, Z => n189);
   U6 : BUF_X1 port map( A => n205, Z => n208);
   U7 : BUF_X1 port map( A => n205, Z => n209);
   U8 : BUF_X1 port map( A => n299, Z => n186);
   U9 : BUF_X1 port map( A => n299, Z => n187);
   U10 : BUF_X1 port map( A => n204, Z => n207);
   U11 : BUF_X1 port map( A => n204, Z => n206);
   U12 : BUF_X1 port map( A => n199, Z => n202);
   U13 : BUF_X1 port map( A => n193, Z => n196);
   U14 : BUF_X1 port map( A => n199, Z => n203);
   U15 : BUF_X1 port map( A => n193, Z => n197);
   U16 : BUF_X1 port map( A => n93, Z => n205);
   U17 : INV_X1 port map( A => n184, ZN => n299);
   U18 : BUF_X1 port map( A => n198, Z => n201);
   U19 : BUF_X1 port map( A => n192, Z => n195);
   U20 : BUF_X1 port map( A => n93, Z => n204);
   U21 : BUF_X1 port map( A => n198, Z => n200);
   U22 : BUF_X1 port map( A => n192, Z => n194);
   U23 : INV_X1 port map( A => n112, ZN => O_45_port);
   U24 : AOI221_X1 port map( B1 => n203, B2 => A_s(43), C1 => n197, C2 => 
                           A_ns(43), A => n237, ZN => n112);
   U25 : INV_X1 port map( A => n113, ZN => n237);
   U26 : INV_X1 port map( A => n114, ZN => O_44_port);
   U27 : AOI221_X1 port map( B1 => n206, B2 => A_ns(43), C1 => n188, C2 => 
                           A_s(43), A => n235, ZN => n114);
   U28 : INV_X1 port map( A => n115, ZN => n235);
   U29 : NAND2_X1 port map( A1 => n185, A2 => n300, ZN => n184);
   U30 : BUF_X1 port map( A => n96, Z => n193);
   U31 : BUF_X1 port map( A => n95, Z => n199);
   U32 : AND2_X1 port map( A1 => n185, A2 => n184, ZN => n93);
   U33 : AOI22_X1 port map( A1 => A_ns(44), A2 => n206, B1 => A_s(44), B2 => 
                           n188, ZN => n113);
   U34 : BUF_X1 port map( A => n96, Z => n192);
   U35 : BUF_X1 port map( A => n95, Z => n198);
   U36 : INV_X1 port map( A => n116, ZN => O_43_port);
   U37 : AOI221_X1 port map( B1 => n206, B2 => A_ns(42), C1 => n188, C2 => 
                           A_s(42), A => n239, ZN => n116);
   U38 : INV_X1 port map( A => n117, ZN => n239);
   U39 : INV_X1 port map( A => n118, ZN => O_42_port);
   U40 : AOI221_X1 port map( B1 => n206, B2 => A_ns(41), C1 => n189, C2 => 
                           A_s(41), A => n241, ZN => n118);
   U41 : INV_X1 port map( A => n119, ZN => n241);
   U42 : INV_X1 port map( A => n120, ZN => O_41_port);
   U43 : AOI221_X1 port map( B1 => n206, B2 => A_ns(40), C1 => n189, C2 => 
                           A_s(40), A => n243, ZN => n120);
   U44 : INV_X1 port map( A => n121, ZN => n243);
   U45 : INV_X1 port map( A => n122, ZN => O_40_port);
   U46 : AOI221_X1 port map( B1 => n206, B2 => A_ns(39), C1 => n189, C2 => 
                           A_s(39), A => n245, ZN => n122);
   U47 : INV_X1 port map( A => n123, ZN => n245);
   U48 : INV_X1 port map( A => n126, ZN => O_38_port);
   U49 : AOI221_X1 port map( B1 => n207, B2 => A_ns(37), C1 => n189, C2 => 
                           A_s(37), A => n249, ZN => n126);
   U50 : INV_X1 port map( A => n127, ZN => n249);
   U51 : INV_X1 port map( A => n128, ZN => O_37_port);
   U52 : AOI221_X1 port map( B1 => n207, B2 => A_ns(36), C1 => n189, C2 => 
                           A_s(36), A => n251, ZN => n128);
   U53 : INV_X1 port map( A => n129, ZN => n251);
   U54 : INV_X1 port map( A => n174, ZN => O_15_port);
   U55 : AOI221_X1 port map( B1 => n209, B2 => A_ns(14), C1 => n191, C2 => 
                           A_s(14), A => n295, ZN => n174);
   U56 : INV_X1 port map( A => n175, ZN => n295);
   U57 : INV_X1 port map( A => n172, ZN => O_16_port);
   U58 : AOI221_X1 port map( B1 => n208, B2 => A_ns(15), C1 => n191, C2 => 
                           A_s(15), A => n293, ZN => n172);
   U59 : INV_X1 port map( A => n173, ZN => n293);
   U60 : INV_X1 port map( A => n170, ZN => O_17_port);
   U61 : AOI221_X1 port map( B1 => n208, B2 => A_ns(16), C1 => n191, C2 => 
                           A_s(16), A => n291, ZN => n170);
   U62 : INV_X1 port map( A => n171, ZN => n291);
   U63 : INV_X1 port map( A => n168, ZN => O_18_port);
   U64 : AOI221_X1 port map( B1 => n208, B2 => A_ns(17), C1 => n191, C2 => 
                           A_s(17), A => n289, ZN => n168);
   U65 : INV_X1 port map( A => n169, ZN => n289);
   U66 : INV_X1 port map( A => n166, ZN => O_19_port);
   U67 : AOI221_X1 port map( B1 => n208, B2 => A_ns(18), C1 => n190, C2 => 
                           A_s(18), A => n287, ZN => n166);
   U68 : INV_X1 port map( A => n167, ZN => n287);
   U69 : INV_X1 port map( A => n164, ZN => O_20_port);
   U70 : AOI221_X1 port map( B1 => n208, B2 => A_ns(19), C1 => n190, C2 => 
                           A_s(19), A => n285, ZN => n164);
   U71 : INV_X1 port map( A => n165, ZN => n285);
   U72 : INV_X1 port map( A => n162, ZN => O_21_port);
   U73 : AOI221_X1 port map( B1 => n208, B2 => A_ns(20), C1 => n190, C2 => 
                           A_s(20), A => n283, ZN => n162);
   U74 : INV_X1 port map( A => n163, ZN => n283);
   U75 : INV_X1 port map( A => n160, ZN => O_22_port);
   U76 : AOI221_X1 port map( B1 => n208, B2 => A_ns(21), C1 => n190, C2 => 
                           A_s(21), A => n281, ZN => n160);
   U77 : INV_X1 port map( A => n161, ZN => n281);
   U78 : INV_X1 port map( A => n158, ZN => O_23_port);
   U79 : AOI221_X1 port map( B1 => n208, B2 => A_ns(22), C1 => n190, C2 => 
                           A_s(22), A => n279, ZN => n158);
   U80 : INV_X1 port map( A => n159, ZN => n279);
   U81 : INV_X1 port map( A => n156, ZN => O_24_port);
   U82 : AOI221_X1 port map( B1 => n208, B2 => A_ns(23), C1 => n190, C2 => 
                           A_s(23), A => n277, ZN => n156);
   U83 : INV_X1 port map( A => n157, ZN => n277);
   U84 : INV_X1 port map( A => n154, ZN => O_25_port);
   U85 : AOI221_X1 port map( B1 => n208, B2 => A_ns(24), C1 => n190, C2 => 
                           A_s(24), A => n275, ZN => n154);
   U86 : INV_X1 port map( A => n155, ZN => n275);
   U87 : INV_X1 port map( A => n152, ZN => O_26_port);
   U88 : AOI221_X1 port map( B1 => n208, B2 => A_ns(25), C1 => n190, C2 => 
                           A_s(25), A => n273, ZN => n152);
   U89 : INV_X1 port map( A => n153, ZN => n273);
   U90 : INV_X1 port map( A => n150, ZN => O_27_port);
   U91 : AOI221_X1 port map( B1 => n208, B2 => A_ns(26), C1 => n190, C2 => 
                           A_s(26), A => n271, ZN => n150);
   U92 : INV_X1 port map( A => n151, ZN => n271);
   U93 : INV_X1 port map( A => n148, ZN => O_28_port);
   U94 : AOI221_X1 port map( B1 => n208, B2 => A_ns(27), C1 => n190, C2 => 
                           A_s(27), A => n269, ZN => n148);
   U95 : INV_X1 port map( A => n149, ZN => n269);
   U96 : INV_X1 port map( A => n146, ZN => O_29_port);
   U97 : AOI221_X1 port map( B1 => n207, B2 => A_ns(28), C1 => n190, C2 => 
                           A_s(28), A => n267, ZN => n146);
   U98 : INV_X1 port map( A => n147, ZN => n267);
   U99 : INV_X1 port map( A => n142, ZN => O_30_port);
   U100 : AOI221_X1 port map( B1 => n207, B2 => A_ns(29), C1 => n190, C2 => 
                           A_s(29), A => n265, ZN => n142);
   U101 : INV_X1 port map( A => n143, ZN => n265);
   U102 : INV_X1 port map( A => n140, ZN => O_31_port);
   U103 : AOI221_X1 port map( B1 => n207, B2 => A_ns(30), C1 => n189, C2 => 
                           A_s(30), A => n263, ZN => n140);
   U104 : INV_X1 port map( A => n141, ZN => n263);
   U105 : INV_X1 port map( A => n138, ZN => O_32_port);
   U106 : AOI221_X1 port map( B1 => n207, B2 => A_ns(31), C1 => n189, C2 => 
                           A_s(31), A => n261, ZN => n138);
   U107 : INV_X1 port map( A => n139, ZN => n261);
   U108 : INV_X1 port map( A => n136, ZN => O_33_port);
   U109 : AOI221_X1 port map( B1 => n207, B2 => A_ns(32), C1 => n189, C2 => 
                           A_s(32), A => n259, ZN => n136);
   U110 : INV_X1 port map( A => n137, ZN => n259);
   U111 : INV_X1 port map( A => n134, ZN => O_34_port);
   U112 : AOI221_X1 port map( B1 => n207, B2 => A_ns(33), C1 => n189, C2 => 
                           A_s(33), A => n257, ZN => n134);
   U113 : INV_X1 port map( A => n135, ZN => n257);
   U114 : INV_X1 port map( A => n124, ZN => O_39_port);
   U115 : AOI221_X1 port map( B1 => n207, B2 => A_ns(38), C1 => n189, C2 => 
                           A_s(38), A => n247, ZN => n124);
   U116 : INV_X1 port map( A => n125, ZN => n247);
   U117 : INV_X1 port map( A => n130, ZN => O_36_port);
   U118 : AOI221_X1 port map( B1 => n207, B2 => A_ns(35), C1 => n189, C2 => 
                           A_s(35), A => n253, ZN => n130);
   U119 : INV_X1 port map( A => n131, ZN => n253);
   U120 : INV_X1 port map( A => n132, ZN => O_35_port);
   U121 : AOI221_X1 port map( B1 => n207, B2 => A_ns(34), C1 => n189, C2 => 
                           A_s(34), A => n255, ZN => n132);
   U122 : INV_X1 port map( A => n133, ZN => n255);
   U123 : INV_X1 port map( A => n176, ZN => O_14_port);
   U124 : AOI221_X1 port map( B1 => n209, B2 => A_ns(13), C1 => n191, C2 => 
                           A_s(13), A => n297, ZN => n176);
   U125 : INV_X1 port map( A => n177, ZN => n297);
   U126 : INV_X1 port map( A => n178, ZN => O_13_port);
   U127 : INV_X1 port map( A => n179, ZN => n298);
   U128 : INV_X1 port map( A => n180, ZN => O_12_port);
   U129 : INV_X1 port map( A => n181, ZN => n232);
   U130 : AOI22_X1 port map( A1 => A_s(17), A2 => n203, B1 => A_ns(17), B2 => 
                           n197, ZN => n167);
   U131 : AOI22_X1 port map( A1 => A_s(19), A2 => n202, B1 => A_ns(19), B2 => 
                           n196, ZN => n163);
   U132 : AOI22_X1 port map( A1 => A_s(20), A2 => n202, B1 => A_ns(20), B2 => 
                           n196, ZN => n161);
   U133 : AOI22_X1 port map( A1 => A_s(21), A2 => n202, B1 => A_ns(21), B2 => 
                           n196, ZN => n159);
   U134 : AOI22_X1 port map( A1 => A_s(22), A2 => n202, B1 => A_ns(22), B2 => 
                           n196, ZN => n157);
   U135 : AOI22_X1 port map( A1 => A_s(23), A2 => n202, B1 => A_ns(23), B2 => 
                           n196, ZN => n155);
   U136 : AOI22_X1 port map( A1 => A_s(24), A2 => n202, B1 => A_ns(24), B2 => 
                           n196, ZN => n153);
   U137 : AOI22_X1 port map( A1 => A_s(25), A2 => n202, B1 => A_ns(25), B2 => 
                           n196, ZN => n151);
   U138 : AOI22_X1 port map( A1 => A_s(26), A2 => n202, B1 => A_ns(26), B2 => 
                           n196, ZN => n149);
   U139 : AOI22_X1 port map( A1 => A_s(27), A2 => n202, B1 => A_ns(27), B2 => 
                           n196, ZN => n147);
   U140 : AOI22_X1 port map( A1 => A_s(13), A2 => n203, B1 => A_ns(13), B2 => 
                           n197, ZN => n175);
   U141 : AOI22_X1 port map( A1 => A_s(14), A2 => n202, B1 => A_ns(14), B2 => 
                           n196, ZN => n173);
   U142 : AOI22_X1 port map( A1 => A_s(16), A2 => n203, B1 => A_ns(16), B2 => 
                           n197, ZN => n169);
   U143 : AOI22_X1 port map( A1 => A_s(18), A2 => n202, B1 => A_ns(18), B2 => 
                           n196, ZN => n165);
   U144 : AOI22_X1 port map( A1 => A_s(28), A2 => n201, B1 => A_ns(28), B2 => 
                           n195, ZN => n143);
   U145 : AOI22_X1 port map( A1 => A_s(29), A2 => n201, B1 => A_ns(29), B2 => 
                           n195, ZN => n141);
   U146 : AOI22_X1 port map( A1 => A_s(15), A2 => n203, B1 => A_ns(15), B2 => 
                           n197, ZN => n171);
   U147 : NOR3_X1 port map( A1 => B(11), A2 => B(12), A3 => n300, ZN => n96);
   U148 : INV_X1 port map( A => B(13), ZN => n300);
   U149 : AND3_X1 port map( A1 => B(11), A2 => n300, A3 => B(12), ZN => n95);
   U150 : AOI22_X1 port map( A1 => A_s(39), A2 => n200, B1 => A_ns(39), B2 => 
                           n194, ZN => n121);
   U151 : AOI22_X1 port map( A1 => A_s(40), A2 => n200, B1 => A_ns(40), B2 => 
                           n194, ZN => n119);
   U152 : AOI22_X1 port map( A1 => A_s(41), A2 => n200, B1 => A_ns(41), B2 => 
                           n194, ZN => n117);
   U153 : AOI22_X1 port map( A1 => A_s(42), A2 => n200, B1 => A_ns(42), B2 => 
                           n194, ZN => n115);
   U154 : AOI22_X1 port map( A1 => A_s(30), A2 => n201, B1 => A_ns(30), B2 => 
                           n195, ZN => n139);
   U155 : AOI22_X1 port map( A1 => A_s(31), A2 => n201, B1 => A_ns(31), B2 => 
                           n195, ZN => n137);
   U156 : AOI22_X1 port map( A1 => A_s(32), A2 => n201, B1 => A_ns(32), B2 => 
                           n195, ZN => n135);
   U157 : AOI22_X1 port map( A1 => A_s(33), A2 => n201, B1 => A_ns(33), B2 => 
                           n195, ZN => n133);
   U158 : AOI22_X1 port map( A1 => A_s(34), A2 => n201, B1 => A_ns(34), B2 => 
                           n195, ZN => n131);
   U159 : AOI22_X1 port map( A1 => A_s(35), A2 => n201, B1 => A_ns(35), B2 => 
                           n195, ZN => n129);
   U160 : AOI22_X1 port map( A1 => A_s(36), A2 => n201, B1 => A_ns(36), B2 => 
                           n195, ZN => n127);
   U161 : AOI22_X1 port map( A1 => A_s(37), A2 => n201, B1 => A_ns(37), B2 => 
                           n195, ZN => n125);
   U162 : AOI22_X1 port map( A1 => A_s(38), A2 => n201, B1 => A_ns(38), B2 => 
                           n195, ZN => n123);
   U163 : INV_X1 port map( A => n106, ZN => O_8_port);
   U164 : AOI221_X1 port map( B1 => n206, B2 => A_ns(7), C1 => n188, C2 => 
                           A_s(7), A => n224, ZN => n106);
   U165 : INV_X1 port map( A => n107, ZN => n224);
   U166 : INV_X1 port map( A => n97, ZN => O_9_port);
   U167 : AOI221_X1 port map( B1 => n206, B2 => A_ns(8), C1 => n188, C2 => 
                           A_s(8), A => n226, ZN => n97);
   U168 : INV_X1 port map( A => n98, ZN => n226);
   U169 : INV_X1 port map( A => n182, ZN => O_10_port);
   U170 : AOI221_X1 port map( B1 => A_ns(9), B2 => n209, C1 => A_s(9), C2 => 
                           n188, A => n228, ZN => n182);
   U171 : INV_X1 port map( A => n183, ZN => n228);
   U172 : INV_X1 port map( A => n92, ZN => O_11_port);
   U173 : AOI221_X1 port map( B1 => n207, B2 => A_ns(10), C1 => n189, C2 => 
                           A_s(10), A => n230, ZN => n92);
   U174 : INV_X1 port map( A => n94, ZN => n230);
   U175 : INV_X1 port map( A => n105, ZN => O_1_port);
   U176 : AOI22_X1 port map( A1 => n188, A2 => A_s(0), B1 => n209, B2 => 
                           A_ns(0), ZN => n105);
   U177 : INV_X1 port map( A => n144, ZN => O_2_port);
   U178 : AOI221_X1 port map( B1 => n207, B2 => A_ns(1), C1 => n190, C2 => 
                           A_s(1), A => n211, ZN => n144);
   U179 : INV_X1 port map( A => n145, ZN => n211);
   U180 : INV_X1 port map( A => n103, ZN => O_3_port);
   U181 : AOI221_X1 port map( B1 => n206, B2 => A_ns(2), C1 => n188, C2 => 
                           A_s(2), A => n214, ZN => n103);
   U182 : INV_X1 port map( A => n104, ZN => n214);
   U183 : INV_X1 port map( A => n110, ZN => O_4_port);
   U184 : AOI221_X1 port map( B1 => n206, B2 => A_ns(3), C1 => n188, C2 => 
                           A_s(3), A => n216, ZN => n110);
   U185 : INV_X1 port map( A => n111, ZN => n216);
   U187 : INV_X1 port map( A => n101, ZN => O_5_port);
   U188 : AOI221_X1 port map( B1 => n206, B2 => A_ns(4), C1 => n188, C2 => 
                           A_s(4), A => n218, ZN => n101);
   U189 : INV_X1 port map( A => n102, ZN => n218);
   U190 : INV_X1 port map( A => n108, ZN => O_6_port);
   U191 : AOI221_X1 port map( B1 => n206, B2 => A_ns(5), C1 => n188, C2 => 
                           A_s(5), A => n220, ZN => n108);
   U192 : INV_X1 port map( A => n109, ZN => n220);
   U193 : INV_X1 port map( A => n99, ZN => O_7_port);
   U194 : AOI221_X1 port map( B1 => n206, B2 => A_ns(6), C1 => n188, C2 => 
                           A_s(6), A => n222, ZN => n99);
   U195 : INV_X1 port map( A => n100, ZN => n222);
   U196 : AOI22_X1 port map( A1 => A_s(0), A2 => n202, B1 => A_ns(0), B2 => 
                           n196, ZN => n145);
   U197 : AOI22_X1 port map( A1 => A_s(1), A2 => n200, B1 => A_ns(1), B2 => 
                           n194, ZN => n104);
   U198 : AOI22_X1 port map( A1 => A_s(2), A2 => n200, B1 => A_ns(2), B2 => 
                           n194, ZN => n111);
   U199 : AOI22_X1 port map( A1 => A_s(3), A2 => n200, B1 => A_ns(3), B2 => 
                           n194, ZN => n102);
   U200 : AOI22_X1 port map( A1 => A_s(4), A2 => n200, B1 => A_ns(4), B2 => 
                           n194, ZN => n109);
   U201 : AOI22_X1 port map( A1 => A_s(5), A2 => n200, B1 => A_ns(5), B2 => 
                           n194, ZN => n100);
   U202 : AOI22_X1 port map( A1 => A_s(6), A2 => n200, B1 => A_ns(6), B2 => 
                           n194, ZN => n107);
   U203 : AOI22_X1 port map( A1 => A_s(7), A2 => n200, B1 => A_ns(7), B2 => 
                           n194, ZN => n98);
   U204 : AOI22_X1 port map( A1 => A_s(8), A2 => n200, B1 => A_ns(8), B2 => 
                           n194, ZN => n183);
   U205 : AOI22_X1 port map( A1 => A_s(9), A2 => n201, B1 => A_ns(9), B2 => 
                           n195, ZN => n94);
   U206 : AOI22_X1 port map( A1 => A_s(10), A2 => n203, B1 => A_ns(10), B2 => 
                           n197, ZN => n181);
   U207 : AOI221_X1 port map( B1 => n209, B2 => A_ns(12), C1 => n191, C2 => 
                           A_s(12), A => n298, ZN => n178);
   U208 : AOI22_X1 port map( A1 => A_s(12), A2 => n203, B1 => A_ns(12), B2 => 
                           n197, ZN => n177);
   U209 : AOI221_X1 port map( B1 => n209, B2 => A_ns(11), C1 => n188, C2 => 
                           A_s(11), A => n232, ZN => n180);
   U210 : AOI22_X1 port map( A1 => A_s(11), A2 => n203, B1 => A_ns(11), B2 => 
                           n197, ZN => n179);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT44_i10 is

   port( A_s, A_ns, B : in std_logic_vector (43 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (43 downto 0));

end BOOTHENC_NBIT44_i10;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT44_i10 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
      n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, 
      n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, 
      n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, 
      n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, O_2_port, n203, O_1_port, 
      O_3_port, n206, O_4_port, n208, O_5_port, n210, O_6_port, n212, O_7_port,
      n214, O_8_port, n216, O_9_port, n218, O_10_port, n220, O_41_port, 
      O_42_port, n223, O_43_port, n225, O_40_port, n227, O_39_port, n229, 
      O_38_port, n231, O_37_port, n233, O_36_port, n235, O_35_port, n237, 
      O_34_port, n239, O_33_port, n241, O_32_port, n243, O_31_port, n245, 
      O_30_port, n247, O_29_port, n249, O_28_port, n251, O_27_port, n253, 
      O_26_port, n255, O_25_port, n257, O_24_port, n259, O_23_port, n261, 
      O_22_port, n263, O_21_port, n265, O_20_port, n267, O_19_port, n269, 
      O_18_port, n271, O_17_port, n273, O_16_port, n275, O_15_port, n277, 
      O_14_port, n279, O_13_port, n281, O_12_port, n283, O_11_port, n285, n286,
      n287, n288 : std_logic;

begin
   O <= ( O_43_port, O_42_port, O_41_port, O_40_port, O_39_port, O_38_port, 
      O_37_port, O_36_port, O_35_port, O_34_port, O_33_port, O_32_port, 
      O_31_port, O_30_port, O_29_port, O_28_port, O_27_port, O_26_port, 
      O_25_port, O_24_port, O_23_port, O_22_port, O_21_port, O_20_port, 
      O_19_port, O_18_port, O_17_port, O_16_port, O_15_port, O_14_port, 
      O_13_port, O_12_port, O_11_port, O_10_port, O_9_port, O_8_port, O_7_port,
      O_6_port, O_5_port, O_4_port, O_3_port, O_2_port, O_1_port, X_Logic0_port
      );
   A_so <= ( A_s(41), A_s(40), A_s(39), A_s(38), A_s(37), A_s(36), A_s(35), 
      A_s(34), A_s(33), A_s(32), A_s(31), A_s(30), A_s(29), A_s(28), A_s(27), 
      A_s(26), A_s(25), A_s(24), A_s(23), A_s(22), A_s(21), A_s(20), A_s(19), 
      A_s(18), A_s(17), A_s(16), A_s(15), A_s(14), A_s(13), A_s(12), A_s(11), 
      A_s(10), A_s(9), A_s(8), A_s(7), A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), 
      A_s(1), A_s(0), X_Logic0_port, X_Logic0_port );
   A_nso <= ( A_ns(41), A_ns(40), A_ns(39), A_ns(38), A_ns(37), A_ns(36), 
      A_ns(35), A_ns(34), A_ns(33), A_ns(32), A_ns(31), A_ns(30), A_ns(29), 
      A_ns(28), A_ns(27), A_ns(26), A_ns(25), A_ns(24), A_ns(23), A_ns(22), 
      A_ns(21), A_ns(20), A_ns(19), A_ns(18), A_ns(17), A_ns(16), A_ns(15), 
      A_ns(14), A_ns(13), A_ns(12), A_ns(11), A_ns(10), A_ns(9), A_ns(8), 
      A_ns(7), A_ns(6), A_ns(5), A_ns(4), A_ns(3), A_ns(2), A_ns(1), A_ns(0), 
      X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U178 : XOR2_X1 port map( A => B(10), B => B(9), Z => n177);
   U2 : BUF_X1 port map( A => n196, Z => n198);
   U3 : BUF_X1 port map( A => n178, Z => n180);
   U4 : CLKBUF_X1 port map( A => n178, Z => n181);
   U5 : CLKBUF_X1 port map( A => n196, Z => n199);
   U6 : CLKBUF_X1 port map( A => n287, Z => n179);
   U7 : CLKBUF_X1 port map( A => n89, Z => n197);
   U8 : BUF_X1 port map( A => n179, Z => n182);
   U9 : BUF_X1 port map( A => n179, Z => n183);
   U10 : BUF_X1 port map( A => n197, Z => n200);
   U11 : BUF_X1 port map( A => n197, Z => n201);
   U12 : BUF_X1 port map( A => n287, Z => n178);
   U13 : BUF_X1 port map( A => n191, Z => n194);
   U14 : BUF_X1 port map( A => n185, Z => n188);
   U15 : BUF_X1 port map( A => n191, Z => n195);
   U16 : BUF_X1 port map( A => n185, Z => n189);
   U17 : BUF_X1 port map( A => n89, Z => n196);
   U18 : INV_X1 port map( A => n176, ZN => n287);
   U19 : BUF_X1 port map( A => n190, Z => n193);
   U20 : BUF_X1 port map( A => n184, Z => n187);
   U21 : BUF_X1 port map( A => n190, Z => n192);
   U22 : BUF_X1 port map( A => n184, Z => n186);
   U23 : INV_X1 port map( A => n106, ZN => O_43_port);
   U24 : AOI221_X1 port map( B1 => n195, B2 => A_s(41), C1 => n189, C2 => 
                           A_ns(41), A => n225, ZN => n106);
   U25 : INV_X1 port map( A => n107, ZN => n225);
   U26 : INV_X1 port map( A => n108, ZN => O_42_port);
   U27 : AOI221_X1 port map( B1 => n198, B2 => A_ns(41), C1 => n180, C2 => 
                           A_s(41), A => n223, ZN => n108);
   U28 : INV_X1 port map( A => n109, ZN => n223);
   U29 : NAND2_X1 port map( A1 => n177, A2 => n288, ZN => n176);
   U30 : BUF_X1 port map( A => n92, Z => n185);
   U31 : BUF_X1 port map( A => n91, Z => n191);
   U32 : AND2_X1 port map( A1 => n177, A2 => n176, ZN => n89);
   U33 : AOI22_X1 port map( A1 => A_ns(42), A2 => n198, B1 => A_s(42), B2 => 
                           n180, ZN => n107);
   U34 : BUF_X1 port map( A => n92, Z => n184);
   U35 : BUF_X1 port map( A => n91, Z => n190);
   U36 : INV_X1 port map( A => n110, ZN => O_41_port);
   U37 : AOI221_X1 port map( B1 => n198, B2 => A_ns(40), C1 => n180, C2 => 
                           A_s(40), A => n227, ZN => n110);
   U38 : INV_X1 port map( A => n111, ZN => n227);
   U39 : INV_X1 port map( A => n112, ZN => O_40_port);
   U40 : AOI221_X1 port map( B1 => n198, B2 => A_ns(39), C1 => n180, C2 => 
                           A_s(39), A => n229, ZN => n112);
   U41 : INV_X1 port map( A => n113, ZN => n229);
   U42 : INV_X1 port map( A => n114, ZN => O_39_port);
   U43 : AOI221_X1 port map( B1 => n198, B2 => A_ns(38), C1 => n180, C2 => 
                           A_s(38), A => n231, ZN => n114);
   U44 : INV_X1 port map( A => n115, ZN => n231);
   U45 : INV_X1 port map( A => n116, ZN => O_38_port);
   U46 : AOI221_X1 port map( B1 => n198, B2 => A_ns(37), C1 => n181, C2 => 
                           A_s(37), A => n233, ZN => n116);
   U47 : INV_X1 port map( A => n117, ZN => n233);
   U48 : INV_X1 port map( A => n118, ZN => O_37_port);
   U49 : AOI221_X1 port map( B1 => n198, B2 => A_ns(36), C1 => n181, C2 => 
                           A_s(36), A => n235, ZN => n118);
   U50 : INV_X1 port map( A => n119, ZN => n235);
   U51 : INV_X1 port map( A => n120, ZN => O_36_port);
   U52 : AOI221_X1 port map( B1 => n199, B2 => A_ns(35), C1 => n181, C2 => 
                           A_s(35), A => n237, ZN => n120);
   U53 : INV_X1 port map( A => n121, ZN => n237);
   U54 : INV_X1 port map( A => n122, ZN => O_35_port);
   U55 : AOI221_X1 port map( B1 => n199, B2 => A_ns(34), C1 => n181, C2 => 
                           A_s(34), A => n239, ZN => n122);
   U56 : INV_X1 port map( A => n123, ZN => n239);
   U57 : INV_X1 port map( A => n124, ZN => O_34_port);
   U58 : AOI221_X1 port map( B1 => n199, B2 => A_ns(33), C1 => n181, C2 => 
                           A_s(33), A => n241, ZN => n124);
   U59 : INV_X1 port map( A => n125, ZN => n241);
   U60 : INV_X1 port map( A => n126, ZN => O_33_port);
   U61 : AOI221_X1 port map( B1 => n199, B2 => A_ns(32), C1 => n181, C2 => 
                           A_s(32), A => n243, ZN => n126);
   U62 : INV_X1 port map( A => n127, ZN => n243);
   U63 : INV_X1 port map( A => n164, ZN => O_15_port);
   U64 : AOI221_X1 port map( B1 => n200, B2 => A_ns(14), C1 => n182, C2 => 
                           A_s(14), A => n279, ZN => n164);
   U65 : INV_X1 port map( A => n165, ZN => n279);
   U66 : INV_X1 port map( A => n162, ZN => O_16_port);
   U67 : AOI221_X1 port map( B1 => n200, B2 => A_ns(15), C1 => n182, C2 => 
                           A_s(15), A => n277, ZN => n162);
   U68 : INV_X1 port map( A => n163, ZN => n277);
   U69 : INV_X1 port map( A => n160, ZN => O_17_port);
   U70 : AOI221_X1 port map( B1 => n200, B2 => A_ns(16), C1 => n182, C2 => 
                           A_s(16), A => n275, ZN => n160);
   U71 : INV_X1 port map( A => n161, ZN => n275);
   U72 : INV_X1 port map( A => n158, ZN => O_18_port);
   U73 : AOI221_X1 port map( B1 => n200, B2 => A_ns(17), C1 => n182, C2 => 
                           A_s(17), A => n273, ZN => n158);
   U74 : INV_X1 port map( A => n159, ZN => n273);
   U75 : INV_X1 port map( A => n156, ZN => O_19_port);
   U76 : AOI221_X1 port map( B1 => n200, B2 => A_ns(18), C1 => n182, C2 => 
                           A_s(18), A => n271, ZN => n156);
   U77 : INV_X1 port map( A => n157, ZN => n271);
   U78 : INV_X1 port map( A => n154, ZN => O_20_port);
   U79 : AOI221_X1 port map( B1 => n200, B2 => A_ns(19), C1 => n182, C2 => 
                           A_s(19), A => n269, ZN => n154);
   U80 : INV_X1 port map( A => n155, ZN => n269);
   U81 : INV_X1 port map( A => n152, ZN => O_21_port);
   U82 : AOI221_X1 port map( B1 => n200, B2 => A_ns(20), C1 => n182, C2 => 
                           A_s(20), A => n267, ZN => n152);
   U83 : INV_X1 port map( A => n153, ZN => n267);
   U84 : INV_X1 port map( A => n150, ZN => O_22_port);
   U85 : AOI221_X1 port map( B1 => n200, B2 => A_ns(21), C1 => n182, C2 => 
                           A_s(21), A => n265, ZN => n150);
   U86 : INV_X1 port map( A => n151, ZN => n265);
   U87 : INV_X1 port map( A => n148, ZN => O_23_port);
   U88 : AOI221_X1 port map( B1 => n200, B2 => A_ns(22), C1 => n182, C2 => 
                           A_s(22), A => n263, ZN => n148);
   U89 : INV_X1 port map( A => n149, ZN => n263);
   U90 : INV_X1 port map( A => n146, ZN => O_24_port);
   U91 : AOI221_X1 port map( B1 => n200, B2 => A_ns(23), C1 => n182, C2 => 
                           A_s(23), A => n261, ZN => n146);
   U92 : INV_X1 port map( A => n147, ZN => n261);
   U93 : INV_X1 port map( A => n144, ZN => O_25_port);
   U94 : AOI221_X1 port map( B1 => n200, B2 => A_ns(24), C1 => n182, C2 => 
                           A_s(24), A => n259, ZN => n144);
   U95 : INV_X1 port map( A => n145, ZN => n259);
   U96 : INV_X1 port map( A => n142, ZN => O_26_port);
   U97 : AOI221_X1 port map( B1 => n199, B2 => A_ns(25), C1 => n182, C2 => 
                           A_s(25), A => n257, ZN => n142);
   U98 : INV_X1 port map( A => n143, ZN => n257);
   U99 : INV_X1 port map( A => n140, ZN => O_27_port);
   U100 : AOI221_X1 port map( B1 => n199, B2 => A_ns(26), C1 => n182, C2 => 
                           A_s(26), A => n255, ZN => n140);
   U101 : INV_X1 port map( A => n141, ZN => n255);
   U102 : INV_X1 port map( A => n138, ZN => O_28_port);
   U103 : AOI221_X1 port map( B1 => n199, B2 => A_ns(27), C1 => n181, C2 => 
                           A_s(27), A => n253, ZN => n138);
   U104 : INV_X1 port map( A => n139, ZN => n253);
   U105 : INV_X1 port map( A => n136, ZN => O_29_port);
   U106 : AOI221_X1 port map( B1 => n199, B2 => A_ns(28), C1 => n181, C2 => 
                           A_s(28), A => n251, ZN => n136);
   U107 : INV_X1 port map( A => n137, ZN => n251);
   U108 : INV_X1 port map( A => n132, ZN => O_30_port);
   U109 : AOI221_X1 port map( B1 => n199, B2 => A_ns(29), C1 => n181, C2 => 
                           A_s(29), A => n249, ZN => n132);
   U110 : INV_X1 port map( A => n133, ZN => n249);
   U111 : INV_X1 port map( A => n130, ZN => O_31_port);
   U112 : AOI221_X1 port map( B1 => n199, B2 => A_ns(30), C1 => n181, C2 => 
                           A_s(30), A => n247, ZN => n130);
   U113 : INV_X1 port map( A => n131, ZN => n247);
   U114 : INV_X1 port map( A => n128, ZN => O_32_port);
   U115 : AOI221_X1 port map( B1 => n199, B2 => A_ns(31), C1 => n181, C2 => 
                           A_s(31), A => n245, ZN => n128);
   U116 : INV_X1 port map( A => n129, ZN => n245);
   U117 : INV_X1 port map( A => n168, ZN => O_13_port);
   U118 : AOI221_X1 port map( B1 => n201, B2 => A_ns(12), C1 => n183, C2 => 
                           A_s(12), A => n283, ZN => n168);
   U119 : INV_X1 port map( A => n169, ZN => n283);
   U120 : INV_X1 port map( A => n166, ZN => O_14_port);
   U121 : AOI221_X1 port map( B1 => n200, B2 => A_ns(13), C1 => n183, C2 => 
                           A_s(13), A => n281, ZN => n166);
   U122 : INV_X1 port map( A => n167, ZN => n281);
   U123 : INV_X1 port map( A => n170, ZN => O_12_port);
   U124 : AOI221_X1 port map( B1 => n201, B2 => A_ns(11), C1 => n183, C2 => 
                           A_s(11), A => n285, ZN => n170);
   U125 : INV_X1 port map( A => n171, ZN => n285);
   U126 : INV_X1 port map( A => n172, ZN => O_11_port);
   U127 : INV_X1 port map( A => n173, ZN => n286);
   U128 : INV_X1 port map( A => n174, ZN => O_10_port);
   U129 : INV_X1 port map( A => n175, ZN => n220);
   U130 : AOI22_X1 port map( A1 => A_s(15), A2 => n194, B1 => A_ns(15), B2 => 
                           n188, ZN => n161);
   U131 : AOI22_X1 port map( A1 => A_s(17), A2 => n194, B1 => A_ns(17), B2 => 
                           n188, ZN => n157);
   U132 : AOI22_X1 port map( A1 => A_s(18), A2 => n194, B1 => A_ns(18), B2 => 
                           n188, ZN => n155);
   U133 : AOI22_X1 port map( A1 => A_s(19), A2 => n194, B1 => A_ns(19), B2 => 
                           n188, ZN => n153);
   U134 : AOI22_X1 port map( A1 => A_s(20), A2 => n194, B1 => A_ns(20), B2 => 
                           n188, ZN => n151);
   U135 : AOI22_X1 port map( A1 => A_s(21), A2 => n194, B1 => A_ns(21), B2 => 
                           n188, ZN => n149);
   U136 : AOI22_X1 port map( A1 => A_s(22), A2 => n194, B1 => A_ns(22), B2 => 
                           n188, ZN => n147);
   U137 : AOI22_X1 port map( A1 => A_s(23), A2 => n194, B1 => A_ns(23), B2 => 
                           n188, ZN => n145);
   U138 : AOI22_X1 port map( A1 => A_s(24), A2 => n194, B1 => A_ns(24), B2 => 
                           n188, ZN => n143);
   U139 : AOI22_X1 port map( A1 => A_s(25), A2 => n194, B1 => A_ns(25), B2 => 
                           n188, ZN => n141);
   U140 : AOI22_X1 port map( A1 => A_s(11), A2 => n195, B1 => A_ns(11), B2 => 
                           n189, ZN => n169);
   U141 : AOI22_X1 port map( A1 => A_s(12), A2 => n195, B1 => A_ns(12), B2 => 
                           n189, ZN => n167);
   U142 : AOI22_X1 port map( A1 => A_s(14), A2 => n194, B1 => A_ns(14), B2 => 
                           n188, ZN => n163);
   U143 : AOI22_X1 port map( A1 => A_s(16), A2 => n194, B1 => A_ns(16), B2 => 
                           n188, ZN => n159);
   U144 : AOI22_X1 port map( A1 => A_s(28), A2 => n193, B1 => A_ns(28), B2 => 
                           n187, ZN => n133);
   U145 : AOI22_X1 port map( A1 => A_s(26), A2 => n193, B1 => A_ns(26), B2 => 
                           n187, ZN => n139);
   U146 : AOI22_X1 port map( A1 => A_s(27), A2 => n193, B1 => A_ns(27), B2 => 
                           n187, ZN => n137);
   U147 : AOI22_X1 port map( A1 => A_s(29), A2 => n193, B1 => A_ns(29), B2 => 
                           n187, ZN => n131);
   U148 : AOI22_X1 port map( A1 => A_s(30), A2 => n193, B1 => A_ns(30), B2 => 
                           n187, ZN => n129);
   U149 : AOI22_X1 port map( A1 => A_s(31), A2 => n193, B1 => A_ns(31), B2 => 
                           n187, ZN => n127);
   U150 : AOI22_X1 port map( A1 => A_s(32), A2 => n193, B1 => A_ns(32), B2 => 
                           n187, ZN => n125);
   U151 : AOI22_X1 port map( A1 => A_s(33), A2 => n193, B1 => A_ns(33), B2 => 
                           n187, ZN => n123);
   U152 : AOI22_X1 port map( A1 => A_s(34), A2 => n193, B1 => A_ns(34), B2 => 
                           n187, ZN => n121);
   U153 : AOI22_X1 port map( A1 => A_s(35), A2 => n193, B1 => A_ns(35), B2 => 
                           n187, ZN => n119);
   U154 : AOI22_X1 port map( A1 => A_s(13), A2 => n195, B1 => A_ns(13), B2 => 
                           n189, ZN => n165);
   U155 : NOR3_X1 port map( A1 => B(10), A2 => B(9), A3 => n288, ZN => n92);
   U156 : INV_X1 port map( A => B(11), ZN => n288);
   U157 : AND3_X1 port map( A1 => B(10), A2 => n288, A3 => B(9), ZN => n91);
   U158 : AOI22_X1 port map( A1 => A_s(37), A2 => n192, B1 => A_ns(37), B2 => 
                           n186, ZN => n115);
   U159 : AOI22_X1 port map( A1 => A_s(38), A2 => n192, B1 => A_ns(38), B2 => 
                           n186, ZN => n113);
   U160 : AOI22_X1 port map( A1 => A_s(39), A2 => n192, B1 => A_ns(39), B2 => 
                           n186, ZN => n111);
   U161 : AOI22_X1 port map( A1 => A_s(40), A2 => n192, B1 => A_ns(40), B2 => 
                           n186, ZN => n109);
   U162 : AOI22_X1 port map( A1 => A_s(36), A2 => n192, B1 => A_ns(36), B2 => 
                           n186, ZN => n117);
   U163 : INV_X1 port map( A => n100, ZN => O_8_port);
   U164 : AOI221_X1 port map( B1 => A_ns(7), B2 => n201, C1 => A_s(7), C2 => 
                           n180, A => n216, ZN => n100);
   U165 : INV_X1 port map( A => n101, ZN => n216);
   U166 : INV_X1 port map( A => n88, ZN => O_9_port);
   U167 : AOI221_X1 port map( B1 => n199, B2 => A_ns(8), C1 => n181, C2 => 
                           A_s(8), A => n218, ZN => n88);
   U168 : INV_X1 port map( A => n90, ZN => n218);
   U169 : INV_X1 port map( A => n99, ZN => O_1_port);
   U170 : AOI22_X1 port map( A1 => n180, A2 => A_s(0), B1 => n201, B2 => 
                           A_ns(0), ZN => n99);
   U171 : INV_X1 port map( A => n134, ZN => O_2_port);
   U172 : AOI221_X1 port map( B1 => n199, B2 => A_ns(1), C1 => n181, C2 => 
                           A_s(1), A => n203, ZN => n134);
   U173 : INV_X1 port map( A => n135, ZN => n203);
   U174 : INV_X1 port map( A => n97, ZN => O_3_port);
   U175 : AOI221_X1 port map( B1 => n198, B2 => A_ns(2), C1 => n180, C2 => 
                           A_s(2), A => n206, ZN => n97);
   U176 : INV_X1 port map( A => n98, ZN => n206);
   U177 : INV_X1 port map( A => n104, ZN => O_4_port);
   U179 : AOI221_X1 port map( B1 => n198, B2 => A_ns(3), C1 => n180, C2 => 
                           A_s(3), A => n208, ZN => n104);
   U180 : INV_X1 port map( A => n105, ZN => n208);
   U181 : INV_X1 port map( A => n95, ZN => O_5_port);
   U182 : AOI221_X1 port map( B1 => n198, B2 => A_ns(4), C1 => n180, C2 => 
                           A_s(4), A => n210, ZN => n95);
   U183 : INV_X1 port map( A => n96, ZN => n210);
   U184 : INV_X1 port map( A => n102, ZN => O_6_port);
   U185 : AOI221_X1 port map( B1 => n198, B2 => A_ns(5), C1 => n180, C2 => 
                           A_s(5), A => n212, ZN => n102);
   U186 : INV_X1 port map( A => n103, ZN => n212);
   U187 : INV_X1 port map( A => n93, ZN => O_7_port);
   U188 : AOI221_X1 port map( B1 => n198, B2 => A_ns(6), C1 => n180, C2 => 
                           A_s(6), A => n214, ZN => n93);
   U189 : INV_X1 port map( A => n94, ZN => n214);
   U190 : AOI22_X1 port map( A1 => A_s(0), A2 => n193, B1 => A_ns(0), B2 => 
                           n187, ZN => n135);
   U191 : AOI22_X1 port map( A1 => A_s(1), A2 => n192, B1 => A_ns(1), B2 => 
                           n186, ZN => n98);
   U192 : AOI22_X1 port map( A1 => A_s(2), A2 => n192, B1 => A_ns(2), B2 => 
                           n186, ZN => n105);
   U193 : AOI22_X1 port map( A1 => A_s(3), A2 => n192, B1 => A_ns(3), B2 => 
                           n186, ZN => n96);
   U194 : AOI22_X1 port map( A1 => A_s(4), A2 => n192, B1 => A_ns(4), B2 => 
                           n186, ZN => n103);
   U195 : AOI22_X1 port map( A1 => A_s(5), A2 => n192, B1 => A_ns(5), B2 => 
                           n186, ZN => n94);
   U196 : AOI22_X1 port map( A1 => A_s(6), A2 => n192, B1 => A_ns(6), B2 => 
                           n186, ZN => n101);
   U197 : AOI22_X1 port map( A1 => A_s(7), A2 => n193, B1 => A_ns(7), B2 => 
                           n187, ZN => n90);
   U198 : AOI22_X1 port map( A1 => A_s(8), A2 => n192, B1 => A_ns(8), B2 => 
                           n186, ZN => n175);
   U199 : AOI221_X1 port map( B1 => n200, B2 => A_ns(10), C1 => n183, C2 => 
                           A_s(10), A => n286, ZN => n172);
   U200 : AOI22_X1 port map( A1 => A_s(10), A2 => n195, B1 => A_ns(10), B2 => 
                           n189, ZN => n171);
   U201 : AOI221_X1 port map( B1 => n198, B2 => A_ns(9), C1 => n180, C2 => 
                           A_s(9), A => n220, ZN => n174);
   U202 : AOI22_X1 port map( A1 => A_s(9), A2 => n195, B1 => A_ns(9), B2 => 
                           n189, ZN => n173);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT42_i8 is

   port( A_s, A_ns, B : in std_logic_vector (41 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (41 downto 0));

end BOOTHENC_NBIT42_i8;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT42_i8 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
      n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, 
      n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, 
      n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, 
      n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, 
      n192, n193, O_2_port, n195, O_1_port, O_3_port, n198, O_4_port, n200, 
      O_5_port, n202, O_6_port, n204, O_7_port, n206, O_8_port, n208, O_39_port
      , O_40_port, n211, O_41_port, n213, O_38_port, n215, O_37_port, n217, 
      O_36_port, n219, O_35_port, n221, O_34_port, n223, O_33_port, n225, 
      O_32_port, n227, O_31_port, n229, O_30_port, n231, O_29_port, n233, 
      O_28_port, n235, O_27_port, n237, O_26_port, n239, O_25_port, n241, 
      O_24_port, n243, O_23_port, n245, O_22_port, n247, O_21_port, n249, 
      O_20_port, n251, O_19_port, n253, O_18_port, n255, O_17_port, n257, 
      O_16_port, n259, O_15_port, n261, O_14_port, n263, O_13_port, n265, 
      O_12_port, n267, O_11_port, n269, O_10_port, n271, n272, O_9_port, n274, 
      n275, n276 : std_logic;

begin
   O <= ( O_41_port, O_40_port, O_39_port, O_38_port, O_37_port, O_36_port, 
      O_35_port, O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, 
      O_29_port, O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, 
      O_23_port, O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, 
      O_17_port, O_16_port, O_15_port, O_14_port, O_13_port, O_12_port, 
      O_11_port, O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, 
      O_4_port, O_3_port, O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(39), A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), 
      A_s(32), A_s(31), A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), 
      A_s(24), A_s(23), A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), 
      A_s(16), A_s(15), A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), 
      A_s(8), A_s(7), A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), 
      X_Logic0_port, X_Logic0_port );
   A_nso <= ( A_ns(39), A_ns(38), A_ns(37), A_ns(36), A_ns(35), A_ns(34), 
      A_ns(33), A_ns(32), A_ns(31), A_ns(30), A_ns(29), A_ns(28), A_ns(27), 
      A_ns(26), A_ns(25), A_ns(24), A_ns(23), A_ns(22), A_ns(21), A_ns(20), 
      A_ns(19), A_ns(18), A_ns(17), A_ns(16), A_ns(15), A_ns(14), A_ns(13), 
      A_ns(12), A_ns(11), A_ns(10), A_ns(9), A_ns(8), A_ns(7), A_ns(6), A_ns(5)
      , A_ns(4), A_ns(3), A_ns(2), A_ns(1), A_ns(0), X_Logic0_port, 
      X_Logic0_port );
   
   X_Logic0_port <= '0';
   U170 : XOR2_X1 port map( A => B(7), B => B(8), Z => n169);
   U2 : INV_X1 port map( A => n166, ZN => O_10_port);
   U3 : CLKBUF_X1 port map( A => n189, Z => n193);
   U4 : CLKBUF_X1 port map( A => n170, Z => n173);
   U5 : CLKBUF_X1 port map( A => n275, Z => n171);
   U6 : CLKBUF_X1 port map( A => n188, Z => n191);
   U7 : CLKBUF_X1 port map( A => n85, Z => n189);
   U8 : CLKBUF_X1 port map( A => n182, Z => n185);
   U9 : CLKBUF_X1 port map( A => n176, Z => n179);
   U10 : CLKBUF_X1 port map( A => n88, Z => n177);
   U11 : CLKBUF_X1 port map( A => n87, Z => n183);
   U12 : BUF_X1 port map( A => n171, Z => n174);
   U13 : BUF_X1 port map( A => n170, Z => n172);
   U14 : BUF_X1 port map( A => n171, Z => n175);
   U15 : BUF_X1 port map( A => n189, Z => n192);
   U16 : BUF_X1 port map( A => n188, Z => n190);
   U17 : BUF_X1 port map( A => n275, Z => n170);
   U18 : BUF_X1 port map( A => n183, Z => n186);
   U19 : BUF_X1 port map( A => n177, Z => n180);
   U20 : BUF_X1 port map( A => n182, Z => n184);
   U21 : BUF_X1 port map( A => n176, Z => n178);
   U22 : BUF_X1 port map( A => n183, Z => n187);
   U23 : BUF_X1 port map( A => n177, Z => n181);
   U24 : BUF_X1 port map( A => n85, Z => n188);
   U25 : INV_X1 port map( A => n168, ZN => n275);
   U26 : INV_X1 port map( A => n102, ZN => O_41_port);
   U27 : AOI221_X1 port map( B1 => n187, B2 => A_s(39), C1 => n181, C2 => 
                           A_ns(39), A => n213, ZN => n102);
   U28 : INV_X1 port map( A => n103, ZN => n213);
   U29 : INV_X1 port map( A => n104, ZN => O_40_port);
   U30 : AOI221_X1 port map( B1 => n190, B2 => A_ns(39), C1 => n172, C2 => 
                           A_s(39), A => n211, ZN => n104);
   U31 : INV_X1 port map( A => n105, ZN => n211);
   U32 : AOI22_X1 port map( A1 => A_ns(40), A2 => n190, B1 => A_s(40), B2 => 
                           n172, ZN => n103);
   U33 : NAND2_X1 port map( A1 => n169, A2 => n276, ZN => n168);
   U34 : BUF_X1 port map( A => n88, Z => n176);
   U35 : BUF_X1 port map( A => n87, Z => n182);
   U36 : AND2_X1 port map( A1 => n169, A2 => n168, ZN => n85);
   U37 : INV_X1 port map( A => n106, ZN => O_39_port);
   U38 : AOI221_X1 port map( B1 => n190, B2 => A_ns(38), C1 => n172, C2 => 
                           A_s(38), A => n215, ZN => n106);
   U39 : INV_X1 port map( A => n107, ZN => n215);
   U40 : INV_X1 port map( A => n108, ZN => O_38_port);
   U41 : AOI221_X1 port map( B1 => n190, B2 => A_ns(37), C1 => n172, C2 => 
                           A_s(37), A => n217, ZN => n108);
   U42 : INV_X1 port map( A => n109, ZN => n217);
   U43 : INV_X1 port map( A => n110, ZN => O_37_port);
   U44 : AOI221_X1 port map( B1 => n190, B2 => A_ns(36), C1 => n172, C2 => 
                           A_s(36), A => n219, ZN => n110);
   U45 : INV_X1 port map( A => n111, ZN => n219);
   U46 : INV_X1 port map( A => n112, ZN => O_36_port);
   U47 : AOI221_X1 port map( B1 => n190, B2 => A_ns(35), C1 => n173, C2 => 
                           A_s(35), A => n221, ZN => n112);
   U48 : INV_X1 port map( A => n113, ZN => n221);
   U49 : INV_X1 port map( A => n116, ZN => O_34_port);
   U50 : AOI221_X1 port map( B1 => n191, B2 => A_ns(33), C1 => n173, C2 => 
                           A_s(33), A => n225, ZN => n116);
   U51 : INV_X1 port map( A => n117, ZN => n225);
   U52 : INV_X1 port map( A => n118, ZN => O_33_port);
   U53 : AOI221_X1 port map( B1 => n191, B2 => A_ns(32), C1 => n173, C2 => 
                           A_s(32), A => n227, ZN => n118);
   U54 : INV_X1 port map( A => n119, ZN => n227);
   U55 : INV_X1 port map( A => n164, ZN => O_11_port);
   U56 : AOI221_X1 port map( B1 => n192, B2 => A_ns(10), C1 => n175, C2 => 
                           A_s(10), A => n271, ZN => n164);
   U57 : INV_X1 port map( A => n165, ZN => n271);
   U58 : INV_X1 port map( A => n162, ZN => O_12_port);
   U59 : AOI221_X1 port map( B1 => n192, B2 => A_ns(11), C1 => n175, C2 => 
                           A_s(11), A => n269, ZN => n162);
   U60 : INV_X1 port map( A => n163, ZN => n269);
   U61 : INV_X1 port map( A => n160, ZN => O_13_port);
   U62 : AOI221_X1 port map( B1 => n192, B2 => A_ns(12), C1 => n174, C2 => 
                           A_s(12), A => n267, ZN => n160);
   U63 : INV_X1 port map( A => n161, ZN => n267);
   U64 : INV_X1 port map( A => n158, ZN => O_14_port);
   U65 : AOI221_X1 port map( B1 => n192, B2 => A_ns(13), C1 => n174, C2 => 
                           A_s(13), A => n265, ZN => n158);
   U66 : INV_X1 port map( A => n159, ZN => n265);
   U67 : INV_X1 port map( A => n156, ZN => O_15_port);
   U68 : AOI221_X1 port map( B1 => n192, B2 => A_ns(14), C1 => n174, C2 => 
                           A_s(14), A => n263, ZN => n156);
   U69 : INV_X1 port map( A => n157, ZN => n263);
   U70 : INV_X1 port map( A => n154, ZN => O_16_port);
   U71 : AOI221_X1 port map( B1 => n192, B2 => A_ns(15), C1 => n174, C2 => 
                           A_s(15), A => n261, ZN => n154);
   U72 : INV_X1 port map( A => n155, ZN => n261);
   U73 : INV_X1 port map( A => n152, ZN => O_17_port);
   U74 : AOI221_X1 port map( B1 => n192, B2 => A_ns(16), C1 => n174, C2 => 
                           A_s(16), A => n259, ZN => n152);
   U75 : INV_X1 port map( A => n153, ZN => n259);
   U76 : INV_X1 port map( A => n150, ZN => O_18_port);
   U77 : AOI221_X1 port map( B1 => n192, B2 => A_ns(17), C1 => n174, C2 => 
                           A_s(17), A => n257, ZN => n150);
   U78 : INV_X1 port map( A => n151, ZN => n257);
   U79 : INV_X1 port map( A => n148, ZN => O_19_port);
   U80 : AOI221_X1 port map( B1 => n192, B2 => A_ns(18), C1 => n174, C2 => 
                           A_s(18), A => n255, ZN => n148);
   U81 : INV_X1 port map( A => n149, ZN => n255);
   U82 : INV_X1 port map( A => n146, ZN => O_20_port);
   U83 : AOI221_X1 port map( B1 => n192, B2 => A_ns(19), C1 => n174, C2 => 
                           A_s(19), A => n253, ZN => n146);
   U84 : INV_X1 port map( A => n147, ZN => n253);
   U85 : INV_X1 port map( A => n144, ZN => O_21_port);
   U86 : AOI221_X1 port map( B1 => n192, B2 => A_ns(20), C1 => n174, C2 => 
                           A_s(20), A => n251, ZN => n144);
   U87 : INV_X1 port map( A => n145, ZN => n251);
   U88 : INV_X1 port map( A => n142, ZN => O_22_port);
   U89 : AOI221_X1 port map( B1 => n192, B2 => A_ns(21), C1 => n174, C2 => 
                           A_s(21), A => n249, ZN => n142);
   U90 : INV_X1 port map( A => n143, ZN => n249);
   U91 : INV_X1 port map( A => n140, ZN => O_23_port);
   U92 : AOI221_X1 port map( B1 => n192, B2 => A_ns(22), C1 => n174, C2 => 
                           A_s(22), A => n247, ZN => n140);
   U93 : INV_X1 port map( A => n141, ZN => n247);
   U94 : INV_X1 port map( A => n138, ZN => O_24_port);
   U95 : AOI221_X1 port map( B1 => n191, B2 => A_ns(23), C1 => n174, C2 => 
                           A_s(23), A => n245, ZN => n138);
   U96 : INV_X1 port map( A => n139, ZN => n245);
   U97 : INV_X1 port map( A => n136, ZN => O_25_port);
   U98 : AOI221_X1 port map( B1 => n191, B2 => A_ns(24), C1 => n174, C2 => 
                           A_s(24), A => n243, ZN => n136);
   U99 : INV_X1 port map( A => n137, ZN => n243);
   U100 : INV_X1 port map( A => n134, ZN => O_26_port);
   U101 : AOI221_X1 port map( B1 => n191, B2 => A_ns(25), C1 => n173, C2 => 
                           A_s(25), A => n241, ZN => n134);
   U102 : INV_X1 port map( A => n135, ZN => n241);
   U103 : INV_X1 port map( A => n132, ZN => O_27_port);
   U104 : AOI221_X1 port map( B1 => n191, B2 => A_ns(26), C1 => n173, C2 => 
                           A_s(26), A => n239, ZN => n132);
   U105 : INV_X1 port map( A => n133, ZN => n239);
   U106 : INV_X1 port map( A => n130, ZN => O_28_port);
   U107 : AOI221_X1 port map( B1 => n191, B2 => A_ns(27), C1 => n173, C2 => 
                           A_s(27), A => n237, ZN => n130);
   U108 : INV_X1 port map( A => n131, ZN => n237);
   U109 : INV_X1 port map( A => n128, ZN => O_29_port);
   U110 : AOI221_X1 port map( B1 => n191, B2 => A_ns(28), C1 => n173, C2 => 
                           A_s(28), A => n235, ZN => n128);
   U111 : INV_X1 port map( A => n129, ZN => n235);
   U112 : INV_X1 port map( A => n124, ZN => O_30_port);
   U113 : AOI221_X1 port map( B1 => n191, B2 => A_ns(29), C1 => n173, C2 => 
                           A_s(29), A => n233, ZN => n124);
   U114 : INV_X1 port map( A => n125, ZN => n233);
   U115 : INV_X1 port map( A => n122, ZN => O_31_port);
   U116 : AOI221_X1 port map( B1 => n191, B2 => A_ns(30), C1 => n173, C2 => 
                           A_s(30), A => n231, ZN => n122);
   U117 : INV_X1 port map( A => n123, ZN => n231);
   U118 : INV_X1 port map( A => n120, ZN => O_32_port);
   U119 : AOI221_X1 port map( B1 => n191, B2 => A_ns(31), C1 => n173, C2 => 
                           A_s(31), A => n229, ZN => n120);
   U120 : INV_X1 port map( A => n121, ZN => n229);
   U121 : INV_X1 port map( A => n114, ZN => O_35_port);
   U122 : AOI221_X1 port map( B1 => n190, B2 => A_ns(34), C1 => n173, C2 => 
                           A_s(34), A => n223, ZN => n114);
   U123 : INV_X1 port map( A => n115, ZN => n223);
   U124 : AOI221_X1 port map( B1 => n190, B2 => A_ns(9), C1 => n172, C2 => 
                           A_s(9), A => n272, ZN => n166);
   U125 : INV_X1 port map( A => n167, ZN => n272);
   U126 : INV_X1 port map( A => n94, ZN => O_9_port);
   U127 : INV_X1 port map( A => n95, ZN => n274);
   U128 : INV_X1 port map( A => n96, ZN => O_8_port);
   U129 : INV_X1 port map( A => n97, ZN => n208);
   U130 : AOI22_X1 port map( A1 => A_s(17), A2 => n186, B1 => A_ns(17), B2 => 
                           n180, ZN => n149);
   U131 : AOI22_X1 port map( A1 => A_s(18), A2 => n186, B1 => A_ns(18), B2 => 
                           n180, ZN => n147);
   U132 : AOI22_X1 port map( A1 => A_s(19), A2 => n186, B1 => A_ns(19), B2 => 
                           n180, ZN => n145);
   U133 : AOI22_X1 port map( A1 => A_s(20), A2 => n186, B1 => A_ns(20), B2 => 
                           n180, ZN => n143);
   U134 : AOI22_X1 port map( A1 => A_s(21), A2 => n186, B1 => A_ns(21), B2 => 
                           n180, ZN => n141);
   U135 : AOI22_X1 port map( A1 => A_s(13), A2 => n186, B1 => A_ns(13), B2 => 
                           n180, ZN => n157);
   U136 : AOI22_X1 port map( A1 => A_s(15), A2 => n186, B1 => A_ns(15), B2 => 
                           n180, ZN => n153);
   U137 : AOI22_X1 port map( A1 => A_s(16), A2 => n186, B1 => A_ns(16), B2 => 
                           n180, ZN => n151);
   U138 : AOI22_X1 port map( A1 => A_s(22), A2 => n186, B1 => A_ns(22), B2 => 
                           n180, ZN => n139);
   U139 : AOI22_X1 port map( A1 => A_s(23), A2 => n186, B1 => A_ns(23), B2 => 
                           n180, ZN => n137);
   U140 : AOI22_X1 port map( A1 => A_s(9), A2 => n187, B1 => A_ns(9), B2 => 
                           n181, ZN => n165);
   U141 : AOI22_X1 port map( A1 => A_s(10), A2 => n187, B1 => A_ns(10), B2 => 
                           n181, ZN => n163);
   U142 : AOI22_X1 port map( A1 => A_s(12), A2 => n186, B1 => A_ns(12), B2 => 
                           n180, ZN => n159);
   U143 : AOI22_X1 port map( A1 => A_s(14), A2 => n186, B1 => A_ns(14), B2 => 
                           n180, ZN => n155);
   U144 : AOI22_X1 port map( A1 => A_s(35), A2 => n184, B1 => A_ns(35), B2 => 
                           n178, ZN => n111);
   U145 : AOI22_X1 port map( A1 => A_s(36), A2 => n184, B1 => A_ns(36), B2 => 
                           n178, ZN => n109);
   U146 : AOI22_X1 port map( A1 => A_s(37), A2 => n184, B1 => A_ns(37), B2 => 
                           n178, ZN => n107);
   U147 : AOI22_X1 port map( A1 => A_s(38), A2 => n184, B1 => A_ns(38), B2 => 
                           n178, ZN => n105);
   U148 : AOI22_X1 port map( A1 => A_s(26), A2 => n185, B1 => A_ns(26), B2 => 
                           n179, ZN => n131);
   U149 : AOI22_X1 port map( A1 => A_s(24), A2 => n185, B1 => A_ns(24), B2 => 
                           n179, ZN => n135);
   U150 : AOI22_X1 port map( A1 => A_s(25), A2 => n185, B1 => A_ns(25), B2 => 
                           n179, ZN => n133);
   U151 : AOI22_X1 port map( A1 => A_s(27), A2 => n185, B1 => A_ns(27), B2 => 
                           n179, ZN => n129);
   U152 : AOI22_X1 port map( A1 => A_s(28), A2 => n185, B1 => A_ns(28), B2 => 
                           n179, ZN => n125);
   U153 : AOI22_X1 port map( A1 => A_s(29), A2 => n185, B1 => A_ns(29), B2 => 
                           n179, ZN => n123);
   U154 : AOI22_X1 port map( A1 => A_s(30), A2 => n185, B1 => A_ns(30), B2 => 
                           n179, ZN => n121);
   U155 : AOI22_X1 port map( A1 => A_s(31), A2 => n185, B1 => A_ns(31), B2 => 
                           n179, ZN => n119);
   U156 : AOI22_X1 port map( A1 => A_s(32), A2 => n185, B1 => A_ns(32), B2 => 
                           n179, ZN => n117);
   U157 : AOI22_X1 port map( A1 => A_s(33), A2 => n185, B1 => A_ns(33), B2 => 
                           n179, ZN => n115);
   U158 : AOI22_X1 port map( A1 => A_s(11), A2 => n187, B1 => A_ns(11), B2 => 
                           n181, ZN => n161);
   U159 : AOI22_X1 port map( A1 => A_s(34), A2 => n184, B1 => A_ns(34), B2 => 
                           n178, ZN => n113);
   U160 : NOR3_X1 port map( A1 => B(7), A2 => B(8), A3 => n276, ZN => n88);
   U161 : INV_X1 port map( A => B(9), ZN => n276);
   U162 : AND3_X1 port map( A1 => B(7), A2 => n276, A3 => B(8), ZN => n87);
   U163 : INV_X1 port map( A => n93, ZN => O_1_port);
   U164 : AOI22_X1 port map( A1 => n172, A2 => A_s(0), B1 => n193, B2 => 
                           A_ns(0), ZN => n93);
   U165 : INV_X1 port map( A => n126, ZN => O_2_port);
   U166 : AOI221_X1 port map( B1 => n191, B2 => A_ns(1), C1 => n173, C2 => 
                           A_s(1), A => n195, ZN => n126);
   U167 : INV_X1 port map( A => n127, ZN => n195);
   U168 : INV_X1 port map( A => n91, ZN => O_3_port);
   U169 : AOI221_X1 port map( B1 => n190, B2 => A_ns(2), C1 => n172, C2 => 
                           A_s(2), A => n198, ZN => n91);
   U171 : INV_X1 port map( A => n92, ZN => n198);
   U172 : INV_X1 port map( A => n100, ZN => O_4_port);
   U173 : AOI221_X1 port map( B1 => n190, B2 => A_ns(3), C1 => n172, C2 => 
                           A_s(3), A => n200, ZN => n100);
   U174 : INV_X1 port map( A => n101, ZN => n200);
   U175 : INV_X1 port map( A => n89, ZN => O_5_port);
   U176 : AOI221_X1 port map( B1 => n190, B2 => A_ns(4), C1 => n172, C2 => 
                           A_s(4), A => n202, ZN => n89);
   U177 : INV_X1 port map( A => n90, ZN => n202);
   U178 : INV_X1 port map( A => n98, ZN => O_6_port);
   U179 : AOI221_X1 port map( B1 => A_ns(5), B2 => n193, C1 => A_s(5), C2 => 
                           n172, A => n204, ZN => n98);
   U180 : INV_X1 port map( A => n99, ZN => n204);
   U181 : INV_X1 port map( A => n84, ZN => O_7_port);
   U182 : AOI221_X1 port map( B1 => n191, B2 => A_ns(6), C1 => n173, C2 => 
                           A_s(6), A => n206, ZN => n84);
   U183 : INV_X1 port map( A => n86, ZN => n206);
   U184 : AOI22_X1 port map( A1 => A_s(0), A2 => n185, B1 => A_ns(0), B2 => 
                           n179, ZN => n127);
   U185 : AOI22_X1 port map( A1 => A_s(1), A2 => n184, B1 => A_ns(1), B2 => 
                           n178, ZN => n92);
   U186 : AOI22_X1 port map( A1 => A_s(2), A2 => n184, B1 => A_ns(2), B2 => 
                           n178, ZN => n101);
   U187 : AOI22_X1 port map( A1 => A_s(3), A2 => n184, B1 => A_ns(3), B2 => 
                           n178, ZN => n90);
   U188 : AOI22_X1 port map( A1 => A_s(4), A2 => n184, B1 => A_ns(4), B2 => 
                           n178, ZN => n99);
   U189 : AOI22_X1 port map( A1 => A_s(5), A2 => n185, B1 => A_ns(5), B2 => 
                           n179, ZN => n86);
   U190 : AOI22_X1 port map( A1 => A_s(6), A2 => n184, B1 => A_ns(6), B2 => 
                           n178, ZN => n97);
   U191 : AOI221_X1 port map( B1 => n190, B2 => A_ns(8), C1 => n172, C2 => 
                           A_s(8), A => n274, ZN => n94);
   U192 : AOI22_X1 port map( A1 => A_s(8), A2 => n184, B1 => A_ns(8), B2 => 
                           n178, ZN => n167);
   U193 : AOI221_X1 port map( B1 => n190, B2 => A_ns(7), C1 => n172, C2 => 
                           A_s(7), A => n208, ZN => n96);
   U194 : AOI22_X1 port map( A1 => A_s(7), A2 => n184, B1 => A_ns(7), B2 => 
                           n178, ZN => n95);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT40_i6 is

   port( A_s, A_ns, B : in std_logic_vector (39 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (39 downto 0));

end BOOTHENC_NBIT40_i6;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT40_i6 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
      n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104
      , n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
      n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, 
      n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, 
      n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, 
      n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, 
      n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, 
      n177, n178, n179, A_nso_39_port, O_2_port, n182, O_1_port, O_3_port, n185
      , O_4_port, n187, O_5_port, n189, O_6_port, n191, O_37_port, O_38_port, 
      n194, O_39_port, n196, O_36_port, n198, O_35_port, n200, O_34_port, n202,
      O_33_port, n204, O_32_port, n206, O_31_port, n208, O_30_port, n210, 
      O_29_port, n212, O_28_port, n214, O_27_port, n216, O_26_port, n218, 
      O_25_port, n220, O_24_port, n222, O_23_port, n224, O_22_port, n226, 
      O_21_port, n228, O_20_port, n230, O_19_port, n232, O_18_port, n234, 
      O_17_port, n236, O_16_port, n238, O_15_port, n240, O_14_port, n242, 
      O_13_port, n244, O_12_port, n246, O_11_port, n248, O_10_port, n250, n251,
      O_9_port, O_8_port, n254, O_7_port, n256, n257, n258, n259 : std_logic;

begin
   O <= ( O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, 
      O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, 
      O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, 
      O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, O_16_port, 
      O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, O_10_port, 
      O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, O_3_port, 
      O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   A_nso <= ( A_nso_39_port, A_ns(36), A_ns(35), A_ns(34), A_ns(33), A_ns(32), 
      A_ns(31), A_ns(30), A_ns(29), A_ns(28), A_ns(27), A_ns(26), A_ns(25), 
      A_ns(24), A_ns(23), A_ns(22), A_ns(21), A_ns(20), A_ns(19), A_ns(18), 
      A_ns(17), A_ns(16), A_ns(15), A_ns(14), A_ns(13), A_ns(12), A_ns(11), 
      A_ns(10), A_ns(9), A_ns(8), A_ns(7), A_ns(6), A_ns(5), A_ns(4), A_ns(3), 
      A_ns(2), A_ns(1), A_ns(0), X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U162 : XOR2_X1 port map( A => B(5), B => B(6), Z => n161);
   U2 : AND2_X1 port map( A1 => n161, A2 => n160, ZN => n81);
   U3 : BUF_X1 port map( A => n258, Z => n162);
   U4 : CLKBUF_X1 port map( A => n258, Z => n164);
   U5 : CLKBUF_X1 port map( A => n258, Z => n163);
   U6 : CLKBUF_X1 port map( A => n81, Z => n179);
   U7 : CLKBUF_X1 port map( A => n81, Z => n178);
   U8 : CLKBUF_X1 port map( A => n171, Z => n174);
   U9 : CLKBUF_X1 port map( A => n165, Z => n168);
   U10 : CLKBUF_X1 port map( A => n84, Z => n166);
   U11 : CLKBUF_X1 port map( A => n83, Z => n172);
   U12 : BUF_X1 port map( A => A_ns(37), Z => A_nso_39_port);
   U13 : BUF_X1 port map( A => n172, Z => n175);
   U14 : BUF_X1 port map( A => n166, Z => n169);
   U15 : BUF_X2 port map( A => n81, Z => n177);
   U16 : BUF_X1 port map( A => n171, Z => n173);
   U17 : BUF_X1 port map( A => n165, Z => n167);
   U18 : INV_X1 port map( A => n160, ZN => n258);
   U19 : BUF_X1 port map( A => n172, Z => n176);
   U20 : BUF_X1 port map( A => n166, Z => n170);
   U21 : INV_X1 port map( A => n98, ZN => O_39_port);
   U22 : AOI221_X1 port map( B1 => n176, B2 => A_s(37), C1 => n170, C2 => 
                           A_nso_39_port, A => n196, ZN => n98);
   U23 : INV_X1 port map( A => n99, ZN => n196);
   U24 : INV_X1 port map( A => n100, ZN => O_38_port);
   U25 : AOI221_X1 port map( B1 => n177, B2 => A_nso_39_port, C1 => n162, C2 =>
                           A_s(37), A => n194, ZN => n100);
   U26 : INV_X1 port map( A => n101, ZN => n194);
   U27 : AOI22_X1 port map( A1 => A_ns(38), A2 => n177, B1 => A_s(38), B2 => 
                           n162, ZN => n99);
   U28 : NAND2_X1 port map( A1 => n161, A2 => n259, ZN => n160);
   U29 : BUF_X1 port map( A => n84, Z => n165);
   U30 : BUF_X1 port map( A => n83, Z => n171);
   U31 : INV_X1 port map( A => n102, ZN => O_37_port);
   U32 : AOI221_X1 port map( B1 => n177, B2 => A_ns(36), C1 => n162, C2 => 
                           A_s(36), A => n198, ZN => n102);
   U33 : INV_X1 port map( A => n103, ZN => n198);
   U34 : INV_X1 port map( A => n104, ZN => O_36_port);
   U35 : AOI221_X1 port map( B1 => n177, B2 => A_ns(35), C1 => n162, C2 => 
                           A_s(35), A => n200, ZN => n104);
   U36 : INV_X1 port map( A => n105, ZN => n200);
   U37 : INV_X1 port map( A => n106, ZN => O_35_port);
   U38 : AOI221_X1 port map( B1 => n177, B2 => A_ns(34), C1 => n162, C2 => 
                           A_s(34), A => n202, ZN => n106);
   U39 : INV_X1 port map( A => n107, ZN => n202);
   U40 : INV_X1 port map( A => n108, ZN => O_34_port);
   U41 : AOI221_X1 port map( B1 => n177, B2 => A_ns(33), C1 => n163, C2 => 
                           A_s(33), A => n204, ZN => n108);
   U42 : INV_X1 port map( A => n109, ZN => n204);
   U43 : INV_X1 port map( A => n110, ZN => O_33_port);
   U44 : AOI221_X1 port map( B1 => n177, B2 => A_ns(32), C1 => n163, C2 => 
                           A_s(32), A => n206, ZN => n110);
   U45 : INV_X1 port map( A => n111, ZN => n206);
   U46 : INV_X1 port map( A => n112, ZN => O_32_port);
   U47 : AOI221_X1 port map( B1 => n178, B2 => A_ns(31), C1 => n163, C2 => 
                           A_s(31), A => n208, ZN => n112);
   U48 : INV_X1 port map( A => n113, ZN => n208);
   U49 : INV_X1 port map( A => n156, ZN => O_11_port);
   U50 : AOI221_X1 port map( B1 => n179, B2 => A_ns(10), C1 => n164, C2 => 
                           A_s(10), A => n250, ZN => n156);
   U51 : INV_X1 port map( A => n157, ZN => n250);
   U52 : INV_X1 port map( A => n154, ZN => O_12_port);
   U53 : AOI221_X1 port map( B1 => n179, B2 => A_ns(11), C1 => n164, C2 => 
                           A_s(11), A => n248, ZN => n154);
   U54 : INV_X1 port map( A => n155, ZN => n248);
   U55 : INV_X1 port map( A => n152, ZN => O_13_port);
   U56 : AOI221_X1 port map( B1 => n179, B2 => A_ns(12), C1 => n164, C2 => 
                           A_s(12), A => n246, ZN => n152);
   U57 : INV_X1 port map( A => n153, ZN => n246);
   U58 : INV_X1 port map( A => n150, ZN => O_14_port);
   U59 : AOI221_X1 port map( B1 => n179, B2 => A_ns(13), C1 => n164, C2 => 
                           A_s(13), A => n244, ZN => n150);
   U60 : INV_X1 port map( A => n151, ZN => n244);
   U61 : INV_X1 port map( A => n148, ZN => O_15_port);
   U62 : AOI221_X1 port map( B1 => n179, B2 => A_ns(14), C1 => n164, C2 => 
                           A_s(14), A => n242, ZN => n148);
   U63 : INV_X1 port map( A => n149, ZN => n242);
   U64 : INV_X1 port map( A => n146, ZN => O_16_port);
   U65 : AOI221_X1 port map( B1 => n179, B2 => A_ns(15), C1 => n164, C2 => 
                           A_s(15), A => n240, ZN => n146);
   U66 : INV_X1 port map( A => n147, ZN => n240);
   U67 : INV_X1 port map( A => n144, ZN => O_17_port);
   U68 : AOI221_X1 port map( B1 => n179, B2 => A_ns(16), C1 => n164, C2 => 
                           A_s(16), A => n238, ZN => n144);
   U69 : INV_X1 port map( A => n145, ZN => n238);
   U70 : INV_X1 port map( A => n142, ZN => O_18_port);
   U71 : AOI221_X1 port map( B1 => n179, B2 => A_ns(17), C1 => n164, C2 => 
                           A_s(17), A => n236, ZN => n142);
   U72 : INV_X1 port map( A => n143, ZN => n236);
   U73 : INV_X1 port map( A => n140, ZN => O_19_port);
   U74 : AOI221_X1 port map( B1 => n179, B2 => A_ns(18), C1 => n164, C2 => 
                           A_s(18), A => n234, ZN => n140);
   U75 : INV_X1 port map( A => n141, ZN => n234);
   U76 : INV_X1 port map( A => n138, ZN => O_20_port);
   U77 : AOI221_X1 port map( B1 => n179, B2 => A_ns(19), C1 => n164, C2 => 
                           A_s(19), A => n232, ZN => n138);
   U78 : INV_X1 port map( A => n139, ZN => n232);
   U79 : INV_X1 port map( A => n136, ZN => O_21_port);
   U80 : AOI221_X1 port map( B1 => n179, B2 => A_ns(20), C1 => n164, C2 => 
                           A_s(20), A => n230, ZN => n136);
   U81 : INV_X1 port map( A => n137, ZN => n230);
   U82 : INV_X1 port map( A => n134, ZN => O_22_port);
   U83 : AOI221_X1 port map( B1 => n178, B2 => A_ns(21), C1 => n164, C2 => 
                           A_s(21), A => n228, ZN => n134);
   U84 : INV_X1 port map( A => n135, ZN => n228);
   U85 : INV_X1 port map( A => n132, ZN => O_23_port);
   U86 : AOI221_X1 port map( B1 => n178, B2 => A_ns(22), C1 => n164, C2 => 
                           A_s(22), A => n226, ZN => n132);
   U87 : INV_X1 port map( A => n133, ZN => n226);
   U88 : INV_X1 port map( A => n130, ZN => O_24_port);
   U89 : AOI221_X1 port map( B1 => n178, B2 => A_ns(23), C1 => n163, C2 => 
                           A_s(23), A => n224, ZN => n130);
   U90 : INV_X1 port map( A => n131, ZN => n224);
   U91 : INV_X1 port map( A => n128, ZN => O_25_port);
   U92 : AOI221_X1 port map( B1 => n178, B2 => A_ns(24), C1 => n163, C2 => 
                           A_s(24), A => n222, ZN => n128);
   U93 : INV_X1 port map( A => n129, ZN => n222);
   U94 : INV_X1 port map( A => n126, ZN => O_26_port);
   U95 : AOI221_X1 port map( B1 => n178, B2 => A_ns(25), C1 => n163, C2 => 
                           A_s(25), A => n220, ZN => n126);
   U96 : INV_X1 port map( A => n127, ZN => n220);
   U97 : INV_X1 port map( A => n124, ZN => O_27_port);
   U98 : AOI221_X1 port map( B1 => n178, B2 => A_ns(26), C1 => n163, C2 => 
                           A_s(26), A => n218, ZN => n124);
   U99 : INV_X1 port map( A => n125, ZN => n218);
   U100 : INV_X1 port map( A => n122, ZN => O_28_port);
   U101 : AOI221_X1 port map( B1 => n178, B2 => A_ns(27), C1 => n163, C2 => 
                           A_s(27), A => n216, ZN => n122);
   U102 : INV_X1 port map( A => n123, ZN => n216);
   U103 : INV_X1 port map( A => n120, ZN => O_29_port);
   U104 : AOI221_X1 port map( B1 => n178, B2 => A_ns(28), C1 => n163, C2 => 
                           A_s(28), A => n214, ZN => n120);
   U105 : INV_X1 port map( A => n121, ZN => n214);
   U106 : INV_X1 port map( A => n116, ZN => O_30_port);
   U107 : AOI221_X1 port map( B1 => n178, B2 => A_ns(29), C1 => n163, C2 => 
                           A_s(29), A => n212, ZN => n116);
   U108 : INV_X1 port map( A => n117, ZN => n212);
   U109 : INV_X1 port map( A => n114, ZN => O_31_port);
   U110 : AOI221_X1 port map( B1 => n178, B2 => A_ns(30), C1 => n163, C2 => 
                           A_s(30), A => n210, ZN => n114);
   U111 : INV_X1 port map( A => n115, ZN => n210);
   U112 : INV_X1 port map( A => n88, ZN => O_9_port);
   U113 : AOI221_X1 port map( B1 => n177, B2 => A_ns(8), C1 => n162, C2 => 
                           A_s(8), A => n254, ZN => n88);
   U114 : INV_X1 port map( A => n89, ZN => n254);
   U115 : INV_X1 port map( A => n158, ZN => O_10_port);
   U116 : AOI221_X1 port map( B1 => n177, B2 => A_ns(9), C1 => n162, C2 => 
                           A_s(9), A => n251, ZN => n158);
   U117 : INV_X1 port map( A => n159, ZN => n251);
   U118 : INV_X1 port map( A => n90, ZN => O_8_port);
   U119 : AOI221_X1 port map( B1 => n177, B2 => A_ns(7), C1 => n162, C2 => 
                           A_s(7), A => n256, ZN => n90);
   U120 : INV_X1 port map( A => n91, ZN => n256);
   U121 : INV_X1 port map( A => n92, ZN => O_7_port);
   U122 : INV_X1 port map( A => n93, ZN => n257);
   U123 : INV_X1 port map( A => n94, ZN => O_6_port);
   U124 : INV_X1 port map( A => n95, ZN => n191);
   U125 : AOI22_X1 port map( A1 => A_s(11), A2 => n175, B1 => A_ns(11), B2 => 
                           n169, ZN => n153);
   U126 : AOI22_X1 port map( A1 => A_s(13), A2 => n175, B1 => A_ns(13), B2 => 
                           n169, ZN => n149);
   U127 : AOI22_X1 port map( A1 => A_s(14), A2 => n175, B1 => A_ns(14), B2 => 
                           n169, ZN => n147);
   U128 : AOI22_X1 port map( A1 => A_s(15), A2 => n175, B1 => A_ns(15), B2 => 
                           n169, ZN => n145);
   U129 : AOI22_X1 port map( A1 => A_s(16), A2 => n175, B1 => A_ns(16), B2 => 
                           n169, ZN => n143);
   U130 : AOI22_X1 port map( A1 => A_s(17), A2 => n175, B1 => A_ns(17), B2 => 
                           n169, ZN => n141);
   U131 : AOI22_X1 port map( A1 => A_s(18), A2 => n175, B1 => A_ns(18), B2 => 
                           n169, ZN => n139);
   U132 : AOI22_X1 port map( A1 => A_s(19), A2 => n175, B1 => A_ns(19), B2 => 
                           n169, ZN => n137);
   U133 : AOI22_X1 port map( A1 => A_s(20), A2 => n175, B1 => A_ns(20), B2 => 
                           n169, ZN => n135);
   U134 : AOI22_X1 port map( A1 => A_s(21), A2 => n175, B1 => A_ns(21), B2 => 
                           n169, ZN => n133);
   U135 : AOI22_X1 port map( A1 => A_s(7), A2 => n173, B1 => A_ns(7), B2 => 
                           n167, ZN => n89);
   U136 : AOI22_X1 port map( A1 => A_s(8), A2 => n173, B1 => A_ns(8), B2 => 
                           n167, ZN => n159);
   U137 : AOI22_X1 port map( A1 => A_s(10), A2 => n175, B1 => A_ns(10), B2 => 
                           n169, ZN => n155);
   U138 : AOI22_X1 port map( A1 => A_s(12), A2 => n175, B1 => A_ns(12), B2 => 
                           n169, ZN => n151);
   U139 : AOI22_X1 port map( A1 => A_s(33), A2 => n173, B1 => A_ns(33), B2 => 
                           n167, ZN => n107);
   U140 : AOI22_X1 port map( A1 => A_s(34), A2 => n173, B1 => A_ns(34), B2 => 
                           n167, ZN => n105);
   U141 : AOI22_X1 port map( A1 => A_s(35), A2 => n173, B1 => A_ns(35), B2 => 
                           n167, ZN => n103);
   U142 : AOI22_X1 port map( A1 => A_s(36), A2 => n173, B1 => A_ns(36), B2 => 
                           n167, ZN => n101);
   U143 : AOI22_X1 port map( A1 => A_s(24), A2 => n174, B1 => A_ns(24), B2 => 
                           n168, ZN => n127);
   U144 : AOI22_X1 port map( A1 => A_s(23), A2 => n174, B1 => A_ns(23), B2 => 
                           n168, ZN => n129);
   U145 : AOI22_X1 port map( A1 => A_s(25), A2 => n174, B1 => A_ns(25), B2 => 
                           n168, ZN => n125);
   U146 : AOI22_X1 port map( A1 => A_s(26), A2 => n174, B1 => A_ns(26), B2 => 
                           n168, ZN => n123);
   U147 : AOI22_X1 port map( A1 => A_s(27), A2 => n174, B1 => A_ns(27), B2 => 
                           n168, ZN => n121);
   U148 : AOI22_X1 port map( A1 => A_s(28), A2 => n174, B1 => A_ns(28), B2 => 
                           n168, ZN => n117);
   U149 : AOI22_X1 port map( A1 => A_s(22), A2 => n174, B1 => A_ns(22), B2 => 
                           n168, ZN => n131);
   U150 : AOI22_X1 port map( A1 => A_s(29), A2 => n174, B1 => A_ns(29), B2 => 
                           n168, ZN => n115);
   U151 : AOI22_X1 port map( A1 => A_s(30), A2 => n174, B1 => A_ns(30), B2 => 
                           n168, ZN => n113);
   U152 : AOI22_X1 port map( A1 => A_s(31), A2 => n174, B1 => A_ns(31), B2 => 
                           n168, ZN => n111);
   U153 : AOI22_X1 port map( A1 => A_s(9), A2 => n176, B1 => A_ns(9), B2 => 
                           n170, ZN => n157);
   U154 : AOI22_X1 port map( A1 => A_s(32), A2 => n173, B1 => A_ns(32), B2 => 
                           n167, ZN => n109);
   U155 : NOR3_X1 port map( A1 => B(5), A2 => B(6), A3 => n259, ZN => n84);
   U156 : INV_X1 port map( A => B(7), ZN => n259);
   U157 : AND3_X1 port map( A1 => B(5), A2 => n259, A3 => B(6), ZN => n83);
   U158 : INV_X1 port map( A => n87, ZN => O_1_port);
   U159 : AOI22_X1 port map( A1 => n162, A2 => A_s(0), B1 => n179, B2 => 
                           A_ns(0), ZN => n87);
   U160 : INV_X1 port map( A => n118, ZN => O_2_port);
   U161 : AOI221_X1 port map( B1 => n178, B2 => A_ns(1), C1 => n163, C2 => 
                           A_s(1), A => n182, ZN => n118);
   U163 : INV_X1 port map( A => n119, ZN => n182);
   U164 : INV_X1 port map( A => n85, ZN => O_3_port);
   U165 : AOI221_X1 port map( B1 => n177, B2 => A_ns(2), C1 => n162, C2 => 
                           A_s(2), A => n185, ZN => n85);
   U166 : INV_X1 port map( A => n86, ZN => n185);
   U167 : INV_X1 port map( A => n96, ZN => O_4_port);
   U168 : AOI221_X1 port map( B1 => A_ns(3), B2 => n179, C1 => A_s(3), C2 => 
                           n162, A => n187, ZN => n96);
   U169 : INV_X1 port map( A => n97, ZN => n187);
   U170 : INV_X1 port map( A => n80, ZN => O_5_port);
   U171 : AOI221_X1 port map( B1 => n178, B2 => A_ns(4), C1 => n163, C2 => 
                           A_s(4), A => n189, ZN => n80);
   U172 : INV_X1 port map( A => n82, ZN => n189);
   U173 : AOI22_X1 port map( A1 => A_s(0), A2 => n174, B1 => A_ns(0), B2 => 
                           n168, ZN => n119);
   U174 : AOI22_X1 port map( A1 => A_s(1), A2 => n173, B1 => A_ns(1), B2 => 
                           n167, ZN => n86);
   U175 : AOI22_X1 port map( A1 => A_s(2), A2 => n173, B1 => A_ns(2), B2 => 
                           n167, ZN => n97);
   U176 : AOI22_X1 port map( A1 => A_s(3), A2 => n174, B1 => A_ns(3), B2 => 
                           n168, ZN => n82);
   U177 : AOI22_X1 port map( A1 => A_s(4), A2 => n173, B1 => A_ns(4), B2 => 
                           n167, ZN => n95);
   U178 : AOI221_X1 port map( B1 => n177, B2 => A_ns(6), C1 => n162, C2 => 
                           A_s(6), A => n257, ZN => n92);
   U179 : AOI22_X1 port map( A1 => A_s(6), A2 => n173, B1 => A_ns(6), B2 => 
                           n167, ZN => n91);
   U180 : AOI221_X1 port map( B1 => n177, B2 => A_ns(5), C1 => n162, C2 => 
                           A_s(5), A => n191, ZN => n94);
   U181 : AOI22_X1 port map( A1 => A_s(5), A2 => n173, B1 => A_ns(5), B2 => 
                           n167, ZN => n93);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT38_i4 is

   port( A_s, A_ns, B : in std_logic_vector (37 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (37 downto 0));

end BOOTHENC_NBIT38_i4;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT38_i4 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic0_port, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
      n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, 
      n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, 
      n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, 
      n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, 
      n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, 
      n149, n150, n151, n152, n153, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, O_2_port, n168, O_1_port, O_3_port, n171, 
      O_4_port, n173, O_35_port, O_36_port, n176, O_37_port, n178, O_34_port, 
      n180, O_33_port, n182, O_32_port, n184, O_31_port, n186, O_30_port, n188,
      O_29_port, n190, O_28_port, n192, O_27_port, n194, O_26_port, n196, 
      O_25_port, n198, O_24_port, n200, O_23_port, n202, O_22_port, n204, 
      O_21_port, n206, O_20_port, n208, O_19_port, n210, O_18_port, n212, 
      O_17_port, n214, O_16_port, n216, O_15_port, n218, O_14_port, n220, 
      O_13_port, n222, O_12_port, n224, O_11_port, n226, O_10_port, n228, n229,
      O_9_port, O_8_port, n232, O_7_port, n234, O_6_port, n236, O_5_port, n238,
      n239, n240, n241 : std_logic;

begin
   O <= ( O_37_port, O_36_port, O_35_port, O_34_port, O_33_port, O_32_port, 
      O_31_port, O_30_port, O_29_port, O_28_port, O_27_port, O_26_port, 
      O_25_port, O_24_port, O_23_port, O_22_port, O_21_port, O_20_port, 
      O_19_port, O_18_port, O_17_port, O_16_port, O_15_port, O_14_port, 
      O_13_port, O_12_port, O_11_port, O_10_port, O_9_port, O_8_port, O_7_port,
      O_6_port, O_5_port, O_4_port, O_3_port, O_2_port, O_1_port, X_Logic0_port
      );
   A_so <= ( A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), A_s(30), A_s(29), 
      A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), A_s(22), A_s(21), 
      A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), A_s(14), A_s(13), 
      A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), A_s(6), A_s(5), A_s(4)
      , A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, X_Logic0_port );
   A_nso <= ( A_ns(35), A_ns(34), A_ns(33), A_ns(32), A_ns(31), A_ns(30), 
      A_ns(29), A_ns(28), A_ns(27), A_ns(26), A_ns(25), A_ns(24), A_ns(23), 
      A_ns(22), A_ns(21), A_ns(20), A_ns(19), A_ns(18), A_ns(17), A_ns(16), 
      A_ns(15), A_ns(14), A_ns(13), A_ns(12), A_ns(11), A_ns(10), A_ns(9), 
      A_ns(8), A_ns(7), A_ns(6), A_ns(5), A_ns(4), A_ns(3), A_ns(2), A_ns(1), 
      A_ns(0), X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U154 : XOR2_X1 port map( A => B(3), B => B(4), Z => n153);
   U2 : INV_X2 port map( A => n128, ZN => O_21_port);
   U3 : INV_X1 port map( A => n142, ZN => O_14_port);
   U4 : AND2_X1 port map( A1 => n153, A2 => n152, ZN => n77);
   U5 : CLKBUF_X1 port map( A => n80, Z => n160);
   U6 : BUF_X2 port map( A => n240, Z => n155);
   U7 : CLKBUF_X1 port map( A => n240, Z => n156);
   U8 : CLKBUF_X1 port map( A => n240, Z => n157);
   U9 : BUF_X2 port map( A => n79, Z => n161);
   U10 : CLKBUF_X1 port map( A => n79, Z => n162);
   U11 : CLKBUF_X1 port map( A => n79, Z => n163);
   U12 : BUF_X2 port map( A => n80, Z => n158);
   U13 : CLKBUF_X1 port map( A => n80, Z => n159);
   U14 : BUF_X2 port map( A => n77, Z => n164);
   U15 : INV_X1 port map( A => n152, ZN => n240);
   U16 : CLKBUF_X1 port map( A => n77, Z => n165);
   U17 : CLKBUF_X1 port map( A => n77, Z => n166);
   U18 : NAND2_X1 port map( A1 => n153, A2 => n241, ZN => n152);
   U19 : INV_X1 port map( A => n94, ZN => O_37_port);
   U20 : AOI221_X1 port map( B1 => n163, B2 => A_s(35), C1 => n160, C2 => 
                           A_ns(35), A => n178, ZN => n94);
   U21 : INV_X1 port map( A => n95, ZN => n178);
   U22 : INV_X1 port map( A => n98, ZN => O_35_port);
   U23 : AOI221_X1 port map( B1 => n164, B2 => A_ns(34), C1 => n155, C2 => 
                           A_s(34), A => n180, ZN => n98);
   U24 : INV_X1 port map( A => n99, ZN => n180);
   U25 : INV_X1 port map( A => n100, ZN => O_34_port);
   U26 : AOI221_X1 port map( B1 => n164, B2 => A_ns(33), C1 => n155, C2 => 
                           A_s(33), A => n182, ZN => n100);
   U27 : INV_X1 port map( A => n101, ZN => n182);
   U28 : INV_X1 port map( A => n102, ZN => O_33_port);
   U29 : AOI221_X1 port map( B1 => n164, B2 => A_ns(32), C1 => n156, C2 => 
                           A_s(32), A => n184, ZN => n102);
   U30 : INV_X1 port map( A => n103, ZN => n184);
   U31 : INV_X1 port map( A => n86, ZN => O_7_port);
   U32 : AOI221_X1 port map( B1 => n164, B2 => A_ns(6), C1 => n155, C2 => 
                           A_s(6), A => n236, ZN => n86);
   U33 : INV_X1 port map( A => n87, ZN => n236);
   U34 : INV_X1 port map( A => n84, ZN => O_8_port);
   U35 : AOI221_X1 port map( B1 => n164, B2 => A_ns(7), C1 => n155, C2 => 
                           A_s(7), A => n234, ZN => n84);
   U36 : INV_X1 port map( A => n85, ZN => n234);
   U37 : INV_X1 port map( A => n82, ZN => O_9_port);
   U38 : AOI221_X1 port map( B1 => n164, B2 => A_ns(8), C1 => n155, C2 => 
                           A_s(8), A => n232, ZN => n82);
   U39 : INV_X1 port map( A => n83, ZN => n232);
   U40 : INV_X1 port map( A => n150, ZN => O_10_port);
   U41 : AOI221_X1 port map( B1 => n164, B2 => A_ns(9), C1 => n155, C2 => 
                           A_s(9), A => n229, ZN => n150);
   U42 : INV_X1 port map( A => n151, ZN => n229);
   U43 : INV_X1 port map( A => n148, ZN => O_11_port);
   U44 : AOI221_X1 port map( B1 => n166, B2 => A_ns(10), C1 => n157, C2 => 
                           A_s(10), A => n228, ZN => n148);
   U45 : INV_X1 port map( A => n149, ZN => n228);
   U46 : INV_X1 port map( A => n146, ZN => O_12_port);
   U47 : AOI221_X1 port map( B1 => n166, B2 => A_ns(11), C1 => n157, C2 => 
                           A_s(11), A => n226, ZN => n146);
   U48 : INV_X1 port map( A => n147, ZN => n226);
   U49 : INV_X1 port map( A => n144, ZN => O_13_port);
   U50 : AOI221_X1 port map( B1 => n166, B2 => A_ns(12), C1 => n157, C2 => 
                           A_s(12), A => n224, ZN => n144);
   U51 : INV_X1 port map( A => n145, ZN => n224);
   U52 : AOI221_X1 port map( B1 => n166, B2 => A_ns(13), C1 => n157, C2 => 
                           A_s(13), A => n222, ZN => n142);
   U53 : INV_X1 port map( A => n143, ZN => n222);
   U54 : INV_X1 port map( A => n140, ZN => O_15_port);
   U55 : AOI221_X1 port map( B1 => n166, B2 => A_ns(14), C1 => n157, C2 => 
                           A_s(14), A => n220, ZN => n140);
   U56 : INV_X1 port map( A => n141, ZN => n220);
   U57 : INV_X1 port map( A => n138, ZN => O_16_port);
   U58 : AOI221_X1 port map( B1 => n166, B2 => A_ns(15), C1 => n157, C2 => 
                           A_s(15), A => n218, ZN => n138);
   U59 : INV_X1 port map( A => n139, ZN => n218);
   U60 : INV_X1 port map( A => n136, ZN => O_17_port);
   U61 : AOI221_X1 port map( B1 => n166, B2 => A_ns(16), C1 => n157, C2 => 
                           A_s(16), A => n216, ZN => n136);
   U62 : INV_X1 port map( A => n137, ZN => n216);
   U63 : INV_X1 port map( A => n134, ZN => O_18_port);
   U64 : AOI221_X1 port map( B1 => n165, B2 => A_ns(17), C1 => n157, C2 => 
                           A_s(17), A => n214, ZN => n134);
   U65 : INV_X1 port map( A => n135, ZN => n214);
   U66 : INV_X1 port map( A => n132, ZN => O_19_port);
   U67 : AOI221_X1 port map( B1 => n166, B2 => A_ns(18), C1 => n157, C2 => 
                           A_s(18), A => n212, ZN => n132);
   U68 : INV_X1 port map( A => n133, ZN => n212);
   U69 : INV_X1 port map( A => n130, ZN => O_20_port);
   U70 : AOI221_X1 port map( B1 => n166, B2 => A_ns(19), C1 => n157, C2 => 
                           A_s(19), A => n210, ZN => n130);
   U71 : INV_X1 port map( A => n131, ZN => n210);
   U72 : AOI221_X1 port map( B1 => n165, B2 => A_ns(20), C1 => n157, C2 => 
                           A_s(20), A => n208, ZN => n128);
   U73 : INV_X1 port map( A => n129, ZN => n208);
   U74 : INV_X1 port map( A => n126, ZN => O_22_port);
   U75 : AOI221_X1 port map( B1 => n165, B2 => A_ns(21), C1 => n156, C2 => 
                           A_s(21), A => n206, ZN => n126);
   U76 : INV_X1 port map( A => n127, ZN => n206);
   U77 : INV_X1 port map( A => n124, ZN => O_23_port);
   U78 : AOI221_X1 port map( B1 => n165, B2 => A_ns(22), C1 => n156, C2 => 
                           A_s(22), A => n204, ZN => n124);
   U79 : INV_X1 port map( A => n125, ZN => n204);
   U80 : INV_X1 port map( A => n122, ZN => O_24_port);
   U81 : AOI221_X1 port map( B1 => n165, B2 => A_ns(23), C1 => n156, C2 => 
                           A_s(23), A => n202, ZN => n122);
   U82 : INV_X1 port map( A => n123, ZN => n202);
   U83 : INV_X1 port map( A => n120, ZN => O_25_port);
   U84 : AOI221_X1 port map( B1 => n165, B2 => A_ns(24), C1 => n156, C2 => 
                           A_s(24), A => n200, ZN => n120);
   U85 : INV_X1 port map( A => n121, ZN => n200);
   U86 : INV_X1 port map( A => n118, ZN => O_26_port);
   U87 : AOI221_X1 port map( B1 => n165, B2 => A_ns(25), C1 => n156, C2 => 
                           A_s(25), A => n198, ZN => n118);
   U88 : INV_X1 port map( A => n119, ZN => n198);
   U89 : INV_X1 port map( A => n116, ZN => O_27_port);
   U90 : AOI221_X1 port map( B1 => n165, B2 => A_ns(26), C1 => n156, C2 => 
                           A_s(26), A => n196, ZN => n116);
   U91 : INV_X1 port map( A => n117, ZN => n196);
   U92 : INV_X1 port map( A => n114, ZN => O_28_port);
   U93 : AOI221_X1 port map( B1 => n165, B2 => A_ns(27), C1 => n156, C2 => 
                           A_s(27), A => n194, ZN => n114);
   U94 : INV_X1 port map( A => n115, ZN => n194);
   U95 : INV_X1 port map( A => n112, ZN => O_29_port);
   U96 : AOI221_X1 port map( B1 => n165, B2 => A_ns(28), C1 => n156, C2 => 
                           A_s(28), A => n192, ZN => n112);
   U97 : INV_X1 port map( A => n113, ZN => n192);
   U98 : INV_X1 port map( A => n108, ZN => O_30_port);
   U99 : AOI221_X1 port map( B1 => n165, B2 => A_ns(29), C1 => n156, C2 => 
                           A_s(29), A => n190, ZN => n108);
   U100 : INV_X1 port map( A => n109, ZN => n190);
   U101 : INV_X1 port map( A => n106, ZN => O_31_port);
   U102 : AOI221_X1 port map( B1 => n165, B2 => A_ns(30), C1 => n156, C2 => 
                           A_s(30), A => n188, ZN => n106);
   U103 : INV_X1 port map( A => n107, ZN => n188);
   U104 : INV_X1 port map( A => n104, ZN => O_32_port);
   U105 : AOI221_X1 port map( B1 => n164, B2 => A_ns(31), C1 => n156, C2 => 
                           A_s(31), A => n186, ZN => n104);
   U106 : INV_X1 port map( A => n105, ZN => n186);
   U107 : INV_X1 port map( A => n88, ZN => O_6_port);
   U108 : AOI221_X1 port map( B1 => n164, B2 => A_ns(5), C1 => n155, C2 => 
                           A_s(5), A => n238, ZN => n88);
   U109 : INV_X1 port map( A => n89, ZN => n238);
   U110 : INV_X1 port map( A => n96, ZN => O_36_port);
   U111 : AOI221_X1 port map( B1 => n164, B2 => A_ns(35), C1 => n155, C2 => 
                           A_s(35), A => n176, ZN => n96);
   U112 : INV_X1 port map( A => n97, ZN => n176);
   U113 : INV_X1 port map( A => n90, ZN => O_5_port);
   U114 : INV_X1 port map( A => n91, ZN => n239);
   U115 : INV_X1 port map( A => n92, ZN => O_4_port);
   U116 : INV_X1 port map( A => n93, ZN => n173);
   U117 : INV_X1 port map( A => B(5), ZN => n241);
   U118 : NOR3_X1 port map( A1 => B(3), A2 => B(4), A3 => n241, ZN => n80);
   U119 : AOI22_X1 port map( A1 => A_s(9), A2 => n163, B1 => A_ns(9), B2 => 
                           n160, ZN => n149);
   U120 : AOI22_X1 port map( A1 => A_s(11), A2 => n163, B1 => A_ns(11), B2 => 
                           n160, ZN => n145);
   U121 : AOI22_X1 port map( A1 => A_s(12), A2 => n163, B1 => A_ns(12), B2 => 
                           n160, ZN => n143);
   U122 : AOI22_X1 port map( A1 => A_s(13), A2 => n163, B1 => A_ns(13), B2 => 
                           n160, ZN => n141);
   U123 : AOI22_X1 port map( A1 => A_s(14), A2 => n163, B1 => A_ns(14), B2 => 
                           n160, ZN => n139);
   U124 : AOI22_X1 port map( A1 => A_s(15), A2 => n163, B1 => A_ns(15), B2 => 
                           n160, ZN => n137);
   U125 : AOI22_X1 port map( A1 => A_s(16), A2 => n163, B1 => A_ns(16), B2 => 
                           n160, ZN => n135);
   U126 : AOI22_X1 port map( A1 => A_s(17), A2 => n163, B1 => A_ns(17), B2 => 
                           n160, ZN => n133);
   U127 : AOI22_X1 port map( A1 => A_s(18), A2 => n163, B1 => A_ns(18), B2 => 
                           n160, ZN => n131);
   U128 : AOI22_X1 port map( A1 => A_s(19), A2 => n163, B1 => A_ns(19), B2 => 
                           n160, ZN => n129);
   U129 : AOI22_X1 port map( A1 => A_s(34), A2 => n161, B1 => A_ns(34), B2 => 
                           n158, ZN => n97);
   U130 : AOI22_X1 port map( A1 => A_s(5), A2 => n161, B1 => A_ns(5), B2 => 
                           n158, ZN => n87);
   U131 : AOI22_X1 port map( A1 => A_s(6), A2 => n161, B1 => A_ns(6), B2 => 
                           n158, ZN => n85);
   U132 : AOI22_X1 port map( A1 => A_s(8), A2 => n161, B1 => A_ns(8), B2 => 
                           n158, ZN => n151);
   U133 : AOI22_X1 port map( A1 => A_s(10), A2 => n163, B1 => A_ns(10), B2 => 
                           n160, ZN => n147);
   U134 : AOI22_X1 port map( A1 => A_s(31), A2 => n161, B1 => A_ns(31), B2 => 
                           n158, ZN => n103);
   U135 : AOI22_X1 port map( A1 => A_s(32), A2 => n161, B1 => A_ns(32), B2 => 
                           n158, ZN => n101);
   U136 : AOI22_X1 port map( A1 => A_s(33), A2 => n161, B1 => A_ns(33), B2 => 
                           n158, ZN => n99);
   U137 : AOI22_X1 port map( A1 => A_s(22), A2 => n162, B1 => A_ns(22), B2 => 
                           n159, ZN => n123);
   U138 : AOI22_X1 port map( A1 => A_s(20), A2 => n162, B1 => A_ns(20), B2 => 
                           n159, ZN => n127);
   U139 : AOI22_X1 port map( A1 => A_s(21), A2 => n162, B1 => A_ns(21), B2 => 
                           n159, ZN => n125);
   U140 : AOI22_X1 port map( A1 => A_s(23), A2 => n162, B1 => A_ns(23), B2 => 
                           n159, ZN => n121);
   U141 : AOI22_X1 port map( A1 => A_s(24), A2 => n162, B1 => A_ns(24), B2 => 
                           n159, ZN => n119);
   U142 : AOI22_X1 port map( A1 => A_s(25), A2 => n162, B1 => A_ns(25), B2 => 
                           n159, ZN => n117);
   U143 : AOI22_X1 port map( A1 => A_s(26), A2 => n162, B1 => A_ns(26), B2 => 
                           n159, ZN => n115);
   U144 : AOI22_X1 port map( A1 => A_s(27), A2 => n162, B1 => A_ns(27), B2 => 
                           n159, ZN => n113);
   U145 : AOI22_X1 port map( A1 => A_s(28), A2 => n162, B1 => A_ns(28), B2 => 
                           n159, ZN => n109);
   U146 : AOI22_X1 port map( A1 => A_s(29), A2 => n162, B1 => A_ns(29), B2 => 
                           n159, ZN => n107);
   U147 : AOI22_X1 port map( A1 => A_s(7), A2 => n161, B1 => A_ns(7), B2 => 
                           n158, ZN => n83);
   U148 : AOI22_X1 port map( A1 => A_s(30), A2 => n161, B1 => A_ns(30), B2 => 
                           n158, ZN => n105);
   U149 : AOI22_X1 port map( A1 => A_ns(36), A2 => n164, B1 => A_s(36), B2 => 
                           n155, ZN => n95);
   U150 : AND3_X1 port map( A1 => B(3), A2 => n241, A3 => B(4), ZN => n79);
   U151 : INV_X1 port map( A => n81, ZN => O_1_port);
   U152 : AOI22_X1 port map( A1 => n155, A2 => A_s(0), B1 => n166, B2 => 
                           A_ns(0), ZN => n81);
   U153 : INV_X1 port map( A => n110, ZN => O_2_port);
   U155 : AOI221_X1 port map( B1 => A_ns(1), B2 => n166, C1 => A_s(1), C2 => 
                           n155, A => n168, ZN => n110);
   U156 : INV_X1 port map( A => n111, ZN => n168);
   U157 : INV_X1 port map( A => n76, ZN => O_3_port);
   U158 : AOI221_X1 port map( B1 => n165, B2 => A_ns(2), C1 => n156, C2 => 
                           A_s(2), A => n171, ZN => n76);
   U159 : INV_X1 port map( A => n78, ZN => n171);
   U160 : AOI22_X1 port map( A1 => A_s(0), A2 => n162, B1 => A_ns(0), B2 => 
                           n159, ZN => n111);
   U161 : AOI22_X1 port map( A1 => A_s(1), A2 => n162, B1 => A_ns(1), B2 => 
                           n159, ZN => n78);
   U162 : AOI22_X1 port map( A1 => A_s(2), A2 => n161, B1 => A_ns(2), B2 => 
                           n158, ZN => n93);
   U163 : AOI221_X1 port map( B1 => n164, B2 => A_ns(4), C1 => n155, C2 => 
                           A_s(4), A => n239, ZN => n90);
   U164 : AOI22_X1 port map( A1 => A_s(4), A2 => n161, B1 => A_ns(4), B2 => 
                           n158, ZN => n89);
   U165 : AOI221_X1 port map( B1 => n164, B2 => A_ns(3), C1 => n155, C2 => 
                           A_s(3), A => n173, ZN => n92);
   U166 : AOI22_X1 port map( A1 => A_s(3), A2 => n161, B1 => A_ns(3), B2 => 
                           n158, ZN => n91);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT36_i2 is

   port( A_s, A_ns, B : in std_logic_vector (35 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (35 downto 0));

end BOOTHENC_NBIT36_i2;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT36_i2 is

   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, n72, n74, n75, n76, n77, n78, n79, n81, n83, n84, n85,
      n87, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, net35751, net39408, net40332, 
      net40345, net41959, net42029, net43199, net43203, net41985, O_7_port, 
      n149, n150, A_so_3_port, n152, n153, n154, A_nso_7_port, n156, n157, 
      A_nso_8_port, A_nso_5_port, n160, O_6_port, n162, n163, O_3_port, n165, 
      n166, n167, n168, n169, O_4_port, n171, n172, n173, n174, n175, n176, 
      n177, n178, n179, n180, O_2_port, O_1_port, O_33_port, O_34_port, n185, 
      O_35_port, n187, O_32_port, n189, O_31_port, n191, O_30_port, n193, 
      O_29_port, n195, O_28_port, n197, O_27_port, n199, O_26_port, n201, 
      O_25_port, n203, O_24_port, n205, O_23_port, n207, O_22_port, n209, 
      O_21_port, n211, O_20_port, n213, O_19_port, n215, O_18_port, n217, 
      O_17_port, n219, O_16_port, n221, O_15_port, n223, O_14_port, n225, 
      O_13_port, n227, O_12_port, n229, O_11_port, n231, O_10_port, n233, n234,
      O_9_port, O_8_port, n237, n238, n239, O_5_port, n241, n242 : std_logic;

begin
   O <= ( O_35_port, O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, 
      O_29_port, O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, 
      O_23_port, O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, 
      O_17_port, O_16_port, O_15_port, O_14_port, O_13_port, O_12_port, 
      O_11_port, O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, 
      O_4_port, O_3_port, O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(33), A_s(32), A_s(31), A_s(30), A_s(29), A_s(28), A_s(27), 
      A_s(26), A_s(25), A_s(24), A_s(23), A_s(22), A_s(21), A_s(20), A_s(19), 
      A_s(18), A_s(17), A_s(16), A_s(15), A_s(14), A_s(13), A_s(12), A_s(11), 
      A_s(10), A_s(9), A_s(8), A_s(7), A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), 
      A_so_3_port, A_s(0), X_Logic0_port, X_Logic0_port );
   A_nso <= ( A_ns(33), A_ns(32), A_ns(31), A_ns(30), A_ns(29), A_ns(28), 
      A_ns(27), A_ns(26), A_ns(25), A_ns(24), A_ns(23), A_ns(22), A_ns(21), 
      A_ns(20), A_ns(19), A_ns(18), A_ns(17), A_ns(16), A_ns(15), A_ns(14), 
      A_ns(13), A_ns(12), A_ns(11), A_ns(10), A_ns(9), A_ns(8), A_ns(7), 
      A_nso_8_port, A_nso_7_port, A_ns(4), A_nso_5_port, A_ns(2), A_ns(1), 
      A_ns(0), X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : OR3_X2 port map( A1 => n156, A2 => n157, A3 => n239, ZN => O_7_port);
   U3 : BUF_X1 port map( A => n76, Z => n178);
   U4 : BUF_X1 port map( A => A_s(1), Z => A_so_3_port);
   U5 : AND2_X1 port map( A1 => net43199, A2 => net35751, ZN => n149);
   U6 : AND2_X1 port map( A1 => net43199, A2 => net35751, ZN => n150);
   U7 : CLKBUF_X1 port map( A => n150, Z => n177);
   U8 : CLKBUF_X1 port map( A => A_ns(6), Z => n152);
   U9 : AOI22_X1 port map( A1 => A_s(1), A2 => n76, B1 => A_ns(1), B2 => n166, 
                           ZN => n89);
   U10 : OAI211_X1 port map( C1 => n153, C2 => n154, A => n165, B => n89, ZN =>
                           O_3_port);
   U11 : INV_X1 port map( A => A_ns(2), ZN => n153);
   U12 : INV_X1 port map( A => n160, ZN => n154);
   U13 : NAND3_X1 port map( A1 => net43199, A2 => n144, A3 => A_ns(1), ZN => 
                           n174);
   U14 : XOR2_X1 port map( A => B(2), B => B(1), Z => net41985);
   U15 : NAND2_X1 port map( A1 => net41985, A2 => net35751, ZN => n144);
   U16 : BUF_X1 port map( A => B(2), Z => net41959);
   U17 : XOR2_X1 port map( A => B(1), B => B(2), Z => net43199);
   U18 : XNOR2_X1 port map( A => B(1), B => B(2), ZN => net43203);
   U19 : BUF_X2 port map( A => B(1), Z => net40332);
   U20 : BUF_X2 port map( A => A_ns(5), Z => A_nso_7_port);
   U21 : AND2_X1 port map( A1 => net39408, A2 => n152, ZN => n156);
   U22 : AND2_X1 port map( A1 => n176, A2 => A_s(6), ZN => n157);
   U23 : BUF_X2 port map( A => n152, Z => A_nso_8_port);
   U24 : BUF_X2 port map( A => A_ns(3), Z => A_nso_5_port);
   U25 : AND3_X1 port map( A1 => net41959, A2 => net35751, A3 => net40332, ZN 
                           => n76);
   U26 : NOR2_X1 port map( A1 => net43203, A2 => B(3), ZN => net42029);
   U27 : AND2_X1 port map( A1 => n144, A2 => net43199, ZN => n160);
   U28 : BUF_X1 port map( A => n160, Z => net40345);
   U29 : INV_X2 port map( A => B(3), ZN => net35751);
   U30 : OR3_X2 port map( A1 => n162, A2 => n163, A3 => n241, ZN => O_6_port);
   U31 : AND2_X1 port map( A1 => net39408, A2 => A_ns(5), ZN => n162);
   U32 : AND2_X1 port map( A1 => n177, A2 => A_s(5), ZN => n163);
   U33 : BUF_X4 port map( A => n150, Z => n176);
   U34 : NAND2_X1 port map( A1 => n149, A2 => A_s(2), ZN => n165);
   U35 : NOR3_X1 port map( A1 => net40332, A2 => net41959, A3 => net35751, ZN 
                           => n166);
   U36 : BUF_X2 port map( A => n168, Z => n167);
   U37 : BUF_X2 port map( A => n166, Z => n168);
   U38 : BUF_X2 port map( A => n77, Z => n169);
   U39 : NAND3_X1 port map( A1 => n171, A2 => n172, A3 => n87, ZN => O_4_port);
   U40 : NAND2_X1 port map( A1 => n160, A2 => A_ns(3), ZN => n171);
   U41 : NAND2_X1 port map( A1 => n150, A2 => A_s(3), ZN => n172);
   U42 : BUF_X2 port map( A => n76, Z => n180);
   U43 : BUF_X2 port map( A => n160, Z => net39408);
   U44 : NAND2_X1 port map( A1 => n174, A2 => n173, ZN => O_2_port);
   U45 : AND2_X1 port map( A1 => n175, A2 => n103, ZN => n173);
   U46 : NAND2_X1 port map( A1 => net42029, A2 => A_s(1), ZN => n175);
   U47 : CLKBUF_X1 port map( A => n76, Z => n179);
   U48 : INV_X1 port map( A => n83, ZN => n241);
   U49 : AOI22_X1 port map( A1 => n179, A2 => A_s(0), B1 => n167, B2 => A_ns(0)
                           , ZN => n103);
   U50 : AOI221_X1 port map( B1 => net39408, B2 => A_ns(7), C1 => n176, C2 => 
                           A_s(7), A => n238, ZN => n78);
   U51 : INV_X1 port map( A => n79, ZN => n238);
   U52 : AOI221_X1 port map( B1 => net39408, B2 => A_ns(9), C1 => n176, C2 => 
                           A_s(9), A => n234, ZN => n142);
   U53 : INV_X1 port map( A => n143, ZN => n234);
   U54 : AOI221_X1 port map( B1 => net39408, B2 => A_ns(10), C1 => n176, C2 => 
                           A_s(10), A => n233, ZN => n140);
   U55 : INV_X1 port map( A => n141, ZN => n233);
   U56 : AOI22_X1 port map( A1 => A_s(9), A2 => n179, B1 => A_ns(9), B2 => n169
                           , ZN => n141);
   U57 : INV_X1 port map( A => n81, ZN => n239);
   U58 : AOI221_X1 port map( B1 => net39408, B2 => A_ns(8), C1 => n176, C2 => 
                           A_s(8), A => n237, ZN => n74);
   U59 : INV_X1 port map( A => n75, ZN => n237);
   U60 : AOI22_X1 port map( A1 => A_s(7), A2 => n179, B1 => A_ns(7), B2 => n167
                           , ZN => n75);
   U61 : AOI221_X1 port map( B1 => A_ns(4), B2 => net40345, C1 => n150, C2 => 
                           A_s(4), A => n242, ZN => n84);
   U62 : INV_X1 port map( A => n85, ZN => n242);
   U63 : INV_X1 port map( A => n90, ZN => O_35_port);
   U64 : AOI221_X1 port map( B1 => n180, B2 => A_s(33), C1 => n169, C2 => 
                           A_ns(33), A => n187, ZN => n90);
   U65 : INV_X1 port map( A => n91, ZN => n187);
   U66 : INV_X1 port map( A => n92, ZN => O_34_port);
   U67 : AOI221_X1 port map( B1 => net39408, B2 => A_ns(33), C1 => n177, C2 => 
                           A_s(33), A => n185, ZN => n92);
   U68 : INV_X1 port map( A => n93, ZN => n185);
   U69 : INV_X1 port map( A => n94, ZN => O_33_port);
   U70 : AOI221_X1 port map( B1 => net40345, B2 => A_ns(32), C1 => n176, C2 => 
                           A_s(32), A => n189, ZN => n94);
   U71 : INV_X1 port map( A => n95, ZN => n189);
   U72 : INV_X1 port map( A => n96, ZN => O_32_port);
   U73 : INV_X1 port map( A => n98, ZN => O_31_port);
   U74 : INV_X1 port map( A => n100, ZN => O_30_port);
   U75 : INV_X1 port map( A => n78, ZN => O_8_port);
   U76 : INV_X1 port map( A => n74, ZN => O_9_port);
   U77 : INV_X1 port map( A => n142, ZN => O_10_port);
   U78 : INV_X1 port map( A => n140, ZN => O_11_port);
   U79 : INV_X1 port map( A => n138, ZN => O_12_port);
   U80 : INV_X1 port map( A => n136, ZN => O_13_port);
   U81 : INV_X1 port map( A => n134, ZN => O_14_port);
   U82 : INV_X1 port map( A => n132, ZN => O_15_port);
   U83 : INV_X1 port map( A => n130, ZN => O_16_port);
   U84 : INV_X1 port map( A => n128, ZN => O_17_port);
   U85 : INV_X1 port map( A => n126, ZN => O_18_port);
   U86 : INV_X1 port map( A => n124, ZN => O_19_port);
   U87 : INV_X1 port map( A => n122, ZN => O_20_port);
   U88 : INV_X1 port map( A => n120, ZN => O_21_port);
   U89 : INV_X1 port map( A => n118, ZN => O_22_port);
   U90 : INV_X1 port map( A => n116, ZN => O_23_port);
   U91 : INV_X1 port map( A => n114, ZN => O_24_port);
   U92 : INV_X1 port map( A => n112, ZN => O_25_port);
   U93 : INV_X1 port map( A => n110, ZN => O_26_port);
   U94 : INV_X1 port map( A => n108, ZN => O_27_port);
   U95 : INV_X1 port map( A => n106, ZN => O_28_port);
   U96 : INV_X1 port map( A => n104, ZN => O_29_port);
   U97 : INV_X1 port map( A => n125, ZN => n217);
   U98 : AOI22_X1 port map( A1 => A_s(17), A2 => n179, B1 => A_ns(17), B2 => 
                           n168, ZN => n125);
   U99 : INV_X1 port map( A => n111, ZN => n203);
   U100 : AOI22_X1 port map( A1 => A_s(24), A2 => n180, B1 => A_ns(24), B2 => 
                           n169, ZN => n111);
   U101 : INV_X1 port map( A => n109, ZN => n201);
   U102 : AOI22_X1 port map( A1 => A_s(25), A2 => n179, B1 => A_ns(25), B2 => 
                           n167, ZN => n109);
   U103 : INV_X1 port map( A => n107, ZN => n199);
   U104 : AOI22_X1 port map( A1 => A_s(26), A2 => n180, B1 => A_ns(26), B2 => 
                           n168, ZN => n107);
   U105 : INV_X1 port map( A => n105, ZN => n197);
   U106 : AOI22_X1 port map( A1 => A_s(27), A2 => n179, B1 => A_ns(27), B2 => 
                           n169, ZN => n105);
   U107 : AOI221_X1 port map( B1 => net39408, B2 => A_ns(11), C1 => n176, C2 =>
                           A_s(11), A => n231, ZN => n138);
   U108 : INV_X1 port map( A => n139, ZN => n231);
   U109 : AOI22_X1 port map( A1 => A_s(10), A2 => n180, B1 => A_ns(10), B2 => 
                           n167, ZN => n139);
   U110 : AOI221_X1 port map( B1 => net39408, B2 => A_ns(14), C1 => n176, C2 =>
                           A_s(14), A => n225, ZN => n132);
   U111 : INV_X1 port map( A => n133, ZN => n225);
   U112 : AOI22_X1 port map( A1 => A_s(13), A2 => n179, B1 => A_ns(13), B2 => 
                           n167, ZN => n133);
   U113 : AOI221_X1 port map( B1 => net39408, B2 => A_ns(15), C1 => n176, C2 =>
                           A_s(15), A => n223, ZN => n130);
   U114 : INV_X1 port map( A => n131, ZN => n223);
   U115 : AOI22_X1 port map( A1 => A_s(14), A2 => n180, B1 => A_ns(14), B2 => 
                           n168, ZN => n131);
   U116 : AOI221_X1 port map( B1 => net39408, B2 => A_ns(16), C1 => n176, C2 =>
                           A_s(16), A => n221, ZN => n128);
   U117 : INV_X1 port map( A => n129, ZN => n221);
   U118 : AOI22_X1 port map( A1 => A_s(15), A2 => n179, B1 => A_ns(15), B2 => 
                           n169, ZN => n129);
   U119 : AOI221_X1 port map( B1 => net39408, B2 => A_ns(17), C1 => n176, C2 =>
                           A_s(17), A => n219, ZN => n126);
   U120 : INV_X1 port map( A => n127, ZN => n219);
   U121 : AOI22_X1 port map( A1 => A_s(16), A2 => n180, B1 => A_ns(16), B2 => 
                           n167, ZN => n127);
   U122 : AOI221_X1 port map( B1 => net39408, B2 => A_ns(31), C1 => n176, C2 =>
                           A_s(31), A => n191, ZN => n96);
   U123 : INV_X1 port map( A => n97, ZN => n191);
   U124 : AOI221_X1 port map( B1 => net40345, B2 => A_ns(30), C1 => n177, C2 =>
                           A_s(30), A => n193, ZN => n98);
   U125 : INV_X1 port map( A => n99, ZN => n193);
   U126 : AOI221_X1 port map( B1 => net39408, B2 => A_ns(29), C1 => n176, C2 =>
                           A_s(29), A => n195, ZN => n100);
   U127 : INV_X1 port map( A => n101, ZN => n195);
   U128 : AOI221_X1 port map( B1 => net39408, B2 => A_ns(12), C1 => n176, C2 =>
                           A_s(12), A => n229, ZN => n136);
   U129 : INV_X1 port map( A => n137, ZN => n229);
   U130 : AOI22_X1 port map( A1 => A_s(11), A2 => n179, B1 => A_ns(11), B2 => 
                           n168, ZN => n137);
   U131 : INV_X1 port map( A => n119, ZN => n211);
   U132 : AOI22_X1 port map( A1 => A_s(20), A2 => n180, B1 => A_ns(20), B2 => 
                           n168, ZN => n119);
   U133 : INV_X1 port map( A => n123, ZN => n215);
   U134 : AOI22_X1 port map( A1 => A_s(18), A2 => n180, B1 => A_ns(18), B2 => 
                           n169, ZN => n123);
   U135 : INV_X1 port map( A => n117, ZN => n209);
   U136 : AOI22_X1 port map( A1 => A_s(21), A2 => n179, B1 => A_ns(21), B2 => 
                           n169, ZN => n117);
   U137 : INV_X1 port map( A => n115, ZN => n207);
   U138 : AOI22_X1 port map( A1 => A_s(22), A2 => n180, B1 => A_ns(22), B2 => 
                           n167, ZN => n115);
   U139 : INV_X1 port map( A => n113, ZN => n205);
   U140 : AOI22_X1 port map( A1 => A_s(23), A2 => n179, B1 => A_ns(23), B2 => 
                           n168, ZN => n113);
   U141 : AOI22_X1 port map( A1 => A_ns(34), A2 => net40345, B1 => A_s(34), B2 
                           => n176, ZN => n91);
   U142 : AOI221_X1 port map( B1 => net39408, B2 => A_ns(13), C1 => n176, C2 =>
                           A_s(13), A => n227, ZN => n134);
   U143 : INV_X1 port map( A => n135, ZN => n227);
   U144 : AOI22_X1 port map( A1 => A_s(12), A2 => n180, B1 => A_ns(12), B2 => 
                           n169, ZN => n135);
   U145 : AOI221_X1 port map( B1 => net40345, B2 => A_ns(20), C1 => n176, C2 =>
                           A_s(20), A => n213, ZN => n120);
   U146 : INV_X1 port map( A => n121, ZN => n213);
   U147 : AOI22_X1 port map( A1 => A_s(19), A2 => n179, B1 => A_ns(19), B2 => 
                           n167, ZN => n121);
   U148 : INV_X1 port map( A => n72, ZN => O_1_port);
   U149 : AOI22_X1 port map( A1 => n150, A2 => A_s(0), B1 => net40345, B2 => 
                           A_ns(0), ZN => n72);
   U150 : INV_X1 port map( A => n84, ZN => O_5_port);
   U151 : AOI22_X1 port map( A1 => A_s(32), A2 => n180, B1 => A_ns(32), B2 => 
                           n168, ZN => n93);
   U152 : AOI22_X1 port map( A1 => A_s(31), A2 => n179, B1 => A_ns(31), B2 => 
                           n167, ZN => n95);
   U153 : AOI22_X1 port map( A1 => A_s(30), A2 => n180, B1 => A_ns(30), B2 => 
                           n169, ZN => n97);
   U154 : AOI22_X1 port map( A1 => A_s(29), A2 => n179, B1 => A_ns(29), B2 => 
                           n168, ZN => n99);
   U155 : AOI22_X1 port map( A1 => A_s(28), A2 => n180, B1 => A_ns(28), B2 => 
                           n167, ZN => n101);
   U156 : AOI22_X1 port map( A1 => A_s(8), A2 => n180, B1 => A_ns(8), B2 => 
                           n168, ZN => n143);
   U157 : AOI22_X1 port map( A1 => A_s(6), A2 => n180, B1 => A_ns(6), B2 => 
                           n169, ZN => n79);
   U158 : AOI22_X1 port map( A1 => A_s(5), A2 => n179, B1 => A_ns(5), B2 => 
                           n168, ZN => n81);
   U159 : AOI22_X1 port map( A1 => A_s(4), A2 => n180, B1 => A_ns(4), B2 => 
                           n167, ZN => n83);
   U160 : AOI22_X1 port map( A1 => A_s(3), A2 => n178, B1 => A_ns(3), B2 => 
                           n169, ZN => n85);
   U161 : AOI22_X1 port map( A1 => A_s(2), A2 => n178, B1 => A_ns(2), B2 => 
                           n168, ZN => n87);
   U162 : NOR3_X1 port map( A1 => net40332, A2 => net41959, A3 => net35751, ZN 
                           => n77);
   U163 : AOI221_X1 port map( B1 => net40345, B2 => A_ns(28), C1 => n176, C2 =>
                           A_s(28), A => n197, ZN => n104);
   U164 : AOI221_X1 port map( B1 => net39408, B2 => A_ns(27), C1 => n176, C2 =>
                           A_s(27), A => n199, ZN => n106);
   U165 : AOI221_X1 port map( B1 => net40345, B2 => A_ns(26), C1 => n177, C2 =>
                           A_s(26), A => n201, ZN => n108);
   U166 : AOI221_X1 port map( B1 => net39408, B2 => A_ns(25), C1 => n176, C2 =>
                           A_s(25), A => n203, ZN => n110);
   U167 : AOI221_X1 port map( B1 => net40345, B2 => A_ns(24), C1 => n176, C2 =>
                           A_s(24), A => n205, ZN => n112);
   U168 : AOI221_X1 port map( B1 => net39408, B2 => A_ns(23), C1 => n177, C2 =>
                           A_s(23), A => n207, ZN => n114);
   U169 : AOI221_X1 port map( B1 => net40345, B2 => A_ns(22), C1 => n176, C2 =>
                           A_s(22), A => n209, ZN => n116);
   U170 : AOI221_X1 port map( B1 => net39408, B2 => A_ns(21), C1 => n176, C2 =>
                           A_s(21), A => n211, ZN => n118);
   U171 : AOI221_X1 port map( B1 => net39408, B2 => A_ns(19), C1 => n177, C2 =>
                           A_s(19), A => n215, ZN => n122);
   U172 : AOI221_X1 port map( B1 => net40345, B2 => A_ns(18), C1 => n176, C2 =>
                           A_s(18), A => n217, ZN => n124);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT34_i0 is

   port( A_s, A_ns, B : in std_logic_vector (33 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (33 downto 0));

end BOOTHENC_NBIT34_i0;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT34_i0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X4
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n81, n82, A_nso_3_port, n84, n85, A_nso_2_port, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, A_nso_4_port, n99, 
      A_nso_5_port, n101, n102, A_nso_7_port, n104, A_nso_8_port, n106, 
      A_nso_9_port, n108, A_nso_10_port, n110, A_nso_11_port, n112, 
      A_nso_12_port, n114, A_nso_13_port, n116, A_nso_14_port, n118, 
      A_nso_15_port, n120, A_nso_16_port, n122, A_nso_17_port, n124, 
      A_nso_18_port, n126, A_nso_19_port, n128, A_nso_20_port, n130, 
      A_nso_21_port, n132, A_nso_22_port, n134, A_nso_23_port, n136, 
      A_nso_24_port, n138, A_nso_25_port, n140, A_nso_26_port, n142, 
      A_nso_27_port, n144, A_nso_28_port, n146, A_nso_29_port, n148, 
      A_nso_30_port, n150, A_nso_31_port, n152, A_nso_32_port, n154, n155, n156
      , A_nso_1_port, n158, n159, n160 : std_logic;

begin
   A_so <= ( A_s(32), A_s(31), A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), 
      A_s(25), A_s(24), A_s(23), A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), 
      A_s(17), A_s(16), A_s(15), A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), 
      A_s(9), A_s(8), A_s(7), A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), 
      A_s(0), X_Logic0_port );
   A_nso <= ( A_ns(32), A_nso_32_port, A_nso_31_port, A_nso_30_port, 
      A_nso_29_port, A_nso_28_port, A_nso_27_port, A_nso_26_port, A_nso_25_port
      , A_nso_24_port, A_nso_23_port, A_nso_22_port, A_nso_21_port, 
      A_nso_20_port, A_nso_19_port, A_nso_18_port, A_nso_17_port, A_nso_16_port
      , A_nso_15_port, A_nso_14_port, A_nso_13_port, A_nso_12_port, 
      A_nso_11_port, A_nso_10_port, A_nso_9_port, A_nso_8_port, A_nso_7_port, 
      A_ns(5), A_nso_5_port, A_nso_4_port, A_nso_3_port, A_nso_2_port, 
      A_nso_1_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U3 : OAI221_X4 port map( B1 => n80, B2 => n152, C1 => n84, C2 => n154, A => 
                           n49, ZN => O(31));
   U4 : OAI221_X4 port map( B1 => n79, B2 => n140, C1 => n93, C2 => n142, A => 
                           n56, ZN => O(25));
   U5 : OAI221_X4 port map( B1 => n80, B2 => n132, C1 => n84, C2 => n134, A => 
                           n60, ZN => O(21));
   U6 : OAI221_X1 port map( B1 => n79, B2 => n120, C1 => n84, C2 => n122, A => 
                           n67, ZN => O(15));
   U7 : OAI221_X1 port map( B1 => n80, B2 => n106, C1 => n108, C2 => n84, A => 
                           n41, ZN => O(8));
   U8 : OAI221_X1 port map( B1 => n95, B2 => n110, C1 => n85, C2 => n112, A => 
                           n72, ZN => O(10));
   U9 : OAI221_X1 port map( B1 => n94, B2 => n112, C1 => n84, C2 => n114, A => 
                           n71, ZN => O(11));
   U10 : OAI221_X1 port map( B1 => n79, B2 => n102, C1 => n85, C2 => n104, A =>
                           n43, ZN => O(6));
   U11 : OAI221_X1 port map( B1 => n94, B2 => n104, C1 => n84, C2 => n106, A =>
                           n42, ZN => O(7));
   U12 : OAI221_X1 port map( B1 => n79, B2 => n108, C1 => n84, C2 => n110, A =>
                           n40, ZN => O(9));
   U13 : OAI221_X1 port map( B1 => n94, B2 => n122, C1 => n92, C2 => n124, A =>
                           n66, ZN => O(16));
   U14 : OAI221_X1 port map( B1 => n95, B2 => n124, C1 => n93, C2 => n126, A =>
                           n65, ZN => O(17));
   U15 : OAI221_X1 port map( B1 => n79, B2 => n128, C1 => n84, C2 => n130, A =>
                           n63, ZN => O(19));
   U16 : OAI222_X1 port map( A1 => n159, A2 => n76, B1 => n155, B2 => n95, C1 
                           => n156, C2 => n85, ZN => O(33));
   U17 : OAI221_X1 port map( B1 => n79, B2 => n134, C1 => n92, C2 => n136, A =>
                           n59, ZN => O(22));
   U18 : INV_X1 port map( A => A_ns(10), ZN => n112);
   U19 : INV_X1 port map( A => A_ns(14), ZN => n120);
   U20 : INV_X1 port map( A => A_ns(29), ZN => n150);
   U21 : CLKBUF_X1 port map( A => n158, Z => n74);
   U22 : OAI221_X4 port map( B1 => n80, B2 => n118, C1 => n85, C2 => n120, A =>
                           n68, ZN => O(14));
   U23 : OAI221_X1 port map( B1 => n75, B2 => n38, C1 => n99, C2 => n78, A => 
                           n46, ZN => O(3));
   U24 : BUF_X1 port map( A => n97, Z => n75);
   U25 : OAI221_X1 port map( B1 => n96, B2 => n38, C1 => n97, C2 => n39, A => 
                           n51, ZN => O(2));
   U26 : INV_X2 port map( A => n106, ZN => A_nso_8_port);
   U27 : OAI221_X4 port map( B1 => n80, B2 => n126, C1 => n85, C2 => n128, A =>
                           n64, ZN => O(18));
   U28 : BUF_X1 port map( A => n38, Z => n94);
   U29 : BUF_X2 port map( A => n81, Z => n88);
   U30 : OAI221_X4 port map( B1 => n94, B2 => n130, C1 => n85, C2 => n132, A =>
                           n61, ZN => O(20));
   U31 : INV_X1 port map( A => n101, ZN => A_nso_5_port);
   U32 : CLKBUF_X1 port map( A => A_ns(2), Z => A_nso_3_port);
   U33 : INV_X2 port map( A => n158, ZN => A_nso_1_port);
   U34 : INV_X1 port map( A => n88, ZN => n76);
   U35 : AND2_X2 port map( A1 => B(0), A2 => n82, ZN => n81);
   U36 : CLKBUF_X1 port map( A => n81, Z => n90);
   U37 : CLKBUF_X1 port map( A => n81, Z => n91);
   U38 : INV_X2 port map( A => n99, ZN => A_nso_4_port);
   U39 : NAND2_X1 port map( A1 => B(0), A2 => n47, ZN => n77);
   U40 : NAND2_X1 port map( A1 => B(0), A2 => n47, ZN => n78);
   U41 : BUF_X2 port map( A => n38, Z => n79);
   U42 : BUF_X2 port map( A => n38, Z => n80);
   U43 : OAI221_X1 port map( B1 => n79, B2 => n101, C1 => n85, C2 => n102, A =>
                           n44, ZN => O(5));
   U44 : OR2_X2 port map( A1 => n160, A2 => B(0), ZN => n38);
   U45 : OAI221_X1 port map( B1 => n79, B2 => n99, C1 => n101, C2 => n85, A => 
                           n45, ZN => O(4));
   U46 : INV_X1 port map( A => B(1), ZN => n82);
   U47 : CLKBUF_X3 port map( A => n77, Z => n84);
   U48 : CLKBUF_X3 port map( A => n78, Z => n85);
   U49 : BUF_X2 port map( A => A_ns(1), Z => A_nso_2_port);
   U50 : CLKBUF_X1 port map( A => n81, Z => n87);
   U51 : CLKBUF_X1 port map( A => n38, Z => n95);
   U52 : CLKBUF_X1 port map( A => n81, Z => n89);
   U53 : CLKBUF_X1 port map( A => n78, Z => n92);
   U54 : CLKBUF_X1 port map( A => n77, Z => n93);
   U55 : INV_X1 port map( A => A_ns(31), ZN => n154);
   U56 : INV_X1 port map( A => A_ns(32), ZN => n155);
   U57 : OAI221_X1 port map( B1 => n79, B2 => n154, C1 => n84, C2 => n155, A =>
                           n48, ZN => O(32));
   U58 : NAND2_X1 port map( A1 => A_s(32), A2 => n88, ZN => n48);
   U59 : NAND2_X1 port map( A1 => A_s(31), A2 => n87, ZN => n49);
   U60 : OAI221_X1 port map( B1 => n94, B2 => n150, C1 => n85, C2 => n152, A =>
                           n50, ZN => O(30));
   U61 : NAND2_X1 port map( A1 => A_s(30), A2 => n88, ZN => n50);
   U62 : NAND2_X1 port map( A1 => A_s(7), A2 => n88, ZN => n42);
   U63 : NAND2_X1 port map( A1 => A_s(8), A2 => n88, ZN => n41);
   U64 : NAND2_X1 port map( A1 => A_s(9), A2 => n88, ZN => n40);
   U65 : NAND2_X1 port map( A1 => A_s(10), A2 => n88, ZN => n72);
   U66 : NAND2_X1 port map( A1 => A_s(11), A2 => n88, ZN => n71);
   U67 : OAI221_X1 port map( B1 => n80, B2 => n114, C1 => n92, C2 => n116, A =>
                           n70, ZN => O(12));
   U68 : NAND2_X1 port map( A1 => A_s(12), A2 => n88, ZN => n70);
   U69 : OAI221_X1 port map( B1 => n79, B2 => n116, C1 => n93, C2 => n118, A =>
                           n69, ZN => O(13));
   U70 : NAND2_X1 port map( A1 => A_s(13), A2 => n88, ZN => n69);
   U71 : NAND2_X1 port map( A1 => A_s(14), A2 => n88, ZN => n68);
   U72 : NAND2_X1 port map( A1 => A_s(15), A2 => n88, ZN => n67);
   U73 : NAND2_X1 port map( A1 => A_s(16), A2 => n88, ZN => n66);
   U74 : NAND2_X1 port map( A1 => A_s(17), A2 => n88, ZN => n65);
   U75 : NAND2_X1 port map( A1 => A_s(18), A2 => n88, ZN => n64);
   U76 : NAND2_X1 port map( A1 => A_s(19), A2 => n88, ZN => n63);
   U77 : NAND2_X1 port map( A1 => A_s(20), A2 => n87, ZN => n61);
   U78 : NAND2_X1 port map( A1 => A_s(21), A2 => n88, ZN => n60);
   U79 : NAND2_X1 port map( A1 => A_s(22), A2 => n87, ZN => n59);
   U80 : OAI221_X1 port map( B1 => n94, B2 => n136, C1 => n85, C2 => n138, A =>
                           n58, ZN => O(23));
   U81 : NAND2_X1 port map( A1 => A_s(23), A2 => n88, ZN => n58);
   U82 : OAI221_X1 port map( B1 => n80, B2 => n138, C1 => n84, C2 => n140, A =>
                           n57, ZN => O(24));
   U83 : NAND2_X1 port map( A1 => A_s(24), A2 => n87, ZN => n57);
   U84 : NAND2_X1 port map( A1 => A_s(25), A2 => n87, ZN => n56);
   U85 : OAI221_X1 port map( B1 => n94, B2 => n142, C1 => n85, C2 => n144, A =>
                           n55, ZN => O(26));
   U86 : NAND2_X1 port map( A1 => A_s(26), A2 => n88, ZN => n55);
   U87 : OAI221_X1 port map( B1 => n95, B2 => n144, C1 => n84, C2 => n146, A =>
                           n54, ZN => O(27));
   U88 : NAND2_X1 port map( A1 => A_s(27), A2 => n87, ZN => n54);
   U89 : OAI221_X1 port map( B1 => n80, B2 => n146, C1 => n92, C2 => n148, A =>
                           n53, ZN => O(28));
   U90 : NAND2_X1 port map( A1 => A_s(28), A2 => n88, ZN => n53);
   U91 : OAI221_X1 port map( B1 => n79, B2 => n148, C1 => n93, C2 => n150, A =>
                           n52, ZN => O(29));
   U92 : NAND2_X1 port map( A1 => A_s(29), A2 => n87, ZN => n52);
   U93 : NAND2_X1 port map( A1 => A_s(6), A2 => n87, ZN => n43);
   U94 : NAND2_X1 port map( A1 => A_s(5), A2 => n89, ZN => n44);
   U95 : NAND2_X1 port map( A1 => A_s(4), A2 => n91, ZN => n45);
   U96 : NAND2_X1 port map( A1 => A_s(3), A2 => n90, ZN => n46);
   U97 : NAND2_X1 port map( A1 => A_s(2), A2 => n81, ZN => n51);
   U98 : INV_X1 port map( A => A_ns(3), ZN => n99);
   U99 : INV_X1 port map( A => A_ns(5), ZN => n102);
   U100 : INV_X1 port map( A => A_ns(7), ZN => n106);
   U101 : INV_X1 port map( A => A_ns(4), ZN => n101);
   U102 : INV_X1 port map( A => A_ns(0), ZN => n158);
   U103 : INV_X1 port map( A => A_ns(8), ZN => n108);
   U104 : INV_X1 port map( A => A_ns(1), ZN => n96);
   U105 : INV_X1 port map( A => A_ns(2), ZN => n97);
   U106 : INV_X1 port map( A => A_ns(6), ZN => n104);
   U107 : INV_X1 port map( A => A_ns(11), ZN => n114);
   U108 : INV_X1 port map( A => A_ns(21), ZN => n134);
   U109 : INV_X1 port map( A => A_ns(26), ZN => n144);
   U110 : INV_X1 port map( A => A_ns(20), ZN => n132);
   U111 : INV_X1 port map( A => A_ns(24), ZN => n140);
   U112 : INV_X1 port map( A => A_ns(30), ZN => n152);
   U113 : INV_X1 port map( A => A_ns(9), ZN => n110);
   U114 : INV_X1 port map( A => A_ns(13), ZN => n118);
   U115 : INV_X1 port map( A => A_ns(15), ZN => n122);
   U116 : INV_X1 port map( A => A_ns(17), ZN => n126);
   U117 : INV_X1 port map( A => A_ns(18), ZN => n128);
   U118 : INV_X1 port map( A => A_ns(19), ZN => n130);
   U119 : INV_X1 port map( A => A_ns(27), ZN => n146);
   U120 : INV_X1 port map( A => A_ns(23), ZN => n138);
   U121 : INV_X1 port map( A => A_ns(25), ZN => n142);
   U122 : INV_X1 port map( A => A_ns(12), ZN => n116);
   U123 : INV_X1 port map( A => A_ns(16), ZN => n124);
   U124 : INV_X1 port map( A => A_ns(28), ZN => n148);
   U125 : INV_X1 port map( A => A_ns(22), ZN => n136);
   U126 : OAI221_X1 port map( B1 => n94, B2 => n74, C1 => n93, C2 => n96, A => 
                           n62, ZN => O(1));
   U127 : NAND2_X1 port map( A1 => A_s(1), A2 => n87, ZN => n62);
   U128 : OAI21_X1 port map( B1 => n92, B2 => n74, A => n73, ZN => O(0));
   U129 : NAND2_X1 port map( A1 => A_s(0), A2 => n87, ZN => n73);
   U130 : NAND2_X1 port map( A1 => B(0), A2 => n82, ZN => n47);
   U131 : NAND2_X1 port map( A1 => B(0), A2 => n47, ZN => n39);
   U132 : INV_X1 port map( A => B(1), ZN => n160);
   U133 : INV_X1 port map( A => n104, ZN => A_nso_7_port);
   U134 : INV_X1 port map( A => n108, ZN => A_nso_9_port);
   U135 : INV_X1 port map( A => n110, ZN => A_nso_10_port);
   U136 : INV_X1 port map( A => n112, ZN => A_nso_11_port);
   U137 : INV_X1 port map( A => n114, ZN => A_nso_12_port);
   U138 : INV_X1 port map( A => n116, ZN => A_nso_13_port);
   U139 : INV_X1 port map( A => n118, ZN => A_nso_14_port);
   U140 : INV_X1 port map( A => n120, ZN => A_nso_15_port);
   U141 : INV_X1 port map( A => n122, ZN => A_nso_16_port);
   U142 : INV_X1 port map( A => n124, ZN => A_nso_17_port);
   U143 : INV_X1 port map( A => n126, ZN => A_nso_18_port);
   U144 : INV_X1 port map( A => n128, ZN => A_nso_19_port);
   U145 : INV_X1 port map( A => n130, ZN => A_nso_20_port);
   U146 : INV_X1 port map( A => n132, ZN => A_nso_21_port);
   U147 : INV_X1 port map( A => n134, ZN => A_nso_22_port);
   U148 : INV_X1 port map( A => n136, ZN => A_nso_23_port);
   U149 : INV_X1 port map( A => n138, ZN => A_nso_24_port);
   U150 : INV_X1 port map( A => n140, ZN => A_nso_25_port);
   U151 : INV_X1 port map( A => n142, ZN => A_nso_26_port);
   U152 : INV_X1 port map( A => n144, ZN => A_nso_27_port);
   U153 : INV_X1 port map( A => n146, ZN => A_nso_28_port);
   U154 : INV_X1 port map( A => n148, ZN => A_nso_29_port);
   U155 : INV_X1 port map( A => n150, ZN => A_nso_30_port);
   U156 : INV_X1 port map( A => n152, ZN => A_nso_31_port);
   U157 : INV_X1 port map( A => n154, ZN => A_nso_32_port);
   U158 : INV_X1 port map( A => A_ns(33), ZN => n156);
   U159 : INV_X1 port map( A => A_s(33), ZN => n159);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHMUL_NBIT32 is

   port( A, B : in std_logic_vector (31 downto 0);  S : out std_logic_vector 
         (63 downto 0));

end BOOTHMUL_NBIT32;

architecture SYN_BEHAVIOURAL of BOOTHMUL_NBIT32 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BOOTHMUL_NBIT32_DW01_sub_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component RCA_NBIT64
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT62
      port( A, B : in std_logic_vector (61 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (61 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT60
      port( A, B : in std_logic_vector (59 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (59 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT58
      port( A, B : in std_logic_vector (57 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (57 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT56
      port( A, B : in std_logic_vector (55 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (55 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT54
      port( A, B : in std_logic_vector (53 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (53 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT52
      port( A, B : in std_logic_vector (51 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (51 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT50
      port( A, B : in std_logic_vector (49 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (49 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT48
      port( A, B : in std_logic_vector (47 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (47 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT46
      port( A, B : in std_logic_vector (45 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (45 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT44
      port( A, B : in std_logic_vector (43 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (43 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT42
      port( A, B : in std_logic_vector (41 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (41 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT40
      port( A, B : in std_logic_vector (39 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (39 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT38
      port( A, B : in std_logic_vector (37 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (37 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT36
      port( A, B : in std_logic_vector (35 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (35 downto 0);  Co : out std_logic);
   end component;
   
   component BOOTHENC_NBIT64_i30
      port( A_s, A_ns, B : in std_logic_vector (63 downto 0);  O, A_so, A_nso :
            out std_logic_vector (63 downto 0));
   end component;
   
   component BOOTHENC_NBIT62_i28
      port( A_s, A_ns, B : in std_logic_vector (61 downto 0);  O, A_so, A_nso :
            out std_logic_vector (61 downto 0));
   end component;
   
   component BOOTHENC_NBIT60_i26
      port( A_s, A_ns, B : in std_logic_vector (59 downto 0);  O, A_so, A_nso :
            out std_logic_vector (59 downto 0));
   end component;
   
   component BOOTHENC_NBIT58_i24
      port( A_s, A_ns, B : in std_logic_vector (57 downto 0);  O, A_so, A_nso :
            out std_logic_vector (57 downto 0));
   end component;
   
   component BOOTHENC_NBIT56_i22
      port( A_s, A_ns, B : in std_logic_vector (55 downto 0);  O, A_so, A_nso :
            out std_logic_vector (55 downto 0));
   end component;
   
   component BOOTHENC_NBIT54_i20
      port( A_s, A_ns, B : in std_logic_vector (53 downto 0);  O, A_so, A_nso :
            out std_logic_vector (53 downto 0));
   end component;
   
   component BOOTHENC_NBIT52_i18
      port( A_s, A_ns, B : in std_logic_vector (51 downto 0);  O, A_so, A_nso :
            out std_logic_vector (51 downto 0));
   end component;
   
   component BOOTHENC_NBIT50_i16
      port( A_s, A_ns, B : in std_logic_vector (49 downto 0);  O, A_so, A_nso :
            out std_logic_vector (49 downto 0));
   end component;
   
   component BOOTHENC_NBIT48_i14
      port( A_s, A_ns, B : in std_logic_vector (47 downto 0);  O, A_so, A_nso :
            out std_logic_vector (47 downto 0));
   end component;
   
   component BOOTHENC_NBIT46_i12
      port( A_s, A_ns, B : in std_logic_vector (45 downto 0);  O, A_so, A_nso :
            out std_logic_vector (45 downto 0));
   end component;
   
   component BOOTHENC_NBIT44_i10
      port( A_s, A_ns, B : in std_logic_vector (43 downto 0);  O, A_so, A_nso :
            out std_logic_vector (43 downto 0));
   end component;
   
   component BOOTHENC_NBIT42_i8
      port( A_s, A_ns, B : in std_logic_vector (41 downto 0);  O, A_so, A_nso :
            out std_logic_vector (41 downto 0));
   end component;
   
   component BOOTHENC_NBIT40_i6
      port( A_s, A_ns, B : in std_logic_vector (39 downto 0);  O, A_so, A_nso :
            out std_logic_vector (39 downto 0));
   end component;
   
   component BOOTHENC_NBIT38_i4
      port( A_s, A_ns, B : in std_logic_vector (37 downto 0);  O, A_so, A_nso :
            out std_logic_vector (37 downto 0));
   end component;
   
   component BOOTHENC_NBIT36_i2
      port( A_s, A_ns, B : in std_logic_vector (35 downto 0);  O, A_so, A_nso :
            out std_logic_vector (35 downto 0));
   end component;
   
   component BOOTHENC_NBIT34_i0
      port( A_s, A_ns, B : in std_logic_vector (33 downto 0);  O, A_so, A_nso :
            out std_logic_vector (33 downto 0));
   end component;
   
   signal X_Logic0_port, A_n_65, A_n_30_port, A_n_29_port, A_n_28_port, 
      A_n_27_port, A_n_26_port, A_n_25_port, A_n_24_port, A_n_23_port, 
      A_n_22_port, A_n_21_port, A_n_20_port, A_n_19_port, A_n_18_port, 
      A_n_17_port, A_n_16_port, A_n_15_port, A_n_14_port, A_n_13_port, 
      A_n_12_port, A_n_11_port, A_n_10_port, A_n_9_port, A_n_8_port, A_n_7_port
      , A_n_6_port, A_n_5_port, A_n_4_port, A_n_3_port, A_n_2_port, A_n_1_port,
      A_n_0_port, SHIFT_1_31_port, SHIFT_1_30_port, SHIFT_1_29_port, 
      SHIFT_1_28_port, SHIFT_1_27_port, SHIFT_1_26_port, SHIFT_1_25_port, 
      SHIFT_1_24_port, SHIFT_1_23_port, SHIFT_1_22_port, SHIFT_1_21_port, 
      SHIFT_1_20_port, SHIFT_1_19_port, SHIFT_1_18_port, SHIFT_1_17_port, 
      SHIFT_1_16_port, SHIFT_1_15_port, SHIFT_1_14_port, SHIFT_1_13_port, 
      SHIFT_1_12_port, SHIFT_1_11_port, SHIFT_1_10_port, SHIFT_1_9_port, 
      SHIFT_1_8_port, SHIFT_1_7_port, SHIFT_1_6_port, SHIFT_1_5_port, 
      SHIFT_1_4_port, SHIFT_1_3_port, SHIFT_1_2_port, SHIFT_1_1_port, 
      SHIFT_1_0_port, SHIFT_15_61_port, SHIFT_15_60_port, SHIFT_15_59_port, 
      SHIFT_15_58_port, SHIFT_15_57_port, SHIFT_15_56_port, SHIFT_15_55_port, 
      SHIFT_15_54_port, SHIFT_15_53_port, SHIFT_15_52_port, SHIFT_15_51_port, 
      SHIFT_15_50_port, SHIFT_15_49_port, SHIFT_15_48_port, SHIFT_15_47_port, 
      SHIFT_15_46_port, SHIFT_15_45_port, SHIFT_15_44_port, SHIFT_15_43_port, 
      SHIFT_15_42_port, SHIFT_15_41_port, SHIFT_15_40_port, SHIFT_15_39_port, 
      SHIFT_15_38_port, SHIFT_15_37_port, SHIFT_15_36_port, SHIFT_15_35_port, 
      SHIFT_15_34_port, SHIFT_15_33_port, SHIFT_15_32_port, SHIFT_15_31_port, 
      SHIFT_15_30_port, SHIFT_15_29_port, SHIFT_15_28_port, SHIFT_15_27_port, 
      SHIFT_15_26_port, SHIFT_15_25_port, SHIFT_15_24_port, SHIFT_15_23_port, 
      SHIFT_15_22_port, SHIFT_15_21_port, SHIFT_15_20_port, SHIFT_15_19_port, 
      SHIFT_15_18_port, SHIFT_15_17_port, SHIFT_15_16_port, SHIFT_15_15_port, 
      SHIFT_15_14_port, SHIFT_15_13_port, SHIFT_15_12_port, SHIFT_15_11_port, 
      SHIFT_15_10_port, SHIFT_15_9_port, SHIFT_15_8_port, SHIFT_15_7_port, 
      SHIFT_15_6_port, SHIFT_15_5_port, SHIFT_15_4_port, SHIFT_15_3_port, 
      SHIFT_15_2_port, SHIFT_15_1_port, SHIFT_15_0_port, SHIFT_14_59_port, 
      SHIFT_14_58_port, SHIFT_14_57_port, SHIFT_14_56_port, SHIFT_14_55_port, 
      SHIFT_14_54_port, SHIFT_14_53_port, SHIFT_14_52_port, SHIFT_14_51_port, 
      SHIFT_14_50_port, SHIFT_14_49_port, SHIFT_14_48_port, SHIFT_14_47_port, 
      SHIFT_14_46_port, SHIFT_14_45_port, SHIFT_14_44_port, SHIFT_14_43_port, 
      SHIFT_14_42_port, SHIFT_14_41_port, SHIFT_14_40_port, SHIFT_14_39_port, 
      SHIFT_14_38_port, SHIFT_14_37_port, SHIFT_14_36_port, SHIFT_14_35_port, 
      SHIFT_14_34_port, SHIFT_14_33_port, SHIFT_14_32_port, SHIFT_14_31_port, 
      SHIFT_14_30_port, SHIFT_14_29_port, SHIFT_14_28_port, SHIFT_14_27_port, 
      SHIFT_14_26_port, SHIFT_14_25_port, SHIFT_14_24_port, SHIFT_14_23_port, 
      SHIFT_14_22_port, SHIFT_14_21_port, SHIFT_14_20_port, SHIFT_14_19_port, 
      SHIFT_14_18_port, SHIFT_14_17_port, SHIFT_14_16_port, SHIFT_14_15_port, 
      SHIFT_14_14_port, SHIFT_14_13_port, SHIFT_14_12_port, SHIFT_14_11_port, 
      SHIFT_14_10_port, SHIFT_14_9_port, SHIFT_14_8_port, SHIFT_14_7_port, 
      SHIFT_14_6_port, SHIFT_14_5_port, SHIFT_14_4_port, SHIFT_14_3_port, 
      SHIFT_14_2_port, SHIFT_14_1_port, SHIFT_14_0_port, SHIFT_13_57_port, 
      SHIFT_13_56_port, SHIFT_13_55_port, SHIFT_13_54_port, SHIFT_13_53_port, 
      SHIFT_13_52_port, SHIFT_13_51_port, SHIFT_13_50_port, SHIFT_13_49_port, 
      SHIFT_13_48_port, SHIFT_13_47_port, SHIFT_13_46_port, SHIFT_13_45_port, 
      SHIFT_13_44_port, SHIFT_13_43_port, SHIFT_13_42_port, SHIFT_13_41_port, 
      SHIFT_13_40_port, SHIFT_13_39_port, SHIFT_13_38_port, SHIFT_13_37_port, 
      SHIFT_13_36_port, SHIFT_13_35_port, SHIFT_13_34_port, SHIFT_13_33_port, 
      SHIFT_13_32_port, SHIFT_13_31_port, SHIFT_13_30_port, SHIFT_13_29_port, 
      SHIFT_13_28_port, SHIFT_13_27_port, SHIFT_13_26_port, SHIFT_13_25_port, 
      SHIFT_13_24_port, SHIFT_13_23_port, SHIFT_13_22_port, SHIFT_13_21_port, 
      SHIFT_13_20_port, SHIFT_13_19_port, SHIFT_13_18_port, SHIFT_13_17_port, 
      SHIFT_13_16_port, SHIFT_13_15_port, SHIFT_13_14_port, SHIFT_13_13_port, 
      SHIFT_13_12_port, SHIFT_13_11_port, SHIFT_13_10_port, SHIFT_13_9_port, 
      SHIFT_13_8_port, SHIFT_13_7_port, SHIFT_13_6_port, SHIFT_13_5_port, 
      SHIFT_13_4_port, SHIFT_13_3_port, SHIFT_13_2_port, SHIFT_13_1_port, 
      SHIFT_13_0_port, SHIFT_12_55_port, SHIFT_12_54_port, SHIFT_12_53_port, 
      SHIFT_12_52_port, SHIFT_12_51_port, SHIFT_12_50_port, SHIFT_12_49_port, 
      SHIFT_12_48_port, SHIFT_12_47_port, SHIFT_12_46_port, SHIFT_12_45_port, 
      SHIFT_12_44_port, SHIFT_12_43_port, SHIFT_12_42_port, SHIFT_12_41_port, 
      SHIFT_12_40_port, SHIFT_12_39_port, SHIFT_12_38_port, SHIFT_12_37_port, 
      SHIFT_12_36_port, SHIFT_12_35_port, SHIFT_12_34_port, SHIFT_12_33_port, 
      SHIFT_12_32_port, SHIFT_12_31_port, SHIFT_12_30_port, SHIFT_12_29_port, 
      SHIFT_12_28_port, SHIFT_12_27_port, SHIFT_12_26_port, SHIFT_12_25_port, 
      SHIFT_12_24_port, SHIFT_12_23_port, SHIFT_12_22_port, SHIFT_12_21_port, 
      SHIFT_12_20_port, SHIFT_12_19_port, SHIFT_12_18_port, SHIFT_12_17_port, 
      SHIFT_12_16_port, SHIFT_12_15_port, SHIFT_12_14_port, SHIFT_12_13_port, 
      SHIFT_12_12_port, SHIFT_12_11_port, SHIFT_12_10_port, SHIFT_12_9_port, 
      SHIFT_12_8_port, SHIFT_12_7_port, SHIFT_12_6_port, SHIFT_12_5_port, 
      SHIFT_12_4_port, SHIFT_12_3_port, SHIFT_12_2_port, SHIFT_12_1_port, 
      SHIFT_12_0_port, SHIFT_11_53_port, SHIFT_11_52_port, SHIFT_11_51_port, 
      SHIFT_11_50_port, SHIFT_11_49_port, SHIFT_11_48_port, SHIFT_11_47_port, 
      SHIFT_11_46_port, SHIFT_11_45_port, SHIFT_11_44_port, SHIFT_11_43_port, 
      SHIFT_11_42_port, SHIFT_11_41_port, SHIFT_11_40_port, SHIFT_11_39_port, 
      SHIFT_11_38_port, SHIFT_11_37_port, SHIFT_11_36_port, SHIFT_11_35_port, 
      SHIFT_11_34_port, SHIFT_11_33_port, SHIFT_11_32_port, SHIFT_11_31_port, 
      SHIFT_11_30_port, SHIFT_11_29_port, SHIFT_11_28_port, SHIFT_11_27_port, 
      SHIFT_11_26_port, SHIFT_11_25_port, SHIFT_11_24_port, SHIFT_11_23_port, 
      SHIFT_11_22_port, SHIFT_11_21_port, SHIFT_11_20_port, SHIFT_11_19_port, 
      SHIFT_11_18_port, SHIFT_11_17_port, SHIFT_11_16_port, SHIFT_11_15_port, 
      SHIFT_11_14_port, SHIFT_11_13_port, SHIFT_11_12_port, SHIFT_11_11_port, 
      SHIFT_11_10_port, SHIFT_11_9_port, SHIFT_11_8_port, SHIFT_11_7_port, 
      SHIFT_11_6_port, SHIFT_11_5_port, SHIFT_11_4_port, SHIFT_11_3_port, 
      SHIFT_11_2_port, SHIFT_11_1_port, SHIFT_11_0_port, SHIFT_10_51_port, 
      SHIFT_10_50_port, SHIFT_10_49_port, SHIFT_10_48_port, SHIFT_10_47_port, 
      SHIFT_10_46_port, SHIFT_10_45_port, SHIFT_10_44_port, SHIFT_10_43_port, 
      SHIFT_10_42_port, SHIFT_10_41_port, SHIFT_10_40_port, SHIFT_10_39_port, 
      SHIFT_10_38_port, SHIFT_10_37_port, SHIFT_10_36_port, SHIFT_10_35_port, 
      SHIFT_10_34_port, SHIFT_10_33_port, SHIFT_10_32_port, SHIFT_10_31_port, 
      SHIFT_10_30_port, SHIFT_10_29_port, SHIFT_10_28_port, SHIFT_10_27_port, 
      SHIFT_10_26_port, SHIFT_10_25_port, SHIFT_10_24_port, SHIFT_10_23_port, 
      SHIFT_10_22_port, SHIFT_10_21_port, SHIFT_10_20_port, SHIFT_10_19_port, 
      SHIFT_10_18_port, SHIFT_10_17_port, SHIFT_10_16_port, SHIFT_10_15_port, 
      SHIFT_10_14_port, SHIFT_10_13_port, SHIFT_10_12_port, SHIFT_10_11_port, 
      SHIFT_10_10_port, SHIFT_10_9_port, SHIFT_10_8_port, SHIFT_10_7_port, 
      SHIFT_10_6_port, SHIFT_10_5_port, SHIFT_10_4_port, SHIFT_10_3_port, 
      SHIFT_10_2_port, SHIFT_10_1_port, SHIFT_10_0_port, SHIFT_9_49_port, 
      SHIFT_9_48_port, SHIFT_9_47_port, SHIFT_9_46_port, SHIFT_9_45_port, 
      SHIFT_9_44_port, SHIFT_9_43_port, SHIFT_9_42_port, SHIFT_9_41_port, 
      SHIFT_9_40_port, SHIFT_9_39_port, SHIFT_9_38_port, SHIFT_9_37_port, 
      SHIFT_9_36_port, SHIFT_9_35_port, SHIFT_9_34_port, SHIFT_9_33_port, 
      SHIFT_9_32_port, SHIFT_9_31_port, SHIFT_9_30_port, SHIFT_9_29_port, 
      SHIFT_9_28_port, SHIFT_9_27_port, SHIFT_9_26_port, SHIFT_9_25_port, 
      SHIFT_9_24_port, SHIFT_9_23_port, SHIFT_9_22_port, SHIFT_9_21_port, 
      SHIFT_9_20_port, SHIFT_9_19_port, SHIFT_9_18_port, SHIFT_9_17_port, 
      SHIFT_9_16_port, SHIFT_9_15_port, SHIFT_9_14_port, SHIFT_9_13_port, 
      SHIFT_9_12_port, SHIFT_9_11_port, SHIFT_9_10_port, SHIFT_9_9_port, 
      SHIFT_9_8_port, SHIFT_9_7_port, SHIFT_9_6_port, SHIFT_9_5_port, 
      SHIFT_9_4_port, SHIFT_9_3_port, SHIFT_9_2_port, SHIFT_9_1_port, 
      SHIFT_9_0_port, SHIFT_8_47_port, SHIFT_8_46_port, SHIFT_8_45_port, 
      SHIFT_8_44_port, SHIFT_8_43_port, SHIFT_8_42_port, SHIFT_8_41_port, 
      SHIFT_8_40_port, SHIFT_8_39_port, SHIFT_8_38_port, SHIFT_8_37_port, 
      SHIFT_8_36_port, SHIFT_8_35_port, SHIFT_8_34_port, SHIFT_8_33_port, 
      SHIFT_8_32_port, SHIFT_8_31_port, SHIFT_8_30_port, SHIFT_8_29_port, 
      SHIFT_8_28_port, SHIFT_8_27_port, SHIFT_8_26_port, SHIFT_8_25_port, 
      SHIFT_8_24_port, SHIFT_8_23_port, SHIFT_8_22_port, SHIFT_8_21_port, 
      SHIFT_8_20_port, SHIFT_8_19_port, SHIFT_8_18_port, SHIFT_8_17_port, 
      SHIFT_8_16_port, SHIFT_8_15_port, SHIFT_8_14_port, SHIFT_8_13_port, 
      SHIFT_8_12_port, SHIFT_8_11_port, SHIFT_8_10_port, SHIFT_8_9_port, 
      SHIFT_8_8_port, SHIFT_8_7_port, SHIFT_8_6_port, SHIFT_8_5_port, 
      SHIFT_8_4_port, SHIFT_8_3_port, SHIFT_8_2_port, SHIFT_8_1_port, 
      SHIFT_8_0_port, SHIFT_7_45_port, SHIFT_7_44_port, SHIFT_7_43_port, 
      SHIFT_7_42_port, SHIFT_7_41_port, SHIFT_7_40_port, SHIFT_7_39_port, 
      SHIFT_7_38_port, SHIFT_7_37_port, SHIFT_7_36_port, SHIFT_7_35_port, 
      SHIFT_7_34_port, SHIFT_7_33_port, SHIFT_7_32_port, SHIFT_7_31_port, 
      SHIFT_7_30_port, SHIFT_7_29_port, SHIFT_7_28_port, SHIFT_7_27_port, 
      SHIFT_7_26_port, SHIFT_7_25_port, SHIFT_7_24_port, SHIFT_7_23_port, 
      SHIFT_7_22_port, SHIFT_7_21_port, SHIFT_7_20_port, SHIFT_7_19_port, 
      SHIFT_7_18_port, SHIFT_7_17_port, SHIFT_7_16_port, SHIFT_7_15_port, 
      SHIFT_7_14_port, SHIFT_7_13_port, SHIFT_7_12_port, SHIFT_7_11_port, 
      SHIFT_7_10_port, SHIFT_7_9_port, SHIFT_7_8_port, SHIFT_7_7_port, 
      SHIFT_7_6_port, SHIFT_7_5_port, SHIFT_7_4_port, SHIFT_7_3_port, 
      SHIFT_7_2_port, SHIFT_7_1_port, SHIFT_7_0_port, SHIFT_6_43_port, 
      SHIFT_6_42_port, SHIFT_6_41_port, SHIFT_6_40_port, SHIFT_6_39_port, 
      SHIFT_6_38_port, SHIFT_6_37_port, SHIFT_6_36_port, SHIFT_6_35_port, 
      SHIFT_6_34_port, SHIFT_6_33_port, SHIFT_6_32_port, SHIFT_6_31_port, 
      SHIFT_6_30_port, SHIFT_6_29_port, SHIFT_6_28_port, SHIFT_6_27_port, 
      SHIFT_6_26_port, SHIFT_6_25_port, SHIFT_6_24_port, SHIFT_6_23_port, 
      SHIFT_6_22_port, SHIFT_6_21_port, SHIFT_6_20_port, SHIFT_6_19_port, 
      SHIFT_6_18_port, SHIFT_6_17_port, SHIFT_6_16_port, SHIFT_6_15_port, 
      SHIFT_6_14_port, SHIFT_6_13_port, SHIFT_6_12_port, SHIFT_6_11_port, 
      SHIFT_6_10_port, SHIFT_6_9_port, SHIFT_6_8_port, SHIFT_6_7_port, 
      SHIFT_6_6_port, SHIFT_6_5_port, SHIFT_6_4_port, SHIFT_6_3_port, 
      SHIFT_6_2_port, SHIFT_6_1_port, SHIFT_6_0_port, SHIFT_5_41_port, 
      SHIFT_5_40_port, SHIFT_5_39_port, SHIFT_5_38_port, SHIFT_5_37_port, 
      SHIFT_5_36_port, SHIFT_5_35_port, SHIFT_5_34_port, SHIFT_5_33_port, 
      SHIFT_5_32_port, SHIFT_5_31_port, SHIFT_5_30_port, SHIFT_5_29_port, 
      SHIFT_5_28_port, SHIFT_5_27_port, SHIFT_5_26_port, SHIFT_5_25_port, 
      SHIFT_5_24_port, SHIFT_5_23_port, SHIFT_5_22_port, SHIFT_5_21_port, 
      SHIFT_5_20_port, SHIFT_5_19_port, SHIFT_5_18_port, SHIFT_5_17_port, 
      SHIFT_5_16_port, SHIFT_5_15_port, SHIFT_5_14_port, SHIFT_5_13_port, 
      SHIFT_5_12_port, SHIFT_5_11_port, SHIFT_5_10_port, SHIFT_5_9_port, 
      SHIFT_5_8_port, SHIFT_5_7_port, SHIFT_5_6_port, SHIFT_5_5_port, 
      SHIFT_5_4_port, SHIFT_5_3_port, SHIFT_5_2_port, SHIFT_5_1_port, 
      SHIFT_5_0_port, SHIFT_4_39_port, SHIFT_4_38_port, SHIFT_4_37_port, 
      SHIFT_4_36_port, SHIFT_4_35_port, SHIFT_4_34_port, SHIFT_4_33_port, 
      SHIFT_4_32_port, SHIFT_4_31_port, SHIFT_4_30_port, SHIFT_4_29_port, 
      SHIFT_4_28_port, SHIFT_4_27_port, SHIFT_4_26_port, SHIFT_4_25_port, 
      SHIFT_4_24_port, SHIFT_4_23_port, SHIFT_4_22_port, SHIFT_4_21_port, 
      SHIFT_4_20_port, SHIFT_4_19_port, SHIFT_4_18_port, SHIFT_4_17_port, 
      SHIFT_4_16_port, SHIFT_4_15_port, SHIFT_4_14_port, SHIFT_4_13_port, 
      SHIFT_4_12_port, SHIFT_4_11_port, SHIFT_4_10_port, SHIFT_4_9_port, 
      SHIFT_4_8_port, SHIFT_4_7_port, SHIFT_4_6_port, SHIFT_4_5_port, 
      SHIFT_4_4_port, SHIFT_4_3_port, SHIFT_4_2_port, SHIFT_4_1_port, 
      SHIFT_4_0_port, SHIFT_3_37_port, SHIFT_3_36_port, SHIFT_3_35_port, 
      SHIFT_3_34_port, SHIFT_3_33_port, SHIFT_3_32_port, SHIFT_3_31_port, 
      SHIFT_3_30_port, SHIFT_3_29_port, SHIFT_3_28_port, SHIFT_3_27_port, 
      SHIFT_3_26_port, SHIFT_3_25_port, SHIFT_3_24_port, SHIFT_3_23_port, 
      SHIFT_3_22_port, SHIFT_3_21_port, SHIFT_3_20_port, SHIFT_3_19_port, 
      SHIFT_3_18_port, SHIFT_3_17_port, SHIFT_3_16_port, SHIFT_3_15_port, 
      SHIFT_3_14_port, SHIFT_3_13_port, SHIFT_3_12_port, SHIFT_3_11_port, 
      SHIFT_3_10_port, SHIFT_3_9_port, SHIFT_3_8_port, SHIFT_3_7_port, 
      SHIFT_3_6_port, SHIFT_3_5_port, SHIFT_3_4_port, SHIFT_3_3_port, 
      SHIFT_3_2_port, SHIFT_3_1_port, SHIFT_3_0_port, SHIFT_2_35_port, 
      SHIFT_2_34_port, SHIFT_2_33_port, SHIFT_2_32_port, SHIFT_2_31_port, 
      SHIFT_2_30_port, SHIFT_2_29_port, SHIFT_2_28_port, SHIFT_2_27_port, 
      SHIFT_2_26_port, SHIFT_2_25_port, SHIFT_2_24_port, SHIFT_2_23_port, 
      SHIFT_2_22_port, SHIFT_2_21_port, SHIFT_2_20_port, SHIFT_2_19_port, 
      SHIFT_2_18_port, SHIFT_2_17_port, SHIFT_2_16_port, SHIFT_2_15_port, 
      SHIFT_2_14_port, SHIFT_2_13_port, SHIFT_2_12_port, SHIFT_2_11_port, 
      SHIFT_2_10_port, SHIFT_2_9_port, SHIFT_2_8_port, SHIFT_2_7_port, 
      SHIFT_2_6_port, SHIFT_2_5_port, SHIFT_2_4_port, SHIFT_2_3_port, 
      SHIFT_2_2_port, SHIFT_2_1_port, SHIFT_2_0_port, SHIFT_1_33_port, 
      SHIFT_1_32_port, SHIFT_n_1_31_port, SHIFT_n_1_30_port, SHIFT_n_1_29_port,
      SHIFT_n_1_28_port, SHIFT_n_1_27_port, SHIFT_n_1_26_port, 
      SHIFT_n_1_25_port, SHIFT_n_1_24_port, SHIFT_n_1_23_port, 
      SHIFT_n_1_22_port, SHIFT_n_1_21_port, SHIFT_n_1_20_port, 
      SHIFT_n_1_19_port, SHIFT_n_1_18_port, SHIFT_n_1_17_port, 
      SHIFT_n_1_16_port, SHIFT_n_1_15_port, SHIFT_n_1_14_port, 
      SHIFT_n_1_13_port, SHIFT_n_1_12_port, SHIFT_n_1_11_port, 
      SHIFT_n_1_10_port, SHIFT_n_1_9_port, SHIFT_n_1_8_port, SHIFT_n_1_7_port, 
      SHIFT_n_1_6_port, SHIFT_n_1_5_port, SHIFT_n_1_4_port, SHIFT_n_1_3_port, 
      SHIFT_n_1_2_port, SHIFT_n_1_1_port, SHIFT_n_1_0_port, SHIFT_n_15_61_port,
      SHIFT_n_15_60_port, SHIFT_n_15_59_port, SHIFT_n_15_58_port, 
      SHIFT_n_15_57_port, SHIFT_n_15_56_port, SHIFT_n_15_55_port, 
      SHIFT_n_15_54_port, SHIFT_n_15_53_port, SHIFT_n_15_52_port, 
      SHIFT_n_15_51_port, SHIFT_n_15_50_port, SHIFT_n_15_49_port, 
      SHIFT_n_15_48_port, SHIFT_n_15_47_port, SHIFT_n_15_46_port, 
      SHIFT_n_15_45_port, SHIFT_n_15_44_port, SHIFT_n_15_43_port, 
      SHIFT_n_15_42_port, SHIFT_n_15_41_port, SHIFT_n_15_40_port, 
      SHIFT_n_15_39_port, SHIFT_n_15_38_port, SHIFT_n_15_37_port, 
      SHIFT_n_15_36_port, SHIFT_n_15_35_port, SHIFT_n_15_34_port, 
      SHIFT_n_15_33_port, SHIFT_n_15_32_port, SHIFT_n_15_31_port, 
      SHIFT_n_15_30_port, SHIFT_n_15_29_port, SHIFT_n_15_28_port, 
      SHIFT_n_15_27_port, SHIFT_n_15_26_port, SHIFT_n_15_25_port, 
      SHIFT_n_15_24_port, SHIFT_n_15_23_port, SHIFT_n_15_22_port, 
      SHIFT_n_15_21_port, SHIFT_n_15_20_port, SHIFT_n_15_19_port, 
      SHIFT_n_15_18_port, SHIFT_n_15_17_port, SHIFT_n_15_16_port, 
      SHIFT_n_15_15_port, SHIFT_n_15_14_port, SHIFT_n_15_13_port, 
      SHIFT_n_15_12_port, SHIFT_n_15_11_port, SHIFT_n_15_10_port, 
      SHIFT_n_15_9_port, SHIFT_n_15_8_port, SHIFT_n_15_7_port, 
      SHIFT_n_15_6_port, SHIFT_n_15_5_port, SHIFT_n_15_4_port, 
      SHIFT_n_15_3_port, SHIFT_n_15_2_port, SHIFT_n_15_1_port, 
      SHIFT_n_15_0_port, SHIFT_n_14_59_port, SHIFT_n_14_58_port, 
      SHIFT_n_14_57_port, SHIFT_n_14_56_port, SHIFT_n_14_55_port, 
      SHIFT_n_14_54_port, SHIFT_n_14_53_port, SHIFT_n_14_52_port, 
      SHIFT_n_14_51_port, SHIFT_n_14_50_port, SHIFT_n_14_49_port, 
      SHIFT_n_14_48_port, SHIFT_n_14_47_port, SHIFT_n_14_46_port, 
      SHIFT_n_14_45_port, SHIFT_n_14_44_port, SHIFT_n_14_43_port, 
      SHIFT_n_14_42_port, SHIFT_n_14_41_port, SHIFT_n_14_40_port, 
      SHIFT_n_14_39_port, SHIFT_n_14_38_port, SHIFT_n_14_37_port, 
      SHIFT_n_14_36_port, SHIFT_n_14_35_port, SHIFT_n_14_34_port, 
      SHIFT_n_14_33_port, SHIFT_n_14_32_port, SHIFT_n_14_31_port, 
      SHIFT_n_14_30_port, SHIFT_n_14_29_port, SHIFT_n_14_28_port, 
      SHIFT_n_14_27_port, SHIFT_n_14_26_port, SHIFT_n_14_25_port, 
      SHIFT_n_14_24_port, SHIFT_n_14_23_port, SHIFT_n_14_22_port, 
      SHIFT_n_14_21_port, SHIFT_n_14_20_port, SHIFT_n_14_19_port, 
      SHIFT_n_14_18_port, SHIFT_n_14_17_port, SHIFT_n_14_16_port, 
      SHIFT_n_14_15_port, SHIFT_n_14_14_port, SHIFT_n_14_13_port, 
      SHIFT_n_14_12_port, SHIFT_n_14_11_port, SHIFT_n_14_10_port, 
      SHIFT_n_14_9_port, SHIFT_n_14_8_port, SHIFT_n_14_7_port, 
      SHIFT_n_14_6_port, SHIFT_n_14_5_port, SHIFT_n_14_4_port, 
      SHIFT_n_14_3_port, SHIFT_n_14_2_port, SHIFT_n_14_1_port, 
      SHIFT_n_14_0_port, SHIFT_n_13_57_port, SHIFT_n_13_56_port, 
      SHIFT_n_13_55_port, SHIFT_n_13_54_port, SHIFT_n_13_53_port, 
      SHIFT_n_13_52_port, SHIFT_n_13_51_port, SHIFT_n_13_50_port, 
      SHIFT_n_13_49_port, SHIFT_n_13_48_port, SHIFT_n_13_47_port, 
      SHIFT_n_13_46_port, SHIFT_n_13_45_port, SHIFT_n_13_44_port, 
      SHIFT_n_13_43_port, SHIFT_n_13_42_port, SHIFT_n_13_41_port, 
      SHIFT_n_13_40_port, SHIFT_n_13_39_port, SHIFT_n_13_38_port, 
      SHIFT_n_13_37_port, SHIFT_n_13_36_port, SHIFT_n_13_35_port, 
      SHIFT_n_13_34_port, SHIFT_n_13_33_port, SHIFT_n_13_32_port, 
      SHIFT_n_13_31_port, SHIFT_n_13_30_port, SHIFT_n_13_29_port, 
      SHIFT_n_13_28_port, SHIFT_n_13_27_port, SHIFT_n_13_26_port, 
      SHIFT_n_13_25_port, SHIFT_n_13_24_port, SHIFT_n_13_23_port, 
      SHIFT_n_13_22_port, SHIFT_n_13_21_port, SHIFT_n_13_20_port, 
      SHIFT_n_13_19_port, SHIFT_n_13_18_port, SHIFT_n_13_17_port, 
      SHIFT_n_13_16_port, SHIFT_n_13_15_port, SHIFT_n_13_14_port, 
      SHIFT_n_13_13_port, SHIFT_n_13_12_port, SHIFT_n_13_11_port, 
      SHIFT_n_13_10_port, SHIFT_n_13_9_port, SHIFT_n_13_8_port, 
      SHIFT_n_13_7_port, SHIFT_n_13_6_port, SHIFT_n_13_5_port, 
      SHIFT_n_13_4_port, SHIFT_n_13_3_port, SHIFT_n_13_2_port, 
      SHIFT_n_13_1_port, SHIFT_n_13_0_port, SHIFT_n_12_55_port, 
      SHIFT_n_12_54_port, SHIFT_n_12_53_port, SHIFT_n_12_52_port, 
      SHIFT_n_12_51_port, SHIFT_n_12_50_port, SHIFT_n_12_49_port, 
      SHIFT_n_12_48_port, SHIFT_n_12_47_port, SHIFT_n_12_46_port, 
      SHIFT_n_12_45_port, SHIFT_n_12_44_port, SHIFT_n_12_43_port, 
      SHIFT_n_12_42_port, SHIFT_n_12_41_port, SHIFT_n_12_40_port, 
      SHIFT_n_12_39_port, SHIFT_n_12_38_port, SHIFT_n_12_37_port, 
      SHIFT_n_12_36_port, SHIFT_n_12_35_port, SHIFT_n_12_34_port, 
      SHIFT_n_12_33_port, SHIFT_n_12_32_port, SHIFT_n_12_31_port, 
      SHIFT_n_12_30_port, SHIFT_n_12_29_port, SHIFT_n_12_28_port, 
      SHIFT_n_12_27_port, SHIFT_n_12_26_port, SHIFT_n_12_25_port, 
      SHIFT_n_12_24_port, SHIFT_n_12_23_port, SHIFT_n_12_22_port, 
      SHIFT_n_12_21_port, SHIFT_n_12_20_port, SHIFT_n_12_19_port, 
      SHIFT_n_12_18_port, SHIFT_n_12_17_port, SHIFT_n_12_16_port, 
      SHIFT_n_12_15_port, SHIFT_n_12_14_port, SHIFT_n_12_13_port, 
      SHIFT_n_12_12_port, SHIFT_n_12_11_port, SHIFT_n_12_10_port, 
      SHIFT_n_12_9_port, SHIFT_n_12_8_port, SHIFT_n_12_7_port, 
      SHIFT_n_12_6_port, SHIFT_n_12_5_port, SHIFT_n_12_4_port, 
      SHIFT_n_12_3_port, SHIFT_n_12_2_port, SHIFT_n_12_1_port, 
      SHIFT_n_12_0_port, SHIFT_n_11_53_port, SHIFT_n_11_52_port, 
      SHIFT_n_11_51_port, SHIFT_n_11_50_port, SHIFT_n_11_49_port, 
      SHIFT_n_11_48_port, SHIFT_n_11_47_port, SHIFT_n_11_46_port, 
      SHIFT_n_11_45_port, SHIFT_n_11_44_port, SHIFT_n_11_43_port, 
      SHIFT_n_11_42_port, SHIFT_n_11_41_port, SHIFT_n_11_40_port, 
      SHIFT_n_11_39_port, SHIFT_n_11_38_port, SHIFT_n_11_37_port, 
      SHIFT_n_11_36_port, SHIFT_n_11_35_port, SHIFT_n_11_34_port, 
      SHIFT_n_11_33_port, SHIFT_n_11_32_port, SHIFT_n_11_31_port, 
      SHIFT_n_11_30_port, SHIFT_n_11_29_port, SHIFT_n_11_28_port, 
      SHIFT_n_11_27_port, SHIFT_n_11_26_port, SHIFT_n_11_25_port, 
      SHIFT_n_11_24_port, SHIFT_n_11_23_port, SHIFT_n_11_22_port, 
      SHIFT_n_11_21_port, SHIFT_n_11_20_port, SHIFT_n_11_19_port, 
      SHIFT_n_11_18_port, SHIFT_n_11_17_port, SHIFT_n_11_16_port, 
      SHIFT_n_11_15_port, SHIFT_n_11_14_port, SHIFT_n_11_13_port, 
      SHIFT_n_11_12_port, SHIFT_n_11_11_port, SHIFT_n_11_10_port, 
      SHIFT_n_11_9_port, SHIFT_n_11_8_port, SHIFT_n_11_7_port, 
      SHIFT_n_11_6_port, SHIFT_n_11_5_port, SHIFT_n_11_4_port, 
      SHIFT_n_11_3_port, SHIFT_n_11_2_port, SHIFT_n_11_1_port, 
      SHIFT_n_11_0_port, SHIFT_n_10_51_port, SHIFT_n_10_50_port, 
      SHIFT_n_10_49_port, SHIFT_n_10_48_port, SHIFT_n_10_47_port, 
      SHIFT_n_10_46_port, SHIFT_n_10_45_port, SHIFT_n_10_44_port, 
      SHIFT_n_10_43_port, SHIFT_n_10_42_port, SHIFT_n_10_41_port, 
      SHIFT_n_10_40_port, SHIFT_n_10_39_port, SHIFT_n_10_38_port, 
      SHIFT_n_10_37_port, SHIFT_n_10_36_port, SHIFT_n_10_35_port, 
      SHIFT_n_10_34_port, SHIFT_n_10_33_port, SHIFT_n_10_32_port, 
      SHIFT_n_10_31_port, SHIFT_n_10_30_port, SHIFT_n_10_29_port, 
      SHIFT_n_10_28_port, SHIFT_n_10_27_port, SHIFT_n_10_26_port, 
      SHIFT_n_10_25_port, SHIFT_n_10_24_port, SHIFT_n_10_23_port, 
      SHIFT_n_10_22_port, SHIFT_n_10_21_port, SHIFT_n_10_20_port, 
      SHIFT_n_10_19_port, SHIFT_n_10_18_port, SHIFT_n_10_17_port, 
      SHIFT_n_10_16_port, SHIFT_n_10_15_port, SHIFT_n_10_14_port, 
      SHIFT_n_10_13_port, SHIFT_n_10_12_port, SHIFT_n_10_11_port, 
      SHIFT_n_10_10_port, SHIFT_n_10_9_port, SHIFT_n_10_8_port, 
      SHIFT_n_10_7_port, SHIFT_n_10_6_port, SHIFT_n_10_5_port, 
      SHIFT_n_10_4_port, SHIFT_n_10_3_port, SHIFT_n_10_2_port, 
      SHIFT_n_10_1_port, SHIFT_n_10_0_port, SHIFT_n_9_49_port, 
      SHIFT_n_9_48_port, SHIFT_n_9_47_port, SHIFT_n_9_46_port, 
      SHIFT_n_9_45_port, SHIFT_n_9_44_port, SHIFT_n_9_43_port, 
      SHIFT_n_9_42_port, SHIFT_n_9_41_port, SHIFT_n_9_40_port, 
      SHIFT_n_9_39_port, SHIFT_n_9_38_port, SHIFT_n_9_37_port, 
      SHIFT_n_9_36_port, SHIFT_n_9_35_port, SHIFT_n_9_34_port, 
      SHIFT_n_9_33_port, SHIFT_n_9_32_port, SHIFT_n_9_31_port, 
      SHIFT_n_9_30_port, SHIFT_n_9_29_port, SHIFT_n_9_28_port, 
      SHIFT_n_9_27_port, SHIFT_n_9_26_port, SHIFT_n_9_25_port, 
      SHIFT_n_9_24_port, SHIFT_n_9_23_port, SHIFT_n_9_22_port, 
      SHIFT_n_9_21_port, SHIFT_n_9_20_port, SHIFT_n_9_19_port, 
      SHIFT_n_9_18_port, SHIFT_n_9_17_port, SHIFT_n_9_16_port, 
      SHIFT_n_9_15_port, SHIFT_n_9_14_port, SHIFT_n_9_13_port, 
      SHIFT_n_9_12_port, SHIFT_n_9_11_port, SHIFT_n_9_10_port, SHIFT_n_9_9_port
      , SHIFT_n_9_8_port, SHIFT_n_9_7_port, SHIFT_n_9_6_port, SHIFT_n_9_5_port,
      SHIFT_n_9_4_port, SHIFT_n_9_3_port, SHIFT_n_9_2_port, SHIFT_n_9_1_port, 
      SHIFT_n_9_0_port, SHIFT_n_8_47_port, SHIFT_n_8_46_port, SHIFT_n_8_45_port
      , SHIFT_n_8_44_port, SHIFT_n_8_43_port, SHIFT_n_8_42_port, 
      SHIFT_n_8_41_port, SHIFT_n_8_40_port, SHIFT_n_8_39_port, 
      SHIFT_n_8_38_port, SHIFT_n_8_37_port, SHIFT_n_8_36_port, 
      SHIFT_n_8_35_port, SHIFT_n_8_34_port, SHIFT_n_8_33_port, 
      SHIFT_n_8_32_port, SHIFT_n_8_31_port, SHIFT_n_8_30_port, 
      SHIFT_n_8_29_port, SHIFT_n_8_28_port, SHIFT_n_8_27_port, 
      SHIFT_n_8_26_port, SHIFT_n_8_25_port, SHIFT_n_8_24_port, 
      SHIFT_n_8_23_port, SHIFT_n_8_22_port, SHIFT_n_8_21_port, 
      SHIFT_n_8_20_port, SHIFT_n_8_19_port, SHIFT_n_8_18_port, 
      SHIFT_n_8_17_port, SHIFT_n_8_16_port, SHIFT_n_8_15_port, 
      SHIFT_n_8_14_port, SHIFT_n_8_13_port, SHIFT_n_8_12_port, 
      SHIFT_n_8_11_port, SHIFT_n_8_10_port, SHIFT_n_8_9_port, SHIFT_n_8_8_port,
      SHIFT_n_8_7_port, SHIFT_n_8_6_port, SHIFT_n_8_5_port, SHIFT_n_8_4_port, 
      SHIFT_n_8_3_port, SHIFT_n_8_2_port, SHIFT_n_8_1_port, SHIFT_n_8_0_port, 
      SHIFT_n_7_45_port, SHIFT_n_7_44_port, SHIFT_n_7_43_port, 
      SHIFT_n_7_42_port, SHIFT_n_7_41_port, SHIFT_n_7_40_port, 
      SHIFT_n_7_39_port, SHIFT_n_7_38_port, SHIFT_n_7_37_port, 
      SHIFT_n_7_36_port, SHIFT_n_7_35_port, SHIFT_n_7_34_port, 
      SHIFT_n_7_33_port, SHIFT_n_7_32_port, SHIFT_n_7_31_port, 
      SHIFT_n_7_30_port, SHIFT_n_7_29_port, SHIFT_n_7_28_port, 
      SHIFT_n_7_27_port, SHIFT_n_7_26_port, SHIFT_n_7_25_port, 
      SHIFT_n_7_24_port, SHIFT_n_7_23_port, SHIFT_n_7_22_port, 
      SHIFT_n_7_21_port, SHIFT_n_7_20_port, SHIFT_n_7_19_port, 
      SHIFT_n_7_18_port, SHIFT_n_7_17_port, SHIFT_n_7_16_port, 
      SHIFT_n_7_15_port, SHIFT_n_7_14_port, SHIFT_n_7_13_port, 
      SHIFT_n_7_12_port, SHIFT_n_7_11_port, SHIFT_n_7_10_port, SHIFT_n_7_9_port
      , SHIFT_n_7_8_port, SHIFT_n_7_7_port, SHIFT_n_7_6_port, SHIFT_n_7_5_port,
      SHIFT_n_7_4_port, SHIFT_n_7_3_port, SHIFT_n_7_2_port, SHIFT_n_7_1_port, 
      SHIFT_n_7_0_port, SHIFT_n_6_43_port, SHIFT_n_6_42_port, SHIFT_n_6_41_port
      , SHIFT_n_6_40_port, SHIFT_n_6_39_port, SHIFT_n_6_38_port, 
      SHIFT_n_6_37_port, SHIFT_n_6_36_port, SHIFT_n_6_35_port, 
      SHIFT_n_6_34_port, SHIFT_n_6_33_port, SHIFT_n_6_32_port, 
      SHIFT_n_6_31_port, SHIFT_n_6_30_port, SHIFT_n_6_29_port, 
      SHIFT_n_6_28_port, SHIFT_n_6_27_port, SHIFT_n_6_26_port, 
      SHIFT_n_6_25_port, SHIFT_n_6_24_port, SHIFT_n_6_23_port, 
      SHIFT_n_6_22_port, SHIFT_n_6_21_port, SHIFT_n_6_20_port, 
      SHIFT_n_6_19_port, SHIFT_n_6_18_port, SHIFT_n_6_17_port, 
      SHIFT_n_6_16_port, SHIFT_n_6_15_port, SHIFT_n_6_14_port, 
      SHIFT_n_6_13_port, SHIFT_n_6_12_port, SHIFT_n_6_11_port, 
      SHIFT_n_6_10_port, SHIFT_n_6_9_port, SHIFT_n_6_8_port, SHIFT_n_6_7_port, 
      SHIFT_n_6_6_port, SHIFT_n_6_5_port, SHIFT_n_6_4_port, SHIFT_n_6_3_port, 
      SHIFT_n_6_2_port, SHIFT_n_6_1_port, SHIFT_n_6_0_port, SHIFT_n_5_41_port, 
      SHIFT_n_5_40_port, SHIFT_n_5_39_port, SHIFT_n_5_38_port, 
      SHIFT_n_5_37_port, SHIFT_n_5_36_port, SHIFT_n_5_35_port, 
      SHIFT_n_5_34_port, SHIFT_n_5_33_port, SHIFT_n_5_32_port, 
      SHIFT_n_5_31_port, SHIFT_n_5_30_port, SHIFT_n_5_29_port, 
      SHIFT_n_5_28_port, SHIFT_n_5_27_port, SHIFT_n_5_26_port, 
      SHIFT_n_5_25_port, SHIFT_n_5_24_port, SHIFT_n_5_23_port, 
      SHIFT_n_5_22_port, SHIFT_n_5_21_port, SHIFT_n_5_20_port, 
      SHIFT_n_5_19_port, SHIFT_n_5_18_port, SHIFT_n_5_17_port, 
      SHIFT_n_5_16_port, SHIFT_n_5_15_port, SHIFT_n_5_14_port, 
      SHIFT_n_5_13_port, SHIFT_n_5_12_port, SHIFT_n_5_11_port, 
      SHIFT_n_5_10_port, SHIFT_n_5_9_port, SHIFT_n_5_8_port, SHIFT_n_5_7_port, 
      SHIFT_n_5_6_port, SHIFT_n_5_5_port, SHIFT_n_5_4_port, SHIFT_n_5_3_port, 
      SHIFT_n_5_2_port, SHIFT_n_5_1_port, SHIFT_n_5_0_port, SHIFT_n_4_39_port, 
      SHIFT_n_4_38_port, SHIFT_n_4_37_port, SHIFT_n_4_36_port, 
      SHIFT_n_4_35_port, SHIFT_n_4_34_port, SHIFT_n_4_33_port, 
      SHIFT_n_4_32_port, SHIFT_n_4_31_port, SHIFT_n_4_30_port, 
      SHIFT_n_4_29_port, SHIFT_n_4_28_port, SHIFT_n_4_27_port, 
      SHIFT_n_4_26_port, SHIFT_n_4_25_port, SHIFT_n_4_24_port, 
      SHIFT_n_4_23_port, SHIFT_n_4_22_port, SHIFT_n_4_21_port, 
      SHIFT_n_4_20_port, SHIFT_n_4_19_port, SHIFT_n_4_18_port, 
      SHIFT_n_4_17_port, SHIFT_n_4_16_port, SHIFT_n_4_15_port, 
      SHIFT_n_4_14_port, SHIFT_n_4_13_port, SHIFT_n_4_12_port, 
      SHIFT_n_4_11_port, SHIFT_n_4_10_port, SHIFT_n_4_9_port, SHIFT_n_4_8_port,
      SHIFT_n_4_7_port, SHIFT_n_4_6_port, SHIFT_n_4_5_port, SHIFT_n_4_4_port, 
      SHIFT_n_4_3_port, SHIFT_n_4_2_port, SHIFT_n_4_1_port, SHIFT_n_4_0_port, 
      SHIFT_n_3_37_port, SHIFT_n_3_36_port, SHIFT_n_3_35_port, 
      SHIFT_n_3_34_port, SHIFT_n_3_33_port, SHIFT_n_3_32_port, 
      SHIFT_n_3_31_port, SHIFT_n_3_30_port, SHIFT_n_3_29_port, 
      SHIFT_n_3_28_port, SHIFT_n_3_27_port, SHIFT_n_3_26_port, 
      SHIFT_n_3_25_port, SHIFT_n_3_24_port, SHIFT_n_3_23_port, 
      SHIFT_n_3_22_port, SHIFT_n_3_21_port, SHIFT_n_3_20_port, 
      SHIFT_n_3_19_port, SHIFT_n_3_18_port, SHIFT_n_3_17_port, 
      SHIFT_n_3_16_port, SHIFT_n_3_15_port, SHIFT_n_3_14_port, 
      SHIFT_n_3_13_port, SHIFT_n_3_12_port, SHIFT_n_3_11_port, 
      SHIFT_n_3_10_port, SHIFT_n_3_9_port, SHIFT_n_3_8_port, SHIFT_n_3_7_port, 
      SHIFT_n_3_6_port, SHIFT_n_3_5_port, SHIFT_n_3_4_port, SHIFT_n_3_3_port, 
      SHIFT_n_3_2_port, SHIFT_n_3_1_port, SHIFT_n_3_0_port, SHIFT_n_2_35_port, 
      SHIFT_n_2_34_port, SHIFT_n_2_33_port, SHIFT_n_2_32_port, 
      SHIFT_n_2_31_port, SHIFT_n_2_30_port, SHIFT_n_2_29_port, 
      SHIFT_n_2_28_port, SHIFT_n_2_27_port, SHIFT_n_2_26_port, 
      SHIFT_n_2_25_port, SHIFT_n_2_24_port, SHIFT_n_2_23_port, 
      SHIFT_n_2_22_port, SHIFT_n_2_21_port, SHIFT_n_2_20_port, 
      SHIFT_n_2_19_port, SHIFT_n_2_18_port, SHIFT_n_2_17_port, 
      SHIFT_n_2_16_port, SHIFT_n_2_15_port, SHIFT_n_2_14_port, 
      SHIFT_n_2_13_port, SHIFT_n_2_12_port, SHIFT_n_2_11_port, 
      SHIFT_n_2_10_port, SHIFT_n_2_9_port, SHIFT_n_2_8_port, SHIFT_n_2_7_port, 
      SHIFT_n_2_6_port, SHIFT_n_2_5_port, SHIFT_n_2_4_port, SHIFT_n_2_3_port, 
      SHIFT_n_2_2_port, SHIFT_n_2_1_port, SHIFT_n_2_0_port, SHIFT_n_1_33_port, 
      SHIFT_n_1_32_port, OTMP_8_15_port, OTMP_8_14_port, OTMP_8_13_port, 
      OTMP_8_12_port, OTMP_8_11_port, OTMP_8_10_port, OTMP_8_9_port, 
      OTMP_8_8_port, OTMP_8_7_port, OTMP_8_6_port, OTMP_8_5_port, OTMP_8_4_port
      , OTMP_8_3_port, OTMP_8_2_port, OTMP_8_1_port, OTMP_8_0_port, 
      OTMP_7_47_port, OTMP_7_46_port, OTMP_7_45_port, OTMP_7_44_port, 
      OTMP_7_43_port, OTMP_7_42_port, OTMP_7_41_port, OTMP_7_40_port, 
      OTMP_7_39_port, OTMP_7_38_port, OTMP_7_37_port, OTMP_7_36_port, 
      OTMP_7_35_port, OTMP_7_34_port, OTMP_7_33_port, OTMP_7_32_port, 
      OTMP_7_31_port, OTMP_7_30_port, OTMP_7_29_port, OTMP_7_28_port, 
      OTMP_7_27_port, OTMP_7_26_port, OTMP_7_25_port, OTMP_7_24_port, 
      OTMP_7_23_port, OTMP_7_22_port, OTMP_7_21_port, OTMP_7_20_port, 
      OTMP_7_19_port, OTMP_7_18_port, OTMP_7_17_port, OTMP_7_16_port, 
      OTMP_7_15_port, OTMP_7_14_port, OTMP_7_13_port, OTMP_7_12_port, 
      OTMP_7_11_port, OTMP_7_10_port, OTMP_7_9_port, OTMP_7_8_port, 
      OTMP_7_7_port, OTMP_7_6_port, OTMP_7_5_port, OTMP_7_4_port, OTMP_7_3_port
      , OTMP_7_2_port, OTMP_7_1_port, OTMP_7_0_port, OTMP_6_45_port, 
      OTMP_6_44_port, OTMP_6_43_port, OTMP_6_42_port, OTMP_6_41_port, 
      OTMP_6_40_port, OTMP_6_39_port, OTMP_6_38_port, OTMP_6_37_port, 
      OTMP_6_36_port, OTMP_6_35_port, OTMP_6_34_port, OTMP_6_33_port, 
      OTMP_6_32_port, OTMP_6_31_port, OTMP_6_30_port, OTMP_6_29_port, 
      OTMP_6_28_port, OTMP_6_27_port, OTMP_6_26_port, OTMP_6_25_port, 
      OTMP_6_24_port, OTMP_6_23_port, OTMP_6_22_port, OTMP_6_21_port, 
      OTMP_6_20_port, OTMP_6_19_port, OTMP_6_18_port, OTMP_6_17_port, 
      OTMP_6_16_port, OTMP_6_15_port, OTMP_6_14_port, OTMP_6_13_port, 
      OTMP_6_12_port, OTMP_6_11_port, OTMP_6_10_port, OTMP_6_9_port, 
      OTMP_6_8_port, OTMP_6_7_port, OTMP_6_6_port, OTMP_6_5_port, OTMP_6_4_port
      , OTMP_6_3_port, OTMP_6_2_port, OTMP_6_1_port, OTMP_6_0_port, 
      OTMP_5_43_port, OTMP_5_42_port, OTMP_5_41_port, OTMP_5_40_port, 
      OTMP_5_39_port, OTMP_5_38_port, OTMP_5_37_port, OTMP_5_36_port, 
      OTMP_5_35_port, OTMP_5_34_port, OTMP_5_33_port, OTMP_5_32_port, 
      OTMP_5_31_port, OTMP_5_30_port, OTMP_5_29_port, OTMP_5_28_port, 
      OTMP_5_27_port, OTMP_5_26_port, OTMP_5_25_port, OTMP_5_24_port, 
      OTMP_5_23_port, OTMP_5_22_port, OTMP_5_21_port, OTMP_5_20_port, 
      OTMP_5_19_port, OTMP_5_18_port, OTMP_5_17_port, OTMP_5_16_port, 
      OTMP_5_15_port, OTMP_5_14_port, OTMP_5_13_port, OTMP_5_12_port, 
      OTMP_5_11_port, OTMP_5_10_port, OTMP_5_9_port, OTMP_5_8_port, 
      OTMP_5_7_port, OTMP_5_6_port, OTMP_5_5_port, OTMP_5_4_port, OTMP_5_3_port
      , OTMP_5_2_port, OTMP_5_1_port, OTMP_5_0_port, OTMP_4_41_port, 
      OTMP_4_40_port, OTMP_4_39_port, OTMP_4_38_port, OTMP_4_37_port, 
      OTMP_4_36_port, OTMP_4_35_port, OTMP_4_34_port, OTMP_4_33_port, 
      OTMP_4_32_port, OTMP_4_31_port, OTMP_4_30_port, OTMP_4_29_port, 
      OTMP_4_28_port, OTMP_4_27_port, OTMP_4_26_port, OTMP_4_25_port, 
      OTMP_4_24_port, OTMP_4_23_port, OTMP_4_22_port, OTMP_4_21_port, 
      OTMP_4_20_port, OTMP_4_19_port, OTMP_4_18_port, OTMP_4_17_port, 
      OTMP_4_16_port, OTMP_4_15_port, OTMP_4_14_port, OTMP_4_13_port, 
      OTMP_4_12_port, OTMP_4_11_port, OTMP_4_10_port, OTMP_4_9_port, 
      OTMP_4_8_port, OTMP_4_7_port, OTMP_4_6_port, OTMP_4_5_port, OTMP_4_4_port
      , OTMP_4_3_port, OTMP_4_2_port, OTMP_4_1_port, OTMP_4_0_port, 
      OTMP_3_39_port, OTMP_3_38_port, OTMP_3_37_port, OTMP_3_36_port, 
      OTMP_3_35_port, OTMP_3_34_port, OTMP_3_33_port, OTMP_3_32_port, 
      OTMP_3_31_port, OTMP_3_30_port, OTMP_3_29_port, OTMP_3_28_port, 
      OTMP_3_27_port, OTMP_3_26_port, OTMP_3_25_port, OTMP_3_24_port, 
      OTMP_3_23_port, OTMP_3_22_port, OTMP_3_21_port, OTMP_3_20_port, 
      OTMP_3_19_port, OTMP_3_18_port, OTMP_3_17_port, OTMP_3_16_port, 
      OTMP_3_15_port, OTMP_3_14_port, OTMP_3_13_port, OTMP_3_12_port, 
      OTMP_3_11_port, OTMP_3_10_port, OTMP_3_9_port, OTMP_3_8_port, 
      OTMP_3_7_port, OTMP_3_6_port, OTMP_3_5_port, OTMP_3_4_port, OTMP_3_3_port
      , OTMP_3_2_port, OTMP_3_1_port, OTMP_3_0_port, OTMP_2_37_port, 
      OTMP_2_36_port, OTMP_2_35_port, OTMP_2_34_port, OTMP_2_33_port, 
      OTMP_2_32_port, OTMP_2_31_port, OTMP_2_30_port, OTMP_2_29_port, 
      OTMP_2_28_port, OTMP_2_27_port, OTMP_2_26_port, OTMP_2_25_port, 
      OTMP_2_24_port, OTMP_2_23_port, OTMP_2_22_port, OTMP_2_21_port, 
      OTMP_2_20_port, OTMP_2_19_port, OTMP_2_18_port, OTMP_2_17_port, 
      OTMP_2_16_port, OTMP_2_15_port, OTMP_2_14_port, OTMP_2_13_port, 
      OTMP_2_12_port, OTMP_2_11_port, OTMP_2_10_port, OTMP_2_9_port, 
      OTMP_2_8_port, OTMP_2_7_port, OTMP_2_6_port, OTMP_2_5_port, OTMP_2_4_port
      , OTMP_2_3_port, OTMP_2_2_port, OTMP_2_1_port, OTMP_2_0_port, 
      OTMP_1_35_port, OTMP_1_34_port, OTMP_1_33_port, OTMP_1_32_port, 
      OTMP_1_31_port, OTMP_1_30_port, OTMP_1_29_port, OTMP_1_28_port, 
      OTMP_1_27_port, OTMP_1_26_port, OTMP_1_25_port, OTMP_1_24_port, 
      OTMP_1_23_port, OTMP_1_22_port, OTMP_1_21_port, OTMP_1_20_port, 
      OTMP_1_19_port, OTMP_1_18_port, OTMP_1_17_port, OTMP_1_16_port, 
      OTMP_1_15_port, OTMP_1_14_port, OTMP_1_13_port, OTMP_1_12_port, 
      OTMP_1_11_port, OTMP_1_10_port, OTMP_1_9_port, OTMP_1_8_port, 
      OTMP_1_7_port, OTMP_1_6_port, OTMP_1_5_port, OTMP_1_4_port, OTMP_1_3_port
      , OTMP_1_2_port, OTMP_1_1_port, OTMP_1_0_port, OTMP_0_34_port, 
      OTMP_0_32_port, OTMP_0_31_port, OTMP_0_30_port, OTMP_0_29_port, 
      OTMP_0_28_port, OTMP_0_27_port, OTMP_0_26_port, OTMP_0_25_port, 
      OTMP_0_24_port, OTMP_0_23_port, OTMP_0_22_port, OTMP_0_21_port, 
      OTMP_0_20_port, OTMP_0_19_port, OTMP_0_18_port, OTMP_0_17_port, 
      OTMP_0_16_port, OTMP_0_15_port, OTMP_0_14_port, OTMP_0_13_port, 
      OTMP_0_12_port, OTMP_0_11_port, OTMP_0_10_port, OTMP_0_9_port, 
      OTMP_0_8_port, OTMP_0_7_port, OTMP_0_6_port, OTMP_0_5_port, OTMP_0_4_port
      , OTMP_0_3_port, OTMP_0_2_port, OTMP_0_1_port, OTMP_0_0_port, 
      OTMP_15_63_port, OTMP_15_62_port, OTMP_15_61_port, OTMP_15_60_port, 
      OTMP_15_59_port, OTMP_15_58_port, OTMP_15_57_port, OTMP_15_56_port, 
      OTMP_15_55_port, OTMP_15_54_port, OTMP_15_53_port, OTMP_15_52_port, 
      OTMP_15_51_port, OTMP_15_50_port, OTMP_15_49_port, OTMP_15_48_port, 
      OTMP_15_47_port, OTMP_15_46_port, OTMP_15_45_port, OTMP_15_44_port, 
      OTMP_15_43_port, OTMP_15_42_port, OTMP_15_41_port, OTMP_15_40_port, 
      OTMP_15_39_port, OTMP_15_38_port, OTMP_15_37_port, OTMP_15_36_port, 
      OTMP_15_35_port, OTMP_15_34_port, OTMP_15_33_port, OTMP_15_32_port, 
      OTMP_15_31_port, OTMP_15_30_port, OTMP_15_29_port, OTMP_15_28_port, 
      OTMP_15_27_port, OTMP_15_26_port, OTMP_15_25_port, OTMP_15_24_port, 
      OTMP_15_23_port, OTMP_15_22_port, OTMP_15_21_port, OTMP_15_20_port, 
      OTMP_15_19_port, OTMP_15_18_port, OTMP_15_17_port, OTMP_15_16_port, 
      OTMP_15_15_port, OTMP_15_14_port, OTMP_15_13_port, OTMP_15_12_port, 
      OTMP_15_11_port, OTMP_15_10_port, OTMP_15_9_port, OTMP_15_8_port, 
      OTMP_15_7_port, OTMP_15_6_port, OTMP_15_5_port, OTMP_15_4_port, 
      OTMP_15_3_port, OTMP_15_2_port, OTMP_15_1_port, OTMP_15_0_port, 
      OTMP_14_61_port, OTMP_14_60_port, OTMP_14_59_port, OTMP_14_58_port, 
      OTMP_14_57_port, OTMP_14_56_port, OTMP_14_55_port, OTMP_14_54_port, 
      OTMP_14_53_port, OTMP_14_52_port, OTMP_14_51_port, OTMP_14_50_port, 
      OTMP_14_49_port, OTMP_14_48_port, OTMP_14_47_port, OTMP_14_46_port, 
      OTMP_14_45_port, OTMP_14_44_port, OTMP_14_43_port, OTMP_14_42_port, 
      OTMP_14_41_port, OTMP_14_40_port, OTMP_14_39_port, OTMP_14_38_port, 
      OTMP_14_37_port, OTMP_14_36_port, OTMP_14_35_port, OTMP_14_34_port, 
      OTMP_14_33_port, OTMP_14_32_port, OTMP_14_31_port, OTMP_14_30_port, 
      OTMP_14_29_port, OTMP_14_28_port, OTMP_14_27_port, OTMP_14_26_port, 
      OTMP_14_25_port, OTMP_14_24_port, OTMP_14_23_port, OTMP_14_22_port, 
      OTMP_14_21_port, OTMP_14_20_port, OTMP_14_19_port, OTMP_14_18_port, 
      OTMP_14_17_port, OTMP_14_16_port, OTMP_14_15_port, OTMP_14_14_port, 
      OTMP_14_13_port, OTMP_14_12_port, OTMP_14_11_port, OTMP_14_10_port, 
      OTMP_14_9_port, OTMP_14_8_port, OTMP_14_7_port, OTMP_14_6_port, 
      OTMP_14_5_port, OTMP_14_4_port, OTMP_14_3_port, OTMP_14_2_port, 
      OTMP_14_1_port, OTMP_14_0_port, OTMP_13_59_port, OTMP_13_58_port, 
      OTMP_13_57_port, OTMP_13_56_port, OTMP_13_55_port, OTMP_13_54_port, 
      OTMP_13_53_port, OTMP_13_52_port, OTMP_13_51_port, OTMP_13_50_port, 
      OTMP_13_49_port, OTMP_13_48_port, OTMP_13_47_port, OTMP_13_46_port, 
      OTMP_13_45_port, OTMP_13_44_port, OTMP_13_43_port, OTMP_13_42_port, 
      OTMP_13_41_port, OTMP_13_40_port, OTMP_13_39_port, OTMP_13_38_port, 
      OTMP_13_37_port, OTMP_13_36_port, OTMP_13_35_port, OTMP_13_34_port, 
      OTMP_13_33_port, OTMP_13_32_port, OTMP_13_31_port, OTMP_13_30_port, 
      OTMP_13_29_port, OTMP_13_28_port, OTMP_13_27_port, OTMP_13_26_port, 
      OTMP_13_25_port, OTMP_13_24_port, OTMP_13_23_port, OTMP_13_22_port, 
      OTMP_13_21_port, OTMP_13_20_port, OTMP_13_19_port, OTMP_13_18_port, 
      OTMP_13_17_port, OTMP_13_16_port, OTMP_13_15_port, OTMP_13_14_port, 
      OTMP_13_13_port, OTMP_13_12_port, OTMP_13_11_port, OTMP_13_10_port, 
      OTMP_13_9_port, OTMP_13_8_port, OTMP_13_7_port, OTMP_13_6_port, 
      OTMP_13_5_port, OTMP_13_4_port, OTMP_13_3_port, OTMP_13_2_port, 
      OTMP_13_1_port, OTMP_13_0_port, OTMP_12_57_port, OTMP_12_56_port, 
      OTMP_12_55_port, OTMP_12_54_port, OTMP_12_53_port, OTMP_12_52_port, 
      OTMP_12_51_port, OTMP_12_50_port, OTMP_12_49_port, OTMP_12_48_port, 
      OTMP_12_47_port, OTMP_12_46_port, OTMP_12_45_port, OTMP_12_44_port, 
      OTMP_12_43_port, OTMP_12_42_port, OTMP_12_41_port, OTMP_12_40_port, 
      OTMP_12_39_port, OTMP_12_38_port, OTMP_12_37_port, OTMP_12_36_port, 
      OTMP_12_35_port, OTMP_12_34_port, OTMP_12_33_port, OTMP_12_32_port, 
      OTMP_12_31_port, OTMP_12_30_port, OTMP_12_29_port, OTMP_12_28_port, 
      OTMP_12_27_port, OTMP_12_26_port, OTMP_12_25_port, OTMP_12_24_port, 
      OTMP_12_23_port, OTMP_12_22_port, OTMP_12_21_port, OTMP_12_20_port, 
      OTMP_12_19_port, OTMP_12_18_port, OTMP_12_17_port, OTMP_12_16_port, 
      OTMP_12_15_port, OTMP_12_14_port, OTMP_12_13_port, OTMP_12_12_port, 
      OTMP_12_11_port, OTMP_12_10_port, OTMP_12_9_port, OTMP_12_8_port, 
      OTMP_12_7_port, OTMP_12_6_port, OTMP_12_5_port, OTMP_12_4_port, 
      OTMP_12_3_port, OTMP_12_2_port, OTMP_12_1_port, OTMP_12_0_port, 
      OTMP_11_55_port, OTMP_11_54_port, OTMP_11_53_port, OTMP_11_52_port, 
      OTMP_11_51_port, OTMP_11_50_port, OTMP_11_49_port, OTMP_11_48_port, 
      OTMP_11_47_port, OTMP_11_46_port, OTMP_11_45_port, OTMP_11_44_port, 
      OTMP_11_43_port, OTMP_11_42_port, OTMP_11_41_port, OTMP_11_40_port, 
      OTMP_11_39_port, OTMP_11_38_port, OTMP_11_37_port, OTMP_11_36_port, 
      OTMP_11_35_port, OTMP_11_34_port, OTMP_11_33_port, OTMP_11_32_port, 
      OTMP_11_31_port, OTMP_11_30_port, OTMP_11_29_port, OTMP_11_28_port, 
      OTMP_11_27_port, OTMP_11_26_port, OTMP_11_25_port, OTMP_11_24_port, 
      OTMP_11_23_port, OTMP_11_22_port, OTMP_11_21_port, OTMP_11_20_port, 
      OTMP_11_19_port, OTMP_11_18_port, OTMP_11_17_port, OTMP_11_16_port, 
      OTMP_11_15_port, OTMP_11_14_port, OTMP_11_13_port, OTMP_11_12_port, 
      OTMP_11_11_port, OTMP_11_10_port, OTMP_11_9_port, OTMP_11_8_port, 
      OTMP_11_7_port, OTMP_11_6_port, OTMP_11_5_port, OTMP_11_4_port, 
      OTMP_11_3_port, OTMP_11_2_port, OTMP_11_1_port, OTMP_11_0_port, 
      OTMP_10_53_port, OTMP_10_52_port, OTMP_10_51_port, OTMP_10_50_port, 
      OTMP_10_49_port, OTMP_10_48_port, OTMP_10_47_port, OTMP_10_46_port, 
      OTMP_10_45_port, OTMP_10_44_port, OTMP_10_43_port, OTMP_10_42_port, 
      OTMP_10_41_port, OTMP_10_40_port, OTMP_10_39_port, OTMP_10_38_port, 
      OTMP_10_37_port, OTMP_10_36_port, OTMP_10_35_port, OTMP_10_34_port, 
      OTMP_10_33_port, OTMP_10_32_port, OTMP_10_31_port, OTMP_10_30_port, 
      OTMP_10_29_port, OTMP_10_28_port, OTMP_10_27_port, OTMP_10_26_port, 
      OTMP_10_25_port, OTMP_10_24_port, OTMP_10_23_port, OTMP_10_22_port, 
      OTMP_10_21_port, OTMP_10_20_port, OTMP_10_19_port, OTMP_10_18_port, 
      OTMP_10_17_port, OTMP_10_16_port, OTMP_10_15_port, OTMP_10_14_port, 
      OTMP_10_13_port, OTMP_10_12_port, OTMP_10_11_port, OTMP_10_10_port, 
      OTMP_10_9_port, OTMP_10_8_port, OTMP_10_7_port, OTMP_10_6_port, 
      OTMP_10_5_port, OTMP_10_4_port, OTMP_10_3_port, OTMP_10_2_port, 
      OTMP_10_1_port, OTMP_10_0_port, OTMP_9_51_port, OTMP_9_50_port, 
      OTMP_9_49_port, OTMP_9_48_port, OTMP_9_47_port, OTMP_9_46_port, 
      OTMP_9_45_port, OTMP_9_44_port, OTMP_9_43_port, OTMP_9_42_port, 
      OTMP_9_41_port, OTMP_9_40_port, OTMP_9_39_port, OTMP_9_38_port, 
      OTMP_9_37_port, OTMP_9_36_port, OTMP_9_35_port, OTMP_9_34_port, 
      OTMP_9_33_port, OTMP_9_32_port, OTMP_9_31_port, OTMP_9_30_port, 
      OTMP_9_29_port, OTMP_9_28_port, OTMP_9_27_port, OTMP_9_26_port, 
      OTMP_9_25_port, OTMP_9_24_port, OTMP_9_23_port, OTMP_9_22_port, 
      OTMP_9_21_port, OTMP_9_20_port, OTMP_9_19_port, OTMP_9_18_port, 
      OTMP_9_17_port, OTMP_9_16_port, OTMP_9_15_port, OTMP_9_14_port, 
      OTMP_9_13_port, OTMP_9_12_port, OTMP_9_11_port, OTMP_9_10_port, 
      OTMP_9_9_port, OTMP_9_8_port, OTMP_9_7_port, OTMP_9_6_port, OTMP_9_5_port
      , OTMP_9_4_port, OTMP_9_3_port, OTMP_9_2_port, OTMP_9_1_port, 
      OTMP_9_0_port, OTMP_8_49_port, OTMP_8_48_port, OTMP_8_47_port, 
      OTMP_8_46_port, OTMP_8_45_port, OTMP_8_44_port, OTMP_8_43_port, 
      OTMP_8_42_port, OTMP_8_41_port, OTMP_8_40_port, OTMP_8_39_port, 
      OTMP_8_38_port, OTMP_8_37_port, OTMP_8_36_port, OTMP_8_35_port, 
      OTMP_8_34_port, OTMP_8_33_port, OTMP_8_32_port, OTMP_8_31_port, 
      OTMP_8_30_port, OTMP_8_29_port, OTMP_8_28_port, OTMP_8_27_port, 
      OTMP_8_26_port, OTMP_8_25_port, OTMP_8_24_port, OTMP_8_23_port, 
      OTMP_8_22_port, OTMP_8_21_port, OTMP_8_20_port, OTMP_8_19_port, 
      OTMP_8_18_port, OTMP_8_17_port, OTMP_8_16_port, PTMP_8_15_port, 
      PTMP_8_14_port, PTMP_8_13_port, PTMP_8_12_port, PTMP_8_11_port, 
      PTMP_8_10_port, PTMP_8_9_port, PTMP_8_8_port, PTMP_8_7_port, 
      PTMP_8_6_port, PTMP_8_5_port, PTMP_8_4_port, PTMP_8_3_port, PTMP_8_2_port
      , PTMP_8_1_port, PTMP_8_0_port, PTMP_7_49_port, PTMP_7_48_port, 
      PTMP_7_47_port, PTMP_7_46_port, PTMP_7_45_port, PTMP_7_44_port, 
      PTMP_7_43_port, PTMP_7_42_port, PTMP_7_41_port, PTMP_7_40_port, 
      PTMP_7_39_port, PTMP_7_38_port, PTMP_7_37_port, PTMP_7_36_port, 
      PTMP_7_35_port, PTMP_7_34_port, PTMP_7_33_port, PTMP_7_32_port, 
      PTMP_7_31_port, PTMP_7_30_port, PTMP_7_29_port, PTMP_7_28_port, 
      PTMP_7_27_port, PTMP_7_26_port, PTMP_7_25_port, PTMP_7_24_port, 
      PTMP_7_23_port, PTMP_7_22_port, PTMP_7_21_port, PTMP_7_20_port, 
      PTMP_7_19_port, PTMP_7_18_port, PTMP_7_17_port, PTMP_7_16_port, 
      PTMP_7_15_port, PTMP_7_14_port, PTMP_7_13_port, PTMP_7_12_port, 
      PTMP_7_11_port, PTMP_7_10_port, PTMP_7_9_port, PTMP_7_8_port, 
      PTMP_7_7_port, PTMP_7_6_port, PTMP_7_5_port, PTMP_7_4_port, PTMP_7_3_port
      , PTMP_7_2_port, PTMP_7_1_port, PTMP_7_0_port, PTMP_6_47_port, 
      PTMP_6_46_port, PTMP_6_45_port, PTMP_6_44_port, PTMP_6_43_port, 
      PTMP_6_42_port, PTMP_6_41_port, PTMP_6_40_port, PTMP_6_39_port, 
      PTMP_6_38_port, PTMP_6_37_port, PTMP_6_36_port, PTMP_6_35_port, 
      PTMP_6_34_port, PTMP_6_33_port, PTMP_6_32_port, PTMP_6_31_port, 
      PTMP_6_30_port, PTMP_6_29_port, PTMP_6_28_port, PTMP_6_27_port, 
      PTMP_6_26_port, PTMP_6_25_port, PTMP_6_24_port, PTMP_6_23_port, 
      PTMP_6_22_port, PTMP_6_21_port, PTMP_6_20_port, PTMP_6_19_port, 
      PTMP_6_18_port, PTMP_6_17_port, PTMP_6_16_port, PTMP_6_15_port, 
      PTMP_6_14_port, PTMP_6_13_port, PTMP_6_12_port, PTMP_6_11_port, 
      PTMP_6_10_port, PTMP_6_9_port, PTMP_6_8_port, PTMP_6_7_port, 
      PTMP_6_6_port, PTMP_6_5_port, PTMP_6_4_port, PTMP_6_3_port, PTMP_6_2_port
      , PTMP_6_1_port, PTMP_6_0_port, PTMP_5_45_port, PTMP_5_44_port, 
      PTMP_5_43_port, PTMP_5_42_port, PTMP_5_41_port, PTMP_5_40_port, 
      PTMP_5_39_port, PTMP_5_38_port, PTMP_5_37_port, PTMP_5_36_port, 
      PTMP_5_35_port, PTMP_5_34_port, PTMP_5_33_port, PTMP_5_32_port, 
      PTMP_5_31_port, PTMP_5_30_port, PTMP_5_29_port, PTMP_5_28_port, 
      PTMP_5_27_port, PTMP_5_26_port, PTMP_5_25_port, PTMP_5_24_port, 
      PTMP_5_23_port, PTMP_5_22_port, PTMP_5_21_port, PTMP_5_20_port, 
      PTMP_5_19_port, PTMP_5_18_port, PTMP_5_17_port, PTMP_5_16_port, 
      PTMP_5_15_port, PTMP_5_14_port, PTMP_5_13_port, PTMP_5_12_port, 
      PTMP_5_11_port, PTMP_5_10_port, PTMP_5_9_port, PTMP_5_8_port, 
      PTMP_5_7_port, PTMP_5_6_port, PTMP_5_5_port, PTMP_5_4_port, PTMP_5_3_port
      , PTMP_5_2_port, PTMP_5_1_port, PTMP_5_0_port, PTMP_4_43_port, 
      PTMP_4_42_port, PTMP_4_41_port, PTMP_4_40_port, PTMP_4_39_port, 
      PTMP_4_38_port, PTMP_4_37_port, PTMP_4_36_port, PTMP_4_35_port, 
      PTMP_4_34_port, PTMP_4_33_port, PTMP_4_32_port, PTMP_4_31_port, 
      PTMP_4_30_port, PTMP_4_29_port, PTMP_4_28_port, PTMP_4_27_port, 
      PTMP_4_26_port, PTMP_4_25_port, PTMP_4_24_port, PTMP_4_23_port, 
      PTMP_4_22_port, PTMP_4_21_port, PTMP_4_20_port, PTMP_4_19_port, 
      PTMP_4_18_port, PTMP_4_17_port, PTMP_4_16_port, PTMP_4_15_port, 
      PTMP_4_14_port, PTMP_4_13_port, PTMP_4_12_port, PTMP_4_11_port, 
      PTMP_4_10_port, PTMP_4_9_port, PTMP_4_8_port, PTMP_4_7_port, 
      PTMP_4_6_port, PTMP_4_5_port, PTMP_4_4_port, PTMP_4_3_port, PTMP_4_2_port
      , PTMP_4_1_port, PTMP_4_0_port, PTMP_3_41_port, PTMP_3_40_port, 
      PTMP_3_39_port, PTMP_3_38_port, PTMP_3_37_port, PTMP_3_36_port, 
      PTMP_3_35_port, PTMP_3_34_port, PTMP_3_33_port, PTMP_3_32_port, 
      PTMP_3_31_port, PTMP_3_30_port, PTMP_3_29_port, PTMP_3_28_port, 
      PTMP_3_27_port, PTMP_3_26_port, PTMP_3_25_port, PTMP_3_24_port, 
      PTMP_3_23_port, PTMP_3_22_port, PTMP_3_21_port, PTMP_3_20_port, 
      PTMP_3_19_port, PTMP_3_18_port, PTMP_3_17_port, PTMP_3_16_port, 
      PTMP_3_15_port, PTMP_3_14_port, PTMP_3_13_port, PTMP_3_12_port, 
      PTMP_3_11_port, PTMP_3_10_port, PTMP_3_9_port, PTMP_3_8_port, 
      PTMP_3_7_port, PTMP_3_6_port, PTMP_3_5_port, PTMP_3_4_port, PTMP_3_3_port
      , PTMP_3_2_port, PTMP_3_1_port, PTMP_3_0_port, PTMP_2_39_port, 
      PTMP_2_38_port, PTMP_2_37_port, PTMP_2_36_port, PTMP_2_35_port, 
      PTMP_2_34_port, PTMP_2_33_port, PTMP_2_32_port, PTMP_2_31_port, 
      PTMP_2_30_port, PTMP_2_29_port, PTMP_2_28_port, PTMP_2_27_port, 
      PTMP_2_26_port, PTMP_2_25_port, PTMP_2_24_port, PTMP_2_23_port, 
      PTMP_2_22_port, PTMP_2_21_port, PTMP_2_20_port, PTMP_2_19_port, 
      PTMP_2_18_port, PTMP_2_17_port, PTMP_2_16_port, PTMP_2_15_port, 
      PTMP_2_14_port, PTMP_2_13_port, PTMP_2_12_port, PTMP_2_11_port, 
      PTMP_2_10_port, PTMP_2_9_port, PTMP_2_8_port, PTMP_2_7_port, 
      PTMP_2_6_port, PTMP_2_5_port, PTMP_2_4_port, PTMP_2_3_port, PTMP_2_2_port
      , PTMP_2_1_port, PTMP_2_0_port, PTMP_1_37_port, PTMP_1_36_port, 
      PTMP_1_35_port, PTMP_1_34_port, PTMP_1_33_port, PTMP_1_32_port, 
      PTMP_1_31_port, PTMP_1_30_port, PTMP_1_29_port, PTMP_1_28_port, 
      PTMP_1_27_port, PTMP_1_26_port, PTMP_1_25_port, PTMP_1_24_port, 
      PTMP_1_23_port, PTMP_1_22_port, PTMP_1_21_port, PTMP_1_20_port, 
      PTMP_1_19_port, PTMP_1_18_port, PTMP_1_17_port, PTMP_1_16_port, 
      PTMP_1_15_port, PTMP_1_14_port, PTMP_1_13_port, PTMP_1_12_port, 
      PTMP_1_11_port, PTMP_1_10_port, PTMP_1_9_port, PTMP_1_8_port, 
      PTMP_1_7_port, PTMP_1_6_port, PTMP_1_5_port, PTMP_1_4_port, PTMP_1_3_port
      , PTMP_1_2_port, PTMP_1_1_port, PTMP_1_0_port, PTMP_0_36_port, 
      PTMP_0_34_port, PTMP_0_33_port, PTMP_0_32_port, PTMP_0_31_port, 
      PTMP_0_30_port, PTMP_0_29_port, PTMP_0_28_port, PTMP_0_27_port, 
      PTMP_0_26_port, PTMP_0_25_port, PTMP_0_24_port, PTMP_0_23_port, 
      PTMP_0_22_port, PTMP_0_21_port, PTMP_0_20_port, PTMP_0_19_port, 
      PTMP_0_18_port, PTMP_0_17_port, PTMP_0_16_port, PTMP_0_15_port, 
      PTMP_0_14_port, PTMP_0_13_port, PTMP_0_12_port, PTMP_0_11_port, 
      PTMP_0_10_port, PTMP_0_9_port, PTMP_0_8_port, PTMP_0_7_port, 
      PTMP_0_6_port, PTMP_0_5_port, PTMP_0_4_port, PTMP_0_3_port, PTMP_0_2_port
      , PTMP_0_1_port, PTMP_0_0_port, PTMP_13_61_port, PTMP_13_60_port, 
      PTMP_13_59_port, PTMP_13_58_port, PTMP_13_57_port, PTMP_13_56_port, 
      PTMP_13_55_port, PTMP_13_54_port, PTMP_13_53_port, PTMP_13_52_port, 
      PTMP_13_51_port, PTMP_13_50_port, PTMP_13_49_port, PTMP_13_48_port, 
      PTMP_13_47_port, PTMP_13_46_port, PTMP_13_45_port, PTMP_13_44_port, 
      PTMP_13_43_port, PTMP_13_42_port, PTMP_13_41_port, PTMP_13_40_port, 
      PTMP_13_39_port, PTMP_13_38_port, PTMP_13_37_port, PTMP_13_36_port, 
      PTMP_13_35_port, PTMP_13_34_port, PTMP_13_33_port, PTMP_13_32_port, 
      PTMP_13_31_port, PTMP_13_30_port, PTMP_13_29_port, PTMP_13_28_port, 
      PTMP_13_27_port, PTMP_13_26_port, PTMP_13_25_port, PTMP_13_24_port, 
      PTMP_13_23_port, PTMP_13_22_port, PTMP_13_21_port, PTMP_13_20_port, 
      PTMP_13_19_port, PTMP_13_18_port, PTMP_13_17_port, PTMP_13_16_port, 
      PTMP_13_15_port, PTMP_13_14_port, PTMP_13_13_port, PTMP_13_12_port, 
      PTMP_13_11_port, PTMP_13_10_port, PTMP_13_9_port, PTMP_13_8_port, 
      PTMP_13_7_port, PTMP_13_6_port, PTMP_13_5_port, PTMP_13_4_port, 
      PTMP_13_3_port, PTMP_13_2_port, PTMP_13_1_port, PTMP_13_0_port, 
      PTMP_12_59_port, PTMP_12_58_port, PTMP_12_57_port, PTMP_12_56_port, 
      PTMP_12_55_port, PTMP_12_54_port, PTMP_12_53_port, PTMP_12_52_port, 
      PTMP_12_51_port, PTMP_12_50_port, PTMP_12_49_port, PTMP_12_48_port, 
      PTMP_12_47_port, PTMP_12_46_port, PTMP_12_45_port, PTMP_12_44_port, 
      PTMP_12_43_port, PTMP_12_42_port, PTMP_12_41_port, PTMP_12_40_port, 
      PTMP_12_39_port, PTMP_12_38_port, PTMP_12_37_port, PTMP_12_36_port, 
      PTMP_12_35_port, PTMP_12_34_port, PTMP_12_33_port, PTMP_12_32_port, 
      PTMP_12_31_port, PTMP_12_30_port, PTMP_12_29_port, PTMP_12_28_port, 
      PTMP_12_27_port, PTMP_12_26_port, PTMP_12_25_port, PTMP_12_24_port, 
      PTMP_12_23_port, PTMP_12_22_port, PTMP_12_21_port, PTMP_12_20_port, 
      PTMP_12_19_port, PTMP_12_18_port, PTMP_12_17_port, PTMP_12_16_port, 
      PTMP_12_15_port, PTMP_12_14_port, PTMP_12_13_port, PTMP_12_12_port, 
      PTMP_12_11_port, PTMP_12_10_port, PTMP_12_9_port, PTMP_12_8_port, 
      PTMP_12_7_port, PTMP_12_6_port, PTMP_12_5_port, PTMP_12_4_port, 
      PTMP_12_3_port, PTMP_12_2_port, PTMP_12_1_port, PTMP_12_0_port, 
      PTMP_11_57_port, PTMP_11_56_port, PTMP_11_55_port, PTMP_11_54_port, 
      PTMP_11_53_port, PTMP_11_52_port, PTMP_11_51_port, PTMP_11_50_port, 
      PTMP_11_49_port, PTMP_11_48_port, PTMP_11_47_port, PTMP_11_46_port, 
      PTMP_11_45_port, PTMP_11_44_port, PTMP_11_43_port, PTMP_11_42_port, 
      PTMP_11_41_port, PTMP_11_40_port, PTMP_11_39_port, PTMP_11_38_port, 
      PTMP_11_37_port, PTMP_11_36_port, PTMP_11_35_port, PTMP_11_34_port, 
      PTMP_11_33_port, PTMP_11_32_port, PTMP_11_31_port, PTMP_11_30_port, 
      PTMP_11_29_port, PTMP_11_28_port, PTMP_11_27_port, PTMP_11_26_port, 
      PTMP_11_25_port, PTMP_11_24_port, PTMP_11_23_port, PTMP_11_22_port, 
      PTMP_11_21_port, PTMP_11_20_port, PTMP_11_19_port, PTMP_11_18_port, 
      PTMP_11_17_port, PTMP_11_16_port, PTMP_11_15_port, PTMP_11_14_port, 
      PTMP_11_13_port, PTMP_11_12_port, PTMP_11_11_port, PTMP_11_10_port, 
      PTMP_11_9_port, PTMP_11_8_port, PTMP_11_7_port, PTMP_11_6_port, 
      PTMP_11_5_port, PTMP_11_4_port, PTMP_11_3_port, PTMP_11_2_port, 
      PTMP_11_1_port, PTMP_11_0_port, PTMP_10_55_port, PTMP_10_54_port, 
      PTMP_10_53_port, PTMP_10_52_port, PTMP_10_51_port, PTMP_10_50_port, 
      PTMP_10_49_port, PTMP_10_48_port, PTMP_10_47_port, PTMP_10_46_port, 
      PTMP_10_45_port, PTMP_10_44_port, PTMP_10_43_port, PTMP_10_42_port, 
      PTMP_10_41_port, PTMP_10_40_port, PTMP_10_39_port, PTMP_10_38_port, 
      PTMP_10_37_port, PTMP_10_36_port, PTMP_10_35_port, PTMP_10_34_port, 
      PTMP_10_33_port, PTMP_10_32_port, PTMP_10_31_port, PTMP_10_30_port, 
      PTMP_10_29_port, PTMP_10_28_port, PTMP_10_27_port, PTMP_10_26_port, 
      PTMP_10_25_port, PTMP_10_24_port, PTMP_10_23_port, PTMP_10_22_port, 
      PTMP_10_21_port, PTMP_10_20_port, PTMP_10_19_port, PTMP_10_18_port, 
      PTMP_10_17_port, PTMP_10_16_port, PTMP_10_15_port, PTMP_10_14_port, 
      PTMP_10_13_port, PTMP_10_12_port, PTMP_10_11_port, PTMP_10_10_port, 
      PTMP_10_9_port, PTMP_10_8_port, PTMP_10_7_port, PTMP_10_6_port, 
      PTMP_10_5_port, PTMP_10_4_port, PTMP_10_3_port, PTMP_10_2_port, 
      PTMP_10_1_port, PTMP_10_0_port, PTMP_9_53_port, PTMP_9_52_port, 
      PTMP_9_51_port, PTMP_9_50_port, PTMP_9_49_port, PTMP_9_48_port, 
      PTMP_9_47_port, PTMP_9_46_port, PTMP_9_45_port, PTMP_9_44_port, 
      PTMP_9_43_port, PTMP_9_42_port, PTMP_9_41_port, PTMP_9_40_port, 
      PTMP_9_39_port, PTMP_9_38_port, PTMP_9_37_port, PTMP_9_36_port, 
      PTMP_9_35_port, PTMP_9_34_port, PTMP_9_33_port, PTMP_9_32_port, 
      PTMP_9_31_port, PTMP_9_30_port, PTMP_9_29_port, PTMP_9_28_port, 
      PTMP_9_27_port, PTMP_9_26_port, PTMP_9_25_port, PTMP_9_24_port, 
      PTMP_9_23_port, PTMP_9_22_port, PTMP_9_21_port, PTMP_9_20_port, 
      PTMP_9_19_port, PTMP_9_18_port, PTMP_9_17_port, PTMP_9_16_port, 
      PTMP_9_15_port, PTMP_9_14_port, PTMP_9_13_port, PTMP_9_12_port, 
      PTMP_9_11_port, PTMP_9_10_port, PTMP_9_9_port, PTMP_9_8_port, 
      PTMP_9_7_port, PTMP_9_6_port, PTMP_9_5_port, PTMP_9_4_port, PTMP_9_3_port
      , PTMP_9_2_port, PTMP_9_1_port, PTMP_9_0_port, PTMP_8_51_port, 
      PTMP_8_50_port, PTMP_8_49_port, PTMP_8_48_port, PTMP_8_47_port, 
      PTMP_8_46_port, PTMP_8_45_port, PTMP_8_44_port, PTMP_8_43_port, 
      PTMP_8_42_port, PTMP_8_41_port, PTMP_8_40_port, PTMP_8_39_port, 
      PTMP_8_38_port, PTMP_8_37_port, PTMP_8_36_port, PTMP_8_35_port, 
      PTMP_8_34_port, PTMP_8_33_port, PTMP_8_32_port, PTMP_8_31_port, 
      PTMP_8_30_port, PTMP_8_29_port, PTMP_8_28_port, PTMP_8_27_port, 
      PTMP_8_26_port, PTMP_8_25_port, PTMP_8_24_port, PTMP_8_23_port, 
      PTMP_8_22_port, PTMP_8_21_port, PTMP_8_20_port, PTMP_8_19_port, 
      PTMP_8_18_port, PTMP_8_17_port, PTMP_8_16_port, n4, n5, n6, n7, n8, n9, 
      n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n_1080, 
      n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, 
      n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, 
      n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, 
      n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, 
      n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, 
      n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, 
      n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, 
      n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, 
      n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, 
      n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, 
      n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, 
      n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, 
      n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, 
      n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, 
      n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, 
      n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, 
      n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, 
      n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, 
      n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, 
      n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, 
      n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, 
      n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, 
      n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, 
      n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296 : 
      std_logic;

begin
   
   X_Logic0_port <= '0';
   OTMP_15_0_port <= '0';
   SHIFT_n_15_0_port <= '0';
   SHIFT_n_15_1_port <= '0';
   SHIFT_15_0_port <= '0';
   SHIFT_15_1_port <= '0';
   OTMP_14_0_port <= '0';
   SHIFT_n_14_0_port <= '0';
   SHIFT_n_14_1_port <= '0';
   SHIFT_14_0_port <= '0';
   SHIFT_14_1_port <= '0';
   OTMP_13_0_port <= '0';
   SHIFT_n_13_0_port <= '0';
   SHIFT_n_13_1_port <= '0';
   SHIFT_13_0_port <= '0';
   SHIFT_13_1_port <= '0';
   OTMP_12_0_port <= '0';
   SHIFT_n_12_0_port <= '0';
   SHIFT_n_12_1_port <= '0';
   SHIFT_12_0_port <= '0';
   SHIFT_12_1_port <= '0';
   OTMP_11_0_port <= '0';
   SHIFT_n_11_0_port <= '0';
   SHIFT_n_11_1_port <= '0';
   SHIFT_11_0_port <= '0';
   SHIFT_11_1_port <= '0';
   OTMP_10_0_port <= '0';
   SHIFT_n_10_0_port <= '0';
   SHIFT_n_10_1_port <= '0';
   SHIFT_10_0_port <= '0';
   SHIFT_10_1_port <= '0';
   OTMP_9_0_port <= '0';
   SHIFT_n_9_0_port <= '0';
   SHIFT_n_9_1_port <= '0';
   SHIFT_9_0_port <= '0';
   SHIFT_9_1_port <= '0';
   OTMP_8_0_port <= '0';
   SHIFT_n_8_0_port <= '0';
   SHIFT_n_8_1_port <= '0';
   SHIFT_8_0_port <= '0';
   SHIFT_8_1_port <= '0';
   OTMP_7_0_port <= '0';
   SHIFT_n_7_0_port <= '0';
   SHIFT_n_7_1_port <= '0';
   SHIFT_7_0_port <= '0';
   SHIFT_7_1_port <= '0';
   OTMP_6_0_port <= '0';
   SHIFT_n_6_0_port <= '0';
   SHIFT_n_6_1_port <= '0';
   SHIFT_6_0_port <= '0';
   SHIFT_6_1_port <= '0';
   OTMP_5_0_port <= '0';
   SHIFT_n_5_0_port <= '0';
   SHIFT_n_5_1_port <= '0';
   SHIFT_5_0_port <= '0';
   SHIFT_5_1_port <= '0';
   OTMP_4_0_port <= '0';
   SHIFT_n_4_0_port <= '0';
   SHIFT_n_4_1_port <= '0';
   SHIFT_4_0_port <= '0';
   SHIFT_4_1_port <= '0';
   OTMP_3_0_port <= '0';
   SHIFT_n_3_0_port <= '0';
   SHIFT_n_3_1_port <= '0';
   SHIFT_3_0_port <= '0';
   SHIFT_3_1_port <= '0';
   OTMP_2_0_port <= '0';
   SHIFT_n_2_0_port <= '0';
   SHIFT_n_2_1_port <= '0';
   SHIFT_2_0_port <= '0';
   SHIFT_2_1_port <= '0';
   OTMP_1_0_port <= '0';
   SHIFT_n_1_0_port <= '0';
   SHIFT_1_0_port <= '0';
   n4 <= '0';
   n5 <= '0';
   ENC1 : BOOTHENC_NBIT34_i0 port map( A_s(33) => A(31), A_s(32) => A(31), 
                           A_s(31) => A(31), A_s(30) => A(30), A_s(29) => A(29)
                           , A_s(28) => A(28), A_s(27) => A(27), A_s(26) => 
                           A(26), A_s(25) => A(25), A_s(24) => A(24), A_s(23) 
                           => A(23), A_s(22) => A(22), A_s(21) => A(21), 
                           A_s(20) => A(20), A_s(19) => A(19), A_s(18) => A(18)
                           , A_s(17) => A(17), A_s(16) => A(16), A_s(15) => 
                           A(15), A_s(14) => A(14), A_s(13) => A(13), A_s(12) 
                           => A(12), A_s(11) => A(11), A_s(10) => A(10), A_s(9)
                           => A(9), A_s(8) => A(8), A_s(7) => A(7), A_s(6) => 
                           A(6), A_s(5) => A(5), A_s(4) => A(4), A_s(3) => A(3)
                           , A_s(2) => n7, A_s(1) => n8, A_s(0) => n9, A_ns(33)
                           => A_n_65, A_ns(32) => A_n_65, A_ns(31) => A_n_65, 
                           A_ns(30) => A_n_30_port, A_ns(29) => A_n_29_port, 
                           A_ns(28) => A_n_28_port, A_ns(27) => A_n_27_port, 
                           A_ns(26) => A_n_26_port, A_ns(25) => A_n_25_port, 
                           A_ns(24) => A_n_24_port, A_ns(23) => A_n_23_port, 
                           A_ns(22) => A_n_22_port, A_ns(21) => A_n_21_port, 
                           A_ns(20) => A_n_20_port, A_ns(19) => A_n_19_port, 
                           A_ns(18) => A_n_18_port, A_ns(17) => A_n_17_port, 
                           A_ns(16) => A_n_16_port, A_ns(15) => A_n_15_port, 
                           A_ns(14) => A_n_14_port, A_ns(13) => A_n_13_port, 
                           A_ns(12) => A_n_12_port, A_ns(11) => A_n_11_port, 
                           A_ns(10) => A_n_10_port, A_ns(9) => A_n_9_port, 
                           A_ns(8) => A_n_8_port, A_ns(7) => A_n_7_port, 
                           A_ns(6) => A_n_6_port, A_ns(5) => A_n_5_port, 
                           A_ns(4) => A_n_4_port, A_ns(3) => A_n_3_port, 
                           A_ns(2) => A_n_2_port, A_ns(1) => A_n_1_port, 
                           A_ns(0) => A_n_0_port, B(33) => B(31), B(32) => 
                           B(31), B(31) => B(31), B(30) => B(30), B(29) => 
                           B(29), B(28) => B(28), B(27) => B(27), B(26) => 
                           B(26), B(25) => B(25), B(24) => B(24), B(23) => 
                           B(23), B(22) => B(22), B(21) => B(21), B(20) => 
                           B(20), B(19) => B(19), B(18) => B(18), B(17) => 
                           B(17), B(16) => B(16), B(15) => B(15), B(14) => 
                           B(14), B(13) => B(13), B(12) => B(12), B(11) => 
                           B(11), B(10) => B(10), B(9) => B(9), B(8) => B(8), 
                           B(7) => B(7), B(6) => B(6), B(5) => B(5), B(4) => 
                           B(4), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), O(33) => OTMP_0_34_port, O(32) => 
                           OTMP_0_32_port, O(31) => OTMP_0_31_port, O(30) => 
                           OTMP_0_30_port, O(29) => OTMP_0_29_port, O(28) => 
                           OTMP_0_28_port, O(27) => OTMP_0_27_port, O(26) => 
                           OTMP_0_26_port, O(25) => OTMP_0_25_port, O(24) => 
                           OTMP_0_24_port, O(23) => OTMP_0_23_port, O(22) => 
                           OTMP_0_22_port, O(21) => OTMP_0_21_port, O(20) => 
                           OTMP_0_20_port, O(19) => OTMP_0_19_port, O(18) => 
                           OTMP_0_18_port, O(17) => OTMP_0_17_port, O(16) => 
                           OTMP_0_16_port, O(15) => OTMP_0_15_port, O(14) => 
                           OTMP_0_14_port, O(13) => OTMP_0_13_port, O(12) => 
                           OTMP_0_12_port, O(11) => OTMP_0_11_port, O(10) => 
                           OTMP_0_10_port, O(9) => OTMP_0_9_port, O(8) => 
                           OTMP_0_8_port, O(7) => OTMP_0_7_port, O(6) => 
                           OTMP_0_6_port, O(5) => OTMP_0_5_port, O(4) => 
                           OTMP_0_4_port, O(3) => OTMP_0_3_port, O(2) => 
                           OTMP_0_2_port, O(1) => OTMP_0_1_port, O(0) => 
                           OTMP_0_0_port, A_so(33) => SHIFT_1_33_port, A_so(32)
                           => SHIFT_1_32_port, A_so(31) => SHIFT_1_31_port, 
                           A_so(30) => SHIFT_1_30_port, A_so(29) => 
                           SHIFT_1_29_port, A_so(28) => SHIFT_1_28_port, 
                           A_so(27) => SHIFT_1_27_port, A_so(26) => 
                           SHIFT_1_26_port, A_so(25) => SHIFT_1_25_port, 
                           A_so(24) => SHIFT_1_24_port, A_so(23) => 
                           SHIFT_1_23_port, A_so(22) => SHIFT_1_22_port, 
                           A_so(21) => SHIFT_1_21_port, A_so(20) => 
                           SHIFT_1_20_port, A_so(19) => SHIFT_1_19_port, 
                           A_so(18) => SHIFT_1_18_port, A_so(17) => 
                           SHIFT_1_17_port, A_so(16) => SHIFT_1_16_port, 
                           A_so(15) => SHIFT_1_15_port, A_so(14) => 
                           SHIFT_1_14_port, A_so(13) => SHIFT_1_13_port, 
                           A_so(12) => SHIFT_1_12_port, A_so(11) => 
                           SHIFT_1_11_port, A_so(10) => SHIFT_1_10_port, 
                           A_so(9) => SHIFT_1_9_port, A_so(8) => SHIFT_1_8_port
                           , A_so(7) => SHIFT_1_7_port, A_so(6) => 
                           SHIFT_1_6_port, A_so(5) => SHIFT_1_5_port, A_so(4) 
                           => SHIFT_1_4_port, A_so(3) => SHIFT_1_3_port, 
                           A_so(2) => SHIFT_1_2_port, A_so(1) => SHIFT_1_1_port
                           , A_so(0) => n_1080, A_nso(33) => SHIFT_n_1_33_port,
                           A_nso(32) => SHIFT_n_1_32_port, A_nso(31) => 
                           SHIFT_n_1_31_port, A_nso(30) => SHIFT_n_1_30_port, 
                           A_nso(29) => SHIFT_n_1_29_port, A_nso(28) => 
                           SHIFT_n_1_28_port, A_nso(27) => SHIFT_n_1_27_port, 
                           A_nso(26) => SHIFT_n_1_26_port, A_nso(25) => 
                           SHIFT_n_1_25_port, A_nso(24) => SHIFT_n_1_24_port, 
                           A_nso(23) => SHIFT_n_1_23_port, A_nso(22) => 
                           SHIFT_n_1_22_port, A_nso(21) => SHIFT_n_1_21_port, 
                           A_nso(20) => SHIFT_n_1_20_port, A_nso(19) => 
                           SHIFT_n_1_19_port, A_nso(18) => SHIFT_n_1_18_port, 
                           A_nso(17) => SHIFT_n_1_17_port, A_nso(16) => 
                           SHIFT_n_1_16_port, A_nso(15) => SHIFT_n_1_15_port, 
                           A_nso(14) => SHIFT_n_1_14_port, A_nso(13) => 
                           SHIFT_n_1_13_port, A_nso(12) => SHIFT_n_1_12_port, 
                           A_nso(11) => SHIFT_n_1_11_port, A_nso(10) => 
                           SHIFT_n_1_10_port, A_nso(9) => SHIFT_n_1_9_port, 
                           A_nso(8) => SHIFT_n_1_8_port, A_nso(7) => 
                           SHIFT_n_1_7_port, A_nso(6) => SHIFT_n_1_6_port, 
                           A_nso(5) => SHIFT_n_1_5_port, A_nso(4) => 
                           SHIFT_n_1_4_port, A_nso(3) => SHIFT_n_1_3_port, 
                           A_nso(2) => SHIFT_n_1_2_port, A_nso(1) => 
                           SHIFT_n_1_1_port, A_nso(0) => n_1081);
   ENC_1 : BOOTHENC_NBIT36_i2 port map( A_s(35) => SHIFT_1_33_port, A_s(34) => 
                           SHIFT_1_33_port, A_s(33) => SHIFT_1_33_port, A_s(32)
                           => SHIFT_1_32_port, A_s(31) => SHIFT_1_31_port, 
                           A_s(30) => SHIFT_1_30_port, A_s(29) => 
                           SHIFT_1_29_port, A_s(28) => SHIFT_1_28_port, A_s(27)
                           => SHIFT_1_27_port, A_s(26) => SHIFT_1_26_port, 
                           A_s(25) => SHIFT_1_25_port, A_s(24) => 
                           SHIFT_1_24_port, A_s(23) => SHIFT_1_23_port, A_s(22)
                           => SHIFT_1_22_port, A_s(21) => SHIFT_1_21_port, 
                           A_s(20) => SHIFT_1_20_port, A_s(19) => 
                           SHIFT_1_19_port, A_s(18) => SHIFT_1_18_port, A_s(17)
                           => SHIFT_1_17_port, A_s(16) => SHIFT_1_16_port, 
                           A_s(15) => SHIFT_1_15_port, A_s(14) => 
                           SHIFT_1_14_port, A_s(13) => SHIFT_1_13_port, A_s(12)
                           => SHIFT_1_12_port, A_s(11) => SHIFT_1_11_port, 
                           A_s(10) => SHIFT_1_10_port, A_s(9) => SHIFT_1_9_port
                           , A_s(8) => SHIFT_1_8_port, A_s(7) => SHIFT_1_7_port
                           , A_s(6) => SHIFT_1_6_port, A_s(5) => SHIFT_1_5_port
                           , A_s(4) => SHIFT_1_4_port, A_s(3) => SHIFT_1_3_port
                           , A_s(2) => SHIFT_1_2_port, A_s(1) => SHIFT_1_1_port
                           , A_s(0) => SHIFT_1_0_port, A_ns(35) => 
                           SHIFT_n_1_33_port, A_ns(34) => SHIFT_n_1_33_port, 
                           A_ns(33) => SHIFT_n_1_33_port, A_ns(32) => 
                           SHIFT_n_1_32_port, A_ns(31) => SHIFT_n_1_31_port, 
                           A_ns(30) => SHIFT_n_1_30_port, A_ns(29) => 
                           SHIFT_n_1_29_port, A_ns(28) => SHIFT_n_1_28_port, 
                           A_ns(27) => SHIFT_n_1_27_port, A_ns(26) => 
                           SHIFT_n_1_26_port, A_ns(25) => SHIFT_n_1_25_port, 
                           A_ns(24) => SHIFT_n_1_24_port, A_ns(23) => 
                           SHIFT_n_1_23_port, A_ns(22) => SHIFT_n_1_22_port, 
                           A_ns(21) => SHIFT_n_1_21_port, A_ns(20) => 
                           SHIFT_n_1_20_port, A_ns(19) => SHIFT_n_1_19_port, 
                           A_ns(18) => SHIFT_n_1_18_port, A_ns(17) => 
                           SHIFT_n_1_17_port, A_ns(16) => SHIFT_n_1_16_port, 
                           A_ns(15) => SHIFT_n_1_15_port, A_ns(14) => 
                           SHIFT_n_1_14_port, A_ns(13) => SHIFT_n_1_13_port, 
                           A_ns(12) => SHIFT_n_1_12_port, A_ns(11) => 
                           SHIFT_n_1_11_port, A_ns(10) => SHIFT_n_1_10_port, 
                           A_ns(9) => SHIFT_n_1_9_port, A_ns(8) => 
                           SHIFT_n_1_8_port, A_ns(7) => SHIFT_n_1_7_port, 
                           A_ns(6) => SHIFT_n_1_6_port, A_ns(5) => 
                           SHIFT_n_1_5_port, A_ns(4) => SHIFT_n_1_4_port, 
                           A_ns(3) => SHIFT_n_1_3_port, A_ns(2) => 
                           SHIFT_n_1_2_port, A_ns(1) => SHIFT_n_1_1_port, 
                           A_ns(0) => SHIFT_n_1_0_port, B(35) => B(31), B(34) 
                           => B(31), B(33) => B(31), B(32) => B(31), B(31) => 
                           B(31), B(30) => B(30), B(29) => B(29), B(28) => 
                           B(28), B(27) => B(27), B(26) => B(26), B(25) => 
                           B(25), B(24) => B(24), B(23) => B(23), B(22) => 
                           B(22), B(21) => B(21), B(20) => B(20), B(19) => 
                           B(19), B(18) => B(18), B(17) => B(17), B(16) => 
                           B(16), B(15) => B(15), B(14) => B(14), B(13) => 
                           B(13), B(12) => B(12), B(11) => B(11), B(10) => 
                           B(10), B(9) => B(9), B(8) => B(8), B(7) => B(7), 
                           B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3) => 
                           B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), 
                           O(35) => OTMP_1_35_port, O(34) => OTMP_1_34_port, 
                           O(33) => OTMP_1_33_port, O(32) => OTMP_1_32_port, 
                           O(31) => OTMP_1_31_port, O(30) => OTMP_1_30_port, 
                           O(29) => OTMP_1_29_port, O(28) => OTMP_1_28_port, 
                           O(27) => OTMP_1_27_port, O(26) => OTMP_1_26_port, 
                           O(25) => OTMP_1_25_port, O(24) => OTMP_1_24_port, 
                           O(23) => OTMP_1_23_port, O(22) => OTMP_1_22_port, 
                           O(21) => OTMP_1_21_port, O(20) => OTMP_1_20_port, 
                           O(19) => OTMP_1_19_port, O(18) => OTMP_1_18_port, 
                           O(17) => OTMP_1_17_port, O(16) => OTMP_1_16_port, 
                           O(15) => OTMP_1_15_port, O(14) => OTMP_1_14_port, 
                           O(13) => OTMP_1_13_port, O(12) => OTMP_1_12_port, 
                           O(11) => OTMP_1_11_port, O(10) => OTMP_1_10_port, 
                           O(9) => OTMP_1_9_port, O(8) => OTMP_1_8_port, O(7) 
                           => OTMP_1_7_port, O(6) => OTMP_1_6_port, O(5) => 
                           OTMP_1_5_port, O(4) => OTMP_1_4_port, O(3) => 
                           OTMP_1_3_port, O(2) => OTMP_1_2_port, O(1) => 
                           OTMP_1_1_port, O(0) => n_1082, A_so(35) => 
                           SHIFT_2_35_port, A_so(34) => SHIFT_2_34_port, 
                           A_so(33) => SHIFT_2_33_port, A_so(32) => 
                           SHIFT_2_32_port, A_so(31) => SHIFT_2_31_port, 
                           A_so(30) => SHIFT_2_30_port, A_so(29) => 
                           SHIFT_2_29_port, A_so(28) => SHIFT_2_28_port, 
                           A_so(27) => SHIFT_2_27_port, A_so(26) => 
                           SHIFT_2_26_port, A_so(25) => SHIFT_2_25_port, 
                           A_so(24) => SHIFT_2_24_port, A_so(23) => 
                           SHIFT_2_23_port, A_so(22) => SHIFT_2_22_port, 
                           A_so(21) => SHIFT_2_21_port, A_so(20) => 
                           SHIFT_2_20_port, A_so(19) => SHIFT_2_19_port, 
                           A_so(18) => SHIFT_2_18_port, A_so(17) => 
                           SHIFT_2_17_port, A_so(16) => SHIFT_2_16_port, 
                           A_so(15) => SHIFT_2_15_port, A_so(14) => 
                           SHIFT_2_14_port, A_so(13) => SHIFT_2_13_port, 
                           A_so(12) => SHIFT_2_12_port, A_so(11) => 
                           SHIFT_2_11_port, A_so(10) => SHIFT_2_10_port, 
                           A_so(9) => SHIFT_2_9_port, A_so(8) => SHIFT_2_8_port
                           , A_so(7) => SHIFT_2_7_port, A_so(6) => 
                           SHIFT_2_6_port, A_so(5) => SHIFT_2_5_port, A_so(4) 
                           => SHIFT_2_4_port, A_so(3) => SHIFT_2_3_port, 
                           A_so(2) => SHIFT_2_2_port, A_so(1) => n_1083, 
                           A_so(0) => n_1084, A_nso(35) => SHIFT_n_2_35_port, 
                           A_nso(34) => SHIFT_n_2_34_port, A_nso(33) => 
                           SHIFT_n_2_33_port, A_nso(32) => SHIFT_n_2_32_port, 
                           A_nso(31) => SHIFT_n_2_31_port, A_nso(30) => 
                           SHIFT_n_2_30_port, A_nso(29) => SHIFT_n_2_29_port, 
                           A_nso(28) => SHIFT_n_2_28_port, A_nso(27) => 
                           SHIFT_n_2_27_port, A_nso(26) => SHIFT_n_2_26_port, 
                           A_nso(25) => SHIFT_n_2_25_port, A_nso(24) => 
                           SHIFT_n_2_24_port, A_nso(23) => SHIFT_n_2_23_port, 
                           A_nso(22) => SHIFT_n_2_22_port, A_nso(21) => 
                           SHIFT_n_2_21_port, A_nso(20) => SHIFT_n_2_20_port, 
                           A_nso(19) => SHIFT_n_2_19_port, A_nso(18) => 
                           SHIFT_n_2_18_port, A_nso(17) => SHIFT_n_2_17_port, 
                           A_nso(16) => SHIFT_n_2_16_port, A_nso(15) => 
                           SHIFT_n_2_15_port, A_nso(14) => SHIFT_n_2_14_port, 
                           A_nso(13) => SHIFT_n_2_13_port, A_nso(12) => 
                           SHIFT_n_2_12_port, A_nso(11) => SHIFT_n_2_11_port, 
                           A_nso(10) => SHIFT_n_2_10_port, A_nso(9) => 
                           SHIFT_n_2_9_port, A_nso(8) => SHIFT_n_2_8_port, 
                           A_nso(7) => SHIFT_n_2_7_port, A_nso(6) => 
                           SHIFT_n_2_6_port, A_nso(5) => SHIFT_n_2_5_port, 
                           A_nso(4) => SHIFT_n_2_4_port, A_nso(3) => 
                           SHIFT_n_2_3_port, A_nso(2) => SHIFT_n_2_2_port, 
                           A_nso(1) => n_1085, A_nso(0) => n_1086);
   ENC_2 : BOOTHENC_NBIT38_i4 port map( A_s(37) => SHIFT_2_35_port, A_s(36) => 
                           SHIFT_2_35_port, A_s(35) => SHIFT_2_35_port, A_s(34)
                           => SHIFT_2_34_port, A_s(33) => SHIFT_2_33_port, 
                           A_s(32) => SHIFT_2_32_port, A_s(31) => 
                           SHIFT_2_31_port, A_s(30) => SHIFT_2_30_port, A_s(29)
                           => SHIFT_2_29_port, A_s(28) => SHIFT_2_28_port, 
                           A_s(27) => SHIFT_2_27_port, A_s(26) => 
                           SHIFT_2_26_port, A_s(25) => SHIFT_2_25_port, A_s(24)
                           => SHIFT_2_24_port, A_s(23) => SHIFT_2_23_port, 
                           A_s(22) => SHIFT_2_22_port, A_s(21) => 
                           SHIFT_2_21_port, A_s(20) => SHIFT_2_20_port, A_s(19)
                           => SHIFT_2_19_port, A_s(18) => SHIFT_2_18_port, 
                           A_s(17) => SHIFT_2_17_port, A_s(16) => 
                           SHIFT_2_16_port, A_s(15) => SHIFT_2_15_port, A_s(14)
                           => SHIFT_2_14_port, A_s(13) => SHIFT_2_13_port, 
                           A_s(12) => SHIFT_2_12_port, A_s(11) => 
                           SHIFT_2_11_port, A_s(10) => SHIFT_2_10_port, A_s(9) 
                           => SHIFT_2_9_port, A_s(8) => SHIFT_2_8_port, A_s(7) 
                           => SHIFT_2_7_port, A_s(6) => SHIFT_2_6_port, A_s(5) 
                           => SHIFT_2_5_port, A_s(4) => SHIFT_2_4_port, A_s(3) 
                           => SHIFT_2_3_port, A_s(2) => SHIFT_2_2_port, A_s(1) 
                           => SHIFT_2_1_port, A_s(0) => SHIFT_2_0_port, 
                           A_ns(37) => SHIFT_n_2_35_port, A_ns(36) => 
                           SHIFT_n_2_35_port, A_ns(35) => SHIFT_n_2_35_port, 
                           A_ns(34) => SHIFT_n_2_34_port, A_ns(33) => 
                           SHIFT_n_2_33_port, A_ns(32) => SHIFT_n_2_32_port, 
                           A_ns(31) => SHIFT_n_2_31_port, A_ns(30) => 
                           SHIFT_n_2_30_port, A_ns(29) => SHIFT_n_2_29_port, 
                           A_ns(28) => SHIFT_n_2_28_port, A_ns(27) => 
                           SHIFT_n_2_27_port, A_ns(26) => SHIFT_n_2_26_port, 
                           A_ns(25) => SHIFT_n_2_25_port, A_ns(24) => 
                           SHIFT_n_2_24_port, A_ns(23) => SHIFT_n_2_23_port, 
                           A_ns(22) => SHIFT_n_2_22_port, A_ns(21) => 
                           SHIFT_n_2_21_port, A_ns(20) => SHIFT_n_2_20_port, 
                           A_ns(19) => SHIFT_n_2_19_port, A_ns(18) => 
                           SHIFT_n_2_18_port, A_ns(17) => SHIFT_n_2_17_port, 
                           A_ns(16) => SHIFT_n_2_16_port, A_ns(15) => 
                           SHIFT_n_2_15_port, A_ns(14) => SHIFT_n_2_14_port, 
                           A_ns(13) => SHIFT_n_2_13_port, A_ns(12) => 
                           SHIFT_n_2_12_port, A_ns(11) => SHIFT_n_2_11_port, 
                           A_ns(10) => SHIFT_n_2_10_port, A_ns(9) => 
                           SHIFT_n_2_9_port, A_ns(8) => SHIFT_n_2_8_port, 
                           A_ns(7) => SHIFT_n_2_7_port, A_ns(6) => 
                           SHIFT_n_2_6_port, A_ns(5) => SHIFT_n_2_5_port, 
                           A_ns(4) => SHIFT_n_2_4_port, A_ns(3) => 
                           SHIFT_n_2_3_port, A_ns(2) => SHIFT_n_2_2_port, 
                           A_ns(1) => SHIFT_n_2_1_port, A_ns(0) => 
                           SHIFT_n_2_0_port, B(37) => B(31), B(36) => B(31), 
                           B(35) => B(31), B(34) => B(31), B(33) => B(31), 
                           B(32) => B(31), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), O(37) => OTMP_2_37_port, O(36) 
                           => OTMP_2_36_port, O(35) => OTMP_2_35_port, O(34) =>
                           OTMP_2_34_port, O(33) => OTMP_2_33_port, O(32) => 
                           OTMP_2_32_port, O(31) => OTMP_2_31_port, O(30) => 
                           OTMP_2_30_port, O(29) => OTMP_2_29_port, O(28) => 
                           OTMP_2_28_port, O(27) => OTMP_2_27_port, O(26) => 
                           OTMP_2_26_port, O(25) => OTMP_2_25_port, O(24) => 
                           OTMP_2_24_port, O(23) => OTMP_2_23_port, O(22) => 
                           OTMP_2_22_port, O(21) => OTMP_2_21_port, O(20) => 
                           OTMP_2_20_port, O(19) => OTMP_2_19_port, O(18) => 
                           OTMP_2_18_port, O(17) => OTMP_2_17_port, O(16) => 
                           OTMP_2_16_port, O(15) => OTMP_2_15_port, O(14) => 
                           OTMP_2_14_port, O(13) => OTMP_2_13_port, O(12) => 
                           OTMP_2_12_port, O(11) => OTMP_2_11_port, O(10) => 
                           OTMP_2_10_port, O(9) => OTMP_2_9_port, O(8) => 
                           OTMP_2_8_port, O(7) => OTMP_2_7_port, O(6) => 
                           OTMP_2_6_port, O(5) => OTMP_2_5_port, O(4) => 
                           OTMP_2_4_port, O(3) => OTMP_2_3_port, O(2) => 
                           OTMP_2_2_port, O(1) => OTMP_2_1_port, O(0) => n_1087
                           , A_so(37) => SHIFT_3_37_port, A_so(36) => 
                           SHIFT_3_36_port, A_so(35) => SHIFT_3_35_port, 
                           A_so(34) => SHIFT_3_34_port, A_so(33) => 
                           SHIFT_3_33_port, A_so(32) => SHIFT_3_32_port, 
                           A_so(31) => SHIFT_3_31_port, A_so(30) => 
                           SHIFT_3_30_port, A_so(29) => SHIFT_3_29_port, 
                           A_so(28) => SHIFT_3_28_port, A_so(27) => 
                           SHIFT_3_27_port, A_so(26) => SHIFT_3_26_port, 
                           A_so(25) => SHIFT_3_25_port, A_so(24) => 
                           SHIFT_3_24_port, A_so(23) => SHIFT_3_23_port, 
                           A_so(22) => SHIFT_3_22_port, A_so(21) => 
                           SHIFT_3_21_port, A_so(20) => SHIFT_3_20_port, 
                           A_so(19) => SHIFT_3_19_port, A_so(18) => 
                           SHIFT_3_18_port, A_so(17) => SHIFT_3_17_port, 
                           A_so(16) => SHIFT_3_16_port, A_so(15) => 
                           SHIFT_3_15_port, A_so(14) => SHIFT_3_14_port, 
                           A_so(13) => SHIFT_3_13_port, A_so(12) => 
                           SHIFT_3_12_port, A_so(11) => SHIFT_3_11_port, 
                           A_so(10) => SHIFT_3_10_port, A_so(9) => 
                           SHIFT_3_9_port, A_so(8) => SHIFT_3_8_port, A_so(7) 
                           => SHIFT_3_7_port, A_so(6) => SHIFT_3_6_port, 
                           A_so(5) => SHIFT_3_5_port, A_so(4) => SHIFT_3_4_port
                           , A_so(3) => SHIFT_3_3_port, A_so(2) => 
                           SHIFT_3_2_port, A_so(1) => n_1088, A_so(0) => n_1089
                           , A_nso(37) => SHIFT_n_3_37_port, A_nso(36) => 
                           SHIFT_n_3_36_port, A_nso(35) => SHIFT_n_3_35_port, 
                           A_nso(34) => SHIFT_n_3_34_port, A_nso(33) => 
                           SHIFT_n_3_33_port, A_nso(32) => SHIFT_n_3_32_port, 
                           A_nso(31) => SHIFT_n_3_31_port, A_nso(30) => 
                           SHIFT_n_3_30_port, A_nso(29) => SHIFT_n_3_29_port, 
                           A_nso(28) => SHIFT_n_3_28_port, A_nso(27) => 
                           SHIFT_n_3_27_port, A_nso(26) => SHIFT_n_3_26_port, 
                           A_nso(25) => SHIFT_n_3_25_port, A_nso(24) => 
                           SHIFT_n_3_24_port, A_nso(23) => SHIFT_n_3_23_port, 
                           A_nso(22) => SHIFT_n_3_22_port, A_nso(21) => 
                           SHIFT_n_3_21_port, A_nso(20) => SHIFT_n_3_20_port, 
                           A_nso(19) => SHIFT_n_3_19_port, A_nso(18) => 
                           SHIFT_n_3_18_port, A_nso(17) => SHIFT_n_3_17_port, 
                           A_nso(16) => SHIFT_n_3_16_port, A_nso(15) => 
                           SHIFT_n_3_15_port, A_nso(14) => SHIFT_n_3_14_port, 
                           A_nso(13) => SHIFT_n_3_13_port, A_nso(12) => 
                           SHIFT_n_3_12_port, A_nso(11) => SHIFT_n_3_11_port, 
                           A_nso(10) => SHIFT_n_3_10_port, A_nso(9) => 
                           SHIFT_n_3_9_port, A_nso(8) => SHIFT_n_3_8_port, 
                           A_nso(7) => SHIFT_n_3_7_port, A_nso(6) => 
                           SHIFT_n_3_6_port, A_nso(5) => SHIFT_n_3_5_port, 
                           A_nso(4) => SHIFT_n_3_4_port, A_nso(3) => 
                           SHIFT_n_3_3_port, A_nso(2) => SHIFT_n_3_2_port, 
                           A_nso(1) => n_1090, A_nso(0) => n_1091);
   ENC_3 : BOOTHENC_NBIT40_i6 port map( A_s(39) => n21, A_s(38) => n21, A_s(37)
                           => n21, A_s(36) => SHIFT_3_36_port, A_s(35) => 
                           SHIFT_3_35_port, A_s(34) => SHIFT_3_34_port, A_s(33)
                           => SHIFT_3_33_port, A_s(32) => SHIFT_3_32_port, 
                           A_s(31) => SHIFT_3_31_port, A_s(30) => 
                           SHIFT_3_30_port, A_s(29) => SHIFT_3_29_port, A_s(28)
                           => SHIFT_3_28_port, A_s(27) => SHIFT_3_27_port, 
                           A_s(26) => SHIFT_3_26_port, A_s(25) => 
                           SHIFT_3_25_port, A_s(24) => SHIFT_3_24_port, A_s(23)
                           => SHIFT_3_23_port, A_s(22) => SHIFT_3_22_port, 
                           A_s(21) => SHIFT_3_21_port, A_s(20) => 
                           SHIFT_3_20_port, A_s(19) => SHIFT_3_19_port, A_s(18)
                           => SHIFT_3_18_port, A_s(17) => SHIFT_3_17_port, 
                           A_s(16) => SHIFT_3_16_port, A_s(15) => 
                           SHIFT_3_15_port, A_s(14) => SHIFT_3_14_port, A_s(13)
                           => SHIFT_3_13_port, A_s(12) => SHIFT_3_12_port, 
                           A_s(11) => SHIFT_3_11_port, A_s(10) => 
                           SHIFT_3_10_port, A_s(9) => SHIFT_3_9_port, A_s(8) =>
                           SHIFT_3_8_port, A_s(7) => SHIFT_3_7_port, A_s(6) => 
                           SHIFT_3_6_port, A_s(5) => SHIFT_3_5_port, A_s(4) => 
                           SHIFT_3_4_port, A_s(3) => SHIFT_3_3_port, A_s(2) => 
                           SHIFT_3_2_port, A_s(1) => SHIFT_3_1_port, A_s(0) => 
                           SHIFT_3_0_port, A_ns(39) => SHIFT_n_3_37_port, 
                           A_ns(38) => SHIFT_n_3_37_port, A_ns(37) => 
                           SHIFT_n_3_37_port, A_ns(36) => SHIFT_n_3_36_port, 
                           A_ns(35) => SHIFT_n_3_35_port, A_ns(34) => 
                           SHIFT_n_3_34_port, A_ns(33) => SHIFT_n_3_33_port, 
                           A_ns(32) => SHIFT_n_3_32_port, A_ns(31) => 
                           SHIFT_n_3_31_port, A_ns(30) => SHIFT_n_3_30_port, 
                           A_ns(29) => SHIFT_n_3_29_port, A_ns(28) => 
                           SHIFT_n_3_28_port, A_ns(27) => SHIFT_n_3_27_port, 
                           A_ns(26) => SHIFT_n_3_26_port, A_ns(25) => 
                           SHIFT_n_3_25_port, A_ns(24) => SHIFT_n_3_24_port, 
                           A_ns(23) => SHIFT_n_3_23_port, A_ns(22) => 
                           SHIFT_n_3_22_port, A_ns(21) => SHIFT_n_3_21_port, 
                           A_ns(20) => SHIFT_n_3_20_port, A_ns(19) => 
                           SHIFT_n_3_19_port, A_ns(18) => SHIFT_n_3_18_port, 
                           A_ns(17) => SHIFT_n_3_17_port, A_ns(16) => 
                           SHIFT_n_3_16_port, A_ns(15) => SHIFT_n_3_15_port, 
                           A_ns(14) => SHIFT_n_3_14_port, A_ns(13) => 
                           SHIFT_n_3_13_port, A_ns(12) => SHIFT_n_3_12_port, 
                           A_ns(11) => SHIFT_n_3_11_port, A_ns(10) => 
                           SHIFT_n_3_10_port, A_ns(9) => SHIFT_n_3_9_port, 
                           A_ns(8) => SHIFT_n_3_8_port, A_ns(7) => 
                           SHIFT_n_3_7_port, A_ns(6) => SHIFT_n_3_6_port, 
                           A_ns(5) => SHIFT_n_3_5_port, A_ns(4) => 
                           SHIFT_n_3_4_port, A_ns(3) => SHIFT_n_3_3_port, 
                           A_ns(2) => SHIFT_n_3_2_port, A_ns(1) => 
                           SHIFT_n_3_1_port, A_ns(0) => SHIFT_n_3_0_port, B(39)
                           => B(31), B(38) => B(31), B(37) => B(31), B(36) => 
                           B(31), B(35) => B(31), B(34) => B(31), B(33) => 
                           B(31), B(32) => B(31), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), O(39) => OTMP_3_39_port, 
                           O(38) => OTMP_3_38_port, O(37) => OTMP_3_37_port, 
                           O(36) => OTMP_3_36_port, O(35) => OTMP_3_35_port, 
                           O(34) => OTMP_3_34_port, O(33) => OTMP_3_33_port, 
                           O(32) => OTMP_3_32_port, O(31) => OTMP_3_31_port, 
                           O(30) => OTMP_3_30_port, O(29) => OTMP_3_29_port, 
                           O(28) => OTMP_3_28_port, O(27) => OTMP_3_27_port, 
                           O(26) => OTMP_3_26_port, O(25) => OTMP_3_25_port, 
                           O(24) => OTMP_3_24_port, O(23) => OTMP_3_23_port, 
                           O(22) => OTMP_3_22_port, O(21) => OTMP_3_21_port, 
                           O(20) => OTMP_3_20_port, O(19) => OTMP_3_19_port, 
                           O(18) => OTMP_3_18_port, O(17) => OTMP_3_17_port, 
                           O(16) => OTMP_3_16_port, O(15) => OTMP_3_15_port, 
                           O(14) => OTMP_3_14_port, O(13) => OTMP_3_13_port, 
                           O(12) => OTMP_3_12_port, O(11) => OTMP_3_11_port, 
                           O(10) => OTMP_3_10_port, O(9) => OTMP_3_9_port, O(8)
                           => OTMP_3_8_port, O(7) => OTMP_3_7_port, O(6) => 
                           OTMP_3_6_port, O(5) => OTMP_3_5_port, O(4) => 
                           OTMP_3_4_port, O(3) => OTMP_3_3_port, O(2) => 
                           OTMP_3_2_port, O(1) => OTMP_3_1_port, O(0) => n_1092
                           , A_so(39) => SHIFT_4_39_port, A_so(38) => 
                           SHIFT_4_38_port, A_so(37) => SHIFT_4_37_port, 
                           A_so(36) => SHIFT_4_36_port, A_so(35) => 
                           SHIFT_4_35_port, A_so(34) => SHIFT_4_34_port, 
                           A_so(33) => SHIFT_4_33_port, A_so(32) => 
                           SHIFT_4_32_port, A_so(31) => SHIFT_4_31_port, 
                           A_so(30) => SHIFT_4_30_port, A_so(29) => 
                           SHIFT_4_29_port, A_so(28) => SHIFT_4_28_port, 
                           A_so(27) => SHIFT_4_27_port, A_so(26) => 
                           SHIFT_4_26_port, A_so(25) => SHIFT_4_25_port, 
                           A_so(24) => SHIFT_4_24_port, A_so(23) => 
                           SHIFT_4_23_port, A_so(22) => SHIFT_4_22_port, 
                           A_so(21) => SHIFT_4_21_port, A_so(20) => 
                           SHIFT_4_20_port, A_so(19) => SHIFT_4_19_port, 
                           A_so(18) => SHIFT_4_18_port, A_so(17) => 
                           SHIFT_4_17_port, A_so(16) => SHIFT_4_16_port, 
                           A_so(15) => SHIFT_4_15_port, A_so(14) => 
                           SHIFT_4_14_port, A_so(13) => SHIFT_4_13_port, 
                           A_so(12) => SHIFT_4_12_port, A_so(11) => 
                           SHIFT_4_11_port, A_so(10) => SHIFT_4_10_port, 
                           A_so(9) => SHIFT_4_9_port, A_so(8) => SHIFT_4_8_port
                           , A_so(7) => SHIFT_4_7_port, A_so(6) => 
                           SHIFT_4_6_port, A_so(5) => SHIFT_4_5_port, A_so(4) 
                           => SHIFT_4_4_port, A_so(3) => SHIFT_4_3_port, 
                           A_so(2) => SHIFT_4_2_port, A_so(1) => n_1093, 
                           A_so(0) => n_1094, A_nso(39) => SHIFT_n_4_39_port, 
                           A_nso(38) => SHIFT_n_4_38_port, A_nso(37) => 
                           SHIFT_n_4_37_port, A_nso(36) => SHIFT_n_4_36_port, 
                           A_nso(35) => SHIFT_n_4_35_port, A_nso(34) => 
                           SHIFT_n_4_34_port, A_nso(33) => SHIFT_n_4_33_port, 
                           A_nso(32) => SHIFT_n_4_32_port, A_nso(31) => 
                           SHIFT_n_4_31_port, A_nso(30) => SHIFT_n_4_30_port, 
                           A_nso(29) => SHIFT_n_4_29_port, A_nso(28) => 
                           SHIFT_n_4_28_port, A_nso(27) => SHIFT_n_4_27_port, 
                           A_nso(26) => SHIFT_n_4_26_port, A_nso(25) => 
                           SHIFT_n_4_25_port, A_nso(24) => SHIFT_n_4_24_port, 
                           A_nso(23) => SHIFT_n_4_23_port, A_nso(22) => 
                           SHIFT_n_4_22_port, A_nso(21) => SHIFT_n_4_21_port, 
                           A_nso(20) => SHIFT_n_4_20_port, A_nso(19) => 
                           SHIFT_n_4_19_port, A_nso(18) => SHIFT_n_4_18_port, 
                           A_nso(17) => SHIFT_n_4_17_port, A_nso(16) => 
                           SHIFT_n_4_16_port, A_nso(15) => SHIFT_n_4_15_port, 
                           A_nso(14) => SHIFT_n_4_14_port, A_nso(13) => 
                           SHIFT_n_4_13_port, A_nso(12) => SHIFT_n_4_12_port, 
                           A_nso(11) => SHIFT_n_4_11_port, A_nso(10) => 
                           SHIFT_n_4_10_port, A_nso(9) => SHIFT_n_4_9_port, 
                           A_nso(8) => SHIFT_n_4_8_port, A_nso(7) => 
                           SHIFT_n_4_7_port, A_nso(6) => SHIFT_n_4_6_port, 
                           A_nso(5) => SHIFT_n_4_5_port, A_nso(4) => 
                           SHIFT_n_4_4_port, A_nso(3) => SHIFT_n_4_3_port, 
                           A_nso(2) => SHIFT_n_4_2_port, A_nso(1) => n_1095, 
                           A_nso(0) => n_1096);
   ENC_4 : BOOTHENC_NBIT42_i8 port map( A_s(41) => SHIFT_4_39_port, A_s(40) => 
                           SHIFT_4_39_port, A_s(39) => SHIFT_4_39_port, A_s(38)
                           => SHIFT_4_38_port, A_s(37) => SHIFT_4_37_port, 
                           A_s(36) => SHIFT_4_36_port, A_s(35) => 
                           SHIFT_4_35_port, A_s(34) => SHIFT_4_34_port, A_s(33)
                           => SHIFT_4_33_port, A_s(32) => SHIFT_4_32_port, 
                           A_s(31) => SHIFT_4_31_port, A_s(30) => 
                           SHIFT_4_30_port, A_s(29) => SHIFT_4_29_port, A_s(28)
                           => SHIFT_4_28_port, A_s(27) => SHIFT_4_27_port, 
                           A_s(26) => SHIFT_4_26_port, A_s(25) => 
                           SHIFT_4_25_port, A_s(24) => SHIFT_4_24_port, A_s(23)
                           => SHIFT_4_23_port, A_s(22) => SHIFT_4_22_port, 
                           A_s(21) => SHIFT_4_21_port, A_s(20) => 
                           SHIFT_4_20_port, A_s(19) => SHIFT_4_19_port, A_s(18)
                           => SHIFT_4_18_port, A_s(17) => SHIFT_4_17_port, 
                           A_s(16) => SHIFT_4_16_port, A_s(15) => 
                           SHIFT_4_15_port, A_s(14) => SHIFT_4_14_port, A_s(13)
                           => SHIFT_4_13_port, A_s(12) => SHIFT_4_12_port, 
                           A_s(11) => SHIFT_4_11_port, A_s(10) => 
                           SHIFT_4_10_port, A_s(9) => SHIFT_4_9_port, A_s(8) =>
                           SHIFT_4_8_port, A_s(7) => SHIFT_4_7_port, A_s(6) => 
                           SHIFT_4_6_port, A_s(5) => SHIFT_4_5_port, A_s(4) => 
                           SHIFT_4_4_port, A_s(3) => SHIFT_4_3_port, A_s(2) => 
                           SHIFT_4_2_port, A_s(1) => SHIFT_4_1_port, A_s(0) => 
                           SHIFT_4_0_port, A_ns(41) => SHIFT_n_4_39_port, 
                           A_ns(40) => SHIFT_n_4_39_port, A_ns(39) => 
                           SHIFT_n_4_39_port, A_ns(38) => SHIFT_n_4_38_port, 
                           A_ns(37) => SHIFT_n_4_37_port, A_ns(36) => 
                           SHIFT_n_4_36_port, A_ns(35) => SHIFT_n_4_35_port, 
                           A_ns(34) => SHIFT_n_4_34_port, A_ns(33) => 
                           SHIFT_n_4_33_port, A_ns(32) => SHIFT_n_4_32_port, 
                           A_ns(31) => SHIFT_n_4_31_port, A_ns(30) => 
                           SHIFT_n_4_30_port, A_ns(29) => SHIFT_n_4_29_port, 
                           A_ns(28) => SHIFT_n_4_28_port, A_ns(27) => 
                           SHIFT_n_4_27_port, A_ns(26) => SHIFT_n_4_26_port, 
                           A_ns(25) => SHIFT_n_4_25_port, A_ns(24) => 
                           SHIFT_n_4_24_port, A_ns(23) => SHIFT_n_4_23_port, 
                           A_ns(22) => SHIFT_n_4_22_port, A_ns(21) => 
                           SHIFT_n_4_21_port, A_ns(20) => SHIFT_n_4_20_port, 
                           A_ns(19) => SHIFT_n_4_19_port, A_ns(18) => 
                           SHIFT_n_4_18_port, A_ns(17) => SHIFT_n_4_17_port, 
                           A_ns(16) => SHIFT_n_4_16_port, A_ns(15) => 
                           SHIFT_n_4_15_port, A_ns(14) => SHIFT_n_4_14_port, 
                           A_ns(13) => SHIFT_n_4_13_port, A_ns(12) => 
                           SHIFT_n_4_12_port, A_ns(11) => SHIFT_n_4_11_port, 
                           A_ns(10) => SHIFT_n_4_10_port, A_ns(9) => 
                           SHIFT_n_4_9_port, A_ns(8) => SHIFT_n_4_8_port, 
                           A_ns(7) => SHIFT_n_4_7_port, A_ns(6) => 
                           SHIFT_n_4_6_port, A_ns(5) => SHIFT_n_4_5_port, 
                           A_ns(4) => SHIFT_n_4_4_port, A_ns(3) => 
                           SHIFT_n_4_3_port, A_ns(2) => SHIFT_n_4_2_port, 
                           A_ns(1) => SHIFT_n_4_1_port, A_ns(0) => 
                           SHIFT_n_4_0_port, B(41) => B(31), B(40) => B(31), 
                           B(39) => B(31), B(38) => B(31), B(37) => B(31), 
                           B(36) => B(31), B(35) => B(31), B(34) => B(31), 
                           B(33) => B(31), B(32) => B(31), B(31) => B(31), 
                           B(30) => B(30), B(29) => B(29), B(28) => B(28), 
                           B(27) => B(27), B(26) => B(26), B(25) => B(25), 
                           B(24) => B(24), B(23) => B(23), B(22) => B(22), 
                           B(21) => B(21), B(20) => B(20), B(19) => B(19), 
                           B(18) => B(18), B(17) => B(17), B(16) => B(16), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => B(0), O(41) => 
                           OTMP_4_41_port, O(40) => OTMP_4_40_port, O(39) => 
                           OTMP_4_39_port, O(38) => OTMP_4_38_port, O(37) => 
                           OTMP_4_37_port, O(36) => OTMP_4_36_port, O(35) => 
                           OTMP_4_35_port, O(34) => OTMP_4_34_port, O(33) => 
                           OTMP_4_33_port, O(32) => OTMP_4_32_port, O(31) => 
                           OTMP_4_31_port, O(30) => OTMP_4_30_port, O(29) => 
                           OTMP_4_29_port, O(28) => OTMP_4_28_port, O(27) => 
                           OTMP_4_27_port, O(26) => OTMP_4_26_port, O(25) => 
                           OTMP_4_25_port, O(24) => OTMP_4_24_port, O(23) => 
                           OTMP_4_23_port, O(22) => OTMP_4_22_port, O(21) => 
                           OTMP_4_21_port, O(20) => OTMP_4_20_port, O(19) => 
                           OTMP_4_19_port, O(18) => OTMP_4_18_port, O(17) => 
                           OTMP_4_17_port, O(16) => OTMP_4_16_port, O(15) => 
                           OTMP_4_15_port, O(14) => OTMP_4_14_port, O(13) => 
                           OTMP_4_13_port, O(12) => OTMP_4_12_port, O(11) => 
                           OTMP_4_11_port, O(10) => OTMP_4_10_port, O(9) => 
                           OTMP_4_9_port, O(8) => OTMP_4_8_port, O(7) => 
                           OTMP_4_7_port, O(6) => OTMP_4_6_port, O(5) => 
                           OTMP_4_5_port, O(4) => OTMP_4_4_port, O(3) => 
                           OTMP_4_3_port, O(2) => OTMP_4_2_port, O(1) => 
                           OTMP_4_1_port, O(0) => n_1097, A_so(41) => 
                           SHIFT_5_41_port, A_so(40) => SHIFT_5_40_port, 
                           A_so(39) => SHIFT_5_39_port, A_so(38) => 
                           SHIFT_5_38_port, A_so(37) => SHIFT_5_37_port, 
                           A_so(36) => SHIFT_5_36_port, A_so(35) => 
                           SHIFT_5_35_port, A_so(34) => SHIFT_5_34_port, 
                           A_so(33) => SHIFT_5_33_port, A_so(32) => 
                           SHIFT_5_32_port, A_so(31) => SHIFT_5_31_port, 
                           A_so(30) => SHIFT_5_30_port, A_so(29) => 
                           SHIFT_5_29_port, A_so(28) => SHIFT_5_28_port, 
                           A_so(27) => SHIFT_5_27_port, A_so(26) => 
                           SHIFT_5_26_port, A_so(25) => SHIFT_5_25_port, 
                           A_so(24) => SHIFT_5_24_port, A_so(23) => 
                           SHIFT_5_23_port, A_so(22) => SHIFT_5_22_port, 
                           A_so(21) => SHIFT_5_21_port, A_so(20) => 
                           SHIFT_5_20_port, A_so(19) => SHIFT_5_19_port, 
                           A_so(18) => SHIFT_5_18_port, A_so(17) => 
                           SHIFT_5_17_port, A_so(16) => SHIFT_5_16_port, 
                           A_so(15) => SHIFT_5_15_port, A_so(14) => 
                           SHIFT_5_14_port, A_so(13) => SHIFT_5_13_port, 
                           A_so(12) => SHIFT_5_12_port, A_so(11) => 
                           SHIFT_5_11_port, A_so(10) => SHIFT_5_10_port, 
                           A_so(9) => SHIFT_5_9_port, A_so(8) => SHIFT_5_8_port
                           , A_so(7) => SHIFT_5_7_port, A_so(6) => 
                           SHIFT_5_6_port, A_so(5) => SHIFT_5_5_port, A_so(4) 
                           => SHIFT_5_4_port, A_so(3) => SHIFT_5_3_port, 
                           A_so(2) => SHIFT_5_2_port, A_so(1) => n_1098, 
                           A_so(0) => n_1099, A_nso(41) => SHIFT_n_5_41_port, 
                           A_nso(40) => SHIFT_n_5_40_port, A_nso(39) => 
                           SHIFT_n_5_39_port, A_nso(38) => SHIFT_n_5_38_port, 
                           A_nso(37) => SHIFT_n_5_37_port, A_nso(36) => 
                           SHIFT_n_5_36_port, A_nso(35) => SHIFT_n_5_35_port, 
                           A_nso(34) => SHIFT_n_5_34_port, A_nso(33) => 
                           SHIFT_n_5_33_port, A_nso(32) => SHIFT_n_5_32_port, 
                           A_nso(31) => SHIFT_n_5_31_port, A_nso(30) => 
                           SHIFT_n_5_30_port, A_nso(29) => SHIFT_n_5_29_port, 
                           A_nso(28) => SHIFT_n_5_28_port, A_nso(27) => 
                           SHIFT_n_5_27_port, A_nso(26) => SHIFT_n_5_26_port, 
                           A_nso(25) => SHIFT_n_5_25_port, A_nso(24) => 
                           SHIFT_n_5_24_port, A_nso(23) => SHIFT_n_5_23_port, 
                           A_nso(22) => SHIFT_n_5_22_port, A_nso(21) => 
                           SHIFT_n_5_21_port, A_nso(20) => SHIFT_n_5_20_port, 
                           A_nso(19) => SHIFT_n_5_19_port, A_nso(18) => 
                           SHIFT_n_5_18_port, A_nso(17) => SHIFT_n_5_17_port, 
                           A_nso(16) => SHIFT_n_5_16_port, A_nso(15) => 
                           SHIFT_n_5_15_port, A_nso(14) => SHIFT_n_5_14_port, 
                           A_nso(13) => SHIFT_n_5_13_port, A_nso(12) => 
                           SHIFT_n_5_12_port, A_nso(11) => SHIFT_n_5_11_port, 
                           A_nso(10) => SHIFT_n_5_10_port, A_nso(9) => 
                           SHIFT_n_5_9_port, A_nso(8) => SHIFT_n_5_8_port, 
                           A_nso(7) => SHIFT_n_5_7_port, A_nso(6) => 
                           SHIFT_n_5_6_port, A_nso(5) => SHIFT_n_5_5_port, 
                           A_nso(4) => SHIFT_n_5_4_port, A_nso(3) => 
                           SHIFT_n_5_3_port, A_nso(2) => SHIFT_n_5_2_port, 
                           A_nso(1) => n_1100, A_nso(0) => n_1101);
   ENC_5 : BOOTHENC_NBIT44_i10 port map( A_s(43) => SHIFT_5_41_port, A_s(42) =>
                           SHIFT_5_41_port, A_s(41) => SHIFT_5_41_port, A_s(40)
                           => SHIFT_5_40_port, A_s(39) => SHIFT_5_39_port, 
                           A_s(38) => SHIFT_5_38_port, A_s(37) => 
                           SHIFT_5_37_port, A_s(36) => SHIFT_5_36_port, A_s(35)
                           => SHIFT_5_35_port, A_s(34) => SHIFT_5_34_port, 
                           A_s(33) => SHIFT_5_33_port, A_s(32) => 
                           SHIFT_5_32_port, A_s(31) => SHIFT_5_31_port, A_s(30)
                           => SHIFT_5_30_port, A_s(29) => SHIFT_5_29_port, 
                           A_s(28) => SHIFT_5_28_port, A_s(27) => 
                           SHIFT_5_27_port, A_s(26) => SHIFT_5_26_port, A_s(25)
                           => SHIFT_5_25_port, A_s(24) => SHIFT_5_24_port, 
                           A_s(23) => SHIFT_5_23_port, A_s(22) => 
                           SHIFT_5_22_port, A_s(21) => SHIFT_5_21_port, A_s(20)
                           => SHIFT_5_20_port, A_s(19) => SHIFT_5_19_port, 
                           A_s(18) => SHIFT_5_18_port, A_s(17) => 
                           SHIFT_5_17_port, A_s(16) => SHIFT_5_16_port, A_s(15)
                           => SHIFT_5_15_port, A_s(14) => SHIFT_5_14_port, 
                           A_s(13) => SHIFT_5_13_port, A_s(12) => 
                           SHIFT_5_12_port, A_s(11) => SHIFT_5_11_port, A_s(10)
                           => SHIFT_5_10_port, A_s(9) => SHIFT_5_9_port, A_s(8)
                           => SHIFT_5_8_port, A_s(7) => SHIFT_5_7_port, A_s(6) 
                           => SHIFT_5_6_port, A_s(5) => SHIFT_5_5_port, A_s(4) 
                           => SHIFT_5_4_port, A_s(3) => SHIFT_5_3_port, A_s(2) 
                           => SHIFT_5_2_port, A_s(1) => SHIFT_5_1_port, A_s(0) 
                           => SHIFT_5_0_port, A_ns(43) => SHIFT_n_5_41_port, 
                           A_ns(42) => SHIFT_n_5_41_port, A_ns(41) => 
                           SHIFT_n_5_41_port, A_ns(40) => SHIFT_n_5_40_port, 
                           A_ns(39) => SHIFT_n_5_39_port, A_ns(38) => 
                           SHIFT_n_5_38_port, A_ns(37) => SHIFT_n_5_37_port, 
                           A_ns(36) => SHIFT_n_5_36_port, A_ns(35) => 
                           SHIFT_n_5_35_port, A_ns(34) => SHIFT_n_5_34_port, 
                           A_ns(33) => SHIFT_n_5_33_port, A_ns(32) => 
                           SHIFT_n_5_32_port, A_ns(31) => SHIFT_n_5_31_port, 
                           A_ns(30) => SHIFT_n_5_30_port, A_ns(29) => 
                           SHIFT_n_5_29_port, A_ns(28) => SHIFT_n_5_28_port, 
                           A_ns(27) => SHIFT_n_5_27_port, A_ns(26) => 
                           SHIFT_n_5_26_port, A_ns(25) => SHIFT_n_5_25_port, 
                           A_ns(24) => SHIFT_n_5_24_port, A_ns(23) => 
                           SHIFT_n_5_23_port, A_ns(22) => SHIFT_n_5_22_port, 
                           A_ns(21) => SHIFT_n_5_21_port, A_ns(20) => 
                           SHIFT_n_5_20_port, A_ns(19) => SHIFT_n_5_19_port, 
                           A_ns(18) => SHIFT_n_5_18_port, A_ns(17) => 
                           SHIFT_n_5_17_port, A_ns(16) => SHIFT_n_5_16_port, 
                           A_ns(15) => SHIFT_n_5_15_port, A_ns(14) => 
                           SHIFT_n_5_14_port, A_ns(13) => SHIFT_n_5_13_port, 
                           A_ns(12) => SHIFT_n_5_12_port, A_ns(11) => 
                           SHIFT_n_5_11_port, A_ns(10) => SHIFT_n_5_10_port, 
                           A_ns(9) => SHIFT_n_5_9_port, A_ns(8) => 
                           SHIFT_n_5_8_port, A_ns(7) => SHIFT_n_5_7_port, 
                           A_ns(6) => SHIFT_n_5_6_port, A_ns(5) => 
                           SHIFT_n_5_5_port, A_ns(4) => SHIFT_n_5_4_port, 
                           A_ns(3) => SHIFT_n_5_3_port, A_ns(2) => 
                           SHIFT_n_5_2_port, A_ns(1) => SHIFT_n_5_1_port, 
                           A_ns(0) => SHIFT_n_5_0_port, B(43) => B(31), B(42) 
                           => B(31), B(41) => B(31), B(40) => B(31), B(39) => 
                           B(31), B(38) => B(31), B(37) => B(31), B(36) => 
                           B(31), B(35) => B(31), B(34) => B(31), B(33) => 
                           B(31), B(32) => B(31), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), O(43) => OTMP_5_43_port, 
                           O(42) => OTMP_5_42_port, O(41) => OTMP_5_41_port, 
                           O(40) => OTMP_5_40_port, O(39) => OTMP_5_39_port, 
                           O(38) => OTMP_5_38_port, O(37) => OTMP_5_37_port, 
                           O(36) => OTMP_5_36_port, O(35) => OTMP_5_35_port, 
                           O(34) => OTMP_5_34_port, O(33) => OTMP_5_33_port, 
                           O(32) => OTMP_5_32_port, O(31) => OTMP_5_31_port, 
                           O(30) => OTMP_5_30_port, O(29) => OTMP_5_29_port, 
                           O(28) => OTMP_5_28_port, O(27) => OTMP_5_27_port, 
                           O(26) => OTMP_5_26_port, O(25) => OTMP_5_25_port, 
                           O(24) => OTMP_5_24_port, O(23) => OTMP_5_23_port, 
                           O(22) => OTMP_5_22_port, O(21) => OTMP_5_21_port, 
                           O(20) => OTMP_5_20_port, O(19) => OTMP_5_19_port, 
                           O(18) => OTMP_5_18_port, O(17) => OTMP_5_17_port, 
                           O(16) => OTMP_5_16_port, O(15) => OTMP_5_15_port, 
                           O(14) => OTMP_5_14_port, O(13) => OTMP_5_13_port, 
                           O(12) => OTMP_5_12_port, O(11) => OTMP_5_11_port, 
                           O(10) => OTMP_5_10_port, O(9) => OTMP_5_9_port, O(8)
                           => OTMP_5_8_port, O(7) => OTMP_5_7_port, O(6) => 
                           OTMP_5_6_port, O(5) => OTMP_5_5_port, O(4) => 
                           OTMP_5_4_port, O(3) => OTMP_5_3_port, O(2) => 
                           OTMP_5_2_port, O(1) => OTMP_5_1_port, O(0) => n_1102
                           , A_so(43) => SHIFT_6_43_port, A_so(42) => 
                           SHIFT_6_42_port, A_so(41) => SHIFT_6_41_port, 
                           A_so(40) => SHIFT_6_40_port, A_so(39) => 
                           SHIFT_6_39_port, A_so(38) => SHIFT_6_38_port, 
                           A_so(37) => SHIFT_6_37_port, A_so(36) => 
                           SHIFT_6_36_port, A_so(35) => SHIFT_6_35_port, 
                           A_so(34) => SHIFT_6_34_port, A_so(33) => 
                           SHIFT_6_33_port, A_so(32) => SHIFT_6_32_port, 
                           A_so(31) => SHIFT_6_31_port, A_so(30) => 
                           SHIFT_6_30_port, A_so(29) => SHIFT_6_29_port, 
                           A_so(28) => SHIFT_6_28_port, A_so(27) => 
                           SHIFT_6_27_port, A_so(26) => SHIFT_6_26_port, 
                           A_so(25) => SHIFT_6_25_port, A_so(24) => 
                           SHIFT_6_24_port, A_so(23) => SHIFT_6_23_port, 
                           A_so(22) => SHIFT_6_22_port, A_so(21) => 
                           SHIFT_6_21_port, A_so(20) => SHIFT_6_20_port, 
                           A_so(19) => SHIFT_6_19_port, A_so(18) => 
                           SHIFT_6_18_port, A_so(17) => SHIFT_6_17_port, 
                           A_so(16) => SHIFT_6_16_port, A_so(15) => 
                           SHIFT_6_15_port, A_so(14) => SHIFT_6_14_port, 
                           A_so(13) => SHIFT_6_13_port, A_so(12) => 
                           SHIFT_6_12_port, A_so(11) => SHIFT_6_11_port, 
                           A_so(10) => SHIFT_6_10_port, A_so(9) => 
                           SHIFT_6_9_port, A_so(8) => SHIFT_6_8_port, A_so(7) 
                           => SHIFT_6_7_port, A_so(6) => SHIFT_6_6_port, 
                           A_so(5) => SHIFT_6_5_port, A_so(4) => SHIFT_6_4_port
                           , A_so(3) => SHIFT_6_3_port, A_so(2) => 
                           SHIFT_6_2_port, A_so(1) => n_1103, A_so(0) => n_1104
                           , A_nso(43) => SHIFT_n_6_43_port, A_nso(42) => 
                           SHIFT_n_6_42_port, A_nso(41) => SHIFT_n_6_41_port, 
                           A_nso(40) => SHIFT_n_6_40_port, A_nso(39) => 
                           SHIFT_n_6_39_port, A_nso(38) => SHIFT_n_6_38_port, 
                           A_nso(37) => SHIFT_n_6_37_port, A_nso(36) => 
                           SHIFT_n_6_36_port, A_nso(35) => SHIFT_n_6_35_port, 
                           A_nso(34) => SHIFT_n_6_34_port, A_nso(33) => 
                           SHIFT_n_6_33_port, A_nso(32) => SHIFT_n_6_32_port, 
                           A_nso(31) => SHIFT_n_6_31_port, A_nso(30) => 
                           SHIFT_n_6_30_port, A_nso(29) => SHIFT_n_6_29_port, 
                           A_nso(28) => SHIFT_n_6_28_port, A_nso(27) => 
                           SHIFT_n_6_27_port, A_nso(26) => SHIFT_n_6_26_port, 
                           A_nso(25) => SHIFT_n_6_25_port, A_nso(24) => 
                           SHIFT_n_6_24_port, A_nso(23) => SHIFT_n_6_23_port, 
                           A_nso(22) => SHIFT_n_6_22_port, A_nso(21) => 
                           SHIFT_n_6_21_port, A_nso(20) => SHIFT_n_6_20_port, 
                           A_nso(19) => SHIFT_n_6_19_port, A_nso(18) => 
                           SHIFT_n_6_18_port, A_nso(17) => SHIFT_n_6_17_port, 
                           A_nso(16) => SHIFT_n_6_16_port, A_nso(15) => 
                           SHIFT_n_6_15_port, A_nso(14) => SHIFT_n_6_14_port, 
                           A_nso(13) => SHIFT_n_6_13_port, A_nso(12) => 
                           SHIFT_n_6_12_port, A_nso(11) => SHIFT_n_6_11_port, 
                           A_nso(10) => SHIFT_n_6_10_port, A_nso(9) => 
                           SHIFT_n_6_9_port, A_nso(8) => SHIFT_n_6_8_port, 
                           A_nso(7) => SHIFT_n_6_7_port, A_nso(6) => 
                           SHIFT_n_6_6_port, A_nso(5) => SHIFT_n_6_5_port, 
                           A_nso(4) => SHIFT_n_6_4_port, A_nso(3) => 
                           SHIFT_n_6_3_port, A_nso(2) => SHIFT_n_6_2_port, 
                           A_nso(1) => n_1105, A_nso(0) => n_1106);
   ENC_6 : BOOTHENC_NBIT46_i12 port map( A_s(45) => SHIFT_6_43_port, A_s(44) =>
                           SHIFT_6_43_port, A_s(43) => SHIFT_6_43_port, A_s(42)
                           => SHIFT_6_42_port, A_s(41) => SHIFT_6_41_port, 
                           A_s(40) => SHIFT_6_40_port, A_s(39) => 
                           SHIFT_6_39_port, A_s(38) => SHIFT_6_38_port, A_s(37)
                           => SHIFT_6_37_port, A_s(36) => SHIFT_6_36_port, 
                           A_s(35) => SHIFT_6_35_port, A_s(34) => 
                           SHIFT_6_34_port, A_s(33) => SHIFT_6_33_port, A_s(32)
                           => SHIFT_6_32_port, A_s(31) => SHIFT_6_31_port, 
                           A_s(30) => SHIFT_6_30_port, A_s(29) => 
                           SHIFT_6_29_port, A_s(28) => SHIFT_6_28_port, A_s(27)
                           => SHIFT_6_27_port, A_s(26) => SHIFT_6_26_port, 
                           A_s(25) => SHIFT_6_25_port, A_s(24) => 
                           SHIFT_6_24_port, A_s(23) => SHIFT_6_23_port, A_s(22)
                           => SHIFT_6_22_port, A_s(21) => SHIFT_6_21_port, 
                           A_s(20) => SHIFT_6_20_port, A_s(19) => 
                           SHIFT_6_19_port, A_s(18) => SHIFT_6_18_port, A_s(17)
                           => SHIFT_6_17_port, A_s(16) => SHIFT_6_16_port, 
                           A_s(15) => SHIFT_6_15_port, A_s(14) => 
                           SHIFT_6_14_port, A_s(13) => SHIFT_6_13_port, A_s(12)
                           => SHIFT_6_12_port, A_s(11) => SHIFT_6_11_port, 
                           A_s(10) => SHIFT_6_10_port, A_s(9) => SHIFT_6_9_port
                           , A_s(8) => SHIFT_6_8_port, A_s(7) => SHIFT_6_7_port
                           , A_s(6) => SHIFT_6_6_port, A_s(5) => SHIFT_6_5_port
                           , A_s(4) => SHIFT_6_4_port, A_s(3) => SHIFT_6_3_port
                           , A_s(2) => SHIFT_6_2_port, A_s(1) => SHIFT_6_1_port
                           , A_s(0) => SHIFT_6_0_port, A_ns(45) => 
                           SHIFT_n_6_43_port, A_ns(44) => SHIFT_n_6_43_port, 
                           A_ns(43) => SHIFT_n_6_43_port, A_ns(42) => 
                           SHIFT_n_6_42_port, A_ns(41) => SHIFT_n_6_41_port, 
                           A_ns(40) => SHIFT_n_6_40_port, A_ns(39) => 
                           SHIFT_n_6_39_port, A_ns(38) => SHIFT_n_6_38_port, 
                           A_ns(37) => SHIFT_n_6_37_port, A_ns(36) => 
                           SHIFT_n_6_36_port, A_ns(35) => SHIFT_n_6_35_port, 
                           A_ns(34) => SHIFT_n_6_34_port, A_ns(33) => 
                           SHIFT_n_6_33_port, A_ns(32) => SHIFT_n_6_32_port, 
                           A_ns(31) => SHIFT_n_6_31_port, A_ns(30) => 
                           SHIFT_n_6_30_port, A_ns(29) => SHIFT_n_6_29_port, 
                           A_ns(28) => SHIFT_n_6_28_port, A_ns(27) => 
                           SHIFT_n_6_27_port, A_ns(26) => SHIFT_n_6_26_port, 
                           A_ns(25) => SHIFT_n_6_25_port, A_ns(24) => 
                           SHIFT_n_6_24_port, A_ns(23) => SHIFT_n_6_23_port, 
                           A_ns(22) => SHIFT_n_6_22_port, A_ns(21) => 
                           SHIFT_n_6_21_port, A_ns(20) => SHIFT_n_6_20_port, 
                           A_ns(19) => SHIFT_n_6_19_port, A_ns(18) => 
                           SHIFT_n_6_18_port, A_ns(17) => SHIFT_n_6_17_port, 
                           A_ns(16) => SHIFT_n_6_16_port, A_ns(15) => 
                           SHIFT_n_6_15_port, A_ns(14) => SHIFT_n_6_14_port, 
                           A_ns(13) => SHIFT_n_6_13_port, A_ns(12) => 
                           SHIFT_n_6_12_port, A_ns(11) => SHIFT_n_6_11_port, 
                           A_ns(10) => SHIFT_n_6_10_port, A_ns(9) => 
                           SHIFT_n_6_9_port, A_ns(8) => SHIFT_n_6_8_port, 
                           A_ns(7) => SHIFT_n_6_7_port, A_ns(6) => 
                           SHIFT_n_6_6_port, A_ns(5) => SHIFT_n_6_5_port, 
                           A_ns(4) => SHIFT_n_6_4_port, A_ns(3) => 
                           SHIFT_n_6_3_port, A_ns(2) => SHIFT_n_6_2_port, 
                           A_ns(1) => SHIFT_n_6_1_port, A_ns(0) => 
                           SHIFT_n_6_0_port, B(45) => B(31), B(44) => B(31), 
                           B(43) => B(31), B(42) => B(31), B(41) => B(31), 
                           B(40) => B(31), B(39) => B(31), B(38) => B(31), 
                           B(37) => B(31), B(36) => B(31), B(35) => B(31), 
                           B(34) => B(31), B(33) => B(31), B(32) => B(31), 
                           B(31) => B(31), B(30) => B(30), B(29) => B(29), 
                           B(28) => B(28), B(27) => B(27), B(26) => B(26), 
                           B(25) => B(25), B(24) => B(24), B(23) => B(23), 
                           B(22) => B(22), B(21) => B(21), B(20) => B(20), 
                           B(19) => B(19), B(18) => B(18), B(17) => B(17), 
                           B(16) => B(16), B(15) => B(15), B(14) => B(14), 
                           B(13) => B(13), B(12) => B(12), B(11) => B(11), 
                           B(10) => B(10), B(9) => B(9), B(8) => B(8), B(7) => 
                           B(7), B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3)
                           => B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), 
                           O(45) => OTMP_6_45_port, O(44) => OTMP_6_44_port, 
                           O(43) => OTMP_6_43_port, O(42) => OTMP_6_42_port, 
                           O(41) => OTMP_6_41_port, O(40) => OTMP_6_40_port, 
                           O(39) => OTMP_6_39_port, O(38) => OTMP_6_38_port, 
                           O(37) => OTMP_6_37_port, O(36) => OTMP_6_36_port, 
                           O(35) => OTMP_6_35_port, O(34) => OTMP_6_34_port, 
                           O(33) => OTMP_6_33_port, O(32) => OTMP_6_32_port, 
                           O(31) => OTMP_6_31_port, O(30) => OTMP_6_30_port, 
                           O(29) => OTMP_6_29_port, O(28) => OTMP_6_28_port, 
                           O(27) => OTMP_6_27_port, O(26) => OTMP_6_26_port, 
                           O(25) => OTMP_6_25_port, O(24) => OTMP_6_24_port, 
                           O(23) => OTMP_6_23_port, O(22) => OTMP_6_22_port, 
                           O(21) => OTMP_6_21_port, O(20) => OTMP_6_20_port, 
                           O(19) => OTMP_6_19_port, O(18) => OTMP_6_18_port, 
                           O(17) => OTMP_6_17_port, O(16) => OTMP_6_16_port, 
                           O(15) => OTMP_6_15_port, O(14) => OTMP_6_14_port, 
                           O(13) => OTMP_6_13_port, O(12) => OTMP_6_12_port, 
                           O(11) => OTMP_6_11_port, O(10) => OTMP_6_10_port, 
                           O(9) => OTMP_6_9_port, O(8) => OTMP_6_8_port, O(7) 
                           => OTMP_6_7_port, O(6) => OTMP_6_6_port, O(5) => 
                           OTMP_6_5_port, O(4) => OTMP_6_4_port, O(3) => 
                           OTMP_6_3_port, O(2) => OTMP_6_2_port, O(1) => 
                           OTMP_6_1_port, O(0) => n_1107, A_so(45) => 
                           SHIFT_7_45_port, A_so(44) => SHIFT_7_44_port, 
                           A_so(43) => SHIFT_7_43_port, A_so(42) => 
                           SHIFT_7_42_port, A_so(41) => SHIFT_7_41_port, 
                           A_so(40) => SHIFT_7_40_port, A_so(39) => 
                           SHIFT_7_39_port, A_so(38) => SHIFT_7_38_port, 
                           A_so(37) => SHIFT_7_37_port, A_so(36) => 
                           SHIFT_7_36_port, A_so(35) => SHIFT_7_35_port, 
                           A_so(34) => SHIFT_7_34_port, A_so(33) => 
                           SHIFT_7_33_port, A_so(32) => SHIFT_7_32_port, 
                           A_so(31) => SHIFT_7_31_port, A_so(30) => 
                           SHIFT_7_30_port, A_so(29) => SHIFT_7_29_port, 
                           A_so(28) => SHIFT_7_28_port, A_so(27) => 
                           SHIFT_7_27_port, A_so(26) => SHIFT_7_26_port, 
                           A_so(25) => SHIFT_7_25_port, A_so(24) => 
                           SHIFT_7_24_port, A_so(23) => SHIFT_7_23_port, 
                           A_so(22) => SHIFT_7_22_port, A_so(21) => 
                           SHIFT_7_21_port, A_so(20) => SHIFT_7_20_port, 
                           A_so(19) => SHIFT_7_19_port, A_so(18) => 
                           SHIFT_7_18_port, A_so(17) => SHIFT_7_17_port, 
                           A_so(16) => SHIFT_7_16_port, A_so(15) => 
                           SHIFT_7_15_port, A_so(14) => SHIFT_7_14_port, 
                           A_so(13) => SHIFT_7_13_port, A_so(12) => 
                           SHIFT_7_12_port, A_so(11) => SHIFT_7_11_port, 
                           A_so(10) => SHIFT_7_10_port, A_so(9) => 
                           SHIFT_7_9_port, A_so(8) => SHIFT_7_8_port, A_so(7) 
                           => SHIFT_7_7_port, A_so(6) => SHIFT_7_6_port, 
                           A_so(5) => SHIFT_7_5_port, A_so(4) => SHIFT_7_4_port
                           , A_so(3) => SHIFT_7_3_port, A_so(2) => 
                           SHIFT_7_2_port, A_so(1) => n_1108, A_so(0) => n_1109
                           , A_nso(45) => SHIFT_n_7_45_port, A_nso(44) => 
                           SHIFT_n_7_44_port, A_nso(43) => SHIFT_n_7_43_port, 
                           A_nso(42) => SHIFT_n_7_42_port, A_nso(41) => 
                           SHIFT_n_7_41_port, A_nso(40) => SHIFT_n_7_40_port, 
                           A_nso(39) => SHIFT_n_7_39_port, A_nso(38) => 
                           SHIFT_n_7_38_port, A_nso(37) => SHIFT_n_7_37_port, 
                           A_nso(36) => SHIFT_n_7_36_port, A_nso(35) => 
                           SHIFT_n_7_35_port, A_nso(34) => SHIFT_n_7_34_port, 
                           A_nso(33) => SHIFT_n_7_33_port, A_nso(32) => 
                           SHIFT_n_7_32_port, A_nso(31) => SHIFT_n_7_31_port, 
                           A_nso(30) => SHIFT_n_7_30_port, A_nso(29) => 
                           SHIFT_n_7_29_port, A_nso(28) => SHIFT_n_7_28_port, 
                           A_nso(27) => SHIFT_n_7_27_port, A_nso(26) => 
                           SHIFT_n_7_26_port, A_nso(25) => SHIFT_n_7_25_port, 
                           A_nso(24) => SHIFT_n_7_24_port, A_nso(23) => 
                           SHIFT_n_7_23_port, A_nso(22) => SHIFT_n_7_22_port, 
                           A_nso(21) => SHIFT_n_7_21_port, A_nso(20) => 
                           SHIFT_n_7_20_port, A_nso(19) => SHIFT_n_7_19_port, 
                           A_nso(18) => SHIFT_n_7_18_port, A_nso(17) => 
                           SHIFT_n_7_17_port, A_nso(16) => SHIFT_n_7_16_port, 
                           A_nso(15) => SHIFT_n_7_15_port, A_nso(14) => 
                           SHIFT_n_7_14_port, A_nso(13) => SHIFT_n_7_13_port, 
                           A_nso(12) => SHIFT_n_7_12_port, A_nso(11) => 
                           SHIFT_n_7_11_port, A_nso(10) => SHIFT_n_7_10_port, 
                           A_nso(9) => SHIFT_n_7_9_port, A_nso(8) => 
                           SHIFT_n_7_8_port, A_nso(7) => SHIFT_n_7_7_port, 
                           A_nso(6) => SHIFT_n_7_6_port, A_nso(5) => 
                           SHIFT_n_7_5_port, A_nso(4) => SHIFT_n_7_4_port, 
                           A_nso(3) => SHIFT_n_7_3_port, A_nso(2) => 
                           SHIFT_n_7_2_port, A_nso(1) => n_1110, A_nso(0) => 
                           n_1111);
   ENC_7 : BOOTHENC_NBIT48_i14 port map( A_s(47) => SHIFT_7_45_port, A_s(46) =>
                           SHIFT_7_45_port, A_s(45) => SHIFT_7_45_port, A_s(44)
                           => SHIFT_7_44_port, A_s(43) => SHIFT_7_43_port, 
                           A_s(42) => SHIFT_7_42_port, A_s(41) => 
                           SHIFT_7_41_port, A_s(40) => SHIFT_7_40_port, A_s(39)
                           => SHIFT_7_39_port, A_s(38) => SHIFT_7_38_port, 
                           A_s(37) => SHIFT_7_37_port, A_s(36) => 
                           SHIFT_7_36_port, A_s(35) => SHIFT_7_35_port, A_s(34)
                           => SHIFT_7_34_port, A_s(33) => SHIFT_7_33_port, 
                           A_s(32) => SHIFT_7_32_port, A_s(31) => 
                           SHIFT_7_31_port, A_s(30) => SHIFT_7_30_port, A_s(29)
                           => SHIFT_7_29_port, A_s(28) => SHIFT_7_28_port, 
                           A_s(27) => SHIFT_7_27_port, A_s(26) => 
                           SHIFT_7_26_port, A_s(25) => SHIFT_7_25_port, A_s(24)
                           => SHIFT_7_24_port, A_s(23) => SHIFT_7_23_port, 
                           A_s(22) => SHIFT_7_22_port, A_s(21) => 
                           SHIFT_7_21_port, A_s(20) => SHIFT_7_20_port, A_s(19)
                           => SHIFT_7_19_port, A_s(18) => SHIFT_7_18_port, 
                           A_s(17) => SHIFT_7_17_port, A_s(16) => 
                           SHIFT_7_16_port, A_s(15) => SHIFT_7_15_port, A_s(14)
                           => SHIFT_7_14_port, A_s(13) => SHIFT_7_13_port, 
                           A_s(12) => SHIFT_7_12_port, A_s(11) => 
                           SHIFT_7_11_port, A_s(10) => SHIFT_7_10_port, A_s(9) 
                           => SHIFT_7_9_port, A_s(8) => SHIFT_7_8_port, A_s(7) 
                           => SHIFT_7_7_port, A_s(6) => SHIFT_7_6_port, A_s(5) 
                           => SHIFT_7_5_port, A_s(4) => SHIFT_7_4_port, A_s(3) 
                           => SHIFT_7_3_port, A_s(2) => SHIFT_7_2_port, A_s(1) 
                           => SHIFT_7_1_port, A_s(0) => SHIFT_7_0_port, 
                           A_ns(47) => SHIFT_n_7_45_port, A_ns(46) => 
                           SHIFT_n_7_45_port, A_ns(45) => SHIFT_n_7_45_port, 
                           A_ns(44) => SHIFT_n_7_44_port, A_ns(43) => 
                           SHIFT_n_7_43_port, A_ns(42) => SHIFT_n_7_42_port, 
                           A_ns(41) => SHIFT_n_7_41_port, A_ns(40) => 
                           SHIFT_n_7_40_port, A_ns(39) => SHIFT_n_7_39_port, 
                           A_ns(38) => SHIFT_n_7_38_port, A_ns(37) => 
                           SHIFT_n_7_37_port, A_ns(36) => SHIFT_n_7_36_port, 
                           A_ns(35) => SHIFT_n_7_35_port, A_ns(34) => 
                           SHIFT_n_7_34_port, A_ns(33) => SHIFT_n_7_33_port, 
                           A_ns(32) => SHIFT_n_7_32_port, A_ns(31) => 
                           SHIFT_n_7_31_port, A_ns(30) => SHIFT_n_7_30_port, 
                           A_ns(29) => SHIFT_n_7_29_port, A_ns(28) => 
                           SHIFT_n_7_28_port, A_ns(27) => SHIFT_n_7_27_port, 
                           A_ns(26) => SHIFT_n_7_26_port, A_ns(25) => 
                           SHIFT_n_7_25_port, A_ns(24) => SHIFT_n_7_24_port, 
                           A_ns(23) => SHIFT_n_7_23_port, A_ns(22) => 
                           SHIFT_n_7_22_port, A_ns(21) => SHIFT_n_7_21_port, 
                           A_ns(20) => SHIFT_n_7_20_port, A_ns(19) => 
                           SHIFT_n_7_19_port, A_ns(18) => SHIFT_n_7_18_port, 
                           A_ns(17) => SHIFT_n_7_17_port, A_ns(16) => 
                           SHIFT_n_7_16_port, A_ns(15) => SHIFT_n_7_15_port, 
                           A_ns(14) => SHIFT_n_7_14_port, A_ns(13) => 
                           SHIFT_n_7_13_port, A_ns(12) => SHIFT_n_7_12_port, 
                           A_ns(11) => SHIFT_n_7_11_port, A_ns(10) => 
                           SHIFT_n_7_10_port, A_ns(9) => SHIFT_n_7_9_port, 
                           A_ns(8) => SHIFT_n_7_8_port, A_ns(7) => 
                           SHIFT_n_7_7_port, A_ns(6) => SHIFT_n_7_6_port, 
                           A_ns(5) => SHIFT_n_7_5_port, A_ns(4) => 
                           SHIFT_n_7_4_port, A_ns(3) => SHIFT_n_7_3_port, 
                           A_ns(2) => SHIFT_n_7_2_port, A_ns(1) => 
                           SHIFT_n_7_1_port, A_ns(0) => SHIFT_n_7_0_port, B(47)
                           => B(31), B(46) => B(31), B(45) => B(31), B(44) => 
                           B(31), B(43) => B(31), B(42) => B(31), B(41) => 
                           B(31), B(40) => B(31), B(39) => B(31), B(38) => 
                           B(31), B(37) => B(31), B(36) => B(31), B(35) => 
                           B(31), B(34) => B(31), B(33) => B(31), B(32) => 
                           B(31), B(31) => B(31), B(30) => B(30), B(29) => 
                           B(29), B(28) => B(28), B(27) => B(27), B(26) => 
                           B(26), B(25) => B(25), B(24) => B(24), B(23) => 
                           B(23), B(22) => B(22), B(21) => B(21), B(20) => 
                           B(20), B(19) => B(19), B(18) => B(18), B(17) => 
                           B(17), B(16) => B(16), B(15) => B(15), B(14) => 
                           B(14), B(13) => B(13), B(12) => B(12), B(11) => 
                           B(11), B(10) => B(10), B(9) => B(9), B(8) => B(8), 
                           B(7) => B(7), B(6) => B(6), B(5) => B(5), B(4) => 
                           B(4), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), O(47) => OTMP_7_47_port, O(46) => 
                           OTMP_7_46_port, O(45) => OTMP_7_45_port, O(44) => 
                           OTMP_7_44_port, O(43) => OTMP_7_43_port, O(42) => 
                           OTMP_7_42_port, O(41) => OTMP_7_41_port, O(40) => 
                           OTMP_7_40_port, O(39) => OTMP_7_39_port, O(38) => 
                           OTMP_7_38_port, O(37) => OTMP_7_37_port, O(36) => 
                           OTMP_7_36_port, O(35) => OTMP_7_35_port, O(34) => 
                           OTMP_7_34_port, O(33) => OTMP_7_33_port, O(32) => 
                           OTMP_7_32_port, O(31) => OTMP_7_31_port, O(30) => 
                           OTMP_7_30_port, O(29) => OTMP_7_29_port, O(28) => 
                           OTMP_7_28_port, O(27) => OTMP_7_27_port, O(26) => 
                           OTMP_7_26_port, O(25) => OTMP_7_25_port, O(24) => 
                           OTMP_7_24_port, O(23) => OTMP_7_23_port, O(22) => 
                           OTMP_7_22_port, O(21) => OTMP_7_21_port, O(20) => 
                           OTMP_7_20_port, O(19) => OTMP_7_19_port, O(18) => 
                           OTMP_7_18_port, O(17) => OTMP_7_17_port, O(16) => 
                           OTMP_7_16_port, O(15) => OTMP_7_15_port, O(14) => 
                           OTMP_7_14_port, O(13) => OTMP_7_13_port, O(12) => 
                           OTMP_7_12_port, O(11) => OTMP_7_11_port, O(10) => 
                           OTMP_7_10_port, O(9) => OTMP_7_9_port, O(8) => 
                           OTMP_7_8_port, O(7) => OTMP_7_7_port, O(6) => 
                           OTMP_7_6_port, O(5) => OTMP_7_5_port, O(4) => 
                           OTMP_7_4_port, O(3) => OTMP_7_3_port, O(2) => 
                           OTMP_7_2_port, O(1) => OTMP_7_1_port, O(0) => n_1112
                           , A_so(47) => SHIFT_8_47_port, A_so(46) => 
                           SHIFT_8_46_port, A_so(45) => SHIFT_8_45_port, 
                           A_so(44) => SHIFT_8_44_port, A_so(43) => 
                           SHIFT_8_43_port, A_so(42) => SHIFT_8_42_port, 
                           A_so(41) => SHIFT_8_41_port, A_so(40) => 
                           SHIFT_8_40_port, A_so(39) => SHIFT_8_39_port, 
                           A_so(38) => SHIFT_8_38_port, A_so(37) => 
                           SHIFT_8_37_port, A_so(36) => SHIFT_8_36_port, 
                           A_so(35) => SHIFT_8_35_port, A_so(34) => 
                           SHIFT_8_34_port, A_so(33) => SHIFT_8_33_port, 
                           A_so(32) => SHIFT_8_32_port, A_so(31) => 
                           SHIFT_8_31_port, A_so(30) => SHIFT_8_30_port, 
                           A_so(29) => SHIFT_8_29_port, A_so(28) => 
                           SHIFT_8_28_port, A_so(27) => SHIFT_8_27_port, 
                           A_so(26) => SHIFT_8_26_port, A_so(25) => 
                           SHIFT_8_25_port, A_so(24) => SHIFT_8_24_port, 
                           A_so(23) => SHIFT_8_23_port, A_so(22) => 
                           SHIFT_8_22_port, A_so(21) => SHIFT_8_21_port, 
                           A_so(20) => SHIFT_8_20_port, A_so(19) => 
                           SHIFT_8_19_port, A_so(18) => SHIFT_8_18_port, 
                           A_so(17) => SHIFT_8_17_port, A_so(16) => 
                           SHIFT_8_16_port, A_so(15) => SHIFT_8_15_port, 
                           A_so(14) => SHIFT_8_14_port, A_so(13) => 
                           SHIFT_8_13_port, A_so(12) => SHIFT_8_12_port, 
                           A_so(11) => SHIFT_8_11_port, A_so(10) => 
                           SHIFT_8_10_port, A_so(9) => SHIFT_8_9_port, A_so(8) 
                           => SHIFT_8_8_port, A_so(7) => SHIFT_8_7_port, 
                           A_so(6) => SHIFT_8_6_port, A_so(5) => SHIFT_8_5_port
                           , A_so(4) => SHIFT_8_4_port, A_so(3) => 
                           SHIFT_8_3_port, A_so(2) => SHIFT_8_2_port, A_so(1) 
                           => n_1113, A_so(0) => n_1114, A_nso(47) => 
                           SHIFT_n_8_47_port, A_nso(46) => SHIFT_n_8_46_port, 
                           A_nso(45) => SHIFT_n_8_45_port, A_nso(44) => 
                           SHIFT_n_8_44_port, A_nso(43) => SHIFT_n_8_43_port, 
                           A_nso(42) => SHIFT_n_8_42_port, A_nso(41) => 
                           SHIFT_n_8_41_port, A_nso(40) => SHIFT_n_8_40_port, 
                           A_nso(39) => SHIFT_n_8_39_port, A_nso(38) => 
                           SHIFT_n_8_38_port, A_nso(37) => SHIFT_n_8_37_port, 
                           A_nso(36) => SHIFT_n_8_36_port, A_nso(35) => 
                           SHIFT_n_8_35_port, A_nso(34) => SHIFT_n_8_34_port, 
                           A_nso(33) => SHIFT_n_8_33_port, A_nso(32) => 
                           SHIFT_n_8_32_port, A_nso(31) => SHIFT_n_8_31_port, 
                           A_nso(30) => SHIFT_n_8_30_port, A_nso(29) => 
                           SHIFT_n_8_29_port, A_nso(28) => SHIFT_n_8_28_port, 
                           A_nso(27) => SHIFT_n_8_27_port, A_nso(26) => 
                           SHIFT_n_8_26_port, A_nso(25) => SHIFT_n_8_25_port, 
                           A_nso(24) => SHIFT_n_8_24_port, A_nso(23) => 
                           SHIFT_n_8_23_port, A_nso(22) => SHIFT_n_8_22_port, 
                           A_nso(21) => SHIFT_n_8_21_port, A_nso(20) => 
                           SHIFT_n_8_20_port, A_nso(19) => SHIFT_n_8_19_port, 
                           A_nso(18) => SHIFT_n_8_18_port, A_nso(17) => 
                           SHIFT_n_8_17_port, A_nso(16) => SHIFT_n_8_16_port, 
                           A_nso(15) => SHIFT_n_8_15_port, A_nso(14) => 
                           SHIFT_n_8_14_port, A_nso(13) => SHIFT_n_8_13_port, 
                           A_nso(12) => SHIFT_n_8_12_port, A_nso(11) => 
                           SHIFT_n_8_11_port, A_nso(10) => SHIFT_n_8_10_port, 
                           A_nso(9) => SHIFT_n_8_9_port, A_nso(8) => 
                           SHIFT_n_8_8_port, A_nso(7) => SHIFT_n_8_7_port, 
                           A_nso(6) => SHIFT_n_8_6_port, A_nso(5) => 
                           SHIFT_n_8_5_port, A_nso(4) => SHIFT_n_8_4_port, 
                           A_nso(3) => SHIFT_n_8_3_port, A_nso(2) => 
                           SHIFT_n_8_2_port, A_nso(1) => n_1115, A_nso(0) => 
                           n_1116);
   ENC_8 : BOOTHENC_NBIT50_i16 port map( A_s(49) => SHIFT_8_47_port, A_s(48) =>
                           SHIFT_8_47_port, A_s(47) => SHIFT_8_47_port, A_s(46)
                           => SHIFT_8_46_port, A_s(45) => SHIFT_8_45_port, 
                           A_s(44) => SHIFT_8_44_port, A_s(43) => 
                           SHIFT_8_43_port, A_s(42) => SHIFT_8_42_port, A_s(41)
                           => SHIFT_8_41_port, A_s(40) => SHIFT_8_40_port, 
                           A_s(39) => SHIFT_8_39_port, A_s(38) => 
                           SHIFT_8_38_port, A_s(37) => SHIFT_8_37_port, A_s(36)
                           => SHIFT_8_36_port, A_s(35) => SHIFT_8_35_port, 
                           A_s(34) => SHIFT_8_34_port, A_s(33) => 
                           SHIFT_8_33_port, A_s(32) => SHIFT_8_32_port, A_s(31)
                           => SHIFT_8_31_port, A_s(30) => SHIFT_8_30_port, 
                           A_s(29) => SHIFT_8_29_port, A_s(28) => 
                           SHIFT_8_28_port, A_s(27) => SHIFT_8_27_port, A_s(26)
                           => SHIFT_8_26_port, A_s(25) => SHIFT_8_25_port, 
                           A_s(24) => SHIFT_8_24_port, A_s(23) => 
                           SHIFT_8_23_port, A_s(22) => SHIFT_8_22_port, A_s(21)
                           => SHIFT_8_21_port, A_s(20) => SHIFT_8_20_port, 
                           A_s(19) => SHIFT_8_19_port, A_s(18) => 
                           SHIFT_8_18_port, A_s(17) => SHIFT_8_17_port, A_s(16)
                           => SHIFT_8_16_port, A_s(15) => SHIFT_8_15_port, 
                           A_s(14) => SHIFT_8_14_port, A_s(13) => 
                           SHIFT_8_13_port, A_s(12) => SHIFT_8_12_port, A_s(11)
                           => SHIFT_8_11_port, A_s(10) => SHIFT_8_10_port, 
                           A_s(9) => SHIFT_8_9_port, A_s(8) => SHIFT_8_8_port, 
                           A_s(7) => SHIFT_8_7_port, A_s(6) => SHIFT_8_6_port, 
                           A_s(5) => SHIFT_8_5_port, A_s(4) => SHIFT_8_4_port, 
                           A_s(3) => SHIFT_8_3_port, A_s(2) => SHIFT_8_2_port, 
                           A_s(1) => SHIFT_8_1_port, A_s(0) => SHIFT_8_0_port, 
                           A_ns(49) => SHIFT_n_8_47_port, A_ns(48) => 
                           SHIFT_n_8_47_port, A_ns(47) => SHIFT_n_8_47_port, 
                           A_ns(46) => SHIFT_n_8_46_port, A_ns(45) => 
                           SHIFT_n_8_45_port, A_ns(44) => SHIFT_n_8_44_port, 
                           A_ns(43) => SHIFT_n_8_43_port, A_ns(42) => 
                           SHIFT_n_8_42_port, A_ns(41) => SHIFT_n_8_41_port, 
                           A_ns(40) => SHIFT_n_8_40_port, A_ns(39) => 
                           SHIFT_n_8_39_port, A_ns(38) => SHIFT_n_8_38_port, 
                           A_ns(37) => SHIFT_n_8_37_port, A_ns(36) => 
                           SHIFT_n_8_36_port, A_ns(35) => SHIFT_n_8_35_port, 
                           A_ns(34) => SHIFT_n_8_34_port, A_ns(33) => 
                           SHIFT_n_8_33_port, A_ns(32) => SHIFT_n_8_32_port, 
                           A_ns(31) => SHIFT_n_8_31_port, A_ns(30) => 
                           SHIFT_n_8_30_port, A_ns(29) => SHIFT_n_8_29_port, 
                           A_ns(28) => SHIFT_n_8_28_port, A_ns(27) => 
                           SHIFT_n_8_27_port, A_ns(26) => SHIFT_n_8_26_port, 
                           A_ns(25) => SHIFT_n_8_25_port, A_ns(24) => 
                           SHIFT_n_8_24_port, A_ns(23) => SHIFT_n_8_23_port, 
                           A_ns(22) => SHIFT_n_8_22_port, A_ns(21) => 
                           SHIFT_n_8_21_port, A_ns(20) => SHIFT_n_8_20_port, 
                           A_ns(19) => SHIFT_n_8_19_port, A_ns(18) => 
                           SHIFT_n_8_18_port, A_ns(17) => SHIFT_n_8_17_port, 
                           A_ns(16) => SHIFT_n_8_16_port, A_ns(15) => 
                           SHIFT_n_8_15_port, A_ns(14) => SHIFT_n_8_14_port, 
                           A_ns(13) => SHIFT_n_8_13_port, A_ns(12) => 
                           SHIFT_n_8_12_port, A_ns(11) => SHIFT_n_8_11_port, 
                           A_ns(10) => SHIFT_n_8_10_port, A_ns(9) => 
                           SHIFT_n_8_9_port, A_ns(8) => SHIFT_n_8_8_port, 
                           A_ns(7) => SHIFT_n_8_7_port, A_ns(6) => 
                           SHIFT_n_8_6_port, A_ns(5) => SHIFT_n_8_5_port, 
                           A_ns(4) => SHIFT_n_8_4_port, A_ns(3) => 
                           SHIFT_n_8_3_port, A_ns(2) => SHIFT_n_8_2_port, 
                           A_ns(1) => SHIFT_n_8_1_port, A_ns(0) => 
                           SHIFT_n_8_0_port, B(49) => B(31), B(48) => B(31), 
                           B(47) => B(31), B(46) => B(31), B(45) => B(31), 
                           B(44) => B(31), B(43) => B(31), B(42) => B(31), 
                           B(41) => B(31), B(40) => B(31), B(39) => B(31), 
                           B(38) => B(31), B(37) => B(31), B(36) => B(31), 
                           B(35) => B(31), B(34) => B(31), B(33) => B(31), 
                           B(32) => B(31), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), O(49) => OTMP_8_49_port, O(48) 
                           => OTMP_8_48_port, O(47) => OTMP_8_47_port, O(46) =>
                           OTMP_8_46_port, O(45) => OTMP_8_45_port, O(44) => 
                           OTMP_8_44_port, O(43) => OTMP_8_43_port, O(42) => 
                           OTMP_8_42_port, O(41) => OTMP_8_41_port, O(40) => 
                           OTMP_8_40_port, O(39) => OTMP_8_39_port, O(38) => 
                           OTMP_8_38_port, O(37) => OTMP_8_37_port, O(36) => 
                           OTMP_8_36_port, O(35) => OTMP_8_35_port, O(34) => 
                           OTMP_8_34_port, O(33) => OTMP_8_33_port, O(32) => 
                           OTMP_8_32_port, O(31) => OTMP_8_31_port, O(30) => 
                           OTMP_8_30_port, O(29) => OTMP_8_29_port, O(28) => 
                           OTMP_8_28_port, O(27) => OTMP_8_27_port, O(26) => 
                           OTMP_8_26_port, O(25) => OTMP_8_25_port, O(24) => 
                           OTMP_8_24_port, O(23) => OTMP_8_23_port, O(22) => 
                           OTMP_8_22_port, O(21) => OTMP_8_21_port, O(20) => 
                           OTMP_8_20_port, O(19) => OTMP_8_19_port, O(18) => 
                           OTMP_8_18_port, O(17) => OTMP_8_17_port, O(16) => 
                           OTMP_8_16_port, O(15) => OTMP_8_15_port, O(14) => 
                           OTMP_8_14_port, O(13) => OTMP_8_13_port, O(12) => 
                           OTMP_8_12_port, O(11) => OTMP_8_11_port, O(10) => 
                           OTMP_8_10_port, O(9) => OTMP_8_9_port, O(8) => 
                           OTMP_8_8_port, O(7) => OTMP_8_7_port, O(6) => 
                           OTMP_8_6_port, O(5) => OTMP_8_5_port, O(4) => 
                           OTMP_8_4_port, O(3) => OTMP_8_3_port, O(2) => 
                           OTMP_8_2_port, O(1) => OTMP_8_1_port, O(0) => n_1117
                           , A_so(49) => SHIFT_9_49_port, A_so(48) => 
                           SHIFT_9_48_port, A_so(47) => SHIFT_9_47_port, 
                           A_so(46) => SHIFT_9_46_port, A_so(45) => 
                           SHIFT_9_45_port, A_so(44) => SHIFT_9_44_port, 
                           A_so(43) => SHIFT_9_43_port, A_so(42) => 
                           SHIFT_9_42_port, A_so(41) => SHIFT_9_41_port, 
                           A_so(40) => SHIFT_9_40_port, A_so(39) => 
                           SHIFT_9_39_port, A_so(38) => SHIFT_9_38_port, 
                           A_so(37) => SHIFT_9_37_port, A_so(36) => 
                           SHIFT_9_36_port, A_so(35) => SHIFT_9_35_port, 
                           A_so(34) => SHIFT_9_34_port, A_so(33) => 
                           SHIFT_9_33_port, A_so(32) => SHIFT_9_32_port, 
                           A_so(31) => SHIFT_9_31_port, A_so(30) => 
                           SHIFT_9_30_port, A_so(29) => SHIFT_9_29_port, 
                           A_so(28) => SHIFT_9_28_port, A_so(27) => 
                           SHIFT_9_27_port, A_so(26) => SHIFT_9_26_port, 
                           A_so(25) => SHIFT_9_25_port, A_so(24) => 
                           SHIFT_9_24_port, A_so(23) => SHIFT_9_23_port, 
                           A_so(22) => SHIFT_9_22_port, A_so(21) => 
                           SHIFT_9_21_port, A_so(20) => SHIFT_9_20_port, 
                           A_so(19) => SHIFT_9_19_port, A_so(18) => 
                           SHIFT_9_18_port, A_so(17) => SHIFT_9_17_port, 
                           A_so(16) => SHIFT_9_16_port, A_so(15) => 
                           SHIFT_9_15_port, A_so(14) => SHIFT_9_14_port, 
                           A_so(13) => SHIFT_9_13_port, A_so(12) => 
                           SHIFT_9_12_port, A_so(11) => SHIFT_9_11_port, 
                           A_so(10) => SHIFT_9_10_port, A_so(9) => 
                           SHIFT_9_9_port, A_so(8) => SHIFT_9_8_port, A_so(7) 
                           => SHIFT_9_7_port, A_so(6) => SHIFT_9_6_port, 
                           A_so(5) => SHIFT_9_5_port, A_so(4) => SHIFT_9_4_port
                           , A_so(3) => SHIFT_9_3_port, A_so(2) => 
                           SHIFT_9_2_port, A_so(1) => n_1118, A_so(0) => n_1119
                           , A_nso(49) => SHIFT_n_9_49_port, A_nso(48) => 
                           SHIFT_n_9_48_port, A_nso(47) => SHIFT_n_9_47_port, 
                           A_nso(46) => SHIFT_n_9_46_port, A_nso(45) => 
                           SHIFT_n_9_45_port, A_nso(44) => SHIFT_n_9_44_port, 
                           A_nso(43) => SHIFT_n_9_43_port, A_nso(42) => 
                           SHIFT_n_9_42_port, A_nso(41) => SHIFT_n_9_41_port, 
                           A_nso(40) => SHIFT_n_9_40_port, A_nso(39) => 
                           SHIFT_n_9_39_port, A_nso(38) => SHIFT_n_9_38_port, 
                           A_nso(37) => SHIFT_n_9_37_port, A_nso(36) => 
                           SHIFT_n_9_36_port, A_nso(35) => SHIFT_n_9_35_port, 
                           A_nso(34) => SHIFT_n_9_34_port, A_nso(33) => 
                           SHIFT_n_9_33_port, A_nso(32) => SHIFT_n_9_32_port, 
                           A_nso(31) => SHIFT_n_9_31_port, A_nso(30) => 
                           SHIFT_n_9_30_port, A_nso(29) => SHIFT_n_9_29_port, 
                           A_nso(28) => SHIFT_n_9_28_port, A_nso(27) => 
                           SHIFT_n_9_27_port, A_nso(26) => SHIFT_n_9_26_port, 
                           A_nso(25) => SHIFT_n_9_25_port, A_nso(24) => 
                           SHIFT_n_9_24_port, A_nso(23) => SHIFT_n_9_23_port, 
                           A_nso(22) => SHIFT_n_9_22_port, A_nso(21) => 
                           SHIFT_n_9_21_port, A_nso(20) => SHIFT_n_9_20_port, 
                           A_nso(19) => SHIFT_n_9_19_port, A_nso(18) => 
                           SHIFT_n_9_18_port, A_nso(17) => SHIFT_n_9_17_port, 
                           A_nso(16) => SHIFT_n_9_16_port, A_nso(15) => 
                           SHIFT_n_9_15_port, A_nso(14) => SHIFT_n_9_14_port, 
                           A_nso(13) => SHIFT_n_9_13_port, A_nso(12) => 
                           SHIFT_n_9_12_port, A_nso(11) => SHIFT_n_9_11_port, 
                           A_nso(10) => SHIFT_n_9_10_port, A_nso(9) => 
                           SHIFT_n_9_9_port, A_nso(8) => SHIFT_n_9_8_port, 
                           A_nso(7) => SHIFT_n_9_7_port, A_nso(6) => 
                           SHIFT_n_9_6_port, A_nso(5) => SHIFT_n_9_5_port, 
                           A_nso(4) => SHIFT_n_9_4_port, A_nso(3) => 
                           SHIFT_n_9_3_port, A_nso(2) => SHIFT_n_9_2_port, 
                           A_nso(1) => n_1120, A_nso(0) => n_1121);
   ENC_9 : BOOTHENC_NBIT52_i18 port map( A_s(51) => SHIFT_9_49_port, A_s(50) =>
                           SHIFT_9_49_port, A_s(49) => SHIFT_9_49_port, A_s(48)
                           => SHIFT_9_48_port, A_s(47) => SHIFT_9_47_port, 
                           A_s(46) => SHIFT_9_46_port, A_s(45) => 
                           SHIFT_9_45_port, A_s(44) => SHIFT_9_44_port, A_s(43)
                           => SHIFT_9_43_port, A_s(42) => SHIFT_9_42_port, 
                           A_s(41) => SHIFT_9_41_port, A_s(40) => 
                           SHIFT_9_40_port, A_s(39) => SHIFT_9_39_port, A_s(38)
                           => SHIFT_9_38_port, A_s(37) => SHIFT_9_37_port, 
                           A_s(36) => SHIFT_9_36_port, A_s(35) => 
                           SHIFT_9_35_port, A_s(34) => SHIFT_9_34_port, A_s(33)
                           => SHIFT_9_33_port, A_s(32) => SHIFT_9_32_port, 
                           A_s(31) => SHIFT_9_31_port, A_s(30) => 
                           SHIFT_9_30_port, A_s(29) => SHIFT_9_29_port, A_s(28)
                           => SHIFT_9_28_port, A_s(27) => SHIFT_9_27_port, 
                           A_s(26) => SHIFT_9_26_port, A_s(25) => 
                           SHIFT_9_25_port, A_s(24) => SHIFT_9_24_port, A_s(23)
                           => SHIFT_9_23_port, A_s(22) => SHIFT_9_22_port, 
                           A_s(21) => SHIFT_9_21_port, A_s(20) => 
                           SHIFT_9_20_port, A_s(19) => SHIFT_9_19_port, A_s(18)
                           => SHIFT_9_18_port, A_s(17) => SHIFT_9_17_port, 
                           A_s(16) => SHIFT_9_16_port, A_s(15) => 
                           SHIFT_9_15_port, A_s(14) => SHIFT_9_14_port, A_s(13)
                           => SHIFT_9_13_port, A_s(12) => SHIFT_9_12_port, 
                           A_s(11) => SHIFT_9_11_port, A_s(10) => 
                           SHIFT_9_10_port, A_s(9) => SHIFT_9_9_port, A_s(8) =>
                           SHIFT_9_8_port, A_s(7) => SHIFT_9_7_port, A_s(6) => 
                           SHIFT_9_6_port, A_s(5) => SHIFT_9_5_port, A_s(4) => 
                           SHIFT_9_4_port, A_s(3) => SHIFT_9_3_port, A_s(2) => 
                           SHIFT_9_2_port, A_s(1) => SHIFT_9_1_port, A_s(0) => 
                           SHIFT_9_0_port, A_ns(51) => SHIFT_n_9_49_port, 
                           A_ns(50) => SHIFT_n_9_49_port, A_ns(49) => 
                           SHIFT_n_9_49_port, A_ns(48) => SHIFT_n_9_48_port, 
                           A_ns(47) => SHIFT_n_9_47_port, A_ns(46) => 
                           SHIFT_n_9_46_port, A_ns(45) => SHIFT_n_9_45_port, 
                           A_ns(44) => SHIFT_n_9_44_port, A_ns(43) => 
                           SHIFT_n_9_43_port, A_ns(42) => SHIFT_n_9_42_port, 
                           A_ns(41) => SHIFT_n_9_41_port, A_ns(40) => 
                           SHIFT_n_9_40_port, A_ns(39) => SHIFT_n_9_39_port, 
                           A_ns(38) => SHIFT_n_9_38_port, A_ns(37) => 
                           SHIFT_n_9_37_port, A_ns(36) => SHIFT_n_9_36_port, 
                           A_ns(35) => SHIFT_n_9_35_port, A_ns(34) => 
                           SHIFT_n_9_34_port, A_ns(33) => SHIFT_n_9_33_port, 
                           A_ns(32) => SHIFT_n_9_32_port, A_ns(31) => 
                           SHIFT_n_9_31_port, A_ns(30) => SHIFT_n_9_30_port, 
                           A_ns(29) => SHIFT_n_9_29_port, A_ns(28) => 
                           SHIFT_n_9_28_port, A_ns(27) => SHIFT_n_9_27_port, 
                           A_ns(26) => SHIFT_n_9_26_port, A_ns(25) => 
                           SHIFT_n_9_25_port, A_ns(24) => SHIFT_n_9_24_port, 
                           A_ns(23) => SHIFT_n_9_23_port, A_ns(22) => 
                           SHIFT_n_9_22_port, A_ns(21) => SHIFT_n_9_21_port, 
                           A_ns(20) => SHIFT_n_9_20_port, A_ns(19) => 
                           SHIFT_n_9_19_port, A_ns(18) => SHIFT_n_9_18_port, 
                           A_ns(17) => SHIFT_n_9_17_port, A_ns(16) => 
                           SHIFT_n_9_16_port, A_ns(15) => SHIFT_n_9_15_port, 
                           A_ns(14) => SHIFT_n_9_14_port, A_ns(13) => 
                           SHIFT_n_9_13_port, A_ns(12) => SHIFT_n_9_12_port, 
                           A_ns(11) => SHIFT_n_9_11_port, A_ns(10) => 
                           SHIFT_n_9_10_port, A_ns(9) => SHIFT_n_9_9_port, 
                           A_ns(8) => SHIFT_n_9_8_port, A_ns(7) => 
                           SHIFT_n_9_7_port, A_ns(6) => SHIFT_n_9_6_port, 
                           A_ns(5) => SHIFT_n_9_5_port, A_ns(4) => 
                           SHIFT_n_9_4_port, A_ns(3) => SHIFT_n_9_3_port, 
                           A_ns(2) => SHIFT_n_9_2_port, A_ns(1) => 
                           SHIFT_n_9_1_port, A_ns(0) => SHIFT_n_9_0_port, B(51)
                           => B(31), B(50) => B(31), B(49) => B(31), B(48) => 
                           B(31), B(47) => B(31), B(46) => B(31), B(45) => 
                           B(31), B(44) => B(31), B(43) => B(31), B(42) => 
                           B(31), B(41) => B(31), B(40) => B(31), B(39) => 
                           B(31), B(38) => B(31), B(37) => B(31), B(36) => 
                           B(31), B(35) => B(31), B(34) => B(31), B(33) => 
                           B(31), B(32) => B(31), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), O(51) => OTMP_9_51_port, 
                           O(50) => OTMP_9_50_port, O(49) => OTMP_9_49_port, 
                           O(48) => OTMP_9_48_port, O(47) => OTMP_9_47_port, 
                           O(46) => OTMP_9_46_port, O(45) => OTMP_9_45_port, 
                           O(44) => OTMP_9_44_port, O(43) => OTMP_9_43_port, 
                           O(42) => OTMP_9_42_port, O(41) => OTMP_9_41_port, 
                           O(40) => OTMP_9_40_port, O(39) => OTMP_9_39_port, 
                           O(38) => OTMP_9_38_port, O(37) => OTMP_9_37_port, 
                           O(36) => OTMP_9_36_port, O(35) => OTMP_9_35_port, 
                           O(34) => OTMP_9_34_port, O(33) => OTMP_9_33_port, 
                           O(32) => OTMP_9_32_port, O(31) => OTMP_9_31_port, 
                           O(30) => OTMP_9_30_port, O(29) => OTMP_9_29_port, 
                           O(28) => OTMP_9_28_port, O(27) => OTMP_9_27_port, 
                           O(26) => OTMP_9_26_port, O(25) => OTMP_9_25_port, 
                           O(24) => OTMP_9_24_port, O(23) => OTMP_9_23_port, 
                           O(22) => OTMP_9_22_port, O(21) => OTMP_9_21_port, 
                           O(20) => OTMP_9_20_port, O(19) => OTMP_9_19_port, 
                           O(18) => OTMP_9_18_port, O(17) => OTMP_9_17_port, 
                           O(16) => OTMP_9_16_port, O(15) => OTMP_9_15_port, 
                           O(14) => OTMP_9_14_port, O(13) => OTMP_9_13_port, 
                           O(12) => OTMP_9_12_port, O(11) => OTMP_9_11_port, 
                           O(10) => OTMP_9_10_port, O(9) => OTMP_9_9_port, O(8)
                           => OTMP_9_8_port, O(7) => OTMP_9_7_port, O(6) => 
                           OTMP_9_6_port, O(5) => OTMP_9_5_port, O(4) => 
                           OTMP_9_4_port, O(3) => OTMP_9_3_port, O(2) => 
                           OTMP_9_2_port, O(1) => OTMP_9_1_port, O(0) => n_1122
                           , A_so(51) => SHIFT_10_51_port, A_so(50) => 
                           SHIFT_10_50_port, A_so(49) => SHIFT_10_49_port, 
                           A_so(48) => SHIFT_10_48_port, A_so(47) => 
                           SHIFT_10_47_port, A_so(46) => SHIFT_10_46_port, 
                           A_so(45) => SHIFT_10_45_port, A_so(44) => 
                           SHIFT_10_44_port, A_so(43) => SHIFT_10_43_port, 
                           A_so(42) => SHIFT_10_42_port, A_so(41) => 
                           SHIFT_10_41_port, A_so(40) => SHIFT_10_40_port, 
                           A_so(39) => SHIFT_10_39_port, A_so(38) => 
                           SHIFT_10_38_port, A_so(37) => SHIFT_10_37_port, 
                           A_so(36) => SHIFT_10_36_port, A_so(35) => 
                           SHIFT_10_35_port, A_so(34) => SHIFT_10_34_port, 
                           A_so(33) => SHIFT_10_33_port, A_so(32) => 
                           SHIFT_10_32_port, A_so(31) => SHIFT_10_31_port, 
                           A_so(30) => SHIFT_10_30_port, A_so(29) => 
                           SHIFT_10_29_port, A_so(28) => SHIFT_10_28_port, 
                           A_so(27) => SHIFT_10_27_port, A_so(26) => 
                           SHIFT_10_26_port, A_so(25) => SHIFT_10_25_port, 
                           A_so(24) => SHIFT_10_24_port, A_so(23) => 
                           SHIFT_10_23_port, A_so(22) => SHIFT_10_22_port, 
                           A_so(21) => SHIFT_10_21_port, A_so(20) => 
                           SHIFT_10_20_port, A_so(19) => SHIFT_10_19_port, 
                           A_so(18) => SHIFT_10_18_port, A_so(17) => 
                           SHIFT_10_17_port, A_so(16) => SHIFT_10_16_port, 
                           A_so(15) => SHIFT_10_15_port, A_so(14) => 
                           SHIFT_10_14_port, A_so(13) => SHIFT_10_13_port, 
                           A_so(12) => SHIFT_10_12_port, A_so(11) => 
                           SHIFT_10_11_port, A_so(10) => SHIFT_10_10_port, 
                           A_so(9) => SHIFT_10_9_port, A_so(8) => 
                           SHIFT_10_8_port, A_so(7) => SHIFT_10_7_port, A_so(6)
                           => SHIFT_10_6_port, A_so(5) => SHIFT_10_5_port, 
                           A_so(4) => SHIFT_10_4_port, A_so(3) => 
                           SHIFT_10_3_port, A_so(2) => SHIFT_10_2_port, A_so(1)
                           => n_1123, A_so(0) => n_1124, A_nso(51) => 
                           SHIFT_n_10_51_port, A_nso(50) => SHIFT_n_10_50_port,
                           A_nso(49) => SHIFT_n_10_49_port, A_nso(48) => 
                           SHIFT_n_10_48_port, A_nso(47) => SHIFT_n_10_47_port,
                           A_nso(46) => SHIFT_n_10_46_port, A_nso(45) => 
                           SHIFT_n_10_45_port, A_nso(44) => SHIFT_n_10_44_port,
                           A_nso(43) => SHIFT_n_10_43_port, A_nso(42) => 
                           SHIFT_n_10_42_port, A_nso(41) => SHIFT_n_10_41_port,
                           A_nso(40) => SHIFT_n_10_40_port, A_nso(39) => 
                           SHIFT_n_10_39_port, A_nso(38) => SHIFT_n_10_38_port,
                           A_nso(37) => SHIFT_n_10_37_port, A_nso(36) => 
                           SHIFT_n_10_36_port, A_nso(35) => SHIFT_n_10_35_port,
                           A_nso(34) => SHIFT_n_10_34_port, A_nso(33) => 
                           SHIFT_n_10_33_port, A_nso(32) => SHIFT_n_10_32_port,
                           A_nso(31) => SHIFT_n_10_31_port, A_nso(30) => 
                           SHIFT_n_10_30_port, A_nso(29) => SHIFT_n_10_29_port,
                           A_nso(28) => SHIFT_n_10_28_port, A_nso(27) => 
                           SHIFT_n_10_27_port, A_nso(26) => SHIFT_n_10_26_port,
                           A_nso(25) => SHIFT_n_10_25_port, A_nso(24) => 
                           SHIFT_n_10_24_port, A_nso(23) => SHIFT_n_10_23_port,
                           A_nso(22) => SHIFT_n_10_22_port, A_nso(21) => 
                           SHIFT_n_10_21_port, A_nso(20) => SHIFT_n_10_20_port,
                           A_nso(19) => SHIFT_n_10_19_port, A_nso(18) => 
                           SHIFT_n_10_18_port, A_nso(17) => SHIFT_n_10_17_port,
                           A_nso(16) => SHIFT_n_10_16_port, A_nso(15) => 
                           SHIFT_n_10_15_port, A_nso(14) => SHIFT_n_10_14_port,
                           A_nso(13) => SHIFT_n_10_13_port, A_nso(12) => 
                           SHIFT_n_10_12_port, A_nso(11) => SHIFT_n_10_11_port,
                           A_nso(10) => SHIFT_n_10_10_port, A_nso(9) => 
                           SHIFT_n_10_9_port, A_nso(8) => SHIFT_n_10_8_port, 
                           A_nso(7) => SHIFT_n_10_7_port, A_nso(6) => 
                           SHIFT_n_10_6_port, A_nso(5) => SHIFT_n_10_5_port, 
                           A_nso(4) => SHIFT_n_10_4_port, A_nso(3) => 
                           SHIFT_n_10_3_port, A_nso(2) => SHIFT_n_10_2_port, 
                           A_nso(1) => n_1125, A_nso(0) => n_1126);
   ENC_10 : BOOTHENC_NBIT54_i20 port map( A_s(53) => SHIFT_10_51_port, A_s(52) 
                           => SHIFT_10_51_port, A_s(51) => SHIFT_10_51_port, 
                           A_s(50) => SHIFT_10_50_port, A_s(49) => 
                           SHIFT_10_49_port, A_s(48) => SHIFT_10_48_port, 
                           A_s(47) => SHIFT_10_47_port, A_s(46) => 
                           SHIFT_10_46_port, A_s(45) => SHIFT_10_45_port, 
                           A_s(44) => SHIFT_10_44_port, A_s(43) => 
                           SHIFT_10_43_port, A_s(42) => SHIFT_10_42_port, 
                           A_s(41) => SHIFT_10_41_port, A_s(40) => 
                           SHIFT_10_40_port, A_s(39) => SHIFT_10_39_port, 
                           A_s(38) => SHIFT_10_38_port, A_s(37) => 
                           SHIFT_10_37_port, A_s(36) => SHIFT_10_36_port, 
                           A_s(35) => SHIFT_10_35_port, A_s(34) => 
                           SHIFT_10_34_port, A_s(33) => SHIFT_10_33_port, 
                           A_s(32) => SHIFT_10_32_port, A_s(31) => 
                           SHIFT_10_31_port, A_s(30) => SHIFT_10_30_port, 
                           A_s(29) => SHIFT_10_29_port, A_s(28) => 
                           SHIFT_10_28_port, A_s(27) => SHIFT_10_27_port, 
                           A_s(26) => SHIFT_10_26_port, A_s(25) => 
                           SHIFT_10_25_port, A_s(24) => SHIFT_10_24_port, 
                           A_s(23) => SHIFT_10_23_port, A_s(22) => 
                           SHIFT_10_22_port, A_s(21) => SHIFT_10_21_port, 
                           A_s(20) => SHIFT_10_20_port, A_s(19) => 
                           SHIFT_10_19_port, A_s(18) => SHIFT_10_18_port, 
                           A_s(17) => SHIFT_10_17_port, A_s(16) => 
                           SHIFT_10_16_port, A_s(15) => SHIFT_10_15_port, 
                           A_s(14) => SHIFT_10_14_port, A_s(13) => 
                           SHIFT_10_13_port, A_s(12) => SHIFT_10_12_port, 
                           A_s(11) => SHIFT_10_11_port, A_s(10) => 
                           SHIFT_10_10_port, A_s(9) => SHIFT_10_9_port, A_s(8) 
                           => SHIFT_10_8_port, A_s(7) => SHIFT_10_7_port, 
                           A_s(6) => SHIFT_10_6_port, A_s(5) => SHIFT_10_5_port
                           , A_s(4) => SHIFT_10_4_port, A_s(3) => 
                           SHIFT_10_3_port, A_s(2) => SHIFT_10_2_port, A_s(1) 
                           => SHIFT_10_1_port, A_s(0) => SHIFT_10_0_port, 
                           A_ns(53) => SHIFT_n_10_51_port, A_ns(52) => 
                           SHIFT_n_10_51_port, A_ns(51) => SHIFT_n_10_51_port, 
                           A_ns(50) => SHIFT_n_10_50_port, A_ns(49) => 
                           SHIFT_n_10_49_port, A_ns(48) => SHIFT_n_10_48_port, 
                           A_ns(47) => SHIFT_n_10_47_port, A_ns(46) => 
                           SHIFT_n_10_46_port, A_ns(45) => SHIFT_n_10_45_port, 
                           A_ns(44) => SHIFT_n_10_44_port, A_ns(43) => 
                           SHIFT_n_10_43_port, A_ns(42) => SHIFT_n_10_42_port, 
                           A_ns(41) => SHIFT_n_10_41_port, A_ns(40) => 
                           SHIFT_n_10_40_port, A_ns(39) => SHIFT_n_10_39_port, 
                           A_ns(38) => SHIFT_n_10_38_port, A_ns(37) => 
                           SHIFT_n_10_37_port, A_ns(36) => SHIFT_n_10_36_port, 
                           A_ns(35) => SHIFT_n_10_35_port, A_ns(34) => 
                           SHIFT_n_10_34_port, A_ns(33) => SHIFT_n_10_33_port, 
                           A_ns(32) => SHIFT_n_10_32_port, A_ns(31) => 
                           SHIFT_n_10_31_port, A_ns(30) => SHIFT_n_10_30_port, 
                           A_ns(29) => SHIFT_n_10_29_port, A_ns(28) => 
                           SHIFT_n_10_28_port, A_ns(27) => SHIFT_n_10_27_port, 
                           A_ns(26) => SHIFT_n_10_26_port, A_ns(25) => 
                           SHIFT_n_10_25_port, A_ns(24) => SHIFT_n_10_24_port, 
                           A_ns(23) => SHIFT_n_10_23_port, A_ns(22) => 
                           SHIFT_n_10_22_port, A_ns(21) => SHIFT_n_10_21_port, 
                           A_ns(20) => SHIFT_n_10_20_port, A_ns(19) => 
                           SHIFT_n_10_19_port, A_ns(18) => SHIFT_n_10_18_port, 
                           A_ns(17) => SHIFT_n_10_17_port, A_ns(16) => 
                           SHIFT_n_10_16_port, A_ns(15) => SHIFT_n_10_15_port, 
                           A_ns(14) => SHIFT_n_10_14_port, A_ns(13) => 
                           SHIFT_n_10_13_port, A_ns(12) => SHIFT_n_10_12_port, 
                           A_ns(11) => SHIFT_n_10_11_port, A_ns(10) => 
                           SHIFT_n_10_10_port, A_ns(9) => SHIFT_n_10_9_port, 
                           A_ns(8) => SHIFT_n_10_8_port, A_ns(7) => 
                           SHIFT_n_10_7_port, A_ns(6) => SHIFT_n_10_6_port, 
                           A_ns(5) => SHIFT_n_10_5_port, A_ns(4) => 
                           SHIFT_n_10_4_port, A_ns(3) => SHIFT_n_10_3_port, 
                           A_ns(2) => SHIFT_n_10_2_port, A_ns(1) => 
                           SHIFT_n_10_1_port, A_ns(0) => SHIFT_n_10_0_port, 
                           B(53) => B(31), B(52) => B(31), B(51) => B(31), 
                           B(50) => B(31), B(49) => B(31), B(48) => B(31), 
                           B(47) => B(31), B(46) => B(31), B(45) => B(31), 
                           B(44) => B(31), B(43) => B(31), B(42) => B(31), 
                           B(41) => B(31), B(40) => B(31), B(39) => B(31), 
                           B(38) => B(31), B(37) => B(31), B(36) => B(31), 
                           B(35) => B(31), B(34) => B(31), B(33) => B(31), 
                           B(32) => B(31), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), O(53) => OTMP_10_53_port, O(52) 
                           => OTMP_10_52_port, O(51) => OTMP_10_51_port, O(50) 
                           => OTMP_10_50_port, O(49) => OTMP_10_49_port, O(48) 
                           => OTMP_10_48_port, O(47) => OTMP_10_47_port, O(46) 
                           => OTMP_10_46_port, O(45) => OTMP_10_45_port, O(44) 
                           => OTMP_10_44_port, O(43) => OTMP_10_43_port, O(42) 
                           => OTMP_10_42_port, O(41) => OTMP_10_41_port, O(40) 
                           => OTMP_10_40_port, O(39) => OTMP_10_39_port, O(38) 
                           => OTMP_10_38_port, O(37) => OTMP_10_37_port, O(36) 
                           => OTMP_10_36_port, O(35) => OTMP_10_35_port, O(34) 
                           => OTMP_10_34_port, O(33) => OTMP_10_33_port, O(32) 
                           => OTMP_10_32_port, O(31) => OTMP_10_31_port, O(30) 
                           => OTMP_10_30_port, O(29) => OTMP_10_29_port, O(28) 
                           => OTMP_10_28_port, O(27) => OTMP_10_27_port, O(26) 
                           => OTMP_10_26_port, O(25) => OTMP_10_25_port, O(24) 
                           => OTMP_10_24_port, O(23) => OTMP_10_23_port, O(22) 
                           => OTMP_10_22_port, O(21) => OTMP_10_21_port, O(20) 
                           => OTMP_10_20_port, O(19) => OTMP_10_19_port, O(18) 
                           => OTMP_10_18_port, O(17) => OTMP_10_17_port, O(16) 
                           => OTMP_10_16_port, O(15) => OTMP_10_15_port, O(14) 
                           => OTMP_10_14_port, O(13) => OTMP_10_13_port, O(12) 
                           => OTMP_10_12_port, O(11) => OTMP_10_11_port, O(10) 
                           => OTMP_10_10_port, O(9) => OTMP_10_9_port, O(8) => 
                           OTMP_10_8_port, O(7) => OTMP_10_7_port, O(6) => 
                           OTMP_10_6_port, O(5) => OTMP_10_5_port, O(4) => 
                           OTMP_10_4_port, O(3) => OTMP_10_3_port, O(2) => 
                           OTMP_10_2_port, O(1) => OTMP_10_1_port, O(0) => 
                           n_1127, A_so(53) => SHIFT_11_53_port, A_so(52) => 
                           SHIFT_11_52_port, A_so(51) => SHIFT_11_51_port, 
                           A_so(50) => SHIFT_11_50_port, A_so(49) => 
                           SHIFT_11_49_port, A_so(48) => SHIFT_11_48_port, 
                           A_so(47) => SHIFT_11_47_port, A_so(46) => 
                           SHIFT_11_46_port, A_so(45) => SHIFT_11_45_port, 
                           A_so(44) => SHIFT_11_44_port, A_so(43) => 
                           SHIFT_11_43_port, A_so(42) => SHIFT_11_42_port, 
                           A_so(41) => SHIFT_11_41_port, A_so(40) => 
                           SHIFT_11_40_port, A_so(39) => SHIFT_11_39_port, 
                           A_so(38) => SHIFT_11_38_port, A_so(37) => 
                           SHIFT_11_37_port, A_so(36) => SHIFT_11_36_port, 
                           A_so(35) => SHIFT_11_35_port, A_so(34) => 
                           SHIFT_11_34_port, A_so(33) => SHIFT_11_33_port, 
                           A_so(32) => SHIFT_11_32_port, A_so(31) => 
                           SHIFT_11_31_port, A_so(30) => SHIFT_11_30_port, 
                           A_so(29) => SHIFT_11_29_port, A_so(28) => 
                           SHIFT_11_28_port, A_so(27) => SHIFT_11_27_port, 
                           A_so(26) => SHIFT_11_26_port, A_so(25) => 
                           SHIFT_11_25_port, A_so(24) => SHIFT_11_24_port, 
                           A_so(23) => SHIFT_11_23_port, A_so(22) => 
                           SHIFT_11_22_port, A_so(21) => SHIFT_11_21_port, 
                           A_so(20) => SHIFT_11_20_port, A_so(19) => 
                           SHIFT_11_19_port, A_so(18) => SHIFT_11_18_port, 
                           A_so(17) => SHIFT_11_17_port, A_so(16) => 
                           SHIFT_11_16_port, A_so(15) => SHIFT_11_15_port, 
                           A_so(14) => SHIFT_11_14_port, A_so(13) => 
                           SHIFT_11_13_port, A_so(12) => SHIFT_11_12_port, 
                           A_so(11) => SHIFT_11_11_port, A_so(10) => 
                           SHIFT_11_10_port, A_so(9) => SHIFT_11_9_port, 
                           A_so(8) => SHIFT_11_8_port, A_so(7) => 
                           SHIFT_11_7_port, A_so(6) => SHIFT_11_6_port, A_so(5)
                           => SHIFT_11_5_port, A_so(4) => SHIFT_11_4_port, 
                           A_so(3) => SHIFT_11_3_port, A_so(2) => 
                           SHIFT_11_2_port, A_so(1) => n_1128, A_so(0) => 
                           n_1129, A_nso(53) => SHIFT_n_11_53_port, A_nso(52) 
                           => SHIFT_n_11_52_port, A_nso(51) => 
                           SHIFT_n_11_51_port, A_nso(50) => SHIFT_n_11_50_port,
                           A_nso(49) => SHIFT_n_11_49_port, A_nso(48) => 
                           SHIFT_n_11_48_port, A_nso(47) => SHIFT_n_11_47_port,
                           A_nso(46) => SHIFT_n_11_46_port, A_nso(45) => 
                           SHIFT_n_11_45_port, A_nso(44) => SHIFT_n_11_44_port,
                           A_nso(43) => SHIFT_n_11_43_port, A_nso(42) => 
                           SHIFT_n_11_42_port, A_nso(41) => SHIFT_n_11_41_port,
                           A_nso(40) => SHIFT_n_11_40_port, A_nso(39) => 
                           SHIFT_n_11_39_port, A_nso(38) => SHIFT_n_11_38_port,
                           A_nso(37) => SHIFT_n_11_37_port, A_nso(36) => 
                           SHIFT_n_11_36_port, A_nso(35) => SHIFT_n_11_35_port,
                           A_nso(34) => SHIFT_n_11_34_port, A_nso(33) => 
                           SHIFT_n_11_33_port, A_nso(32) => SHIFT_n_11_32_port,
                           A_nso(31) => SHIFT_n_11_31_port, A_nso(30) => 
                           SHIFT_n_11_30_port, A_nso(29) => SHIFT_n_11_29_port,
                           A_nso(28) => SHIFT_n_11_28_port, A_nso(27) => 
                           SHIFT_n_11_27_port, A_nso(26) => SHIFT_n_11_26_port,
                           A_nso(25) => SHIFT_n_11_25_port, A_nso(24) => 
                           SHIFT_n_11_24_port, A_nso(23) => SHIFT_n_11_23_port,
                           A_nso(22) => SHIFT_n_11_22_port, A_nso(21) => 
                           SHIFT_n_11_21_port, A_nso(20) => SHIFT_n_11_20_port,
                           A_nso(19) => SHIFT_n_11_19_port, A_nso(18) => 
                           SHIFT_n_11_18_port, A_nso(17) => SHIFT_n_11_17_port,
                           A_nso(16) => SHIFT_n_11_16_port, A_nso(15) => 
                           SHIFT_n_11_15_port, A_nso(14) => SHIFT_n_11_14_port,
                           A_nso(13) => SHIFT_n_11_13_port, A_nso(12) => 
                           SHIFT_n_11_12_port, A_nso(11) => SHIFT_n_11_11_port,
                           A_nso(10) => SHIFT_n_11_10_port, A_nso(9) => 
                           SHIFT_n_11_9_port, A_nso(8) => SHIFT_n_11_8_port, 
                           A_nso(7) => SHIFT_n_11_7_port, A_nso(6) => 
                           SHIFT_n_11_6_port, A_nso(5) => SHIFT_n_11_5_port, 
                           A_nso(4) => SHIFT_n_11_4_port, A_nso(3) => 
                           SHIFT_n_11_3_port, A_nso(2) => SHIFT_n_11_2_port, 
                           A_nso(1) => n_1130, A_nso(0) => n_1131);
   ENC_11 : BOOTHENC_NBIT56_i22 port map( A_s(55) => SHIFT_11_53_port, A_s(54) 
                           => SHIFT_11_53_port, A_s(53) => SHIFT_11_53_port, 
                           A_s(52) => SHIFT_11_52_port, A_s(51) => 
                           SHIFT_11_51_port, A_s(50) => SHIFT_11_50_port, 
                           A_s(49) => SHIFT_11_49_port, A_s(48) => 
                           SHIFT_11_48_port, A_s(47) => SHIFT_11_47_port, 
                           A_s(46) => SHIFT_11_46_port, A_s(45) => 
                           SHIFT_11_45_port, A_s(44) => SHIFT_11_44_port, 
                           A_s(43) => SHIFT_11_43_port, A_s(42) => 
                           SHIFT_11_42_port, A_s(41) => SHIFT_11_41_port, 
                           A_s(40) => SHIFT_11_40_port, A_s(39) => 
                           SHIFT_11_39_port, A_s(38) => SHIFT_11_38_port, 
                           A_s(37) => SHIFT_11_37_port, A_s(36) => 
                           SHIFT_11_36_port, A_s(35) => SHIFT_11_35_port, 
                           A_s(34) => SHIFT_11_34_port, A_s(33) => 
                           SHIFT_11_33_port, A_s(32) => SHIFT_11_32_port, 
                           A_s(31) => SHIFT_11_31_port, A_s(30) => 
                           SHIFT_11_30_port, A_s(29) => SHIFT_11_29_port, 
                           A_s(28) => SHIFT_11_28_port, A_s(27) => 
                           SHIFT_11_27_port, A_s(26) => SHIFT_11_26_port, 
                           A_s(25) => SHIFT_11_25_port, A_s(24) => 
                           SHIFT_11_24_port, A_s(23) => SHIFT_11_23_port, 
                           A_s(22) => SHIFT_11_22_port, A_s(21) => 
                           SHIFT_11_21_port, A_s(20) => SHIFT_11_20_port, 
                           A_s(19) => SHIFT_11_19_port, A_s(18) => 
                           SHIFT_11_18_port, A_s(17) => SHIFT_11_17_port, 
                           A_s(16) => SHIFT_11_16_port, A_s(15) => 
                           SHIFT_11_15_port, A_s(14) => SHIFT_11_14_port, 
                           A_s(13) => SHIFT_11_13_port, A_s(12) => 
                           SHIFT_11_12_port, A_s(11) => SHIFT_11_11_port, 
                           A_s(10) => SHIFT_11_10_port, A_s(9) => 
                           SHIFT_11_9_port, A_s(8) => SHIFT_11_8_port, A_s(7) 
                           => SHIFT_11_7_port, A_s(6) => SHIFT_11_6_port, 
                           A_s(5) => SHIFT_11_5_port, A_s(4) => SHIFT_11_4_port
                           , A_s(3) => SHIFT_11_3_port, A_s(2) => 
                           SHIFT_11_2_port, A_s(1) => SHIFT_11_1_port, A_s(0) 
                           => SHIFT_11_0_port, A_ns(55) => SHIFT_n_11_53_port, 
                           A_ns(54) => SHIFT_n_11_53_port, A_ns(53) => 
                           SHIFT_n_11_53_port, A_ns(52) => SHIFT_n_11_52_port, 
                           A_ns(51) => SHIFT_n_11_51_port, A_ns(50) => 
                           SHIFT_n_11_50_port, A_ns(49) => SHIFT_n_11_49_port, 
                           A_ns(48) => SHIFT_n_11_48_port, A_ns(47) => 
                           SHIFT_n_11_47_port, A_ns(46) => SHIFT_n_11_46_port, 
                           A_ns(45) => SHIFT_n_11_45_port, A_ns(44) => 
                           SHIFT_n_11_44_port, A_ns(43) => SHIFT_n_11_43_port, 
                           A_ns(42) => SHIFT_n_11_42_port, A_ns(41) => 
                           SHIFT_n_11_41_port, A_ns(40) => SHIFT_n_11_40_port, 
                           A_ns(39) => SHIFT_n_11_39_port, A_ns(38) => 
                           SHIFT_n_11_38_port, A_ns(37) => SHIFT_n_11_37_port, 
                           A_ns(36) => SHIFT_n_11_36_port, A_ns(35) => 
                           SHIFT_n_11_35_port, A_ns(34) => SHIFT_n_11_34_port, 
                           A_ns(33) => SHIFT_n_11_33_port, A_ns(32) => 
                           SHIFT_n_11_32_port, A_ns(31) => SHIFT_n_11_31_port, 
                           A_ns(30) => SHIFT_n_11_30_port, A_ns(29) => 
                           SHIFT_n_11_29_port, A_ns(28) => SHIFT_n_11_28_port, 
                           A_ns(27) => SHIFT_n_11_27_port, A_ns(26) => 
                           SHIFT_n_11_26_port, A_ns(25) => SHIFT_n_11_25_port, 
                           A_ns(24) => SHIFT_n_11_24_port, A_ns(23) => 
                           SHIFT_n_11_23_port, A_ns(22) => SHIFT_n_11_22_port, 
                           A_ns(21) => SHIFT_n_11_21_port, A_ns(20) => 
                           SHIFT_n_11_20_port, A_ns(19) => SHIFT_n_11_19_port, 
                           A_ns(18) => SHIFT_n_11_18_port, A_ns(17) => 
                           SHIFT_n_11_17_port, A_ns(16) => SHIFT_n_11_16_port, 
                           A_ns(15) => SHIFT_n_11_15_port, A_ns(14) => 
                           SHIFT_n_11_14_port, A_ns(13) => SHIFT_n_11_13_port, 
                           A_ns(12) => SHIFT_n_11_12_port, A_ns(11) => 
                           SHIFT_n_11_11_port, A_ns(10) => SHIFT_n_11_10_port, 
                           A_ns(9) => SHIFT_n_11_9_port, A_ns(8) => 
                           SHIFT_n_11_8_port, A_ns(7) => SHIFT_n_11_7_port, 
                           A_ns(6) => SHIFT_n_11_6_port, A_ns(5) => 
                           SHIFT_n_11_5_port, A_ns(4) => SHIFT_n_11_4_port, 
                           A_ns(3) => SHIFT_n_11_3_port, A_ns(2) => 
                           SHIFT_n_11_2_port, A_ns(1) => SHIFT_n_11_1_port, 
                           A_ns(0) => SHIFT_n_11_0_port, B(55) => B(31), B(54) 
                           => B(31), B(53) => B(31), B(52) => B(31), B(51) => 
                           B(31), B(50) => B(31), B(49) => B(31), B(48) => 
                           B(31), B(47) => B(31), B(46) => B(31), B(45) => 
                           B(31), B(44) => B(31), B(43) => B(31), B(42) => 
                           B(31), B(41) => B(31), B(40) => B(31), B(39) => 
                           B(31), B(38) => B(31), B(37) => B(31), B(36) => 
                           B(31), B(35) => B(31), B(34) => B(31), B(33) => 
                           B(31), B(32) => B(31), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), O(55) => OTMP_11_55_port, 
                           O(54) => OTMP_11_54_port, O(53) => OTMP_11_53_port, 
                           O(52) => OTMP_11_52_port, O(51) => OTMP_11_51_port, 
                           O(50) => OTMP_11_50_port, O(49) => OTMP_11_49_port, 
                           O(48) => OTMP_11_48_port, O(47) => OTMP_11_47_port, 
                           O(46) => OTMP_11_46_port, O(45) => OTMP_11_45_port, 
                           O(44) => OTMP_11_44_port, O(43) => OTMP_11_43_port, 
                           O(42) => OTMP_11_42_port, O(41) => OTMP_11_41_port, 
                           O(40) => OTMP_11_40_port, O(39) => OTMP_11_39_port, 
                           O(38) => OTMP_11_38_port, O(37) => OTMP_11_37_port, 
                           O(36) => OTMP_11_36_port, O(35) => OTMP_11_35_port, 
                           O(34) => OTMP_11_34_port, O(33) => OTMP_11_33_port, 
                           O(32) => OTMP_11_32_port, O(31) => OTMP_11_31_port, 
                           O(30) => OTMP_11_30_port, O(29) => OTMP_11_29_port, 
                           O(28) => OTMP_11_28_port, O(27) => OTMP_11_27_port, 
                           O(26) => OTMP_11_26_port, O(25) => OTMP_11_25_port, 
                           O(24) => OTMP_11_24_port, O(23) => OTMP_11_23_port, 
                           O(22) => OTMP_11_22_port, O(21) => OTMP_11_21_port, 
                           O(20) => OTMP_11_20_port, O(19) => OTMP_11_19_port, 
                           O(18) => OTMP_11_18_port, O(17) => OTMP_11_17_port, 
                           O(16) => OTMP_11_16_port, O(15) => OTMP_11_15_port, 
                           O(14) => OTMP_11_14_port, O(13) => OTMP_11_13_port, 
                           O(12) => OTMP_11_12_port, O(11) => OTMP_11_11_port, 
                           O(10) => OTMP_11_10_port, O(9) => OTMP_11_9_port, 
                           O(8) => OTMP_11_8_port, O(7) => OTMP_11_7_port, O(6)
                           => OTMP_11_6_port, O(5) => OTMP_11_5_port, O(4) => 
                           OTMP_11_4_port, O(3) => OTMP_11_3_port, O(2) => 
                           OTMP_11_2_port, O(1) => OTMP_11_1_port, O(0) => 
                           n_1132, A_so(55) => SHIFT_12_55_port, A_so(54) => 
                           SHIFT_12_54_port, A_so(53) => SHIFT_12_53_port, 
                           A_so(52) => SHIFT_12_52_port, A_so(51) => 
                           SHIFT_12_51_port, A_so(50) => SHIFT_12_50_port, 
                           A_so(49) => SHIFT_12_49_port, A_so(48) => 
                           SHIFT_12_48_port, A_so(47) => SHIFT_12_47_port, 
                           A_so(46) => SHIFT_12_46_port, A_so(45) => 
                           SHIFT_12_45_port, A_so(44) => SHIFT_12_44_port, 
                           A_so(43) => SHIFT_12_43_port, A_so(42) => 
                           SHIFT_12_42_port, A_so(41) => SHIFT_12_41_port, 
                           A_so(40) => SHIFT_12_40_port, A_so(39) => 
                           SHIFT_12_39_port, A_so(38) => SHIFT_12_38_port, 
                           A_so(37) => SHIFT_12_37_port, A_so(36) => 
                           SHIFT_12_36_port, A_so(35) => SHIFT_12_35_port, 
                           A_so(34) => SHIFT_12_34_port, A_so(33) => 
                           SHIFT_12_33_port, A_so(32) => SHIFT_12_32_port, 
                           A_so(31) => SHIFT_12_31_port, A_so(30) => 
                           SHIFT_12_30_port, A_so(29) => SHIFT_12_29_port, 
                           A_so(28) => SHIFT_12_28_port, A_so(27) => 
                           SHIFT_12_27_port, A_so(26) => SHIFT_12_26_port, 
                           A_so(25) => SHIFT_12_25_port, A_so(24) => 
                           SHIFT_12_24_port, A_so(23) => SHIFT_12_23_port, 
                           A_so(22) => SHIFT_12_22_port, A_so(21) => 
                           SHIFT_12_21_port, A_so(20) => SHIFT_12_20_port, 
                           A_so(19) => SHIFT_12_19_port, A_so(18) => 
                           SHIFT_12_18_port, A_so(17) => SHIFT_12_17_port, 
                           A_so(16) => SHIFT_12_16_port, A_so(15) => 
                           SHIFT_12_15_port, A_so(14) => SHIFT_12_14_port, 
                           A_so(13) => SHIFT_12_13_port, A_so(12) => 
                           SHIFT_12_12_port, A_so(11) => SHIFT_12_11_port, 
                           A_so(10) => SHIFT_12_10_port, A_so(9) => 
                           SHIFT_12_9_port, A_so(8) => SHIFT_12_8_port, A_so(7)
                           => SHIFT_12_7_port, A_so(6) => SHIFT_12_6_port, 
                           A_so(5) => SHIFT_12_5_port, A_so(4) => 
                           SHIFT_12_4_port, A_so(3) => SHIFT_12_3_port, A_so(2)
                           => SHIFT_12_2_port, A_so(1) => n_1133, A_so(0) => 
                           n_1134, A_nso(55) => SHIFT_n_12_55_port, A_nso(54) 
                           => SHIFT_n_12_54_port, A_nso(53) => 
                           SHIFT_n_12_53_port, A_nso(52) => SHIFT_n_12_52_port,
                           A_nso(51) => SHIFT_n_12_51_port, A_nso(50) => 
                           SHIFT_n_12_50_port, A_nso(49) => SHIFT_n_12_49_port,
                           A_nso(48) => SHIFT_n_12_48_port, A_nso(47) => 
                           SHIFT_n_12_47_port, A_nso(46) => SHIFT_n_12_46_port,
                           A_nso(45) => SHIFT_n_12_45_port, A_nso(44) => 
                           SHIFT_n_12_44_port, A_nso(43) => SHIFT_n_12_43_port,
                           A_nso(42) => SHIFT_n_12_42_port, A_nso(41) => 
                           SHIFT_n_12_41_port, A_nso(40) => SHIFT_n_12_40_port,
                           A_nso(39) => SHIFT_n_12_39_port, A_nso(38) => 
                           SHIFT_n_12_38_port, A_nso(37) => SHIFT_n_12_37_port,
                           A_nso(36) => SHIFT_n_12_36_port, A_nso(35) => 
                           SHIFT_n_12_35_port, A_nso(34) => SHIFT_n_12_34_port,
                           A_nso(33) => SHIFT_n_12_33_port, A_nso(32) => 
                           SHIFT_n_12_32_port, A_nso(31) => SHIFT_n_12_31_port,
                           A_nso(30) => SHIFT_n_12_30_port, A_nso(29) => 
                           SHIFT_n_12_29_port, A_nso(28) => SHIFT_n_12_28_port,
                           A_nso(27) => SHIFT_n_12_27_port, A_nso(26) => 
                           SHIFT_n_12_26_port, A_nso(25) => SHIFT_n_12_25_port,
                           A_nso(24) => SHIFT_n_12_24_port, A_nso(23) => 
                           SHIFT_n_12_23_port, A_nso(22) => SHIFT_n_12_22_port,
                           A_nso(21) => SHIFT_n_12_21_port, A_nso(20) => 
                           SHIFT_n_12_20_port, A_nso(19) => SHIFT_n_12_19_port,
                           A_nso(18) => SHIFT_n_12_18_port, A_nso(17) => 
                           SHIFT_n_12_17_port, A_nso(16) => SHIFT_n_12_16_port,
                           A_nso(15) => SHIFT_n_12_15_port, A_nso(14) => 
                           SHIFT_n_12_14_port, A_nso(13) => SHIFT_n_12_13_port,
                           A_nso(12) => SHIFT_n_12_12_port, A_nso(11) => 
                           SHIFT_n_12_11_port, A_nso(10) => SHIFT_n_12_10_port,
                           A_nso(9) => SHIFT_n_12_9_port, A_nso(8) => 
                           SHIFT_n_12_8_port, A_nso(7) => SHIFT_n_12_7_port, 
                           A_nso(6) => SHIFT_n_12_6_port, A_nso(5) => 
                           SHIFT_n_12_5_port, A_nso(4) => SHIFT_n_12_4_port, 
                           A_nso(3) => SHIFT_n_12_3_port, A_nso(2) => 
                           SHIFT_n_12_2_port, A_nso(1) => n_1135, A_nso(0) => 
                           n_1136);
   ENC_12 : BOOTHENC_NBIT58_i24 port map( A_s(57) => SHIFT_12_55_port, A_s(56) 
                           => SHIFT_12_55_port, A_s(55) => SHIFT_12_55_port, 
                           A_s(54) => SHIFT_12_54_port, A_s(53) => 
                           SHIFT_12_53_port, A_s(52) => SHIFT_12_52_port, 
                           A_s(51) => SHIFT_12_51_port, A_s(50) => 
                           SHIFT_12_50_port, A_s(49) => SHIFT_12_49_port, 
                           A_s(48) => SHIFT_12_48_port, A_s(47) => 
                           SHIFT_12_47_port, A_s(46) => SHIFT_12_46_port, 
                           A_s(45) => SHIFT_12_45_port, A_s(44) => 
                           SHIFT_12_44_port, A_s(43) => SHIFT_12_43_port, 
                           A_s(42) => SHIFT_12_42_port, A_s(41) => 
                           SHIFT_12_41_port, A_s(40) => SHIFT_12_40_port, 
                           A_s(39) => SHIFT_12_39_port, A_s(38) => 
                           SHIFT_12_38_port, A_s(37) => SHIFT_12_37_port, 
                           A_s(36) => SHIFT_12_36_port, A_s(35) => 
                           SHIFT_12_35_port, A_s(34) => SHIFT_12_34_port, 
                           A_s(33) => SHIFT_12_33_port, A_s(32) => 
                           SHIFT_12_32_port, A_s(31) => SHIFT_12_31_port, 
                           A_s(30) => SHIFT_12_30_port, A_s(29) => 
                           SHIFT_12_29_port, A_s(28) => SHIFT_12_28_port, 
                           A_s(27) => SHIFT_12_27_port, A_s(26) => 
                           SHIFT_12_26_port, A_s(25) => SHIFT_12_25_port, 
                           A_s(24) => SHIFT_12_24_port, A_s(23) => 
                           SHIFT_12_23_port, A_s(22) => SHIFT_12_22_port, 
                           A_s(21) => SHIFT_12_21_port, A_s(20) => 
                           SHIFT_12_20_port, A_s(19) => SHIFT_12_19_port, 
                           A_s(18) => SHIFT_12_18_port, A_s(17) => 
                           SHIFT_12_17_port, A_s(16) => SHIFT_12_16_port, 
                           A_s(15) => SHIFT_12_15_port, A_s(14) => 
                           SHIFT_12_14_port, A_s(13) => SHIFT_12_13_port, 
                           A_s(12) => SHIFT_12_12_port, A_s(11) => 
                           SHIFT_12_11_port, A_s(10) => SHIFT_12_10_port, 
                           A_s(9) => SHIFT_12_9_port, A_s(8) => SHIFT_12_8_port
                           , A_s(7) => SHIFT_12_7_port, A_s(6) => 
                           SHIFT_12_6_port, A_s(5) => SHIFT_12_5_port, A_s(4) 
                           => SHIFT_12_4_port, A_s(3) => SHIFT_12_3_port, 
                           A_s(2) => SHIFT_12_2_port, A_s(1) => SHIFT_12_1_port
                           , A_s(0) => SHIFT_12_0_port, A_ns(57) => 
                           SHIFT_n_12_55_port, A_ns(56) => SHIFT_n_12_55_port, 
                           A_ns(55) => SHIFT_n_12_55_port, A_ns(54) => 
                           SHIFT_n_12_54_port, A_ns(53) => SHIFT_n_12_53_port, 
                           A_ns(52) => SHIFT_n_12_52_port, A_ns(51) => 
                           SHIFT_n_12_51_port, A_ns(50) => SHIFT_n_12_50_port, 
                           A_ns(49) => SHIFT_n_12_49_port, A_ns(48) => 
                           SHIFT_n_12_48_port, A_ns(47) => SHIFT_n_12_47_port, 
                           A_ns(46) => SHIFT_n_12_46_port, A_ns(45) => 
                           SHIFT_n_12_45_port, A_ns(44) => SHIFT_n_12_44_port, 
                           A_ns(43) => SHIFT_n_12_43_port, A_ns(42) => 
                           SHIFT_n_12_42_port, A_ns(41) => SHIFT_n_12_41_port, 
                           A_ns(40) => SHIFT_n_12_40_port, A_ns(39) => 
                           SHIFT_n_12_39_port, A_ns(38) => SHIFT_n_12_38_port, 
                           A_ns(37) => SHIFT_n_12_37_port, A_ns(36) => 
                           SHIFT_n_12_36_port, A_ns(35) => SHIFT_n_12_35_port, 
                           A_ns(34) => SHIFT_n_12_34_port, A_ns(33) => 
                           SHIFT_n_12_33_port, A_ns(32) => SHIFT_n_12_32_port, 
                           A_ns(31) => SHIFT_n_12_31_port, A_ns(30) => 
                           SHIFT_n_12_30_port, A_ns(29) => SHIFT_n_12_29_port, 
                           A_ns(28) => SHIFT_n_12_28_port, A_ns(27) => 
                           SHIFT_n_12_27_port, A_ns(26) => SHIFT_n_12_26_port, 
                           A_ns(25) => SHIFT_n_12_25_port, A_ns(24) => 
                           SHIFT_n_12_24_port, A_ns(23) => SHIFT_n_12_23_port, 
                           A_ns(22) => SHIFT_n_12_22_port, A_ns(21) => 
                           SHIFT_n_12_21_port, A_ns(20) => SHIFT_n_12_20_port, 
                           A_ns(19) => SHIFT_n_12_19_port, A_ns(18) => 
                           SHIFT_n_12_18_port, A_ns(17) => SHIFT_n_12_17_port, 
                           A_ns(16) => SHIFT_n_12_16_port, A_ns(15) => 
                           SHIFT_n_12_15_port, A_ns(14) => SHIFT_n_12_14_port, 
                           A_ns(13) => SHIFT_n_12_13_port, A_ns(12) => 
                           SHIFT_n_12_12_port, A_ns(11) => SHIFT_n_12_11_port, 
                           A_ns(10) => SHIFT_n_12_10_port, A_ns(9) => 
                           SHIFT_n_12_9_port, A_ns(8) => SHIFT_n_12_8_port, 
                           A_ns(7) => SHIFT_n_12_7_port, A_ns(6) => 
                           SHIFT_n_12_6_port, A_ns(5) => SHIFT_n_12_5_port, 
                           A_ns(4) => SHIFT_n_12_4_port, A_ns(3) => 
                           SHIFT_n_12_3_port, A_ns(2) => SHIFT_n_12_2_port, 
                           A_ns(1) => SHIFT_n_12_1_port, A_ns(0) => 
                           SHIFT_n_12_0_port, B(57) => B(31), B(56) => B(31), 
                           B(55) => B(31), B(54) => B(31), B(53) => B(31), 
                           B(52) => B(31), B(51) => B(31), B(50) => B(31), 
                           B(49) => B(31), B(48) => B(31), B(47) => B(31), 
                           B(46) => B(31), B(45) => B(31), B(44) => B(31), 
                           B(43) => B(31), B(42) => B(31), B(41) => B(31), 
                           B(40) => B(31), B(39) => B(31), B(38) => B(31), 
                           B(37) => B(31), B(36) => B(31), B(35) => B(31), 
                           B(34) => B(31), B(33) => B(31), B(32) => B(31), 
                           B(31) => B(31), B(30) => B(30), B(29) => B(29), 
                           B(28) => B(28), B(27) => B(27), B(26) => B(26), 
                           B(25) => B(25), B(24) => B(24), B(23) => B(23), 
                           B(22) => B(22), B(21) => B(21), B(20) => B(20), 
                           B(19) => B(19), B(18) => B(18), B(17) => B(17), 
                           B(16) => B(16), B(15) => B(15), B(14) => B(14), 
                           B(13) => B(13), B(12) => B(12), B(11) => B(11), 
                           B(10) => B(10), B(9) => B(9), B(8) => B(8), B(7) => 
                           B(7), B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3)
                           => B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), 
                           O(57) => OTMP_12_57_port, O(56) => OTMP_12_56_port, 
                           O(55) => OTMP_12_55_port, O(54) => OTMP_12_54_port, 
                           O(53) => OTMP_12_53_port, O(52) => OTMP_12_52_port, 
                           O(51) => OTMP_12_51_port, O(50) => OTMP_12_50_port, 
                           O(49) => OTMP_12_49_port, O(48) => OTMP_12_48_port, 
                           O(47) => OTMP_12_47_port, O(46) => OTMP_12_46_port, 
                           O(45) => OTMP_12_45_port, O(44) => OTMP_12_44_port, 
                           O(43) => OTMP_12_43_port, O(42) => OTMP_12_42_port, 
                           O(41) => OTMP_12_41_port, O(40) => OTMP_12_40_port, 
                           O(39) => OTMP_12_39_port, O(38) => OTMP_12_38_port, 
                           O(37) => OTMP_12_37_port, O(36) => OTMP_12_36_port, 
                           O(35) => OTMP_12_35_port, O(34) => OTMP_12_34_port, 
                           O(33) => OTMP_12_33_port, O(32) => OTMP_12_32_port, 
                           O(31) => OTMP_12_31_port, O(30) => OTMP_12_30_port, 
                           O(29) => OTMP_12_29_port, O(28) => OTMP_12_28_port, 
                           O(27) => OTMP_12_27_port, O(26) => OTMP_12_26_port, 
                           O(25) => OTMP_12_25_port, O(24) => OTMP_12_24_port, 
                           O(23) => OTMP_12_23_port, O(22) => OTMP_12_22_port, 
                           O(21) => OTMP_12_21_port, O(20) => OTMP_12_20_port, 
                           O(19) => OTMP_12_19_port, O(18) => OTMP_12_18_port, 
                           O(17) => OTMP_12_17_port, O(16) => OTMP_12_16_port, 
                           O(15) => OTMP_12_15_port, O(14) => OTMP_12_14_port, 
                           O(13) => OTMP_12_13_port, O(12) => OTMP_12_12_port, 
                           O(11) => OTMP_12_11_port, O(10) => OTMP_12_10_port, 
                           O(9) => OTMP_12_9_port, O(8) => OTMP_12_8_port, O(7)
                           => OTMP_12_7_port, O(6) => OTMP_12_6_port, O(5) => 
                           OTMP_12_5_port, O(4) => OTMP_12_4_port, O(3) => 
                           OTMP_12_3_port, O(2) => OTMP_12_2_port, O(1) => 
                           OTMP_12_1_port, O(0) => n_1137, A_so(57) => 
                           SHIFT_13_57_port, A_so(56) => SHIFT_13_56_port, 
                           A_so(55) => SHIFT_13_55_port, A_so(54) => 
                           SHIFT_13_54_port, A_so(53) => SHIFT_13_53_port, 
                           A_so(52) => SHIFT_13_52_port, A_so(51) => 
                           SHIFT_13_51_port, A_so(50) => SHIFT_13_50_port, 
                           A_so(49) => SHIFT_13_49_port, A_so(48) => 
                           SHIFT_13_48_port, A_so(47) => SHIFT_13_47_port, 
                           A_so(46) => SHIFT_13_46_port, A_so(45) => 
                           SHIFT_13_45_port, A_so(44) => SHIFT_13_44_port, 
                           A_so(43) => SHIFT_13_43_port, A_so(42) => 
                           SHIFT_13_42_port, A_so(41) => SHIFT_13_41_port, 
                           A_so(40) => SHIFT_13_40_port, A_so(39) => 
                           SHIFT_13_39_port, A_so(38) => SHIFT_13_38_port, 
                           A_so(37) => SHIFT_13_37_port, A_so(36) => 
                           SHIFT_13_36_port, A_so(35) => SHIFT_13_35_port, 
                           A_so(34) => SHIFT_13_34_port, A_so(33) => 
                           SHIFT_13_33_port, A_so(32) => SHIFT_13_32_port, 
                           A_so(31) => SHIFT_13_31_port, A_so(30) => 
                           SHIFT_13_30_port, A_so(29) => SHIFT_13_29_port, 
                           A_so(28) => SHIFT_13_28_port, A_so(27) => 
                           SHIFT_13_27_port, A_so(26) => SHIFT_13_26_port, 
                           A_so(25) => SHIFT_13_25_port, A_so(24) => 
                           SHIFT_13_24_port, A_so(23) => SHIFT_13_23_port, 
                           A_so(22) => SHIFT_13_22_port, A_so(21) => 
                           SHIFT_13_21_port, A_so(20) => SHIFT_13_20_port, 
                           A_so(19) => SHIFT_13_19_port, A_so(18) => 
                           SHIFT_13_18_port, A_so(17) => SHIFT_13_17_port, 
                           A_so(16) => SHIFT_13_16_port, A_so(15) => 
                           SHIFT_13_15_port, A_so(14) => SHIFT_13_14_port, 
                           A_so(13) => SHIFT_13_13_port, A_so(12) => 
                           SHIFT_13_12_port, A_so(11) => SHIFT_13_11_port, 
                           A_so(10) => SHIFT_13_10_port, A_so(9) => 
                           SHIFT_13_9_port, A_so(8) => SHIFT_13_8_port, A_so(7)
                           => SHIFT_13_7_port, A_so(6) => SHIFT_13_6_port, 
                           A_so(5) => SHIFT_13_5_port, A_so(4) => 
                           SHIFT_13_4_port, A_so(3) => SHIFT_13_3_port, A_so(2)
                           => SHIFT_13_2_port, A_so(1) => n_1138, A_so(0) => 
                           n_1139, A_nso(57) => SHIFT_n_13_57_port, A_nso(56) 
                           => SHIFT_n_13_56_port, A_nso(55) => 
                           SHIFT_n_13_55_port, A_nso(54) => SHIFT_n_13_54_port,
                           A_nso(53) => SHIFT_n_13_53_port, A_nso(52) => 
                           SHIFT_n_13_52_port, A_nso(51) => SHIFT_n_13_51_port,
                           A_nso(50) => SHIFT_n_13_50_port, A_nso(49) => 
                           SHIFT_n_13_49_port, A_nso(48) => SHIFT_n_13_48_port,
                           A_nso(47) => SHIFT_n_13_47_port, A_nso(46) => 
                           SHIFT_n_13_46_port, A_nso(45) => SHIFT_n_13_45_port,
                           A_nso(44) => SHIFT_n_13_44_port, A_nso(43) => 
                           SHIFT_n_13_43_port, A_nso(42) => SHIFT_n_13_42_port,
                           A_nso(41) => SHIFT_n_13_41_port, A_nso(40) => 
                           SHIFT_n_13_40_port, A_nso(39) => SHIFT_n_13_39_port,
                           A_nso(38) => SHIFT_n_13_38_port, A_nso(37) => 
                           SHIFT_n_13_37_port, A_nso(36) => SHIFT_n_13_36_port,
                           A_nso(35) => SHIFT_n_13_35_port, A_nso(34) => 
                           SHIFT_n_13_34_port, A_nso(33) => SHIFT_n_13_33_port,
                           A_nso(32) => SHIFT_n_13_32_port, A_nso(31) => 
                           SHIFT_n_13_31_port, A_nso(30) => SHIFT_n_13_30_port,
                           A_nso(29) => SHIFT_n_13_29_port, A_nso(28) => 
                           SHIFT_n_13_28_port, A_nso(27) => SHIFT_n_13_27_port,
                           A_nso(26) => SHIFT_n_13_26_port, A_nso(25) => 
                           SHIFT_n_13_25_port, A_nso(24) => SHIFT_n_13_24_port,
                           A_nso(23) => SHIFT_n_13_23_port, A_nso(22) => 
                           SHIFT_n_13_22_port, A_nso(21) => SHIFT_n_13_21_port,
                           A_nso(20) => SHIFT_n_13_20_port, A_nso(19) => 
                           SHIFT_n_13_19_port, A_nso(18) => SHIFT_n_13_18_port,
                           A_nso(17) => SHIFT_n_13_17_port, A_nso(16) => 
                           SHIFT_n_13_16_port, A_nso(15) => SHIFT_n_13_15_port,
                           A_nso(14) => SHIFT_n_13_14_port, A_nso(13) => 
                           SHIFT_n_13_13_port, A_nso(12) => SHIFT_n_13_12_port,
                           A_nso(11) => SHIFT_n_13_11_port, A_nso(10) => 
                           SHIFT_n_13_10_port, A_nso(9) => SHIFT_n_13_9_port, 
                           A_nso(8) => SHIFT_n_13_8_port, A_nso(7) => 
                           SHIFT_n_13_7_port, A_nso(6) => SHIFT_n_13_6_port, 
                           A_nso(5) => SHIFT_n_13_5_port, A_nso(4) => 
                           SHIFT_n_13_4_port, A_nso(3) => SHIFT_n_13_3_port, 
                           A_nso(2) => SHIFT_n_13_2_port, A_nso(1) => n_1140, 
                           A_nso(0) => n_1141);
   ENC_13 : BOOTHENC_NBIT60_i26 port map( A_s(59) => SHIFT_13_57_port, A_s(58) 
                           => SHIFT_13_57_port, A_s(57) => SHIFT_13_57_port, 
                           A_s(56) => SHIFT_13_56_port, A_s(55) => 
                           SHIFT_13_55_port, A_s(54) => SHIFT_13_54_port, 
                           A_s(53) => SHIFT_13_53_port, A_s(52) => 
                           SHIFT_13_52_port, A_s(51) => SHIFT_13_51_port, 
                           A_s(50) => SHIFT_13_50_port, A_s(49) => 
                           SHIFT_13_49_port, A_s(48) => SHIFT_13_48_port, 
                           A_s(47) => SHIFT_13_47_port, A_s(46) => 
                           SHIFT_13_46_port, A_s(45) => SHIFT_13_45_port, 
                           A_s(44) => SHIFT_13_44_port, A_s(43) => 
                           SHIFT_13_43_port, A_s(42) => SHIFT_13_42_port, 
                           A_s(41) => SHIFT_13_41_port, A_s(40) => 
                           SHIFT_13_40_port, A_s(39) => SHIFT_13_39_port, 
                           A_s(38) => SHIFT_13_38_port, A_s(37) => 
                           SHIFT_13_37_port, A_s(36) => SHIFT_13_36_port, 
                           A_s(35) => SHIFT_13_35_port, A_s(34) => 
                           SHIFT_13_34_port, A_s(33) => SHIFT_13_33_port, 
                           A_s(32) => SHIFT_13_32_port, A_s(31) => 
                           SHIFT_13_31_port, A_s(30) => SHIFT_13_30_port, 
                           A_s(29) => SHIFT_13_29_port, A_s(28) => 
                           SHIFT_13_28_port, A_s(27) => SHIFT_13_27_port, 
                           A_s(26) => SHIFT_13_26_port, A_s(25) => 
                           SHIFT_13_25_port, A_s(24) => SHIFT_13_24_port, 
                           A_s(23) => SHIFT_13_23_port, A_s(22) => 
                           SHIFT_13_22_port, A_s(21) => SHIFT_13_21_port, 
                           A_s(20) => SHIFT_13_20_port, A_s(19) => 
                           SHIFT_13_19_port, A_s(18) => SHIFT_13_18_port, 
                           A_s(17) => SHIFT_13_17_port, A_s(16) => 
                           SHIFT_13_16_port, A_s(15) => SHIFT_13_15_port, 
                           A_s(14) => SHIFT_13_14_port, A_s(13) => 
                           SHIFT_13_13_port, A_s(12) => SHIFT_13_12_port, 
                           A_s(11) => SHIFT_13_11_port, A_s(10) => 
                           SHIFT_13_10_port, A_s(9) => SHIFT_13_9_port, A_s(8) 
                           => SHIFT_13_8_port, A_s(7) => SHIFT_13_7_port, 
                           A_s(6) => SHIFT_13_6_port, A_s(5) => SHIFT_13_5_port
                           , A_s(4) => SHIFT_13_4_port, A_s(3) => 
                           SHIFT_13_3_port, A_s(2) => SHIFT_13_2_port, A_s(1) 
                           => SHIFT_13_1_port, A_s(0) => SHIFT_13_0_port, 
                           A_ns(59) => SHIFT_n_13_57_port, A_ns(58) => 
                           SHIFT_n_13_57_port, A_ns(57) => SHIFT_n_13_57_port, 
                           A_ns(56) => SHIFT_n_13_56_port, A_ns(55) => 
                           SHIFT_n_13_55_port, A_ns(54) => SHIFT_n_13_54_port, 
                           A_ns(53) => SHIFT_n_13_53_port, A_ns(52) => 
                           SHIFT_n_13_52_port, A_ns(51) => SHIFT_n_13_51_port, 
                           A_ns(50) => SHIFT_n_13_50_port, A_ns(49) => 
                           SHIFT_n_13_49_port, A_ns(48) => SHIFT_n_13_48_port, 
                           A_ns(47) => SHIFT_n_13_47_port, A_ns(46) => 
                           SHIFT_n_13_46_port, A_ns(45) => SHIFT_n_13_45_port, 
                           A_ns(44) => SHIFT_n_13_44_port, A_ns(43) => 
                           SHIFT_n_13_43_port, A_ns(42) => SHIFT_n_13_42_port, 
                           A_ns(41) => SHIFT_n_13_41_port, A_ns(40) => 
                           SHIFT_n_13_40_port, A_ns(39) => SHIFT_n_13_39_port, 
                           A_ns(38) => SHIFT_n_13_38_port, A_ns(37) => 
                           SHIFT_n_13_37_port, A_ns(36) => SHIFT_n_13_36_port, 
                           A_ns(35) => SHIFT_n_13_35_port, A_ns(34) => 
                           SHIFT_n_13_34_port, A_ns(33) => SHIFT_n_13_33_port, 
                           A_ns(32) => SHIFT_n_13_32_port, A_ns(31) => 
                           SHIFT_n_13_31_port, A_ns(30) => SHIFT_n_13_30_port, 
                           A_ns(29) => SHIFT_n_13_29_port, A_ns(28) => 
                           SHIFT_n_13_28_port, A_ns(27) => SHIFT_n_13_27_port, 
                           A_ns(26) => SHIFT_n_13_26_port, A_ns(25) => 
                           SHIFT_n_13_25_port, A_ns(24) => SHIFT_n_13_24_port, 
                           A_ns(23) => SHIFT_n_13_23_port, A_ns(22) => 
                           SHIFT_n_13_22_port, A_ns(21) => SHIFT_n_13_21_port, 
                           A_ns(20) => SHIFT_n_13_20_port, A_ns(19) => 
                           SHIFT_n_13_19_port, A_ns(18) => SHIFT_n_13_18_port, 
                           A_ns(17) => SHIFT_n_13_17_port, A_ns(16) => 
                           SHIFT_n_13_16_port, A_ns(15) => SHIFT_n_13_15_port, 
                           A_ns(14) => SHIFT_n_13_14_port, A_ns(13) => 
                           SHIFT_n_13_13_port, A_ns(12) => SHIFT_n_13_12_port, 
                           A_ns(11) => SHIFT_n_13_11_port, A_ns(10) => 
                           SHIFT_n_13_10_port, A_ns(9) => SHIFT_n_13_9_port, 
                           A_ns(8) => SHIFT_n_13_8_port, A_ns(7) => 
                           SHIFT_n_13_7_port, A_ns(6) => SHIFT_n_13_6_port, 
                           A_ns(5) => SHIFT_n_13_5_port, A_ns(4) => 
                           SHIFT_n_13_4_port, A_ns(3) => SHIFT_n_13_3_port, 
                           A_ns(2) => SHIFT_n_13_2_port, A_ns(1) => 
                           SHIFT_n_13_1_port, A_ns(0) => SHIFT_n_13_0_port, 
                           B(59) => B(31), B(58) => B(31), B(57) => B(31), 
                           B(56) => B(31), B(55) => B(31), B(54) => B(31), 
                           B(53) => B(31), B(52) => B(31), B(51) => B(31), 
                           B(50) => B(31), B(49) => B(31), B(48) => B(31), 
                           B(47) => B(31), B(46) => B(31), B(45) => B(31), 
                           B(44) => B(31), B(43) => B(31), B(42) => B(31), 
                           B(41) => B(31), B(40) => B(31), B(39) => B(31), 
                           B(38) => B(31), B(37) => B(31), B(36) => B(31), 
                           B(35) => B(31), B(34) => B(31), B(33) => B(31), 
                           B(32) => B(31), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), O(59) => OTMP_13_59_port, O(58) 
                           => OTMP_13_58_port, O(57) => OTMP_13_57_port, O(56) 
                           => OTMP_13_56_port, O(55) => OTMP_13_55_port, O(54) 
                           => OTMP_13_54_port, O(53) => OTMP_13_53_port, O(52) 
                           => OTMP_13_52_port, O(51) => OTMP_13_51_port, O(50) 
                           => OTMP_13_50_port, O(49) => OTMP_13_49_port, O(48) 
                           => OTMP_13_48_port, O(47) => OTMP_13_47_port, O(46) 
                           => OTMP_13_46_port, O(45) => OTMP_13_45_port, O(44) 
                           => OTMP_13_44_port, O(43) => OTMP_13_43_port, O(42) 
                           => OTMP_13_42_port, O(41) => OTMP_13_41_port, O(40) 
                           => OTMP_13_40_port, O(39) => OTMP_13_39_port, O(38) 
                           => OTMP_13_38_port, O(37) => OTMP_13_37_port, O(36) 
                           => OTMP_13_36_port, O(35) => OTMP_13_35_port, O(34) 
                           => OTMP_13_34_port, O(33) => OTMP_13_33_port, O(32) 
                           => OTMP_13_32_port, O(31) => OTMP_13_31_port, O(30) 
                           => OTMP_13_30_port, O(29) => OTMP_13_29_port, O(28) 
                           => OTMP_13_28_port, O(27) => OTMP_13_27_port, O(26) 
                           => OTMP_13_26_port, O(25) => OTMP_13_25_port, O(24) 
                           => OTMP_13_24_port, O(23) => OTMP_13_23_port, O(22) 
                           => OTMP_13_22_port, O(21) => OTMP_13_21_port, O(20) 
                           => OTMP_13_20_port, O(19) => OTMP_13_19_port, O(18) 
                           => OTMP_13_18_port, O(17) => OTMP_13_17_port, O(16) 
                           => OTMP_13_16_port, O(15) => OTMP_13_15_port, O(14) 
                           => OTMP_13_14_port, O(13) => OTMP_13_13_port, O(12) 
                           => OTMP_13_12_port, O(11) => OTMP_13_11_port, O(10) 
                           => OTMP_13_10_port, O(9) => OTMP_13_9_port, O(8) => 
                           OTMP_13_8_port, O(7) => OTMP_13_7_port, O(6) => 
                           OTMP_13_6_port, O(5) => OTMP_13_5_port, O(4) => 
                           OTMP_13_4_port, O(3) => OTMP_13_3_port, O(2) => 
                           OTMP_13_2_port, O(1) => OTMP_13_1_port, O(0) => 
                           n_1142, A_so(59) => SHIFT_14_59_port, A_so(58) => 
                           SHIFT_14_58_port, A_so(57) => SHIFT_14_57_port, 
                           A_so(56) => SHIFT_14_56_port, A_so(55) => 
                           SHIFT_14_55_port, A_so(54) => SHIFT_14_54_port, 
                           A_so(53) => SHIFT_14_53_port, A_so(52) => 
                           SHIFT_14_52_port, A_so(51) => SHIFT_14_51_port, 
                           A_so(50) => SHIFT_14_50_port, A_so(49) => 
                           SHIFT_14_49_port, A_so(48) => SHIFT_14_48_port, 
                           A_so(47) => SHIFT_14_47_port, A_so(46) => 
                           SHIFT_14_46_port, A_so(45) => SHIFT_14_45_port, 
                           A_so(44) => SHIFT_14_44_port, A_so(43) => 
                           SHIFT_14_43_port, A_so(42) => SHIFT_14_42_port, 
                           A_so(41) => SHIFT_14_41_port, A_so(40) => 
                           SHIFT_14_40_port, A_so(39) => SHIFT_14_39_port, 
                           A_so(38) => SHIFT_14_38_port, A_so(37) => 
                           SHIFT_14_37_port, A_so(36) => SHIFT_14_36_port, 
                           A_so(35) => SHIFT_14_35_port, A_so(34) => 
                           SHIFT_14_34_port, A_so(33) => SHIFT_14_33_port, 
                           A_so(32) => SHIFT_14_32_port, A_so(31) => 
                           SHIFT_14_31_port, A_so(30) => SHIFT_14_30_port, 
                           A_so(29) => SHIFT_14_29_port, A_so(28) => 
                           SHIFT_14_28_port, A_so(27) => SHIFT_14_27_port, 
                           A_so(26) => SHIFT_14_26_port, A_so(25) => 
                           SHIFT_14_25_port, A_so(24) => SHIFT_14_24_port, 
                           A_so(23) => SHIFT_14_23_port, A_so(22) => 
                           SHIFT_14_22_port, A_so(21) => SHIFT_14_21_port, 
                           A_so(20) => SHIFT_14_20_port, A_so(19) => 
                           SHIFT_14_19_port, A_so(18) => SHIFT_14_18_port, 
                           A_so(17) => SHIFT_14_17_port, A_so(16) => 
                           SHIFT_14_16_port, A_so(15) => SHIFT_14_15_port, 
                           A_so(14) => SHIFT_14_14_port, A_so(13) => 
                           SHIFT_14_13_port, A_so(12) => SHIFT_14_12_port, 
                           A_so(11) => SHIFT_14_11_port, A_so(10) => 
                           SHIFT_14_10_port, A_so(9) => SHIFT_14_9_port, 
                           A_so(8) => SHIFT_14_8_port, A_so(7) => 
                           SHIFT_14_7_port, A_so(6) => SHIFT_14_6_port, A_so(5)
                           => SHIFT_14_5_port, A_so(4) => SHIFT_14_4_port, 
                           A_so(3) => SHIFT_14_3_port, A_so(2) => 
                           SHIFT_14_2_port, A_so(1) => n_1143, A_so(0) => 
                           n_1144, A_nso(59) => SHIFT_n_14_59_port, A_nso(58) 
                           => SHIFT_n_14_58_port, A_nso(57) => 
                           SHIFT_n_14_57_port, A_nso(56) => SHIFT_n_14_56_port,
                           A_nso(55) => SHIFT_n_14_55_port, A_nso(54) => 
                           SHIFT_n_14_54_port, A_nso(53) => SHIFT_n_14_53_port,
                           A_nso(52) => SHIFT_n_14_52_port, A_nso(51) => 
                           SHIFT_n_14_51_port, A_nso(50) => SHIFT_n_14_50_port,
                           A_nso(49) => SHIFT_n_14_49_port, A_nso(48) => 
                           SHIFT_n_14_48_port, A_nso(47) => SHIFT_n_14_47_port,
                           A_nso(46) => SHIFT_n_14_46_port, A_nso(45) => 
                           SHIFT_n_14_45_port, A_nso(44) => SHIFT_n_14_44_port,
                           A_nso(43) => SHIFT_n_14_43_port, A_nso(42) => 
                           SHIFT_n_14_42_port, A_nso(41) => SHIFT_n_14_41_port,
                           A_nso(40) => SHIFT_n_14_40_port, A_nso(39) => 
                           SHIFT_n_14_39_port, A_nso(38) => SHIFT_n_14_38_port,
                           A_nso(37) => SHIFT_n_14_37_port, A_nso(36) => 
                           SHIFT_n_14_36_port, A_nso(35) => SHIFT_n_14_35_port,
                           A_nso(34) => SHIFT_n_14_34_port, A_nso(33) => 
                           SHIFT_n_14_33_port, A_nso(32) => SHIFT_n_14_32_port,
                           A_nso(31) => SHIFT_n_14_31_port, A_nso(30) => 
                           SHIFT_n_14_30_port, A_nso(29) => SHIFT_n_14_29_port,
                           A_nso(28) => SHIFT_n_14_28_port, A_nso(27) => 
                           SHIFT_n_14_27_port, A_nso(26) => SHIFT_n_14_26_port,
                           A_nso(25) => SHIFT_n_14_25_port, A_nso(24) => 
                           SHIFT_n_14_24_port, A_nso(23) => SHIFT_n_14_23_port,
                           A_nso(22) => SHIFT_n_14_22_port, A_nso(21) => 
                           SHIFT_n_14_21_port, A_nso(20) => SHIFT_n_14_20_port,
                           A_nso(19) => SHIFT_n_14_19_port, A_nso(18) => 
                           SHIFT_n_14_18_port, A_nso(17) => SHIFT_n_14_17_port,
                           A_nso(16) => SHIFT_n_14_16_port, A_nso(15) => 
                           SHIFT_n_14_15_port, A_nso(14) => SHIFT_n_14_14_port,
                           A_nso(13) => SHIFT_n_14_13_port, A_nso(12) => 
                           SHIFT_n_14_12_port, A_nso(11) => SHIFT_n_14_11_port,
                           A_nso(10) => SHIFT_n_14_10_port, A_nso(9) => 
                           SHIFT_n_14_9_port, A_nso(8) => SHIFT_n_14_8_port, 
                           A_nso(7) => SHIFT_n_14_7_port, A_nso(6) => 
                           SHIFT_n_14_6_port, A_nso(5) => SHIFT_n_14_5_port, 
                           A_nso(4) => SHIFT_n_14_4_port, A_nso(3) => 
                           SHIFT_n_14_3_port, A_nso(2) => SHIFT_n_14_2_port, 
                           A_nso(1) => n_1145, A_nso(0) => n_1146);
   ENC_14 : BOOTHENC_NBIT62_i28 port map( A_s(61) => SHIFT_14_59_port, A_s(60) 
                           => SHIFT_14_59_port, A_s(59) => SHIFT_14_59_port, 
                           A_s(58) => SHIFT_14_58_port, A_s(57) => 
                           SHIFT_14_57_port, A_s(56) => SHIFT_14_56_port, 
                           A_s(55) => SHIFT_14_55_port, A_s(54) => 
                           SHIFT_14_54_port, A_s(53) => SHIFT_14_53_port, 
                           A_s(52) => SHIFT_14_52_port, A_s(51) => 
                           SHIFT_14_51_port, A_s(50) => SHIFT_14_50_port, 
                           A_s(49) => SHIFT_14_49_port, A_s(48) => 
                           SHIFT_14_48_port, A_s(47) => SHIFT_14_47_port, 
                           A_s(46) => SHIFT_14_46_port, A_s(45) => 
                           SHIFT_14_45_port, A_s(44) => SHIFT_14_44_port, 
                           A_s(43) => SHIFT_14_43_port, A_s(42) => 
                           SHIFT_14_42_port, A_s(41) => SHIFT_14_41_port, 
                           A_s(40) => SHIFT_14_40_port, A_s(39) => 
                           SHIFT_14_39_port, A_s(38) => SHIFT_14_38_port, 
                           A_s(37) => SHIFT_14_37_port, A_s(36) => 
                           SHIFT_14_36_port, A_s(35) => SHIFT_14_35_port, 
                           A_s(34) => SHIFT_14_34_port, A_s(33) => 
                           SHIFT_14_33_port, A_s(32) => SHIFT_14_32_port, 
                           A_s(31) => SHIFT_14_31_port, A_s(30) => 
                           SHIFT_14_30_port, A_s(29) => SHIFT_14_29_port, 
                           A_s(28) => SHIFT_14_28_port, A_s(27) => 
                           SHIFT_14_27_port, A_s(26) => SHIFT_14_26_port, 
                           A_s(25) => SHIFT_14_25_port, A_s(24) => 
                           SHIFT_14_24_port, A_s(23) => SHIFT_14_23_port, 
                           A_s(22) => SHIFT_14_22_port, A_s(21) => 
                           SHIFT_14_21_port, A_s(20) => SHIFT_14_20_port, 
                           A_s(19) => SHIFT_14_19_port, A_s(18) => 
                           SHIFT_14_18_port, A_s(17) => SHIFT_14_17_port, 
                           A_s(16) => SHIFT_14_16_port, A_s(15) => 
                           SHIFT_14_15_port, A_s(14) => SHIFT_14_14_port, 
                           A_s(13) => SHIFT_14_13_port, A_s(12) => 
                           SHIFT_14_12_port, A_s(11) => SHIFT_14_11_port, 
                           A_s(10) => SHIFT_14_10_port, A_s(9) => 
                           SHIFT_14_9_port, A_s(8) => SHIFT_14_8_port, A_s(7) 
                           => SHIFT_14_7_port, A_s(6) => SHIFT_14_6_port, 
                           A_s(5) => SHIFT_14_5_port, A_s(4) => SHIFT_14_4_port
                           , A_s(3) => SHIFT_14_3_port, A_s(2) => 
                           SHIFT_14_2_port, A_s(1) => SHIFT_14_1_port, A_s(0) 
                           => SHIFT_14_0_port, A_ns(61) => SHIFT_n_14_59_port, 
                           A_ns(60) => SHIFT_n_14_59_port, A_ns(59) => 
                           SHIFT_n_14_59_port, A_ns(58) => SHIFT_n_14_58_port, 
                           A_ns(57) => SHIFT_n_14_57_port, A_ns(56) => 
                           SHIFT_n_14_56_port, A_ns(55) => SHIFT_n_14_55_port, 
                           A_ns(54) => SHIFT_n_14_54_port, A_ns(53) => 
                           SHIFT_n_14_53_port, A_ns(52) => SHIFT_n_14_52_port, 
                           A_ns(51) => SHIFT_n_14_51_port, A_ns(50) => 
                           SHIFT_n_14_50_port, A_ns(49) => SHIFT_n_14_49_port, 
                           A_ns(48) => SHIFT_n_14_48_port, A_ns(47) => 
                           SHIFT_n_14_47_port, A_ns(46) => SHIFT_n_14_46_port, 
                           A_ns(45) => SHIFT_n_14_45_port, A_ns(44) => 
                           SHIFT_n_14_44_port, A_ns(43) => SHIFT_n_14_43_port, 
                           A_ns(42) => SHIFT_n_14_42_port, A_ns(41) => 
                           SHIFT_n_14_41_port, A_ns(40) => SHIFT_n_14_40_port, 
                           A_ns(39) => SHIFT_n_14_39_port, A_ns(38) => 
                           SHIFT_n_14_38_port, A_ns(37) => SHIFT_n_14_37_port, 
                           A_ns(36) => SHIFT_n_14_36_port, A_ns(35) => 
                           SHIFT_n_14_35_port, A_ns(34) => SHIFT_n_14_34_port, 
                           A_ns(33) => SHIFT_n_14_33_port, A_ns(32) => 
                           SHIFT_n_14_32_port, A_ns(31) => SHIFT_n_14_31_port, 
                           A_ns(30) => SHIFT_n_14_30_port, A_ns(29) => 
                           SHIFT_n_14_29_port, A_ns(28) => SHIFT_n_14_28_port, 
                           A_ns(27) => SHIFT_n_14_27_port, A_ns(26) => 
                           SHIFT_n_14_26_port, A_ns(25) => SHIFT_n_14_25_port, 
                           A_ns(24) => SHIFT_n_14_24_port, A_ns(23) => 
                           SHIFT_n_14_23_port, A_ns(22) => SHIFT_n_14_22_port, 
                           A_ns(21) => SHIFT_n_14_21_port, A_ns(20) => 
                           SHIFT_n_14_20_port, A_ns(19) => SHIFT_n_14_19_port, 
                           A_ns(18) => SHIFT_n_14_18_port, A_ns(17) => 
                           SHIFT_n_14_17_port, A_ns(16) => SHIFT_n_14_16_port, 
                           A_ns(15) => SHIFT_n_14_15_port, A_ns(14) => 
                           SHIFT_n_14_14_port, A_ns(13) => SHIFT_n_14_13_port, 
                           A_ns(12) => SHIFT_n_14_12_port, A_ns(11) => 
                           SHIFT_n_14_11_port, A_ns(10) => SHIFT_n_14_10_port, 
                           A_ns(9) => SHIFT_n_14_9_port, A_ns(8) => 
                           SHIFT_n_14_8_port, A_ns(7) => SHIFT_n_14_7_port, 
                           A_ns(6) => SHIFT_n_14_6_port, A_ns(5) => 
                           SHIFT_n_14_5_port, A_ns(4) => SHIFT_n_14_4_port, 
                           A_ns(3) => SHIFT_n_14_3_port, A_ns(2) => 
                           SHIFT_n_14_2_port, A_ns(1) => SHIFT_n_14_1_port, 
                           A_ns(0) => SHIFT_n_14_0_port, B(61) => B(31), B(60) 
                           => B(31), B(59) => B(31), B(58) => B(31), B(57) => 
                           B(31), B(56) => B(31), B(55) => B(31), B(54) => 
                           B(31), B(53) => B(31), B(52) => B(31), B(51) => 
                           B(31), B(50) => B(31), B(49) => B(31), B(48) => 
                           B(31), B(47) => B(31), B(46) => B(31), B(45) => 
                           B(31), B(44) => B(31), B(43) => B(31), B(42) => 
                           B(31), B(41) => B(31), B(40) => B(31), B(39) => 
                           B(31), B(38) => B(31), B(37) => B(31), B(36) => 
                           B(31), B(35) => B(31), B(34) => B(31), B(33) => 
                           B(31), B(32) => B(31), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), O(61) => OTMP_14_61_port, 
                           O(60) => OTMP_14_60_port, O(59) => OTMP_14_59_port, 
                           O(58) => OTMP_14_58_port, O(57) => OTMP_14_57_port, 
                           O(56) => OTMP_14_56_port, O(55) => OTMP_14_55_port, 
                           O(54) => OTMP_14_54_port, O(53) => OTMP_14_53_port, 
                           O(52) => OTMP_14_52_port, O(51) => OTMP_14_51_port, 
                           O(50) => OTMP_14_50_port, O(49) => OTMP_14_49_port, 
                           O(48) => OTMP_14_48_port, O(47) => OTMP_14_47_port, 
                           O(46) => OTMP_14_46_port, O(45) => OTMP_14_45_port, 
                           O(44) => OTMP_14_44_port, O(43) => OTMP_14_43_port, 
                           O(42) => OTMP_14_42_port, O(41) => OTMP_14_41_port, 
                           O(40) => OTMP_14_40_port, O(39) => OTMP_14_39_port, 
                           O(38) => OTMP_14_38_port, O(37) => OTMP_14_37_port, 
                           O(36) => OTMP_14_36_port, O(35) => OTMP_14_35_port, 
                           O(34) => OTMP_14_34_port, O(33) => OTMP_14_33_port, 
                           O(32) => OTMP_14_32_port, O(31) => OTMP_14_31_port, 
                           O(30) => OTMP_14_30_port, O(29) => OTMP_14_29_port, 
                           O(28) => OTMP_14_28_port, O(27) => OTMP_14_27_port, 
                           O(26) => OTMP_14_26_port, O(25) => OTMP_14_25_port, 
                           O(24) => OTMP_14_24_port, O(23) => OTMP_14_23_port, 
                           O(22) => OTMP_14_22_port, O(21) => OTMP_14_21_port, 
                           O(20) => OTMP_14_20_port, O(19) => OTMP_14_19_port, 
                           O(18) => OTMP_14_18_port, O(17) => OTMP_14_17_port, 
                           O(16) => OTMP_14_16_port, O(15) => OTMP_14_15_port, 
                           O(14) => OTMP_14_14_port, O(13) => OTMP_14_13_port, 
                           O(12) => OTMP_14_12_port, O(11) => OTMP_14_11_port, 
                           O(10) => OTMP_14_10_port, O(9) => OTMP_14_9_port, 
                           O(8) => OTMP_14_8_port, O(7) => OTMP_14_7_port, O(6)
                           => OTMP_14_6_port, O(5) => OTMP_14_5_port, O(4) => 
                           OTMP_14_4_port, O(3) => OTMP_14_3_port, O(2) => 
                           OTMP_14_2_port, O(1) => OTMP_14_1_port, O(0) => 
                           n_1147, A_so(61) => SHIFT_15_61_port, A_so(60) => 
                           SHIFT_15_60_port, A_so(59) => SHIFT_15_59_port, 
                           A_so(58) => SHIFT_15_58_port, A_so(57) => 
                           SHIFT_15_57_port, A_so(56) => SHIFT_15_56_port, 
                           A_so(55) => SHIFT_15_55_port, A_so(54) => 
                           SHIFT_15_54_port, A_so(53) => SHIFT_15_53_port, 
                           A_so(52) => SHIFT_15_52_port, A_so(51) => 
                           SHIFT_15_51_port, A_so(50) => SHIFT_15_50_port, 
                           A_so(49) => SHIFT_15_49_port, A_so(48) => 
                           SHIFT_15_48_port, A_so(47) => SHIFT_15_47_port, 
                           A_so(46) => SHIFT_15_46_port, A_so(45) => 
                           SHIFT_15_45_port, A_so(44) => SHIFT_15_44_port, 
                           A_so(43) => SHIFT_15_43_port, A_so(42) => 
                           SHIFT_15_42_port, A_so(41) => SHIFT_15_41_port, 
                           A_so(40) => SHIFT_15_40_port, A_so(39) => 
                           SHIFT_15_39_port, A_so(38) => SHIFT_15_38_port, 
                           A_so(37) => SHIFT_15_37_port, A_so(36) => 
                           SHIFT_15_36_port, A_so(35) => SHIFT_15_35_port, 
                           A_so(34) => SHIFT_15_34_port, A_so(33) => 
                           SHIFT_15_33_port, A_so(32) => SHIFT_15_32_port, 
                           A_so(31) => SHIFT_15_31_port, A_so(30) => 
                           SHIFT_15_30_port, A_so(29) => SHIFT_15_29_port, 
                           A_so(28) => SHIFT_15_28_port, A_so(27) => 
                           SHIFT_15_27_port, A_so(26) => SHIFT_15_26_port, 
                           A_so(25) => SHIFT_15_25_port, A_so(24) => 
                           SHIFT_15_24_port, A_so(23) => SHIFT_15_23_port, 
                           A_so(22) => SHIFT_15_22_port, A_so(21) => 
                           SHIFT_15_21_port, A_so(20) => SHIFT_15_20_port, 
                           A_so(19) => SHIFT_15_19_port, A_so(18) => 
                           SHIFT_15_18_port, A_so(17) => SHIFT_15_17_port, 
                           A_so(16) => SHIFT_15_16_port, A_so(15) => 
                           SHIFT_15_15_port, A_so(14) => SHIFT_15_14_port, 
                           A_so(13) => SHIFT_15_13_port, A_so(12) => 
                           SHIFT_15_12_port, A_so(11) => SHIFT_15_11_port, 
                           A_so(10) => SHIFT_15_10_port, A_so(9) => 
                           SHIFT_15_9_port, A_so(8) => SHIFT_15_8_port, A_so(7)
                           => SHIFT_15_7_port, A_so(6) => SHIFT_15_6_port, 
                           A_so(5) => SHIFT_15_5_port, A_so(4) => 
                           SHIFT_15_4_port, A_so(3) => SHIFT_15_3_port, A_so(2)
                           => SHIFT_15_2_port, A_so(1) => n_1148, A_so(0) => 
                           n_1149, A_nso(61) => SHIFT_n_15_61_port, A_nso(60) 
                           => SHIFT_n_15_60_port, A_nso(59) => 
                           SHIFT_n_15_59_port, A_nso(58) => SHIFT_n_15_58_port,
                           A_nso(57) => SHIFT_n_15_57_port, A_nso(56) => 
                           SHIFT_n_15_56_port, A_nso(55) => SHIFT_n_15_55_port,
                           A_nso(54) => SHIFT_n_15_54_port, A_nso(53) => 
                           SHIFT_n_15_53_port, A_nso(52) => SHIFT_n_15_52_port,
                           A_nso(51) => SHIFT_n_15_51_port, A_nso(50) => 
                           SHIFT_n_15_50_port, A_nso(49) => SHIFT_n_15_49_port,
                           A_nso(48) => SHIFT_n_15_48_port, A_nso(47) => 
                           SHIFT_n_15_47_port, A_nso(46) => SHIFT_n_15_46_port,
                           A_nso(45) => SHIFT_n_15_45_port, A_nso(44) => 
                           SHIFT_n_15_44_port, A_nso(43) => SHIFT_n_15_43_port,
                           A_nso(42) => SHIFT_n_15_42_port, A_nso(41) => 
                           SHIFT_n_15_41_port, A_nso(40) => SHIFT_n_15_40_port,
                           A_nso(39) => SHIFT_n_15_39_port, A_nso(38) => 
                           SHIFT_n_15_38_port, A_nso(37) => SHIFT_n_15_37_port,
                           A_nso(36) => SHIFT_n_15_36_port, A_nso(35) => 
                           SHIFT_n_15_35_port, A_nso(34) => SHIFT_n_15_34_port,
                           A_nso(33) => SHIFT_n_15_33_port, A_nso(32) => 
                           SHIFT_n_15_32_port, A_nso(31) => SHIFT_n_15_31_port,
                           A_nso(30) => SHIFT_n_15_30_port, A_nso(29) => 
                           SHIFT_n_15_29_port, A_nso(28) => SHIFT_n_15_28_port,
                           A_nso(27) => SHIFT_n_15_27_port, A_nso(26) => 
                           SHIFT_n_15_26_port, A_nso(25) => SHIFT_n_15_25_port,
                           A_nso(24) => SHIFT_n_15_24_port, A_nso(23) => 
                           SHIFT_n_15_23_port, A_nso(22) => SHIFT_n_15_22_port,
                           A_nso(21) => SHIFT_n_15_21_port, A_nso(20) => 
                           SHIFT_n_15_20_port, A_nso(19) => SHIFT_n_15_19_port,
                           A_nso(18) => SHIFT_n_15_18_port, A_nso(17) => 
                           SHIFT_n_15_17_port, A_nso(16) => SHIFT_n_15_16_port,
                           A_nso(15) => SHIFT_n_15_15_port, A_nso(14) => 
                           SHIFT_n_15_14_port, A_nso(13) => SHIFT_n_15_13_port,
                           A_nso(12) => SHIFT_n_15_12_port, A_nso(11) => 
                           SHIFT_n_15_11_port, A_nso(10) => SHIFT_n_15_10_port,
                           A_nso(9) => SHIFT_n_15_9_port, A_nso(8) => 
                           SHIFT_n_15_8_port, A_nso(7) => SHIFT_n_15_7_port, 
                           A_nso(6) => SHIFT_n_15_6_port, A_nso(5) => 
                           SHIFT_n_15_5_port, A_nso(4) => SHIFT_n_15_4_port, 
                           A_nso(3) => SHIFT_n_15_3_port, A_nso(2) => 
                           SHIFT_n_15_2_port, A_nso(1) => n_1150, A_nso(0) => 
                           n_1151);
   ENC_15 : BOOTHENC_NBIT64_i30 port map( A_s(63) => SHIFT_15_61_port, A_s(62) 
                           => SHIFT_15_61_port, A_s(61) => SHIFT_15_61_port, 
                           A_s(60) => SHIFT_15_60_port, A_s(59) => 
                           SHIFT_15_59_port, A_s(58) => SHIFT_15_58_port, 
                           A_s(57) => SHIFT_15_57_port, A_s(56) => 
                           SHIFT_15_56_port, A_s(55) => SHIFT_15_55_port, 
                           A_s(54) => SHIFT_15_54_port, A_s(53) => 
                           SHIFT_15_53_port, A_s(52) => SHIFT_15_52_port, 
                           A_s(51) => SHIFT_15_51_port, A_s(50) => 
                           SHIFT_15_50_port, A_s(49) => SHIFT_15_49_port, 
                           A_s(48) => SHIFT_15_48_port, A_s(47) => 
                           SHIFT_15_47_port, A_s(46) => SHIFT_15_46_port, 
                           A_s(45) => SHIFT_15_45_port, A_s(44) => 
                           SHIFT_15_44_port, A_s(43) => SHIFT_15_43_port, 
                           A_s(42) => SHIFT_15_42_port, A_s(41) => 
                           SHIFT_15_41_port, A_s(40) => SHIFT_15_40_port, 
                           A_s(39) => SHIFT_15_39_port, A_s(38) => 
                           SHIFT_15_38_port, A_s(37) => SHIFT_15_37_port, 
                           A_s(36) => SHIFT_15_36_port, A_s(35) => 
                           SHIFT_15_35_port, A_s(34) => SHIFT_15_34_port, 
                           A_s(33) => SHIFT_15_33_port, A_s(32) => 
                           SHIFT_15_32_port, A_s(31) => SHIFT_15_31_port, 
                           A_s(30) => SHIFT_15_30_port, A_s(29) => 
                           SHIFT_15_29_port, A_s(28) => SHIFT_15_28_port, 
                           A_s(27) => SHIFT_15_27_port, A_s(26) => 
                           SHIFT_15_26_port, A_s(25) => SHIFT_15_25_port, 
                           A_s(24) => SHIFT_15_24_port, A_s(23) => 
                           SHIFT_15_23_port, A_s(22) => SHIFT_15_22_port, 
                           A_s(21) => SHIFT_15_21_port, A_s(20) => 
                           SHIFT_15_20_port, A_s(19) => SHIFT_15_19_port, 
                           A_s(18) => SHIFT_15_18_port, A_s(17) => 
                           SHIFT_15_17_port, A_s(16) => SHIFT_15_16_port, 
                           A_s(15) => SHIFT_15_15_port, A_s(14) => 
                           SHIFT_15_14_port, A_s(13) => SHIFT_15_13_port, 
                           A_s(12) => SHIFT_15_12_port, A_s(11) => 
                           SHIFT_15_11_port, A_s(10) => SHIFT_15_10_port, 
                           A_s(9) => SHIFT_15_9_port, A_s(8) => SHIFT_15_8_port
                           , A_s(7) => SHIFT_15_7_port, A_s(6) => 
                           SHIFT_15_6_port, A_s(5) => SHIFT_15_5_port, A_s(4) 
                           => SHIFT_15_4_port, A_s(3) => SHIFT_15_3_port, 
                           A_s(2) => SHIFT_15_2_port, A_s(1) => SHIFT_15_1_port
                           , A_s(0) => SHIFT_15_0_port, A_ns(63) => 
                           SHIFT_n_15_61_port, A_ns(62) => SHIFT_n_15_61_port, 
                           A_ns(61) => SHIFT_n_15_61_port, A_ns(60) => 
                           SHIFT_n_15_60_port, A_ns(59) => SHIFT_n_15_59_port, 
                           A_ns(58) => SHIFT_n_15_58_port, A_ns(57) => 
                           SHIFT_n_15_57_port, A_ns(56) => SHIFT_n_15_56_port, 
                           A_ns(55) => SHIFT_n_15_55_port, A_ns(54) => 
                           SHIFT_n_15_54_port, A_ns(53) => SHIFT_n_15_53_port, 
                           A_ns(52) => SHIFT_n_15_52_port, A_ns(51) => 
                           SHIFT_n_15_51_port, A_ns(50) => SHIFT_n_15_50_port, 
                           A_ns(49) => SHIFT_n_15_49_port, A_ns(48) => 
                           SHIFT_n_15_48_port, A_ns(47) => SHIFT_n_15_47_port, 
                           A_ns(46) => SHIFT_n_15_46_port, A_ns(45) => 
                           SHIFT_n_15_45_port, A_ns(44) => SHIFT_n_15_44_port, 
                           A_ns(43) => SHIFT_n_15_43_port, A_ns(42) => 
                           SHIFT_n_15_42_port, A_ns(41) => SHIFT_n_15_41_port, 
                           A_ns(40) => SHIFT_n_15_40_port, A_ns(39) => 
                           SHIFT_n_15_39_port, A_ns(38) => SHIFT_n_15_38_port, 
                           A_ns(37) => SHIFT_n_15_37_port, A_ns(36) => 
                           SHIFT_n_15_36_port, A_ns(35) => SHIFT_n_15_35_port, 
                           A_ns(34) => SHIFT_n_15_34_port, A_ns(33) => 
                           SHIFT_n_15_33_port, A_ns(32) => SHIFT_n_15_32_port, 
                           A_ns(31) => SHIFT_n_15_31_port, A_ns(30) => 
                           SHIFT_n_15_30_port, A_ns(29) => SHIFT_n_15_29_port, 
                           A_ns(28) => SHIFT_n_15_28_port, A_ns(27) => 
                           SHIFT_n_15_27_port, A_ns(26) => SHIFT_n_15_26_port, 
                           A_ns(25) => SHIFT_n_15_25_port, A_ns(24) => 
                           SHIFT_n_15_24_port, A_ns(23) => SHIFT_n_15_23_port, 
                           A_ns(22) => SHIFT_n_15_22_port, A_ns(21) => 
                           SHIFT_n_15_21_port, A_ns(20) => SHIFT_n_15_20_port, 
                           A_ns(19) => SHIFT_n_15_19_port, A_ns(18) => 
                           SHIFT_n_15_18_port, A_ns(17) => SHIFT_n_15_17_port, 
                           A_ns(16) => SHIFT_n_15_16_port, A_ns(15) => 
                           SHIFT_n_15_15_port, A_ns(14) => SHIFT_n_15_14_port, 
                           A_ns(13) => SHIFT_n_15_13_port, A_ns(12) => 
                           SHIFT_n_15_12_port, A_ns(11) => SHIFT_n_15_11_port, 
                           A_ns(10) => SHIFT_n_15_10_port, A_ns(9) => 
                           SHIFT_n_15_9_port, A_ns(8) => SHIFT_n_15_8_port, 
                           A_ns(7) => SHIFT_n_15_7_port, A_ns(6) => 
                           SHIFT_n_15_6_port, A_ns(5) => SHIFT_n_15_5_port, 
                           A_ns(4) => SHIFT_n_15_4_port, A_ns(3) => 
                           SHIFT_n_15_3_port, A_ns(2) => SHIFT_n_15_2_port, 
                           A_ns(1) => SHIFT_n_15_1_port, A_ns(0) => 
                           SHIFT_n_15_0_port, B(63) => B(31), B(62) => B(31), 
                           B(61) => B(31), B(60) => B(31), B(59) => B(31), 
                           B(58) => B(31), B(57) => B(31), B(56) => B(31), 
                           B(55) => B(31), B(54) => B(31), B(53) => B(31), 
                           B(52) => B(31), B(51) => B(31), B(50) => B(31), 
                           B(49) => B(31), B(48) => B(31), B(47) => B(31), 
                           B(46) => B(31), B(45) => B(31), B(44) => B(31), 
                           B(43) => B(31), B(42) => B(31), B(41) => B(31), 
                           B(40) => B(31), B(39) => B(31), B(38) => B(31), 
                           B(37) => B(31), B(36) => B(31), B(35) => B(31), 
                           B(34) => B(31), B(33) => B(31), B(32) => B(31), 
                           B(31) => B(31), B(30) => B(30), B(29) => B(29), 
                           B(28) => B(28), B(27) => B(27), B(26) => B(26), 
                           B(25) => B(25), B(24) => B(24), B(23) => B(23), 
                           B(22) => B(22), B(21) => B(21), B(20) => B(20), 
                           B(19) => B(19), B(18) => B(18), B(17) => B(17), 
                           B(16) => B(16), B(15) => B(15), B(14) => B(14), 
                           B(13) => B(13), B(12) => B(12), B(11) => B(11), 
                           B(10) => B(10), B(9) => B(9), B(8) => B(8), B(7) => 
                           B(7), B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3)
                           => B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), 
                           O(63) => OTMP_15_63_port, O(62) => OTMP_15_62_port, 
                           O(61) => OTMP_15_61_port, O(60) => OTMP_15_60_port, 
                           O(59) => OTMP_15_59_port, O(58) => OTMP_15_58_port, 
                           O(57) => OTMP_15_57_port, O(56) => OTMP_15_56_port, 
                           O(55) => OTMP_15_55_port, O(54) => OTMP_15_54_port, 
                           O(53) => OTMP_15_53_port, O(52) => OTMP_15_52_port, 
                           O(51) => OTMP_15_51_port, O(50) => OTMP_15_50_port, 
                           O(49) => OTMP_15_49_port, O(48) => OTMP_15_48_port, 
                           O(47) => OTMP_15_47_port, O(46) => OTMP_15_46_port, 
                           O(45) => OTMP_15_45_port, O(44) => OTMP_15_44_port, 
                           O(43) => OTMP_15_43_port, O(42) => OTMP_15_42_port, 
                           O(41) => OTMP_15_41_port, O(40) => OTMP_15_40_port, 
                           O(39) => OTMP_15_39_port, O(38) => OTMP_15_38_port, 
                           O(37) => OTMP_15_37_port, O(36) => OTMP_15_36_port, 
                           O(35) => OTMP_15_35_port, O(34) => OTMP_15_34_port, 
                           O(33) => OTMP_15_33_port, O(32) => OTMP_15_32_port, 
                           O(31) => OTMP_15_31_port, O(30) => OTMP_15_30_port, 
                           O(29) => OTMP_15_29_port, O(28) => OTMP_15_28_port, 
                           O(27) => OTMP_15_27_port, O(26) => OTMP_15_26_port, 
                           O(25) => OTMP_15_25_port, O(24) => OTMP_15_24_port, 
                           O(23) => OTMP_15_23_port, O(22) => OTMP_15_22_port, 
                           O(21) => OTMP_15_21_port, O(20) => OTMP_15_20_port, 
                           O(19) => OTMP_15_19_port, O(18) => OTMP_15_18_port, 
                           O(17) => OTMP_15_17_port, O(16) => OTMP_15_16_port, 
                           O(15) => OTMP_15_15_port, O(14) => OTMP_15_14_port, 
                           O(13) => OTMP_15_13_port, O(12) => OTMP_15_12_port, 
                           O(11) => OTMP_15_11_port, O(10) => OTMP_15_10_port, 
                           O(9) => OTMP_15_9_port, O(8) => OTMP_15_8_port, O(7)
                           => OTMP_15_7_port, O(6) => OTMP_15_6_port, O(5) => 
                           OTMP_15_5_port, O(4) => OTMP_15_4_port, O(3) => 
                           OTMP_15_3_port, O(2) => OTMP_15_2_port, O(1) => 
                           OTMP_15_1_port, O(0) => n_1152, A_so(63) => n_1153, 
                           A_so(62) => n_1154, A_so(61) => n_1155, A_so(60) => 
                           n_1156, A_so(59) => n_1157, A_so(58) => n_1158, 
                           A_so(57) => n_1159, A_so(56) => n_1160, A_so(55) => 
                           n_1161, A_so(54) => n_1162, A_so(53) => n_1163, 
                           A_so(52) => n_1164, A_so(51) => n_1165, A_so(50) => 
                           n_1166, A_so(49) => n_1167, A_so(48) => n_1168, 
                           A_so(47) => n_1169, A_so(46) => n_1170, A_so(45) => 
                           n_1171, A_so(44) => n_1172, A_so(43) => n_1173, 
                           A_so(42) => n_1174, A_so(41) => n_1175, A_so(40) => 
                           n_1176, A_so(39) => n_1177, A_so(38) => n_1178, 
                           A_so(37) => n_1179, A_so(36) => n_1180, A_so(35) => 
                           n_1181, A_so(34) => n_1182, A_so(33) => n_1183, 
                           A_so(32) => n_1184, A_so(31) => n_1185, A_so(30) => 
                           n_1186, A_so(29) => n_1187, A_so(28) => n_1188, 
                           A_so(27) => n_1189, A_so(26) => n_1190, A_so(25) => 
                           n_1191, A_so(24) => n_1192, A_so(23) => n_1193, 
                           A_so(22) => n_1194, A_so(21) => n_1195, A_so(20) => 
                           n_1196, A_so(19) => n_1197, A_so(18) => n_1198, 
                           A_so(17) => n_1199, A_so(16) => n_1200, A_so(15) => 
                           n_1201, A_so(14) => n_1202, A_so(13) => n_1203, 
                           A_so(12) => n_1204, A_so(11) => n_1205, A_so(10) => 
                           n_1206, A_so(9) => n_1207, A_so(8) => n_1208, 
                           A_so(7) => n_1209, A_so(6) => n_1210, A_so(5) => 
                           n_1211, A_so(4) => n_1212, A_so(3) => n_1213, 
                           A_so(2) => n_1214, A_so(1) => n_1215, A_so(0) => 
                           n_1216, A_nso(63) => n_1217, A_nso(62) => n_1218, 
                           A_nso(61) => n_1219, A_nso(60) => n_1220, A_nso(59) 
                           => n_1221, A_nso(58) => n_1222, A_nso(57) => n_1223,
                           A_nso(56) => n_1224, A_nso(55) => n_1225, A_nso(54) 
                           => n_1226, A_nso(53) => n_1227, A_nso(52) => n_1228,
                           A_nso(51) => n_1229, A_nso(50) => n_1230, A_nso(49) 
                           => n_1231, A_nso(48) => n_1232, A_nso(47) => n_1233,
                           A_nso(46) => n_1234, A_nso(45) => n_1235, A_nso(44) 
                           => n_1236, A_nso(43) => n_1237, A_nso(42) => n_1238,
                           A_nso(41) => n_1239, A_nso(40) => n_1240, A_nso(39) 
                           => n_1241, A_nso(38) => n_1242, A_nso(37) => n_1243,
                           A_nso(36) => n_1244, A_nso(35) => n_1245, A_nso(34) 
                           => n_1246, A_nso(33) => n_1247, A_nso(32) => n_1248,
                           A_nso(31) => n_1249, A_nso(30) => n_1250, A_nso(29) 
                           => n_1251, A_nso(28) => n_1252, A_nso(27) => n_1253,
                           A_nso(26) => n_1254, A_nso(25) => n_1255, A_nso(24) 
                           => n_1256, A_nso(23) => n_1257, A_nso(22) => n_1258,
                           A_nso(21) => n_1259, A_nso(20) => n_1260, A_nso(19) 
                           => n_1261, A_nso(18) => n_1262, A_nso(17) => n_1263,
                           A_nso(16) => n_1264, A_nso(15) => n_1265, A_nso(14) 
                           => n_1266, A_nso(13) => n_1267, A_nso(12) => n_1268,
                           A_nso(11) => n_1269, A_nso(10) => n_1270, A_nso(9) 
                           => n_1271, A_nso(8) => n_1272, A_nso(7) => n_1273, 
                           A_nso(6) => n_1274, A_nso(5) => n_1275, A_nso(4) => 
                           n_1276, A_nso(3) => n_1277, A_nso(2) => n_1278, 
                           A_nso(1) => n_1279, A_nso(0) => n_1280);
   ADDER1 : RCA_NBIT36 port map( A(35) => OTMP_0_34_port, A(34) => 
                           OTMP_0_34_port, A(33) => OTMP_0_34_port, A(32) => 
                           OTMP_0_32_port, A(31) => OTMP_0_31_port, A(30) => 
                           OTMP_0_30_port, A(29) => OTMP_0_29_port, A(28) => 
                           OTMP_0_28_port, A(27) => OTMP_0_27_port, A(26) => 
                           OTMP_0_26_port, A(25) => OTMP_0_25_port, A(24) => 
                           OTMP_0_24_port, A(23) => OTMP_0_23_port, A(22) => 
                           OTMP_0_22_port, A(21) => OTMP_0_21_port, A(20) => 
                           OTMP_0_20_port, A(19) => OTMP_0_19_port, A(18) => 
                           OTMP_0_18_port, A(17) => OTMP_0_17_port, A(16) => 
                           OTMP_0_16_port, A(15) => OTMP_0_15_port, A(14) => 
                           OTMP_0_14_port, A(13) => OTMP_0_13_port, A(12) => 
                           OTMP_0_12_port, A(11) => OTMP_0_11_port, A(10) => 
                           OTMP_0_10_port, A(9) => OTMP_0_9_port, A(8) => 
                           OTMP_0_8_port, A(7) => OTMP_0_7_port, A(6) => 
                           OTMP_0_6_port, A(5) => OTMP_0_5_port, A(4) => 
                           OTMP_0_4_port, A(3) => OTMP_0_3_port, A(2) => 
                           OTMP_0_2_port, A(1) => OTMP_0_1_port, A(0) => 
                           OTMP_0_0_port, B(35) => OTMP_1_35_port, B(34) => 
                           OTMP_1_34_port, B(33) => OTMP_1_33_port, B(32) => 
                           OTMP_1_32_port, B(31) => OTMP_1_31_port, B(30) => 
                           OTMP_1_30_port, B(29) => OTMP_1_29_port, B(28) => 
                           OTMP_1_28_port, B(27) => OTMP_1_27_port, B(26) => 
                           OTMP_1_26_port, B(25) => OTMP_1_25_port, B(24) => 
                           OTMP_1_24_port, B(23) => OTMP_1_23_port, B(22) => 
                           OTMP_1_22_port, B(21) => OTMP_1_21_port, B(20) => 
                           OTMP_1_20_port, B(19) => OTMP_1_19_port, B(18) => 
                           OTMP_1_18_port, B(17) => OTMP_1_17_port, B(16) => 
                           OTMP_1_16_port, B(15) => OTMP_1_15_port, B(14) => 
                           OTMP_1_14_port, B(13) => OTMP_1_13_port, B(12) => 
                           OTMP_1_12_port, B(11) => OTMP_1_11_port, B(10) => 
                           OTMP_1_10_port, B(9) => OTMP_1_9_port, B(8) => 
                           OTMP_1_8_port, B(7) => OTMP_1_7_port, B(6) => 
                           OTMP_1_6_port, B(5) => OTMP_1_5_port, B(4) => 
                           OTMP_1_4_port, B(3) => OTMP_1_3_port, B(2) => 
                           OTMP_1_2_port, B(1) => OTMP_1_1_port, B(0) => 
                           OTMP_1_0_port, Ci => X_Logic0_port, S(35) => 
                           PTMP_0_36_port, S(34) => PTMP_0_34_port, S(33) => 
                           PTMP_0_33_port, S(32) => PTMP_0_32_port, S(31) => 
                           PTMP_0_31_port, S(30) => PTMP_0_30_port, S(29) => 
                           PTMP_0_29_port, S(28) => PTMP_0_28_port, S(27) => 
                           PTMP_0_27_port, S(26) => PTMP_0_26_port, S(25) => 
                           PTMP_0_25_port, S(24) => PTMP_0_24_port, S(23) => 
                           PTMP_0_23_port, S(22) => PTMP_0_22_port, S(21) => 
                           PTMP_0_21_port, S(20) => PTMP_0_20_port, S(19) => 
                           PTMP_0_19_port, S(18) => PTMP_0_18_port, S(17) => 
                           PTMP_0_17_port, S(16) => PTMP_0_16_port, S(15) => 
                           PTMP_0_15_port, S(14) => PTMP_0_14_port, S(13) => 
                           PTMP_0_13_port, S(12) => PTMP_0_12_port, S(11) => 
                           PTMP_0_11_port, S(10) => PTMP_0_10_port, S(9) => 
                           PTMP_0_9_port, S(8) => PTMP_0_8_port, S(7) => 
                           PTMP_0_7_port, S(6) => PTMP_0_6_port, S(5) => 
                           PTMP_0_5_port, S(4) => PTMP_0_4_port, S(3) => 
                           PTMP_0_3_port, S(2) => PTMP_0_2_port, S(1) => 
                           PTMP_0_1_port, S(0) => PTMP_0_0_port, Co => n_1281);
   ADDER_2 : RCA_NBIT38 port map( A(37) => n20, A(36) => n20, A(35) => 
                           PTMP_0_36_port, A(34) => PTMP_0_34_port, A(33) => 
                           PTMP_0_33_port, A(32) => PTMP_0_32_port, A(31) => 
                           PTMP_0_31_port, A(30) => PTMP_0_30_port, A(29) => 
                           PTMP_0_29_port, A(28) => PTMP_0_28_port, A(27) => 
                           PTMP_0_27_port, A(26) => PTMP_0_26_port, A(25) => 
                           PTMP_0_25_port, A(24) => PTMP_0_24_port, A(23) => 
                           PTMP_0_23_port, A(22) => PTMP_0_22_port, A(21) => 
                           PTMP_0_21_port, A(20) => PTMP_0_20_port, A(19) => 
                           PTMP_0_19_port, A(18) => PTMP_0_18_port, A(17) => 
                           PTMP_0_17_port, A(16) => PTMP_0_16_port, A(15) => 
                           PTMP_0_15_port, A(14) => PTMP_0_14_port, A(13) => 
                           PTMP_0_13_port, A(12) => PTMP_0_12_port, A(11) => 
                           PTMP_0_11_port, A(10) => PTMP_0_10_port, A(9) => 
                           PTMP_0_9_port, A(8) => PTMP_0_8_port, A(7) => 
                           PTMP_0_7_port, A(6) => PTMP_0_6_port, A(5) => 
                           PTMP_0_5_port, A(4) => PTMP_0_4_port, A(3) => 
                           PTMP_0_3_port, A(2) => PTMP_0_2_port, A(1) => 
                           PTMP_0_1_port, A(0) => PTMP_0_0_port, B(37) => 
                           OTMP_2_37_port, B(36) => OTMP_2_36_port, B(35) => 
                           OTMP_2_35_port, B(34) => OTMP_2_34_port, B(33) => 
                           OTMP_2_33_port, B(32) => OTMP_2_32_port, B(31) => 
                           OTMP_2_31_port, B(30) => OTMP_2_30_port, B(29) => 
                           OTMP_2_29_port, B(28) => OTMP_2_28_port, B(27) => 
                           OTMP_2_27_port, B(26) => OTMP_2_26_port, B(25) => 
                           OTMP_2_25_port, B(24) => OTMP_2_24_port, B(23) => 
                           OTMP_2_23_port, B(22) => OTMP_2_22_port, B(21) => 
                           OTMP_2_21_port, B(20) => OTMP_2_20_port, B(19) => 
                           OTMP_2_19_port, B(18) => OTMP_2_18_port, B(17) => 
                           OTMP_2_17_port, B(16) => OTMP_2_16_port, B(15) => 
                           OTMP_2_15_port, B(14) => OTMP_2_14_port, B(13) => 
                           OTMP_2_13_port, B(12) => OTMP_2_12_port, B(11) => 
                           OTMP_2_11_port, B(10) => OTMP_2_10_port, B(9) => 
                           OTMP_2_9_port, B(8) => OTMP_2_8_port, B(7) => 
                           OTMP_2_7_port, B(6) => OTMP_2_6_port, B(5) => 
                           OTMP_2_5_port, B(4) => OTMP_2_4_port, B(3) => 
                           OTMP_2_3_port, B(2) => OTMP_2_2_port, B(1) => 
                           OTMP_2_1_port, B(0) => OTMP_2_0_port, Ci => 
                           X_Logic0_port, S(37) => PTMP_1_37_port, S(36) => 
                           PTMP_1_36_port, S(35) => PTMP_1_35_port, S(34) => 
                           PTMP_1_34_port, S(33) => PTMP_1_33_port, S(32) => 
                           PTMP_1_32_port, S(31) => PTMP_1_31_port, S(30) => 
                           PTMP_1_30_port, S(29) => PTMP_1_29_port, S(28) => 
                           PTMP_1_28_port, S(27) => PTMP_1_27_port, S(26) => 
                           PTMP_1_26_port, S(25) => PTMP_1_25_port, S(24) => 
                           PTMP_1_24_port, S(23) => PTMP_1_23_port, S(22) => 
                           PTMP_1_22_port, S(21) => PTMP_1_21_port, S(20) => 
                           PTMP_1_20_port, S(19) => PTMP_1_19_port, S(18) => 
                           PTMP_1_18_port, S(17) => PTMP_1_17_port, S(16) => 
                           PTMP_1_16_port, S(15) => PTMP_1_15_port, S(14) => 
                           PTMP_1_14_port, S(13) => PTMP_1_13_port, S(12) => 
                           PTMP_1_12_port, S(11) => PTMP_1_11_port, S(10) => 
                           PTMP_1_10_port, S(9) => PTMP_1_9_port, S(8) => 
                           PTMP_1_8_port, S(7) => PTMP_1_7_port, S(6) => 
                           PTMP_1_6_port, S(5) => PTMP_1_5_port, S(4) => 
                           PTMP_1_4_port, S(3) => PTMP_1_3_port, S(2) => 
                           PTMP_1_2_port, S(1) => PTMP_1_1_port, S(0) => 
                           PTMP_1_0_port, Co => n_1282);
   ADDER_3 : RCA_NBIT40 port map( A(39) => PTMP_1_37_port, A(38) => 
                           PTMP_1_37_port, A(37) => PTMP_1_37_port, A(36) => 
                           PTMP_1_36_port, A(35) => PTMP_1_35_port, A(34) => 
                           PTMP_1_34_port, A(33) => PTMP_1_33_port, A(32) => 
                           PTMP_1_32_port, A(31) => PTMP_1_31_port, A(30) => 
                           PTMP_1_30_port, A(29) => PTMP_1_29_port, A(28) => 
                           PTMP_1_28_port, A(27) => PTMP_1_27_port, A(26) => 
                           PTMP_1_26_port, A(25) => PTMP_1_25_port, A(24) => 
                           PTMP_1_24_port, A(23) => PTMP_1_23_port, A(22) => 
                           PTMP_1_22_port, A(21) => PTMP_1_21_port, A(20) => 
                           PTMP_1_20_port, A(19) => PTMP_1_19_port, A(18) => 
                           PTMP_1_18_port, A(17) => PTMP_1_17_port, A(16) => 
                           PTMP_1_16_port, A(15) => PTMP_1_15_port, A(14) => 
                           PTMP_1_14_port, A(13) => PTMP_1_13_port, A(12) => 
                           PTMP_1_12_port, A(11) => PTMP_1_11_port, A(10) => 
                           PTMP_1_10_port, A(9) => PTMP_1_9_port, A(8) => 
                           PTMP_1_8_port, A(7) => PTMP_1_7_port, A(6) => 
                           PTMP_1_6_port, A(5) => PTMP_1_5_port, A(4) => 
                           PTMP_1_4_port, A(3) => PTMP_1_3_port, A(2) => 
                           PTMP_1_2_port, A(1) => PTMP_1_1_port, A(0) => 
                           PTMP_1_0_port, B(39) => OTMP_3_39_port, B(38) => 
                           OTMP_3_38_port, B(37) => OTMP_3_37_port, B(36) => 
                           OTMP_3_36_port, B(35) => OTMP_3_35_port, B(34) => 
                           OTMP_3_34_port, B(33) => OTMP_3_33_port, B(32) => 
                           OTMP_3_32_port, B(31) => OTMP_3_31_port, B(30) => 
                           OTMP_3_30_port, B(29) => OTMP_3_29_port, B(28) => 
                           OTMP_3_28_port, B(27) => OTMP_3_27_port, B(26) => 
                           OTMP_3_26_port, B(25) => OTMP_3_25_port, B(24) => 
                           OTMP_3_24_port, B(23) => OTMP_3_23_port, B(22) => 
                           OTMP_3_22_port, B(21) => OTMP_3_21_port, B(20) => 
                           OTMP_3_20_port, B(19) => OTMP_3_19_port, B(18) => 
                           OTMP_3_18_port, B(17) => OTMP_3_17_port, B(16) => 
                           OTMP_3_16_port, B(15) => OTMP_3_15_port, B(14) => 
                           OTMP_3_14_port, B(13) => OTMP_3_13_port, B(12) => 
                           OTMP_3_12_port, B(11) => OTMP_3_11_port, B(10) => 
                           OTMP_3_10_port, B(9) => OTMP_3_9_port, B(8) => 
                           OTMP_3_8_port, B(7) => OTMP_3_7_port, B(6) => 
                           OTMP_3_6_port, B(5) => OTMP_3_5_port, B(4) => 
                           OTMP_3_4_port, B(3) => OTMP_3_3_port, B(2) => 
                           OTMP_3_2_port, B(1) => OTMP_3_1_port, B(0) => 
                           OTMP_3_0_port, Ci => X_Logic0_port, S(39) => 
                           PTMP_2_39_port, S(38) => PTMP_2_38_port, S(37) => 
                           PTMP_2_37_port, S(36) => PTMP_2_36_port, S(35) => 
                           PTMP_2_35_port, S(34) => PTMP_2_34_port, S(33) => 
                           PTMP_2_33_port, S(32) => PTMP_2_32_port, S(31) => 
                           PTMP_2_31_port, S(30) => PTMP_2_30_port, S(29) => 
                           PTMP_2_29_port, S(28) => PTMP_2_28_port, S(27) => 
                           PTMP_2_27_port, S(26) => PTMP_2_26_port, S(25) => 
                           PTMP_2_25_port, S(24) => PTMP_2_24_port, S(23) => 
                           PTMP_2_23_port, S(22) => PTMP_2_22_port, S(21) => 
                           PTMP_2_21_port, S(20) => PTMP_2_20_port, S(19) => 
                           PTMP_2_19_port, S(18) => PTMP_2_18_port, S(17) => 
                           PTMP_2_17_port, S(16) => PTMP_2_16_port, S(15) => 
                           PTMP_2_15_port, S(14) => PTMP_2_14_port, S(13) => 
                           PTMP_2_13_port, S(12) => PTMP_2_12_port, S(11) => 
                           PTMP_2_11_port, S(10) => PTMP_2_10_port, S(9) => 
                           PTMP_2_9_port, S(8) => PTMP_2_8_port, S(7) => 
                           PTMP_2_7_port, S(6) => PTMP_2_6_port, S(5) => 
                           PTMP_2_5_port, S(4) => PTMP_2_4_port, S(3) => 
                           PTMP_2_3_port, S(2) => PTMP_2_2_port, S(1) => 
                           PTMP_2_1_port, S(0) => PTMP_2_0_port, Co => n_1283);
   ADDER_4 : RCA_NBIT42 port map( A(41) => PTMP_2_39_port, A(40) => 
                           PTMP_2_39_port, A(39) => PTMP_2_39_port, A(38) => 
                           PTMP_2_38_port, A(37) => PTMP_2_37_port, A(36) => 
                           PTMP_2_36_port, A(35) => PTMP_2_35_port, A(34) => 
                           PTMP_2_34_port, A(33) => PTMP_2_33_port, A(32) => 
                           PTMP_2_32_port, A(31) => PTMP_2_31_port, A(30) => 
                           PTMP_2_30_port, A(29) => PTMP_2_29_port, A(28) => 
                           PTMP_2_28_port, A(27) => PTMP_2_27_port, A(26) => 
                           PTMP_2_26_port, A(25) => PTMP_2_25_port, A(24) => 
                           PTMP_2_24_port, A(23) => PTMP_2_23_port, A(22) => 
                           PTMP_2_22_port, A(21) => PTMP_2_21_port, A(20) => 
                           PTMP_2_20_port, A(19) => PTMP_2_19_port, A(18) => 
                           PTMP_2_18_port, A(17) => PTMP_2_17_port, A(16) => 
                           PTMP_2_16_port, A(15) => PTMP_2_15_port, A(14) => 
                           PTMP_2_14_port, A(13) => PTMP_2_13_port, A(12) => 
                           PTMP_2_12_port, A(11) => PTMP_2_11_port, A(10) => 
                           PTMP_2_10_port, A(9) => PTMP_2_9_port, A(8) => 
                           PTMP_2_8_port, A(7) => PTMP_2_7_port, A(6) => 
                           PTMP_2_6_port, A(5) => PTMP_2_5_port, A(4) => 
                           PTMP_2_4_port, A(3) => PTMP_2_3_port, A(2) => 
                           PTMP_2_2_port, A(1) => PTMP_2_1_port, A(0) => 
                           PTMP_2_0_port, B(41) => OTMP_4_41_port, B(40) => 
                           OTMP_4_40_port, B(39) => OTMP_4_39_port, B(38) => 
                           OTMP_4_38_port, B(37) => OTMP_4_37_port, B(36) => 
                           OTMP_4_36_port, B(35) => OTMP_4_35_port, B(34) => 
                           OTMP_4_34_port, B(33) => OTMP_4_33_port, B(32) => 
                           OTMP_4_32_port, B(31) => OTMP_4_31_port, B(30) => 
                           OTMP_4_30_port, B(29) => OTMP_4_29_port, B(28) => 
                           OTMP_4_28_port, B(27) => OTMP_4_27_port, B(26) => 
                           OTMP_4_26_port, B(25) => OTMP_4_25_port, B(24) => 
                           OTMP_4_24_port, B(23) => OTMP_4_23_port, B(22) => 
                           OTMP_4_22_port, B(21) => OTMP_4_21_port, B(20) => 
                           OTMP_4_20_port, B(19) => OTMP_4_19_port, B(18) => 
                           OTMP_4_18_port, B(17) => OTMP_4_17_port, B(16) => 
                           OTMP_4_16_port, B(15) => OTMP_4_15_port, B(14) => 
                           OTMP_4_14_port, B(13) => OTMP_4_13_port, B(12) => 
                           OTMP_4_12_port, B(11) => OTMP_4_11_port, B(10) => 
                           OTMP_4_10_port, B(9) => OTMP_4_9_port, B(8) => 
                           OTMP_4_8_port, B(7) => OTMP_4_7_port, B(6) => 
                           OTMP_4_6_port, B(5) => OTMP_4_5_port, B(4) => 
                           OTMP_4_4_port, B(3) => OTMP_4_3_port, B(2) => 
                           OTMP_4_2_port, B(1) => OTMP_4_1_port, B(0) => 
                           OTMP_4_0_port, Ci => X_Logic0_port, S(41) => 
                           PTMP_3_41_port, S(40) => PTMP_3_40_port, S(39) => 
                           PTMP_3_39_port, S(38) => PTMP_3_38_port, S(37) => 
                           PTMP_3_37_port, S(36) => PTMP_3_36_port, S(35) => 
                           PTMP_3_35_port, S(34) => PTMP_3_34_port, S(33) => 
                           PTMP_3_33_port, S(32) => PTMP_3_32_port, S(31) => 
                           PTMP_3_31_port, S(30) => PTMP_3_30_port, S(29) => 
                           PTMP_3_29_port, S(28) => PTMP_3_28_port, S(27) => 
                           PTMP_3_27_port, S(26) => PTMP_3_26_port, S(25) => 
                           PTMP_3_25_port, S(24) => PTMP_3_24_port, S(23) => 
                           PTMP_3_23_port, S(22) => PTMP_3_22_port, S(21) => 
                           PTMP_3_21_port, S(20) => PTMP_3_20_port, S(19) => 
                           PTMP_3_19_port, S(18) => PTMP_3_18_port, S(17) => 
                           PTMP_3_17_port, S(16) => PTMP_3_16_port, S(15) => 
                           PTMP_3_15_port, S(14) => PTMP_3_14_port, S(13) => 
                           PTMP_3_13_port, S(12) => PTMP_3_12_port, S(11) => 
                           PTMP_3_11_port, S(10) => PTMP_3_10_port, S(9) => 
                           PTMP_3_9_port, S(8) => PTMP_3_8_port, S(7) => 
                           PTMP_3_7_port, S(6) => PTMP_3_6_port, S(5) => 
                           PTMP_3_5_port, S(4) => PTMP_3_4_port, S(3) => 
                           PTMP_3_3_port, S(2) => PTMP_3_2_port, S(1) => 
                           PTMP_3_1_port, S(0) => PTMP_3_0_port, Co => n_1284);
   ADDER_5 : RCA_NBIT44 port map( A(43) => n16, A(42) => n16, A(41) => 
                           PTMP_3_41_port, A(40) => PTMP_3_40_port, A(39) => 
                           PTMP_3_39_port, A(38) => PTMP_3_38_port, A(37) => 
                           PTMP_3_37_port, A(36) => PTMP_3_36_port, A(35) => 
                           PTMP_3_35_port, A(34) => PTMP_3_34_port, A(33) => 
                           PTMP_3_33_port, A(32) => PTMP_3_32_port, A(31) => 
                           PTMP_3_31_port, A(30) => PTMP_3_30_port, A(29) => 
                           PTMP_3_29_port, A(28) => PTMP_3_28_port, A(27) => 
                           PTMP_3_27_port, A(26) => PTMP_3_26_port, A(25) => 
                           PTMP_3_25_port, A(24) => PTMP_3_24_port, A(23) => 
                           PTMP_3_23_port, A(22) => PTMP_3_22_port, A(21) => 
                           PTMP_3_21_port, A(20) => PTMP_3_20_port, A(19) => 
                           PTMP_3_19_port, A(18) => PTMP_3_18_port, A(17) => 
                           PTMP_3_17_port, A(16) => PTMP_3_16_port, A(15) => 
                           PTMP_3_15_port, A(14) => PTMP_3_14_port, A(13) => 
                           PTMP_3_13_port, A(12) => PTMP_3_12_port, A(11) => 
                           PTMP_3_11_port, A(10) => PTMP_3_10_port, A(9) => 
                           PTMP_3_9_port, A(8) => PTMP_3_8_port, A(7) => 
                           PTMP_3_7_port, A(6) => PTMP_3_6_port, A(5) => 
                           PTMP_3_5_port, A(4) => PTMP_3_4_port, A(3) => 
                           PTMP_3_3_port, A(2) => PTMP_3_2_port, A(1) => 
                           PTMP_3_1_port, A(0) => PTMP_3_0_port, B(43) => 
                           OTMP_5_43_port, B(42) => OTMP_5_42_port, B(41) => 
                           OTMP_5_41_port, B(40) => OTMP_5_40_port, B(39) => 
                           OTMP_5_39_port, B(38) => OTMP_5_38_port, B(37) => 
                           OTMP_5_37_port, B(36) => OTMP_5_36_port, B(35) => 
                           OTMP_5_35_port, B(34) => OTMP_5_34_port, B(33) => 
                           OTMP_5_33_port, B(32) => OTMP_5_32_port, B(31) => 
                           OTMP_5_31_port, B(30) => OTMP_5_30_port, B(29) => 
                           OTMP_5_29_port, B(28) => OTMP_5_28_port, B(27) => 
                           OTMP_5_27_port, B(26) => OTMP_5_26_port, B(25) => 
                           OTMP_5_25_port, B(24) => OTMP_5_24_port, B(23) => 
                           OTMP_5_23_port, B(22) => OTMP_5_22_port, B(21) => 
                           OTMP_5_21_port, B(20) => OTMP_5_20_port, B(19) => 
                           OTMP_5_19_port, B(18) => OTMP_5_18_port, B(17) => 
                           OTMP_5_17_port, B(16) => OTMP_5_16_port, B(15) => 
                           OTMP_5_15_port, B(14) => OTMP_5_14_port, B(13) => 
                           OTMP_5_13_port, B(12) => OTMP_5_12_port, B(11) => 
                           OTMP_5_11_port, B(10) => OTMP_5_10_port, B(9) => 
                           OTMP_5_9_port, B(8) => OTMP_5_8_port, B(7) => 
                           OTMP_5_7_port, B(6) => OTMP_5_6_port, B(5) => 
                           OTMP_5_5_port, B(4) => OTMP_5_4_port, B(3) => 
                           OTMP_5_3_port, B(2) => OTMP_5_2_port, B(1) => 
                           OTMP_5_1_port, B(0) => OTMP_5_0_port, Ci => 
                           X_Logic0_port, S(43) => PTMP_4_43_port, S(42) => 
                           PTMP_4_42_port, S(41) => PTMP_4_41_port, S(40) => 
                           PTMP_4_40_port, S(39) => PTMP_4_39_port, S(38) => 
                           PTMP_4_38_port, S(37) => PTMP_4_37_port, S(36) => 
                           PTMP_4_36_port, S(35) => PTMP_4_35_port, S(34) => 
                           PTMP_4_34_port, S(33) => PTMP_4_33_port, S(32) => 
                           PTMP_4_32_port, S(31) => PTMP_4_31_port, S(30) => 
                           PTMP_4_30_port, S(29) => PTMP_4_29_port, S(28) => 
                           PTMP_4_28_port, S(27) => PTMP_4_27_port, S(26) => 
                           PTMP_4_26_port, S(25) => PTMP_4_25_port, S(24) => 
                           PTMP_4_24_port, S(23) => PTMP_4_23_port, S(22) => 
                           PTMP_4_22_port, S(21) => PTMP_4_21_port, S(20) => 
                           PTMP_4_20_port, S(19) => PTMP_4_19_port, S(18) => 
                           PTMP_4_18_port, S(17) => PTMP_4_17_port, S(16) => 
                           PTMP_4_16_port, S(15) => PTMP_4_15_port, S(14) => 
                           PTMP_4_14_port, S(13) => PTMP_4_13_port, S(12) => 
                           PTMP_4_12_port, S(11) => PTMP_4_11_port, S(10) => 
                           PTMP_4_10_port, S(9) => PTMP_4_9_port, S(8) => 
                           PTMP_4_8_port, S(7) => PTMP_4_7_port, S(6) => 
                           PTMP_4_6_port, S(5) => PTMP_4_5_port, S(4) => 
                           PTMP_4_4_port, S(3) => PTMP_4_3_port, S(2) => 
                           PTMP_4_2_port, S(1) => PTMP_4_1_port, S(0) => 
                           PTMP_4_0_port, Co => n_1285);
   ADDER_6 : RCA_NBIT46 port map( A(45) => n12, A(44) => n12, A(43) => 
                           PTMP_4_43_port, A(42) => PTMP_4_42_port, A(41) => 
                           PTMP_4_41_port, A(40) => PTMP_4_40_port, A(39) => 
                           PTMP_4_39_port, A(38) => PTMP_4_38_port, A(37) => 
                           PTMP_4_37_port, A(36) => PTMP_4_36_port, A(35) => 
                           PTMP_4_35_port, A(34) => PTMP_4_34_port, A(33) => 
                           PTMP_4_33_port, A(32) => PTMP_4_32_port, A(31) => 
                           PTMP_4_31_port, A(30) => PTMP_4_30_port, A(29) => 
                           PTMP_4_29_port, A(28) => PTMP_4_28_port, A(27) => 
                           PTMP_4_27_port, A(26) => PTMP_4_26_port, A(25) => 
                           PTMP_4_25_port, A(24) => PTMP_4_24_port, A(23) => 
                           PTMP_4_23_port, A(22) => PTMP_4_22_port, A(21) => 
                           PTMP_4_21_port, A(20) => PTMP_4_20_port, A(19) => 
                           PTMP_4_19_port, A(18) => PTMP_4_18_port, A(17) => 
                           PTMP_4_17_port, A(16) => PTMP_4_16_port, A(15) => 
                           PTMP_4_15_port, A(14) => PTMP_4_14_port, A(13) => 
                           PTMP_4_13_port, A(12) => PTMP_4_12_port, A(11) => 
                           PTMP_4_11_port, A(10) => PTMP_4_10_port, A(9) => 
                           PTMP_4_9_port, A(8) => PTMP_4_8_port, A(7) => 
                           PTMP_4_7_port, A(6) => PTMP_4_6_port, A(5) => 
                           PTMP_4_5_port, A(4) => PTMP_4_4_port, A(3) => 
                           PTMP_4_3_port, A(2) => PTMP_4_2_port, A(1) => 
                           PTMP_4_1_port, A(0) => PTMP_4_0_port, B(45) => 
                           OTMP_6_45_port, B(44) => OTMP_6_44_port, B(43) => 
                           OTMP_6_43_port, B(42) => OTMP_6_42_port, B(41) => 
                           OTMP_6_41_port, B(40) => OTMP_6_40_port, B(39) => 
                           OTMP_6_39_port, B(38) => OTMP_6_38_port, B(37) => 
                           OTMP_6_37_port, B(36) => OTMP_6_36_port, B(35) => 
                           OTMP_6_35_port, B(34) => OTMP_6_34_port, B(33) => 
                           OTMP_6_33_port, B(32) => OTMP_6_32_port, B(31) => 
                           OTMP_6_31_port, B(30) => OTMP_6_30_port, B(29) => 
                           OTMP_6_29_port, B(28) => OTMP_6_28_port, B(27) => 
                           OTMP_6_27_port, B(26) => OTMP_6_26_port, B(25) => 
                           OTMP_6_25_port, B(24) => OTMP_6_24_port, B(23) => 
                           OTMP_6_23_port, B(22) => OTMP_6_22_port, B(21) => 
                           OTMP_6_21_port, B(20) => OTMP_6_20_port, B(19) => 
                           OTMP_6_19_port, B(18) => OTMP_6_18_port, B(17) => 
                           OTMP_6_17_port, B(16) => OTMP_6_16_port, B(15) => 
                           OTMP_6_15_port, B(14) => OTMP_6_14_port, B(13) => 
                           OTMP_6_13_port, B(12) => OTMP_6_12_port, B(11) => 
                           OTMP_6_11_port, B(10) => OTMP_6_10_port, B(9) => 
                           OTMP_6_9_port, B(8) => OTMP_6_8_port, B(7) => 
                           OTMP_6_7_port, B(6) => OTMP_6_6_port, B(5) => 
                           OTMP_6_5_port, B(4) => OTMP_6_4_port, B(3) => 
                           OTMP_6_3_port, B(2) => OTMP_6_2_port, B(1) => 
                           OTMP_6_1_port, B(0) => OTMP_6_0_port, Ci => 
                           X_Logic0_port, S(45) => PTMP_5_45_port, S(44) => 
                           PTMP_5_44_port, S(43) => PTMP_5_43_port, S(42) => 
                           PTMP_5_42_port, S(41) => PTMP_5_41_port, S(40) => 
                           PTMP_5_40_port, S(39) => PTMP_5_39_port, S(38) => 
                           PTMP_5_38_port, S(37) => PTMP_5_37_port, S(36) => 
                           PTMP_5_36_port, S(35) => PTMP_5_35_port, S(34) => 
                           PTMP_5_34_port, S(33) => PTMP_5_33_port, S(32) => 
                           PTMP_5_32_port, S(31) => PTMP_5_31_port, S(30) => 
                           PTMP_5_30_port, S(29) => PTMP_5_29_port, S(28) => 
                           PTMP_5_28_port, S(27) => PTMP_5_27_port, S(26) => 
                           PTMP_5_26_port, S(25) => PTMP_5_25_port, S(24) => 
                           PTMP_5_24_port, S(23) => PTMP_5_23_port, S(22) => 
                           PTMP_5_22_port, S(21) => PTMP_5_21_port, S(20) => 
                           PTMP_5_20_port, S(19) => PTMP_5_19_port, S(18) => 
                           PTMP_5_18_port, S(17) => PTMP_5_17_port, S(16) => 
                           PTMP_5_16_port, S(15) => PTMP_5_15_port, S(14) => 
                           PTMP_5_14_port, S(13) => PTMP_5_13_port, S(12) => 
                           PTMP_5_12_port, S(11) => PTMP_5_11_port, S(10) => 
                           PTMP_5_10_port, S(9) => PTMP_5_9_port, S(8) => 
                           PTMP_5_8_port, S(7) => PTMP_5_7_port, S(6) => 
                           PTMP_5_6_port, S(5) => PTMP_5_5_port, S(4) => 
                           PTMP_5_4_port, S(3) => PTMP_5_3_port, S(2) => 
                           PTMP_5_2_port, S(1) => PTMP_5_1_port, S(0) => 
                           PTMP_5_0_port, Co => n_1286);
   ADDER_7 : RCA_NBIT48 port map( A(47) => n15, A(46) => n15, A(45) => 
                           PTMP_5_45_port, A(44) => PTMP_5_44_port, A(43) => 
                           PTMP_5_43_port, A(42) => PTMP_5_42_port, A(41) => 
                           PTMP_5_41_port, A(40) => PTMP_5_40_port, A(39) => 
                           PTMP_5_39_port, A(38) => PTMP_5_38_port, A(37) => 
                           PTMP_5_37_port, A(36) => PTMP_5_36_port, A(35) => 
                           PTMP_5_35_port, A(34) => PTMP_5_34_port, A(33) => 
                           PTMP_5_33_port, A(32) => PTMP_5_32_port, A(31) => 
                           PTMP_5_31_port, A(30) => PTMP_5_30_port, A(29) => 
                           PTMP_5_29_port, A(28) => PTMP_5_28_port, A(27) => 
                           PTMP_5_27_port, A(26) => PTMP_5_26_port, A(25) => 
                           PTMP_5_25_port, A(24) => PTMP_5_24_port, A(23) => 
                           PTMP_5_23_port, A(22) => PTMP_5_22_port, A(21) => 
                           PTMP_5_21_port, A(20) => PTMP_5_20_port, A(19) => 
                           PTMP_5_19_port, A(18) => PTMP_5_18_port, A(17) => 
                           PTMP_5_17_port, A(16) => PTMP_5_16_port, A(15) => 
                           PTMP_5_15_port, A(14) => PTMP_5_14_port, A(13) => 
                           PTMP_5_13_port, A(12) => PTMP_5_12_port, A(11) => 
                           PTMP_5_11_port, A(10) => PTMP_5_10_port, A(9) => 
                           PTMP_5_9_port, A(8) => PTMP_5_8_port, A(7) => 
                           PTMP_5_7_port, A(6) => PTMP_5_6_port, A(5) => 
                           PTMP_5_5_port, A(4) => PTMP_5_4_port, A(3) => 
                           PTMP_5_3_port, A(2) => PTMP_5_2_port, A(1) => 
                           PTMP_5_1_port, A(0) => PTMP_5_0_port, B(47) => 
                           OTMP_7_47_port, B(46) => OTMP_7_46_port, B(45) => 
                           OTMP_7_45_port, B(44) => OTMP_7_44_port, B(43) => 
                           OTMP_7_43_port, B(42) => OTMP_7_42_port, B(41) => 
                           OTMP_7_41_port, B(40) => OTMP_7_40_port, B(39) => 
                           OTMP_7_39_port, B(38) => OTMP_7_38_port, B(37) => 
                           OTMP_7_37_port, B(36) => OTMP_7_36_port, B(35) => 
                           OTMP_7_35_port, B(34) => OTMP_7_34_port, B(33) => 
                           OTMP_7_33_port, B(32) => OTMP_7_32_port, B(31) => 
                           OTMP_7_31_port, B(30) => OTMP_7_30_port, B(29) => 
                           OTMP_7_29_port, B(28) => OTMP_7_28_port, B(27) => 
                           OTMP_7_27_port, B(26) => OTMP_7_26_port, B(25) => 
                           OTMP_7_25_port, B(24) => OTMP_7_24_port, B(23) => 
                           OTMP_7_23_port, B(22) => OTMP_7_22_port, B(21) => 
                           OTMP_7_21_port, B(20) => OTMP_7_20_port, B(19) => 
                           OTMP_7_19_port, B(18) => OTMP_7_18_port, B(17) => 
                           OTMP_7_17_port, B(16) => OTMP_7_16_port, B(15) => 
                           OTMP_7_15_port, B(14) => OTMP_7_14_port, B(13) => 
                           OTMP_7_13_port, B(12) => OTMP_7_12_port, B(11) => 
                           OTMP_7_11_port, B(10) => OTMP_7_10_port, B(9) => 
                           OTMP_7_9_port, B(8) => OTMP_7_8_port, B(7) => 
                           OTMP_7_7_port, B(6) => OTMP_7_6_port, B(5) => 
                           OTMP_7_5_port, B(4) => OTMP_7_4_port, B(3) => 
                           OTMP_7_3_port, B(2) => OTMP_7_2_port, B(1) => 
                           OTMP_7_1_port, B(0) => OTMP_7_0_port, Ci => 
                           X_Logic0_port, S(47) => PTMP_6_47_port, S(46) => 
                           PTMP_6_46_port, S(45) => PTMP_6_45_port, S(44) => 
                           PTMP_6_44_port, S(43) => PTMP_6_43_port, S(42) => 
                           PTMP_6_42_port, S(41) => PTMP_6_41_port, S(40) => 
                           PTMP_6_40_port, S(39) => PTMP_6_39_port, S(38) => 
                           PTMP_6_38_port, S(37) => PTMP_6_37_port, S(36) => 
                           PTMP_6_36_port, S(35) => PTMP_6_35_port, S(34) => 
                           PTMP_6_34_port, S(33) => PTMP_6_33_port, S(32) => 
                           PTMP_6_32_port, S(31) => PTMP_6_31_port, S(30) => 
                           PTMP_6_30_port, S(29) => PTMP_6_29_port, S(28) => 
                           PTMP_6_28_port, S(27) => PTMP_6_27_port, S(26) => 
                           PTMP_6_26_port, S(25) => PTMP_6_25_port, S(24) => 
                           PTMP_6_24_port, S(23) => PTMP_6_23_port, S(22) => 
                           PTMP_6_22_port, S(21) => PTMP_6_21_port, S(20) => 
                           PTMP_6_20_port, S(19) => PTMP_6_19_port, S(18) => 
                           PTMP_6_18_port, S(17) => PTMP_6_17_port, S(16) => 
                           PTMP_6_16_port, S(15) => PTMP_6_15_port, S(14) => 
                           PTMP_6_14_port, S(13) => PTMP_6_13_port, S(12) => 
                           PTMP_6_12_port, S(11) => PTMP_6_11_port, S(10) => 
                           PTMP_6_10_port, S(9) => PTMP_6_9_port, S(8) => 
                           PTMP_6_8_port, S(7) => PTMP_6_7_port, S(6) => 
                           PTMP_6_6_port, S(5) => PTMP_6_5_port, S(4) => 
                           PTMP_6_4_port, S(3) => PTMP_6_3_port, S(2) => 
                           PTMP_6_2_port, S(1) => PTMP_6_1_port, S(0) => 
                           PTMP_6_0_port, Co => n_1287);
   ADDER_8 : RCA_NBIT50 port map( A(49) => n6, A(48) => n6, A(47) => 
                           PTMP_6_47_port, A(46) => PTMP_6_46_port, A(45) => 
                           PTMP_6_45_port, A(44) => PTMP_6_44_port, A(43) => 
                           PTMP_6_43_port, A(42) => PTMP_6_42_port, A(41) => 
                           PTMP_6_41_port, A(40) => PTMP_6_40_port, A(39) => 
                           PTMP_6_39_port, A(38) => PTMP_6_38_port, A(37) => 
                           PTMP_6_37_port, A(36) => PTMP_6_36_port, A(35) => 
                           PTMP_6_35_port, A(34) => PTMP_6_34_port, A(33) => 
                           PTMP_6_33_port, A(32) => PTMP_6_32_port, A(31) => 
                           PTMP_6_31_port, A(30) => PTMP_6_30_port, A(29) => 
                           PTMP_6_29_port, A(28) => PTMP_6_28_port, A(27) => 
                           PTMP_6_27_port, A(26) => PTMP_6_26_port, A(25) => 
                           PTMP_6_25_port, A(24) => PTMP_6_24_port, A(23) => 
                           PTMP_6_23_port, A(22) => PTMP_6_22_port, A(21) => 
                           PTMP_6_21_port, A(20) => PTMP_6_20_port, A(19) => 
                           PTMP_6_19_port, A(18) => PTMP_6_18_port, A(17) => 
                           PTMP_6_17_port, A(16) => PTMP_6_16_port, A(15) => 
                           PTMP_6_15_port, A(14) => PTMP_6_14_port, A(13) => 
                           PTMP_6_13_port, A(12) => PTMP_6_12_port, A(11) => 
                           PTMP_6_11_port, A(10) => PTMP_6_10_port, A(9) => 
                           PTMP_6_9_port, A(8) => PTMP_6_8_port, A(7) => 
                           PTMP_6_7_port, A(6) => PTMP_6_6_port, A(5) => 
                           PTMP_6_5_port, A(4) => PTMP_6_4_port, A(3) => 
                           PTMP_6_3_port, A(2) => PTMP_6_2_port, A(1) => 
                           PTMP_6_1_port, A(0) => PTMP_6_0_port, B(49) => 
                           OTMP_8_49_port, B(48) => OTMP_8_48_port, B(47) => 
                           OTMP_8_47_port, B(46) => OTMP_8_46_port, B(45) => 
                           OTMP_8_45_port, B(44) => OTMP_8_44_port, B(43) => 
                           OTMP_8_43_port, B(42) => OTMP_8_42_port, B(41) => 
                           OTMP_8_41_port, B(40) => OTMP_8_40_port, B(39) => 
                           OTMP_8_39_port, B(38) => OTMP_8_38_port, B(37) => 
                           OTMP_8_37_port, B(36) => OTMP_8_36_port, B(35) => 
                           OTMP_8_35_port, B(34) => OTMP_8_34_port, B(33) => 
                           OTMP_8_33_port, B(32) => OTMP_8_32_port, B(31) => 
                           OTMP_8_31_port, B(30) => OTMP_8_30_port, B(29) => 
                           OTMP_8_29_port, B(28) => OTMP_8_28_port, B(27) => 
                           OTMP_8_27_port, B(26) => OTMP_8_26_port, B(25) => 
                           OTMP_8_25_port, B(24) => OTMP_8_24_port, B(23) => 
                           OTMP_8_23_port, B(22) => OTMP_8_22_port, B(21) => 
                           OTMP_8_21_port, B(20) => OTMP_8_20_port, B(19) => 
                           OTMP_8_19_port, B(18) => OTMP_8_18_port, B(17) => 
                           OTMP_8_17_port, B(16) => OTMP_8_16_port, B(15) => 
                           OTMP_8_15_port, B(14) => OTMP_8_14_port, B(13) => 
                           OTMP_8_13_port, B(12) => OTMP_8_12_port, B(11) => 
                           OTMP_8_11_port, B(10) => OTMP_8_10_port, B(9) => 
                           OTMP_8_9_port, B(8) => OTMP_8_8_port, B(7) => 
                           OTMP_8_7_port, B(6) => OTMP_8_6_port, B(5) => 
                           OTMP_8_5_port, B(4) => OTMP_8_4_port, B(3) => 
                           OTMP_8_3_port, B(2) => OTMP_8_2_port, B(1) => 
                           OTMP_8_1_port, B(0) => OTMP_8_0_port, Ci => 
                           X_Logic0_port, S(49) => PTMP_7_49_port, S(48) => 
                           PTMP_7_48_port, S(47) => PTMP_7_47_port, S(46) => 
                           PTMP_7_46_port, S(45) => PTMP_7_45_port, S(44) => 
                           PTMP_7_44_port, S(43) => PTMP_7_43_port, S(42) => 
                           PTMP_7_42_port, S(41) => PTMP_7_41_port, S(40) => 
                           PTMP_7_40_port, S(39) => PTMP_7_39_port, S(38) => 
                           PTMP_7_38_port, S(37) => PTMP_7_37_port, S(36) => 
                           PTMP_7_36_port, S(35) => PTMP_7_35_port, S(34) => 
                           PTMP_7_34_port, S(33) => PTMP_7_33_port, S(32) => 
                           PTMP_7_32_port, S(31) => PTMP_7_31_port, S(30) => 
                           PTMP_7_30_port, S(29) => PTMP_7_29_port, S(28) => 
                           PTMP_7_28_port, S(27) => PTMP_7_27_port, S(26) => 
                           PTMP_7_26_port, S(25) => PTMP_7_25_port, S(24) => 
                           PTMP_7_24_port, S(23) => PTMP_7_23_port, S(22) => 
                           PTMP_7_22_port, S(21) => PTMP_7_21_port, S(20) => 
                           PTMP_7_20_port, S(19) => PTMP_7_19_port, S(18) => 
                           PTMP_7_18_port, S(17) => PTMP_7_17_port, S(16) => 
                           PTMP_7_16_port, S(15) => PTMP_7_15_port, S(14) => 
                           PTMP_7_14_port, S(13) => PTMP_7_13_port, S(12) => 
                           PTMP_7_12_port, S(11) => PTMP_7_11_port, S(10) => 
                           PTMP_7_10_port, S(9) => PTMP_7_9_port, S(8) => 
                           PTMP_7_8_port, S(7) => PTMP_7_7_port, S(6) => 
                           PTMP_7_6_port, S(5) => PTMP_7_5_port, S(4) => 
                           PTMP_7_4_port, S(3) => PTMP_7_3_port, S(2) => 
                           PTMP_7_2_port, S(1) => PTMP_7_1_port, S(0) => 
                           PTMP_7_0_port, Co => n_1288);
   ADDER_9 : RCA_NBIT52 port map( A(51) => n10, A(50) => n10, A(49) => 
                           PTMP_7_49_port, A(48) => PTMP_7_48_port, A(47) => 
                           PTMP_7_47_port, A(46) => PTMP_7_46_port, A(45) => 
                           PTMP_7_45_port, A(44) => PTMP_7_44_port, A(43) => 
                           PTMP_7_43_port, A(42) => PTMP_7_42_port, A(41) => 
                           PTMP_7_41_port, A(40) => PTMP_7_40_port, A(39) => 
                           PTMP_7_39_port, A(38) => PTMP_7_38_port, A(37) => 
                           PTMP_7_37_port, A(36) => PTMP_7_36_port, A(35) => 
                           PTMP_7_35_port, A(34) => PTMP_7_34_port, A(33) => 
                           PTMP_7_33_port, A(32) => PTMP_7_32_port, A(31) => 
                           PTMP_7_31_port, A(30) => PTMP_7_30_port, A(29) => 
                           PTMP_7_29_port, A(28) => PTMP_7_28_port, A(27) => 
                           PTMP_7_27_port, A(26) => PTMP_7_26_port, A(25) => 
                           PTMP_7_25_port, A(24) => PTMP_7_24_port, A(23) => 
                           PTMP_7_23_port, A(22) => PTMP_7_22_port, A(21) => 
                           PTMP_7_21_port, A(20) => PTMP_7_20_port, A(19) => 
                           PTMP_7_19_port, A(18) => PTMP_7_18_port, A(17) => 
                           PTMP_7_17_port, A(16) => PTMP_7_16_port, A(15) => 
                           PTMP_7_15_port, A(14) => PTMP_7_14_port, A(13) => 
                           PTMP_7_13_port, A(12) => PTMP_7_12_port, A(11) => 
                           PTMP_7_11_port, A(10) => PTMP_7_10_port, A(9) => 
                           PTMP_7_9_port, A(8) => PTMP_7_8_port, A(7) => 
                           PTMP_7_7_port, A(6) => PTMP_7_6_port, A(5) => 
                           PTMP_7_5_port, A(4) => PTMP_7_4_port, A(3) => 
                           PTMP_7_3_port, A(2) => PTMP_7_2_port, A(1) => 
                           PTMP_7_1_port, A(0) => PTMP_7_0_port, B(51) => 
                           OTMP_9_51_port, B(50) => OTMP_9_50_port, B(49) => 
                           OTMP_9_49_port, B(48) => OTMP_9_48_port, B(47) => 
                           OTMP_9_47_port, B(46) => OTMP_9_46_port, B(45) => 
                           OTMP_9_45_port, B(44) => OTMP_9_44_port, B(43) => 
                           OTMP_9_43_port, B(42) => OTMP_9_42_port, B(41) => 
                           OTMP_9_41_port, B(40) => OTMP_9_40_port, B(39) => 
                           OTMP_9_39_port, B(38) => OTMP_9_38_port, B(37) => 
                           OTMP_9_37_port, B(36) => OTMP_9_36_port, B(35) => 
                           OTMP_9_35_port, B(34) => OTMP_9_34_port, B(33) => 
                           OTMP_9_33_port, B(32) => OTMP_9_32_port, B(31) => 
                           OTMP_9_31_port, B(30) => OTMP_9_30_port, B(29) => 
                           OTMP_9_29_port, B(28) => OTMP_9_28_port, B(27) => 
                           OTMP_9_27_port, B(26) => OTMP_9_26_port, B(25) => 
                           OTMP_9_25_port, B(24) => OTMP_9_24_port, B(23) => 
                           OTMP_9_23_port, B(22) => OTMP_9_22_port, B(21) => 
                           OTMP_9_21_port, B(20) => OTMP_9_20_port, B(19) => 
                           OTMP_9_19_port, B(18) => OTMP_9_18_port, B(17) => 
                           OTMP_9_17_port, B(16) => OTMP_9_16_port, B(15) => 
                           OTMP_9_15_port, B(14) => OTMP_9_14_port, B(13) => 
                           OTMP_9_13_port, B(12) => OTMP_9_12_port, B(11) => 
                           OTMP_9_11_port, B(10) => OTMP_9_10_port, B(9) => 
                           OTMP_9_9_port, B(8) => OTMP_9_8_port, B(7) => 
                           OTMP_9_7_port, B(6) => OTMP_9_6_port, B(5) => 
                           OTMP_9_5_port, B(4) => OTMP_9_4_port, B(3) => 
                           OTMP_9_3_port, B(2) => OTMP_9_2_port, B(1) => 
                           OTMP_9_1_port, B(0) => OTMP_9_0_port, Ci => 
                           X_Logic0_port, S(51) => PTMP_8_51_port, S(50) => 
                           PTMP_8_50_port, S(49) => PTMP_8_49_port, S(48) => 
                           PTMP_8_48_port, S(47) => PTMP_8_47_port, S(46) => 
                           PTMP_8_46_port, S(45) => PTMP_8_45_port, S(44) => 
                           PTMP_8_44_port, S(43) => PTMP_8_43_port, S(42) => 
                           PTMP_8_42_port, S(41) => PTMP_8_41_port, S(40) => 
                           PTMP_8_40_port, S(39) => PTMP_8_39_port, S(38) => 
                           PTMP_8_38_port, S(37) => PTMP_8_37_port, S(36) => 
                           PTMP_8_36_port, S(35) => PTMP_8_35_port, S(34) => 
                           PTMP_8_34_port, S(33) => PTMP_8_33_port, S(32) => 
                           PTMP_8_32_port, S(31) => PTMP_8_31_port, S(30) => 
                           PTMP_8_30_port, S(29) => PTMP_8_29_port, S(28) => 
                           PTMP_8_28_port, S(27) => PTMP_8_27_port, S(26) => 
                           PTMP_8_26_port, S(25) => PTMP_8_25_port, S(24) => 
                           PTMP_8_24_port, S(23) => PTMP_8_23_port, S(22) => 
                           PTMP_8_22_port, S(21) => PTMP_8_21_port, S(20) => 
                           PTMP_8_20_port, S(19) => PTMP_8_19_port, S(18) => 
                           PTMP_8_18_port, S(17) => PTMP_8_17_port, S(16) => 
                           PTMP_8_16_port, S(15) => PTMP_8_15_port, S(14) => 
                           PTMP_8_14_port, S(13) => PTMP_8_13_port, S(12) => 
                           PTMP_8_12_port, S(11) => PTMP_8_11_port, S(10) => 
                           PTMP_8_10_port, S(9) => PTMP_8_9_port, S(8) => 
                           PTMP_8_8_port, S(7) => PTMP_8_7_port, S(6) => 
                           PTMP_8_6_port, S(5) => PTMP_8_5_port, S(4) => 
                           PTMP_8_4_port, S(3) => PTMP_8_3_port, S(2) => 
                           PTMP_8_2_port, S(1) => PTMP_8_1_port, S(0) => 
                           PTMP_8_0_port, Co => n_1289);
   ADDER_10 : RCA_NBIT54 port map( A(53) => PTMP_8_51_port, A(52) => 
                           PTMP_8_51_port, A(51) => PTMP_8_51_port, A(50) => 
                           PTMP_8_50_port, A(49) => PTMP_8_49_port, A(48) => 
                           PTMP_8_48_port, A(47) => PTMP_8_47_port, A(46) => 
                           PTMP_8_46_port, A(45) => PTMP_8_45_port, A(44) => 
                           PTMP_8_44_port, A(43) => PTMP_8_43_port, A(42) => 
                           PTMP_8_42_port, A(41) => PTMP_8_41_port, A(40) => 
                           PTMP_8_40_port, A(39) => PTMP_8_39_port, A(38) => 
                           PTMP_8_38_port, A(37) => PTMP_8_37_port, A(36) => 
                           PTMP_8_36_port, A(35) => PTMP_8_35_port, A(34) => 
                           PTMP_8_34_port, A(33) => PTMP_8_33_port, A(32) => 
                           PTMP_8_32_port, A(31) => PTMP_8_31_port, A(30) => 
                           PTMP_8_30_port, A(29) => PTMP_8_29_port, A(28) => 
                           PTMP_8_28_port, A(27) => PTMP_8_27_port, A(26) => 
                           PTMP_8_26_port, A(25) => PTMP_8_25_port, A(24) => 
                           PTMP_8_24_port, A(23) => PTMP_8_23_port, A(22) => 
                           PTMP_8_22_port, A(21) => PTMP_8_21_port, A(20) => 
                           PTMP_8_20_port, A(19) => PTMP_8_19_port, A(18) => 
                           PTMP_8_18_port, A(17) => PTMP_8_17_port, A(16) => 
                           PTMP_8_16_port, A(15) => PTMP_8_15_port, A(14) => 
                           PTMP_8_14_port, A(13) => PTMP_8_13_port, A(12) => 
                           PTMP_8_12_port, A(11) => PTMP_8_11_port, A(10) => 
                           PTMP_8_10_port, A(9) => PTMP_8_9_port, A(8) => 
                           PTMP_8_8_port, A(7) => PTMP_8_7_port, A(6) => 
                           PTMP_8_6_port, A(5) => PTMP_8_5_port, A(4) => 
                           PTMP_8_4_port, A(3) => PTMP_8_3_port, A(2) => 
                           PTMP_8_2_port, A(1) => PTMP_8_1_port, A(0) => 
                           PTMP_8_0_port, B(53) => OTMP_10_53_port, B(52) => 
                           OTMP_10_52_port, B(51) => OTMP_10_51_port, B(50) => 
                           OTMP_10_50_port, B(49) => OTMP_10_49_port, B(48) => 
                           OTMP_10_48_port, B(47) => OTMP_10_47_port, B(46) => 
                           OTMP_10_46_port, B(45) => OTMP_10_45_port, B(44) => 
                           OTMP_10_44_port, B(43) => OTMP_10_43_port, B(42) => 
                           OTMP_10_42_port, B(41) => OTMP_10_41_port, B(40) => 
                           OTMP_10_40_port, B(39) => OTMP_10_39_port, B(38) => 
                           OTMP_10_38_port, B(37) => OTMP_10_37_port, B(36) => 
                           OTMP_10_36_port, B(35) => OTMP_10_35_port, B(34) => 
                           OTMP_10_34_port, B(33) => OTMP_10_33_port, B(32) => 
                           OTMP_10_32_port, B(31) => OTMP_10_31_port, B(30) => 
                           OTMP_10_30_port, B(29) => OTMP_10_29_port, B(28) => 
                           OTMP_10_28_port, B(27) => OTMP_10_27_port, B(26) => 
                           OTMP_10_26_port, B(25) => OTMP_10_25_port, B(24) => 
                           OTMP_10_24_port, B(23) => OTMP_10_23_port, B(22) => 
                           OTMP_10_22_port, B(21) => OTMP_10_21_port, B(20) => 
                           OTMP_10_20_port, B(19) => OTMP_10_19_port, B(18) => 
                           OTMP_10_18_port, B(17) => OTMP_10_17_port, B(16) => 
                           OTMP_10_16_port, B(15) => OTMP_10_15_port, B(14) => 
                           OTMP_10_14_port, B(13) => OTMP_10_13_port, B(12) => 
                           OTMP_10_12_port, B(11) => OTMP_10_11_port, B(10) => 
                           OTMP_10_10_port, B(9) => OTMP_10_9_port, B(8) => 
                           OTMP_10_8_port, B(7) => OTMP_10_7_port, B(6) => 
                           OTMP_10_6_port, B(5) => OTMP_10_5_port, B(4) => 
                           OTMP_10_4_port, B(3) => OTMP_10_3_port, B(2) => 
                           OTMP_10_2_port, B(1) => OTMP_10_1_port, B(0) => 
                           OTMP_10_0_port, Ci => X_Logic0_port, S(53) => 
                           PTMP_9_53_port, S(52) => PTMP_9_52_port, S(51) => 
                           PTMP_9_51_port, S(50) => PTMP_9_50_port, S(49) => 
                           PTMP_9_49_port, S(48) => PTMP_9_48_port, S(47) => 
                           PTMP_9_47_port, S(46) => PTMP_9_46_port, S(45) => 
                           PTMP_9_45_port, S(44) => PTMP_9_44_port, S(43) => 
                           PTMP_9_43_port, S(42) => PTMP_9_42_port, S(41) => 
                           PTMP_9_41_port, S(40) => PTMP_9_40_port, S(39) => 
                           PTMP_9_39_port, S(38) => PTMP_9_38_port, S(37) => 
                           PTMP_9_37_port, S(36) => PTMP_9_36_port, S(35) => 
                           PTMP_9_35_port, S(34) => PTMP_9_34_port, S(33) => 
                           PTMP_9_33_port, S(32) => PTMP_9_32_port, S(31) => 
                           PTMP_9_31_port, S(30) => PTMP_9_30_port, S(29) => 
                           PTMP_9_29_port, S(28) => PTMP_9_28_port, S(27) => 
                           PTMP_9_27_port, S(26) => PTMP_9_26_port, S(25) => 
                           PTMP_9_25_port, S(24) => PTMP_9_24_port, S(23) => 
                           PTMP_9_23_port, S(22) => PTMP_9_22_port, S(21) => 
                           PTMP_9_21_port, S(20) => PTMP_9_20_port, S(19) => 
                           PTMP_9_19_port, S(18) => PTMP_9_18_port, S(17) => 
                           PTMP_9_17_port, S(16) => PTMP_9_16_port, S(15) => 
                           PTMP_9_15_port, S(14) => PTMP_9_14_port, S(13) => 
                           PTMP_9_13_port, S(12) => PTMP_9_12_port, S(11) => 
                           PTMP_9_11_port, S(10) => PTMP_9_10_port, S(9) => 
                           PTMP_9_9_port, S(8) => PTMP_9_8_port, S(7) => 
                           PTMP_9_7_port, S(6) => PTMP_9_6_port, S(5) => 
                           PTMP_9_5_port, S(4) => PTMP_9_4_port, S(3) => 
                           PTMP_9_3_port, S(2) => PTMP_9_2_port, S(1) => 
                           PTMP_9_1_port, S(0) => PTMP_9_0_port, Co => n_1290);
   ADDER_11 : RCA_NBIT56 port map( A(55) => n14, A(54) => n14, A(53) => 
                           PTMP_9_53_port, A(52) => PTMP_9_52_port, A(51) => 
                           PTMP_9_51_port, A(50) => PTMP_9_50_port, A(49) => 
                           PTMP_9_49_port, A(48) => PTMP_9_48_port, A(47) => 
                           PTMP_9_47_port, A(46) => PTMP_9_46_port, A(45) => 
                           PTMP_9_45_port, A(44) => PTMP_9_44_port, A(43) => 
                           PTMP_9_43_port, A(42) => PTMP_9_42_port, A(41) => 
                           PTMP_9_41_port, A(40) => PTMP_9_40_port, A(39) => 
                           PTMP_9_39_port, A(38) => PTMP_9_38_port, A(37) => 
                           PTMP_9_37_port, A(36) => PTMP_9_36_port, A(35) => 
                           PTMP_9_35_port, A(34) => PTMP_9_34_port, A(33) => 
                           PTMP_9_33_port, A(32) => PTMP_9_32_port, A(31) => 
                           PTMP_9_31_port, A(30) => PTMP_9_30_port, A(29) => 
                           PTMP_9_29_port, A(28) => PTMP_9_28_port, A(27) => 
                           PTMP_9_27_port, A(26) => PTMP_9_26_port, A(25) => 
                           PTMP_9_25_port, A(24) => PTMP_9_24_port, A(23) => 
                           PTMP_9_23_port, A(22) => PTMP_9_22_port, A(21) => 
                           PTMP_9_21_port, A(20) => PTMP_9_20_port, A(19) => 
                           PTMP_9_19_port, A(18) => PTMP_9_18_port, A(17) => 
                           PTMP_9_17_port, A(16) => PTMP_9_16_port, A(15) => 
                           PTMP_9_15_port, A(14) => PTMP_9_14_port, A(13) => 
                           PTMP_9_13_port, A(12) => PTMP_9_12_port, A(11) => 
                           PTMP_9_11_port, A(10) => PTMP_9_10_port, A(9) => 
                           PTMP_9_9_port, A(8) => PTMP_9_8_port, A(7) => 
                           PTMP_9_7_port, A(6) => PTMP_9_6_port, A(5) => 
                           PTMP_9_5_port, A(4) => PTMP_9_4_port, A(3) => 
                           PTMP_9_3_port, A(2) => PTMP_9_2_port, A(1) => 
                           PTMP_9_1_port, A(0) => PTMP_9_0_port, B(55) => 
                           OTMP_11_55_port, B(54) => OTMP_11_54_port, B(53) => 
                           OTMP_11_53_port, B(52) => OTMP_11_52_port, B(51) => 
                           OTMP_11_51_port, B(50) => OTMP_11_50_port, B(49) => 
                           OTMP_11_49_port, B(48) => OTMP_11_48_port, B(47) => 
                           OTMP_11_47_port, B(46) => OTMP_11_46_port, B(45) => 
                           OTMP_11_45_port, B(44) => OTMP_11_44_port, B(43) => 
                           OTMP_11_43_port, B(42) => OTMP_11_42_port, B(41) => 
                           OTMP_11_41_port, B(40) => OTMP_11_40_port, B(39) => 
                           OTMP_11_39_port, B(38) => OTMP_11_38_port, B(37) => 
                           OTMP_11_37_port, B(36) => OTMP_11_36_port, B(35) => 
                           OTMP_11_35_port, B(34) => OTMP_11_34_port, B(33) => 
                           OTMP_11_33_port, B(32) => OTMP_11_32_port, B(31) => 
                           OTMP_11_31_port, B(30) => OTMP_11_30_port, B(29) => 
                           OTMP_11_29_port, B(28) => OTMP_11_28_port, B(27) => 
                           OTMP_11_27_port, B(26) => OTMP_11_26_port, B(25) => 
                           OTMP_11_25_port, B(24) => OTMP_11_24_port, B(23) => 
                           OTMP_11_23_port, B(22) => OTMP_11_22_port, B(21) => 
                           OTMP_11_21_port, B(20) => OTMP_11_20_port, B(19) => 
                           OTMP_11_19_port, B(18) => OTMP_11_18_port, B(17) => 
                           OTMP_11_17_port, B(16) => OTMP_11_16_port, B(15) => 
                           OTMP_11_15_port, B(14) => OTMP_11_14_port, B(13) => 
                           OTMP_11_13_port, B(12) => OTMP_11_12_port, B(11) => 
                           OTMP_11_11_port, B(10) => OTMP_11_10_port, B(9) => 
                           OTMP_11_9_port, B(8) => OTMP_11_8_port, B(7) => 
                           OTMP_11_7_port, B(6) => OTMP_11_6_port, B(5) => 
                           OTMP_11_5_port, B(4) => OTMP_11_4_port, B(3) => 
                           OTMP_11_3_port, B(2) => OTMP_11_2_port, B(1) => 
                           OTMP_11_1_port, B(0) => OTMP_11_0_port, Ci => 
                           X_Logic0_port, S(55) => PTMP_10_55_port, S(54) => 
                           PTMP_10_54_port, S(53) => PTMP_10_53_port, S(52) => 
                           PTMP_10_52_port, S(51) => PTMP_10_51_port, S(50) => 
                           PTMP_10_50_port, S(49) => PTMP_10_49_port, S(48) => 
                           PTMP_10_48_port, S(47) => PTMP_10_47_port, S(46) => 
                           PTMP_10_46_port, S(45) => PTMP_10_45_port, S(44) => 
                           PTMP_10_44_port, S(43) => PTMP_10_43_port, S(42) => 
                           PTMP_10_42_port, S(41) => PTMP_10_41_port, S(40) => 
                           PTMP_10_40_port, S(39) => PTMP_10_39_port, S(38) => 
                           PTMP_10_38_port, S(37) => PTMP_10_37_port, S(36) => 
                           PTMP_10_36_port, S(35) => PTMP_10_35_port, S(34) => 
                           PTMP_10_34_port, S(33) => PTMP_10_33_port, S(32) => 
                           PTMP_10_32_port, S(31) => PTMP_10_31_port, S(30) => 
                           PTMP_10_30_port, S(29) => PTMP_10_29_port, S(28) => 
                           PTMP_10_28_port, S(27) => PTMP_10_27_port, S(26) => 
                           PTMP_10_26_port, S(25) => PTMP_10_25_port, S(24) => 
                           PTMP_10_24_port, S(23) => PTMP_10_23_port, S(22) => 
                           PTMP_10_22_port, S(21) => PTMP_10_21_port, S(20) => 
                           PTMP_10_20_port, S(19) => PTMP_10_19_port, S(18) => 
                           PTMP_10_18_port, S(17) => PTMP_10_17_port, S(16) => 
                           PTMP_10_16_port, S(15) => PTMP_10_15_port, S(14) => 
                           PTMP_10_14_port, S(13) => PTMP_10_13_port, S(12) => 
                           PTMP_10_12_port, S(11) => PTMP_10_11_port, S(10) => 
                           PTMP_10_10_port, S(9) => PTMP_10_9_port, S(8) => 
                           PTMP_10_8_port, S(7) => PTMP_10_7_port, S(6) => 
                           PTMP_10_6_port, S(5) => PTMP_10_5_port, S(4) => 
                           PTMP_10_4_port, S(3) => PTMP_10_3_port, S(2) => 
                           PTMP_10_2_port, S(1) => PTMP_10_1_port, S(0) => 
                           PTMP_10_0_port, Co => n_1291);
   ADDER_12 : RCA_NBIT58 port map( A(57) => n19, A(56) => n19, A(55) => 
                           PTMP_10_55_port, A(54) => PTMP_10_54_port, A(53) => 
                           PTMP_10_53_port, A(52) => PTMP_10_52_port, A(51) => 
                           PTMP_10_51_port, A(50) => PTMP_10_50_port, A(49) => 
                           PTMP_10_49_port, A(48) => PTMP_10_48_port, A(47) => 
                           PTMP_10_47_port, A(46) => PTMP_10_46_port, A(45) => 
                           PTMP_10_45_port, A(44) => PTMP_10_44_port, A(43) => 
                           PTMP_10_43_port, A(42) => PTMP_10_42_port, A(41) => 
                           PTMP_10_41_port, A(40) => PTMP_10_40_port, A(39) => 
                           PTMP_10_39_port, A(38) => PTMP_10_38_port, A(37) => 
                           PTMP_10_37_port, A(36) => PTMP_10_36_port, A(35) => 
                           PTMP_10_35_port, A(34) => PTMP_10_34_port, A(33) => 
                           PTMP_10_33_port, A(32) => PTMP_10_32_port, A(31) => 
                           PTMP_10_31_port, A(30) => PTMP_10_30_port, A(29) => 
                           PTMP_10_29_port, A(28) => PTMP_10_28_port, A(27) => 
                           PTMP_10_27_port, A(26) => PTMP_10_26_port, A(25) => 
                           PTMP_10_25_port, A(24) => PTMP_10_24_port, A(23) => 
                           PTMP_10_23_port, A(22) => PTMP_10_22_port, A(21) => 
                           PTMP_10_21_port, A(20) => PTMP_10_20_port, A(19) => 
                           PTMP_10_19_port, A(18) => PTMP_10_18_port, A(17) => 
                           PTMP_10_17_port, A(16) => PTMP_10_16_port, A(15) => 
                           PTMP_10_15_port, A(14) => PTMP_10_14_port, A(13) => 
                           PTMP_10_13_port, A(12) => PTMP_10_12_port, A(11) => 
                           PTMP_10_11_port, A(10) => PTMP_10_10_port, A(9) => 
                           PTMP_10_9_port, A(8) => PTMP_10_8_port, A(7) => 
                           PTMP_10_7_port, A(6) => PTMP_10_6_port, A(5) => 
                           PTMP_10_5_port, A(4) => PTMP_10_4_port, A(3) => 
                           PTMP_10_3_port, A(2) => PTMP_10_2_port, A(1) => 
                           PTMP_10_1_port, A(0) => PTMP_10_0_port, B(57) => 
                           OTMP_12_57_port, B(56) => OTMP_12_56_port, B(55) => 
                           OTMP_12_55_port, B(54) => OTMP_12_54_port, B(53) => 
                           OTMP_12_53_port, B(52) => OTMP_12_52_port, B(51) => 
                           OTMP_12_51_port, B(50) => OTMP_12_50_port, B(49) => 
                           OTMP_12_49_port, B(48) => OTMP_12_48_port, B(47) => 
                           OTMP_12_47_port, B(46) => OTMP_12_46_port, B(45) => 
                           OTMP_12_45_port, B(44) => OTMP_12_44_port, B(43) => 
                           OTMP_12_43_port, B(42) => OTMP_12_42_port, B(41) => 
                           OTMP_12_41_port, B(40) => OTMP_12_40_port, B(39) => 
                           OTMP_12_39_port, B(38) => OTMP_12_38_port, B(37) => 
                           OTMP_12_37_port, B(36) => OTMP_12_36_port, B(35) => 
                           OTMP_12_35_port, B(34) => OTMP_12_34_port, B(33) => 
                           OTMP_12_33_port, B(32) => OTMP_12_32_port, B(31) => 
                           OTMP_12_31_port, B(30) => OTMP_12_30_port, B(29) => 
                           OTMP_12_29_port, B(28) => OTMP_12_28_port, B(27) => 
                           OTMP_12_27_port, B(26) => OTMP_12_26_port, B(25) => 
                           OTMP_12_25_port, B(24) => OTMP_12_24_port, B(23) => 
                           OTMP_12_23_port, B(22) => OTMP_12_22_port, B(21) => 
                           OTMP_12_21_port, B(20) => OTMP_12_20_port, B(19) => 
                           OTMP_12_19_port, B(18) => OTMP_12_18_port, B(17) => 
                           OTMP_12_17_port, B(16) => OTMP_12_16_port, B(15) => 
                           OTMP_12_15_port, B(14) => OTMP_12_14_port, B(13) => 
                           OTMP_12_13_port, B(12) => OTMP_12_12_port, B(11) => 
                           OTMP_12_11_port, B(10) => OTMP_12_10_port, B(9) => 
                           OTMP_12_9_port, B(8) => OTMP_12_8_port, B(7) => 
                           OTMP_12_7_port, B(6) => OTMP_12_6_port, B(5) => 
                           OTMP_12_5_port, B(4) => OTMP_12_4_port, B(3) => 
                           OTMP_12_3_port, B(2) => OTMP_12_2_port, B(1) => 
                           OTMP_12_1_port, B(0) => OTMP_12_0_port, Ci => 
                           X_Logic0_port, S(57) => PTMP_11_57_port, S(56) => 
                           PTMP_11_56_port, S(55) => PTMP_11_55_port, S(54) => 
                           PTMP_11_54_port, S(53) => PTMP_11_53_port, S(52) => 
                           PTMP_11_52_port, S(51) => PTMP_11_51_port, S(50) => 
                           PTMP_11_50_port, S(49) => PTMP_11_49_port, S(48) => 
                           PTMP_11_48_port, S(47) => PTMP_11_47_port, S(46) => 
                           PTMP_11_46_port, S(45) => PTMP_11_45_port, S(44) => 
                           PTMP_11_44_port, S(43) => PTMP_11_43_port, S(42) => 
                           PTMP_11_42_port, S(41) => PTMP_11_41_port, S(40) => 
                           PTMP_11_40_port, S(39) => PTMP_11_39_port, S(38) => 
                           PTMP_11_38_port, S(37) => PTMP_11_37_port, S(36) => 
                           PTMP_11_36_port, S(35) => PTMP_11_35_port, S(34) => 
                           PTMP_11_34_port, S(33) => PTMP_11_33_port, S(32) => 
                           PTMP_11_32_port, S(31) => PTMP_11_31_port, S(30) => 
                           PTMP_11_30_port, S(29) => PTMP_11_29_port, S(28) => 
                           PTMP_11_28_port, S(27) => PTMP_11_27_port, S(26) => 
                           PTMP_11_26_port, S(25) => PTMP_11_25_port, S(24) => 
                           PTMP_11_24_port, S(23) => PTMP_11_23_port, S(22) => 
                           PTMP_11_22_port, S(21) => PTMP_11_21_port, S(20) => 
                           PTMP_11_20_port, S(19) => PTMP_11_19_port, S(18) => 
                           PTMP_11_18_port, S(17) => PTMP_11_17_port, S(16) => 
                           PTMP_11_16_port, S(15) => PTMP_11_15_port, S(14) => 
                           PTMP_11_14_port, S(13) => PTMP_11_13_port, S(12) => 
                           PTMP_11_12_port, S(11) => PTMP_11_11_port, S(10) => 
                           PTMP_11_10_port, S(9) => PTMP_11_9_port, S(8) => 
                           PTMP_11_8_port, S(7) => PTMP_11_7_port, S(6) => 
                           PTMP_11_6_port, S(5) => PTMP_11_5_port, S(4) => 
                           PTMP_11_4_port, S(3) => PTMP_11_3_port, S(2) => 
                           PTMP_11_2_port, S(1) => PTMP_11_1_port, S(0) => 
                           PTMP_11_0_port, Co => n_1292);
   ADDER_13 : RCA_NBIT60 port map( A(59) => n13, A(58) => n13, A(57) => 
                           PTMP_11_57_port, A(56) => PTMP_11_56_port, A(55) => 
                           PTMP_11_55_port, A(54) => PTMP_11_54_port, A(53) => 
                           PTMP_11_53_port, A(52) => PTMP_11_52_port, A(51) => 
                           PTMP_11_51_port, A(50) => PTMP_11_50_port, A(49) => 
                           PTMP_11_49_port, A(48) => PTMP_11_48_port, A(47) => 
                           PTMP_11_47_port, A(46) => PTMP_11_46_port, A(45) => 
                           PTMP_11_45_port, A(44) => PTMP_11_44_port, A(43) => 
                           PTMP_11_43_port, A(42) => PTMP_11_42_port, A(41) => 
                           PTMP_11_41_port, A(40) => PTMP_11_40_port, A(39) => 
                           PTMP_11_39_port, A(38) => PTMP_11_38_port, A(37) => 
                           PTMP_11_37_port, A(36) => PTMP_11_36_port, A(35) => 
                           PTMP_11_35_port, A(34) => PTMP_11_34_port, A(33) => 
                           PTMP_11_33_port, A(32) => PTMP_11_32_port, A(31) => 
                           PTMP_11_31_port, A(30) => PTMP_11_30_port, A(29) => 
                           PTMP_11_29_port, A(28) => PTMP_11_28_port, A(27) => 
                           PTMP_11_27_port, A(26) => PTMP_11_26_port, A(25) => 
                           PTMP_11_25_port, A(24) => PTMP_11_24_port, A(23) => 
                           PTMP_11_23_port, A(22) => PTMP_11_22_port, A(21) => 
                           PTMP_11_21_port, A(20) => PTMP_11_20_port, A(19) => 
                           PTMP_11_19_port, A(18) => PTMP_11_18_port, A(17) => 
                           PTMP_11_17_port, A(16) => PTMP_11_16_port, A(15) => 
                           PTMP_11_15_port, A(14) => PTMP_11_14_port, A(13) => 
                           PTMP_11_13_port, A(12) => PTMP_11_12_port, A(11) => 
                           PTMP_11_11_port, A(10) => PTMP_11_10_port, A(9) => 
                           PTMP_11_9_port, A(8) => PTMP_11_8_port, A(7) => 
                           PTMP_11_7_port, A(6) => PTMP_11_6_port, A(5) => 
                           PTMP_11_5_port, A(4) => PTMP_11_4_port, A(3) => 
                           PTMP_11_3_port, A(2) => PTMP_11_2_port, A(1) => 
                           PTMP_11_1_port, A(0) => PTMP_11_0_port, B(59) => 
                           OTMP_13_59_port, B(58) => OTMP_13_58_port, B(57) => 
                           OTMP_13_57_port, B(56) => OTMP_13_56_port, B(55) => 
                           OTMP_13_55_port, B(54) => OTMP_13_54_port, B(53) => 
                           OTMP_13_53_port, B(52) => OTMP_13_52_port, B(51) => 
                           OTMP_13_51_port, B(50) => OTMP_13_50_port, B(49) => 
                           OTMP_13_49_port, B(48) => OTMP_13_48_port, B(47) => 
                           OTMP_13_47_port, B(46) => OTMP_13_46_port, B(45) => 
                           OTMP_13_45_port, B(44) => OTMP_13_44_port, B(43) => 
                           OTMP_13_43_port, B(42) => OTMP_13_42_port, B(41) => 
                           OTMP_13_41_port, B(40) => OTMP_13_40_port, B(39) => 
                           OTMP_13_39_port, B(38) => OTMP_13_38_port, B(37) => 
                           OTMP_13_37_port, B(36) => OTMP_13_36_port, B(35) => 
                           OTMP_13_35_port, B(34) => OTMP_13_34_port, B(33) => 
                           OTMP_13_33_port, B(32) => OTMP_13_32_port, B(31) => 
                           OTMP_13_31_port, B(30) => OTMP_13_30_port, B(29) => 
                           OTMP_13_29_port, B(28) => OTMP_13_28_port, B(27) => 
                           OTMP_13_27_port, B(26) => OTMP_13_26_port, B(25) => 
                           OTMP_13_25_port, B(24) => OTMP_13_24_port, B(23) => 
                           OTMP_13_23_port, B(22) => OTMP_13_22_port, B(21) => 
                           OTMP_13_21_port, B(20) => OTMP_13_20_port, B(19) => 
                           OTMP_13_19_port, B(18) => OTMP_13_18_port, B(17) => 
                           OTMP_13_17_port, B(16) => OTMP_13_16_port, B(15) => 
                           OTMP_13_15_port, B(14) => OTMP_13_14_port, B(13) => 
                           OTMP_13_13_port, B(12) => OTMP_13_12_port, B(11) => 
                           OTMP_13_11_port, B(10) => OTMP_13_10_port, B(9) => 
                           OTMP_13_9_port, B(8) => OTMP_13_8_port, B(7) => 
                           OTMP_13_7_port, B(6) => OTMP_13_6_port, B(5) => 
                           OTMP_13_5_port, B(4) => OTMP_13_4_port, B(3) => 
                           OTMP_13_3_port, B(2) => OTMP_13_2_port, B(1) => 
                           OTMP_13_1_port, B(0) => OTMP_13_0_port, Ci => 
                           X_Logic0_port, S(59) => PTMP_12_59_port, S(58) => 
                           PTMP_12_58_port, S(57) => PTMP_12_57_port, S(56) => 
                           PTMP_12_56_port, S(55) => PTMP_12_55_port, S(54) => 
                           PTMP_12_54_port, S(53) => PTMP_12_53_port, S(52) => 
                           PTMP_12_52_port, S(51) => PTMP_12_51_port, S(50) => 
                           PTMP_12_50_port, S(49) => PTMP_12_49_port, S(48) => 
                           PTMP_12_48_port, S(47) => PTMP_12_47_port, S(46) => 
                           PTMP_12_46_port, S(45) => PTMP_12_45_port, S(44) => 
                           PTMP_12_44_port, S(43) => PTMP_12_43_port, S(42) => 
                           PTMP_12_42_port, S(41) => PTMP_12_41_port, S(40) => 
                           PTMP_12_40_port, S(39) => PTMP_12_39_port, S(38) => 
                           PTMP_12_38_port, S(37) => PTMP_12_37_port, S(36) => 
                           PTMP_12_36_port, S(35) => PTMP_12_35_port, S(34) => 
                           PTMP_12_34_port, S(33) => PTMP_12_33_port, S(32) => 
                           PTMP_12_32_port, S(31) => PTMP_12_31_port, S(30) => 
                           PTMP_12_30_port, S(29) => PTMP_12_29_port, S(28) => 
                           PTMP_12_28_port, S(27) => PTMP_12_27_port, S(26) => 
                           PTMP_12_26_port, S(25) => PTMP_12_25_port, S(24) => 
                           PTMP_12_24_port, S(23) => PTMP_12_23_port, S(22) => 
                           PTMP_12_22_port, S(21) => PTMP_12_21_port, S(20) => 
                           PTMP_12_20_port, S(19) => PTMP_12_19_port, S(18) => 
                           PTMP_12_18_port, S(17) => PTMP_12_17_port, S(16) => 
                           PTMP_12_16_port, S(15) => PTMP_12_15_port, S(14) => 
                           PTMP_12_14_port, S(13) => PTMP_12_13_port, S(12) => 
                           PTMP_12_12_port, S(11) => PTMP_12_11_port, S(10) => 
                           PTMP_12_10_port, S(9) => PTMP_12_9_port, S(8) => 
                           PTMP_12_8_port, S(7) => PTMP_12_7_port, S(6) => 
                           PTMP_12_6_port, S(5) => PTMP_12_5_port, S(4) => 
                           PTMP_12_4_port, S(3) => PTMP_12_3_port, S(2) => 
                           PTMP_12_2_port, S(1) => PTMP_12_1_port, S(0) => 
                           PTMP_12_0_port, Co => n_1293);
   ADDER_14 : RCA_NBIT62 port map( A(61) => n18, A(60) => n18, A(59) => 
                           PTMP_12_59_port, A(58) => PTMP_12_58_port, A(57) => 
                           PTMP_12_57_port, A(56) => PTMP_12_56_port, A(55) => 
                           PTMP_12_55_port, A(54) => PTMP_12_54_port, A(53) => 
                           PTMP_12_53_port, A(52) => PTMP_12_52_port, A(51) => 
                           PTMP_12_51_port, A(50) => PTMP_12_50_port, A(49) => 
                           PTMP_12_49_port, A(48) => PTMP_12_48_port, A(47) => 
                           PTMP_12_47_port, A(46) => PTMP_12_46_port, A(45) => 
                           PTMP_12_45_port, A(44) => PTMP_12_44_port, A(43) => 
                           PTMP_12_43_port, A(42) => PTMP_12_42_port, A(41) => 
                           PTMP_12_41_port, A(40) => PTMP_12_40_port, A(39) => 
                           PTMP_12_39_port, A(38) => PTMP_12_38_port, A(37) => 
                           PTMP_12_37_port, A(36) => PTMP_12_36_port, A(35) => 
                           PTMP_12_35_port, A(34) => PTMP_12_34_port, A(33) => 
                           PTMP_12_33_port, A(32) => PTMP_12_32_port, A(31) => 
                           PTMP_12_31_port, A(30) => PTMP_12_30_port, A(29) => 
                           PTMP_12_29_port, A(28) => PTMP_12_28_port, A(27) => 
                           PTMP_12_27_port, A(26) => PTMP_12_26_port, A(25) => 
                           PTMP_12_25_port, A(24) => PTMP_12_24_port, A(23) => 
                           PTMP_12_23_port, A(22) => PTMP_12_22_port, A(21) => 
                           PTMP_12_21_port, A(20) => PTMP_12_20_port, A(19) => 
                           PTMP_12_19_port, A(18) => PTMP_12_18_port, A(17) => 
                           PTMP_12_17_port, A(16) => PTMP_12_16_port, A(15) => 
                           PTMP_12_15_port, A(14) => PTMP_12_14_port, A(13) => 
                           PTMP_12_13_port, A(12) => PTMP_12_12_port, A(11) => 
                           PTMP_12_11_port, A(10) => PTMP_12_10_port, A(9) => 
                           PTMP_12_9_port, A(8) => PTMP_12_8_port, A(7) => 
                           PTMP_12_7_port, A(6) => PTMP_12_6_port, A(5) => 
                           PTMP_12_5_port, A(4) => PTMP_12_4_port, A(3) => 
                           PTMP_12_3_port, A(2) => PTMP_12_2_port, A(1) => 
                           PTMP_12_1_port, A(0) => PTMP_12_0_port, B(61) => 
                           OTMP_14_61_port, B(60) => OTMP_14_60_port, B(59) => 
                           OTMP_14_59_port, B(58) => OTMP_14_58_port, B(57) => 
                           OTMP_14_57_port, B(56) => OTMP_14_56_port, B(55) => 
                           OTMP_14_55_port, B(54) => OTMP_14_54_port, B(53) => 
                           OTMP_14_53_port, B(52) => OTMP_14_52_port, B(51) => 
                           OTMP_14_51_port, B(50) => OTMP_14_50_port, B(49) => 
                           OTMP_14_49_port, B(48) => OTMP_14_48_port, B(47) => 
                           OTMP_14_47_port, B(46) => OTMP_14_46_port, B(45) => 
                           OTMP_14_45_port, B(44) => OTMP_14_44_port, B(43) => 
                           OTMP_14_43_port, B(42) => OTMP_14_42_port, B(41) => 
                           OTMP_14_41_port, B(40) => OTMP_14_40_port, B(39) => 
                           OTMP_14_39_port, B(38) => OTMP_14_38_port, B(37) => 
                           OTMP_14_37_port, B(36) => OTMP_14_36_port, B(35) => 
                           OTMP_14_35_port, B(34) => OTMP_14_34_port, B(33) => 
                           OTMP_14_33_port, B(32) => OTMP_14_32_port, B(31) => 
                           OTMP_14_31_port, B(30) => OTMP_14_30_port, B(29) => 
                           OTMP_14_29_port, B(28) => OTMP_14_28_port, B(27) => 
                           OTMP_14_27_port, B(26) => OTMP_14_26_port, B(25) => 
                           OTMP_14_25_port, B(24) => OTMP_14_24_port, B(23) => 
                           OTMP_14_23_port, B(22) => OTMP_14_22_port, B(21) => 
                           OTMP_14_21_port, B(20) => OTMP_14_20_port, B(19) => 
                           OTMP_14_19_port, B(18) => OTMP_14_18_port, B(17) => 
                           OTMP_14_17_port, B(16) => OTMP_14_16_port, B(15) => 
                           OTMP_14_15_port, B(14) => OTMP_14_14_port, B(13) => 
                           OTMP_14_13_port, B(12) => OTMP_14_12_port, B(11) => 
                           OTMP_14_11_port, B(10) => OTMP_14_10_port, B(9) => 
                           OTMP_14_9_port, B(8) => OTMP_14_8_port, B(7) => 
                           OTMP_14_7_port, B(6) => OTMP_14_6_port, B(5) => 
                           OTMP_14_5_port, B(4) => OTMP_14_4_port, B(3) => 
                           OTMP_14_3_port, B(2) => OTMP_14_2_port, B(1) => 
                           OTMP_14_1_port, B(0) => OTMP_14_0_port, Ci => 
                           X_Logic0_port, S(61) => PTMP_13_61_port, S(60) => 
                           PTMP_13_60_port, S(59) => PTMP_13_59_port, S(58) => 
                           PTMP_13_58_port, S(57) => PTMP_13_57_port, S(56) => 
                           PTMP_13_56_port, S(55) => PTMP_13_55_port, S(54) => 
                           PTMP_13_54_port, S(53) => PTMP_13_53_port, S(52) => 
                           PTMP_13_52_port, S(51) => PTMP_13_51_port, S(50) => 
                           PTMP_13_50_port, S(49) => PTMP_13_49_port, S(48) => 
                           PTMP_13_48_port, S(47) => PTMP_13_47_port, S(46) => 
                           PTMP_13_46_port, S(45) => PTMP_13_45_port, S(44) => 
                           PTMP_13_44_port, S(43) => PTMP_13_43_port, S(42) => 
                           PTMP_13_42_port, S(41) => PTMP_13_41_port, S(40) => 
                           PTMP_13_40_port, S(39) => PTMP_13_39_port, S(38) => 
                           PTMP_13_38_port, S(37) => PTMP_13_37_port, S(36) => 
                           PTMP_13_36_port, S(35) => PTMP_13_35_port, S(34) => 
                           PTMP_13_34_port, S(33) => PTMP_13_33_port, S(32) => 
                           PTMP_13_32_port, S(31) => PTMP_13_31_port, S(30) => 
                           PTMP_13_30_port, S(29) => PTMP_13_29_port, S(28) => 
                           PTMP_13_28_port, S(27) => PTMP_13_27_port, S(26) => 
                           PTMP_13_26_port, S(25) => PTMP_13_25_port, S(24) => 
                           PTMP_13_24_port, S(23) => PTMP_13_23_port, S(22) => 
                           PTMP_13_22_port, S(21) => PTMP_13_21_port, S(20) => 
                           PTMP_13_20_port, S(19) => PTMP_13_19_port, S(18) => 
                           PTMP_13_18_port, S(17) => PTMP_13_17_port, S(16) => 
                           PTMP_13_16_port, S(15) => PTMP_13_15_port, S(14) => 
                           PTMP_13_14_port, S(13) => PTMP_13_13_port, S(12) => 
                           PTMP_13_12_port, S(11) => PTMP_13_11_port, S(10) => 
                           PTMP_13_10_port, S(9) => PTMP_13_9_port, S(8) => 
                           PTMP_13_8_port, S(7) => PTMP_13_7_port, S(6) => 
                           PTMP_13_6_port, S(5) => PTMP_13_5_port, S(4) => 
                           PTMP_13_4_port, S(3) => PTMP_13_3_port, S(2) => 
                           PTMP_13_2_port, S(1) => PTMP_13_1_port, S(0) => 
                           PTMP_13_0_port, Co => n_1294);
   ADDER_15 : RCA_NBIT64 port map( A(63) => n17, A(62) => n17, A(61) => 
                           PTMP_13_61_port, A(60) => PTMP_13_60_port, A(59) => 
                           PTMP_13_59_port, A(58) => PTMP_13_58_port, A(57) => 
                           PTMP_13_57_port, A(56) => PTMP_13_56_port, A(55) => 
                           PTMP_13_55_port, A(54) => PTMP_13_54_port, A(53) => 
                           PTMP_13_53_port, A(52) => PTMP_13_52_port, A(51) => 
                           PTMP_13_51_port, A(50) => PTMP_13_50_port, A(49) => 
                           PTMP_13_49_port, A(48) => PTMP_13_48_port, A(47) => 
                           PTMP_13_47_port, A(46) => PTMP_13_46_port, A(45) => 
                           PTMP_13_45_port, A(44) => PTMP_13_44_port, A(43) => 
                           PTMP_13_43_port, A(42) => PTMP_13_42_port, A(41) => 
                           PTMP_13_41_port, A(40) => PTMP_13_40_port, A(39) => 
                           PTMP_13_39_port, A(38) => PTMP_13_38_port, A(37) => 
                           PTMP_13_37_port, A(36) => PTMP_13_36_port, A(35) => 
                           PTMP_13_35_port, A(34) => PTMP_13_34_port, A(33) => 
                           PTMP_13_33_port, A(32) => PTMP_13_32_port, A(31) => 
                           PTMP_13_31_port, A(30) => PTMP_13_30_port, A(29) => 
                           PTMP_13_29_port, A(28) => PTMP_13_28_port, A(27) => 
                           PTMP_13_27_port, A(26) => PTMP_13_26_port, A(25) => 
                           PTMP_13_25_port, A(24) => PTMP_13_24_port, A(23) => 
                           PTMP_13_23_port, A(22) => PTMP_13_22_port, A(21) => 
                           PTMP_13_21_port, A(20) => PTMP_13_20_port, A(19) => 
                           PTMP_13_19_port, A(18) => PTMP_13_18_port, A(17) => 
                           PTMP_13_17_port, A(16) => PTMP_13_16_port, A(15) => 
                           PTMP_13_15_port, A(14) => PTMP_13_14_port, A(13) => 
                           PTMP_13_13_port, A(12) => PTMP_13_12_port, A(11) => 
                           PTMP_13_11_port, A(10) => PTMP_13_10_port, A(9) => 
                           PTMP_13_9_port, A(8) => PTMP_13_8_port, A(7) => 
                           PTMP_13_7_port, A(6) => PTMP_13_6_port, A(5) => 
                           PTMP_13_5_port, A(4) => PTMP_13_4_port, A(3) => 
                           PTMP_13_3_port, A(2) => PTMP_13_2_port, A(1) => 
                           PTMP_13_1_port, A(0) => PTMP_13_0_port, B(63) => 
                           OTMP_15_63_port, B(62) => OTMP_15_62_port, B(61) => 
                           OTMP_15_61_port, B(60) => OTMP_15_60_port, B(59) => 
                           OTMP_15_59_port, B(58) => OTMP_15_58_port, B(57) => 
                           OTMP_15_57_port, B(56) => OTMP_15_56_port, B(55) => 
                           OTMP_15_55_port, B(54) => OTMP_15_54_port, B(53) => 
                           OTMP_15_53_port, B(52) => OTMP_15_52_port, B(51) => 
                           OTMP_15_51_port, B(50) => OTMP_15_50_port, B(49) => 
                           OTMP_15_49_port, B(48) => OTMP_15_48_port, B(47) => 
                           OTMP_15_47_port, B(46) => OTMP_15_46_port, B(45) => 
                           OTMP_15_45_port, B(44) => OTMP_15_44_port, B(43) => 
                           OTMP_15_43_port, B(42) => OTMP_15_42_port, B(41) => 
                           OTMP_15_41_port, B(40) => OTMP_15_40_port, B(39) => 
                           OTMP_15_39_port, B(38) => OTMP_15_38_port, B(37) => 
                           OTMP_15_37_port, B(36) => OTMP_15_36_port, B(35) => 
                           OTMP_15_35_port, B(34) => OTMP_15_34_port, B(33) => 
                           OTMP_15_33_port, B(32) => OTMP_15_32_port, B(31) => 
                           OTMP_15_31_port, B(30) => OTMP_15_30_port, B(29) => 
                           OTMP_15_29_port, B(28) => OTMP_15_28_port, B(27) => 
                           OTMP_15_27_port, B(26) => OTMP_15_26_port, B(25) => 
                           OTMP_15_25_port, B(24) => OTMP_15_24_port, B(23) => 
                           OTMP_15_23_port, B(22) => OTMP_15_22_port, B(21) => 
                           OTMP_15_21_port, B(20) => OTMP_15_20_port, B(19) => 
                           OTMP_15_19_port, B(18) => OTMP_15_18_port, B(17) => 
                           OTMP_15_17_port, B(16) => OTMP_15_16_port, B(15) => 
                           OTMP_15_15_port, B(14) => OTMP_15_14_port, B(13) => 
                           OTMP_15_13_port, B(12) => OTMP_15_12_port, B(11) => 
                           OTMP_15_11_port, B(10) => OTMP_15_10_port, B(9) => 
                           OTMP_15_9_port, B(8) => OTMP_15_8_port, B(7) => 
                           OTMP_15_7_port, B(6) => OTMP_15_6_port, B(5) => 
                           OTMP_15_5_port, B(4) => OTMP_15_4_port, B(3) => 
                           OTMP_15_3_port, B(2) => OTMP_15_2_port, B(1) => 
                           OTMP_15_1_port, B(0) => OTMP_15_0_port, Ci => 
                           X_Logic0_port, S(63) => S(63), S(62) => S(62), S(61)
                           => S(61), S(60) => S(60), S(59) => S(59), S(58) => 
                           S(58), S(57) => S(57), S(56) => S(56), S(55) => 
                           S(55), S(54) => S(54), S(53) => S(53), S(52) => 
                           S(52), S(51) => S(51), S(50) => S(50), S(49) => 
                           S(49), S(48) => S(48), S(47) => S(47), S(46) => 
                           S(46), S(45) => S(45), S(44) => S(44), S(43) => 
                           S(43), S(42) => S(42), S(41) => S(41), S(40) => 
                           S(40), S(39) => S(39), S(38) => S(38), S(37) => 
                           S(37), S(36) => S(36), S(35) => S(35), S(34) => 
                           S(34), S(33) => S(33), S(32) => S(32), S(31) => 
                           S(31), S(30) => S(30), S(29) => S(29), S(28) => 
                           S(28), S(27) => S(27), S(26) => S(26), S(25) => 
                           S(25), S(24) => S(24), S(23) => S(23), S(22) => 
                           S(22), S(21) => S(21), S(20) => S(20), S(19) => 
                           S(19), S(18) => S(18), S(17) => S(17), S(16) => 
                           S(16), S(15) => S(15), S(14) => S(14), S(13) => 
                           S(13), S(12) => S(12), S(11) => S(11), S(10) => 
                           S(10), S(9) => S(9), S(8) => S(8), S(7) => S(7), 
                           S(6) => S(6), S(5) => S(5), S(4) => S(4), S(3) => 
                           S(3), S(2) => S(2), S(1) => S(1), S(0) => S(0), Co 
                           => n_1295);
   sub_101 : BOOTHMUL_NBIT32_DW01_sub_0 port map( A(31) => n4, A(30) => n4, 
                           A(29) => n4, A(28) => n4, A(27) => n4, A(26) => n4, 
                           A(25) => n4, A(24) => n4, A(23) => n4, A(22) => n4, 
                           A(21) => n4, A(20) => n4, A(19) => n4, A(18) => n4, 
                           A(17) => n4, A(16) => n4, A(15) => n4, A(14) => n4, 
                           A(13) => n4, A(12) => n4, A(11) => n4, A(10) => n4, 
                           A(9) => n4, A(8) => n4, A(7) => n4, A(6) => n4, A(5)
                           => n4, A(4) => n4, A(3) => n4, A(2) => n4, A(1) => 
                           n4, A(0) => n4, B(31) => A(31), B(30) => A(30), 
                           B(29) => A(29), B(28) => A(28), B(27) => A(27), 
                           B(26) => A(26), B(25) => A(25), B(24) => A(24), 
                           B(23) => A(23), B(22) => A(22), B(21) => A(21), 
                           B(20) => A(20), B(19) => A(19), B(18) => A(18), 
                           B(17) => A(17), B(16) => A(16), B(15) => A(15), 
                           B(14) => A(14), B(13) => A(13), B(12) => A(12), 
                           B(11) => A(11), B(10) => A(10), B(9) => A(9), B(8) 
                           => A(8), B(7) => A(7), B(6) => A(6), B(5) => A(5), 
                           B(4) => A(4), B(3) => A(3), B(2) => A(2), B(1) => 
                           A(1), B(0) => A(0), CI => n5, DIFF(31) => A_n_65, 
                           DIFF(30) => A_n_30_port, DIFF(29) => A_n_29_port, 
                           DIFF(28) => A_n_28_port, DIFF(27) => A_n_27_port, 
                           DIFF(26) => A_n_26_port, DIFF(25) => A_n_25_port, 
                           DIFF(24) => A_n_24_port, DIFF(23) => A_n_23_port, 
                           DIFF(22) => A_n_22_port, DIFF(21) => A_n_21_port, 
                           DIFF(20) => A_n_20_port, DIFF(19) => A_n_19_port, 
                           DIFF(18) => A_n_18_port, DIFF(17) => A_n_17_port, 
                           DIFF(16) => A_n_16_port, DIFF(15) => A_n_15_port, 
                           DIFF(14) => A_n_14_port, DIFF(13) => A_n_13_port, 
                           DIFF(12) => A_n_12_port, DIFF(11) => A_n_11_port, 
                           DIFF(10) => A_n_10_port, DIFF(9) => A_n_9_port, 
                           DIFF(8) => A_n_8_port, DIFF(7) => A_n_7_port, 
                           DIFF(6) => A_n_6_port, DIFF(5) => A_n_5_port, 
                           DIFF(4) => A_n_4_port, DIFF(3) => A_n_3_port, 
                           DIFF(2) => A_n_2_port, DIFF(1) => A_n_1_port, 
                           DIFF(0) => A_n_0_port, CO => n_1296);
   U80 : BUF_X1 port map( A => PTMP_6_47_port, Z => n6);
   U81 : BUF_X1 port map( A => A(0), Z => n9);
   U82 : CLKBUF_X1 port map( A => PTMP_11_57_port, Z => n13);
   U83 : CLKBUF_X1 port map( A => PTMP_9_53_port, Z => n14);
   U84 : CLKBUF_X1 port map( A => PTMP_7_49_port, Z => n10);
   U85 : BUF_X1 port map( A => PTMP_10_55_port, Z => n19);
   U86 : BUF_X1 port map( A => PTMP_12_59_port, Z => n18);
   U87 : BUF_X1 port map( A => PTMP_13_61_port, Z => n17);
   U88 : BUF_X2 port map( A => A(2), Z => n7);
   U89 : BUF_X2 port map( A => A(1), Z => n8);
   U90 : CLKBUF_X1 port map( A => PTMP_3_41_port, Z => n16);
   U91 : BUF_X1 port map( A => PTMP_5_45_port, Z => n15);
   U92 : BUF_X1 port map( A => SHIFT_3_37_port, Z => n21);
   U93 : INV_X1 port map( A => PTMP_4_43_port, ZN => n11);
   U94 : INV_X1 port map( A => n11, ZN => n12);
   U95 : CLKBUF_X1 port map( A => PTMP_0_36_port, Z => n20);

end SYN_BEHAVIOURAL;
