
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_RF_ADDR_W5_DATA_W32 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_RF_ADDR_W5_DATA_W32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_RF_ADDR_W5_DATA_W32.all;

entity RF_ADDR_W5_DATA_W32 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end RF_ADDR_W5_DATA_W32;

architecture SYN_Behavioural of RF_ADDR_W5_DATA_W32 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
      n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, 
      n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, 
      n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, 
      n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, 
      n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, 
      n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, 
      n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, 
      n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, 
      n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, 
      n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, 
      n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, 
      n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, 
      n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, 
      n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, 
      n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, 
      n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, 
      n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, 
      n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, 
      n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, 
      n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, 
      n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, 
      n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, 
      n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, 
      n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, 
      n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, 
      n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, 
      n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, 
      n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, 
      n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, 
      n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, 
      n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, 
      n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, 
      n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, 
      n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, 
      n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, 
      n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, 
      n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, 
      n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, 
      n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, 
      n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, 
      n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, 
      n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, 
      n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, 
      n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, 
      n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, 
      n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, 
      n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, 
      n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, 
      n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, 
      n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, 
      n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, 
      n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, 
      n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, 
      n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, 
      n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, 
      n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, 
      n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, 
      n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, 
      n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, 
      n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, 
      n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, 
      n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, 
      n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, 
      n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, 
      n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, 
      n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, 
      n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, 
      n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, 
      n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, 
      n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, 
      n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, 
      n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, 
      n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, 
      n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, 
      n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, 
      n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, 
      n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, 
      n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, 
      n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, 
      n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, 
      n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, 
      n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, 
      n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, 
      n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, 
      n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, 
      n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, 
      n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, 
      n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, 
      n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, 
      n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, 
      n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, 
      n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, 
      n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, 
      n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, 
      n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, 
      n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, 
      n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, 
      n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, 
      n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, 
      n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, 
      n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, 
      n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, 
      n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, 
      n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, 
      n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, 
      n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, 
      n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, 
      n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n6568, n6569, 
      n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, 
      n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, 
      n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, 
      n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, 
      n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, 
      n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, 
      n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, 
      n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, 
      n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, 
      n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, 
      n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, 
      n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, 
      n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, 
      n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, 
      n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, 
      n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, 
      n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, 
      n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, 
      n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, 
      n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, 
      n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, 
      n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, 
      n8813, n8814, n8815, n8816, n8817, n8820, n8821, n8822, n8823, n8824, 
      n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8835, n8836, 
      n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, 
      n8847, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, 
      n8859, n8860, n8861, n8862, n8865, n8866, n8867, n8868, n8869, n8870, 
      n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8880, n8881, n8882, 
      n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, 
      n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, 
      n8905, n8906, n8907, n8910, n8911, n8912, n8913, n8914, n8915, n8916, 
      n8917, n8918, n8919, n8920, n8921, n8922, n8925, n8926, n8927, n8928, 
      n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8940, 
      n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, 
      n8951, n8952, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, 
      n8963, n8964, n8965, n8966, n8967, n8970, n8971, n8972, n8973, n8974, 
      n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8985, n8986, 
      n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, 
      n8997, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, 
      n9009, n9010, n9011, n9012, n9015, n9016, n9017, n9018, n9019, n9020, 
      n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9030, n9031, n9032, 
      n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, 
      n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, 
      n9055, n9056, n9057, n9060, n9061, n9062, n9063, n9064, n9065, n9066, 
      n9067, n9068, n9069, n9070, n9071, n9072, n9075, n9076, n9077, n9078, 
      n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9090, 
      n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, 
      n9101, n9102, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, 
      n9113, n9114, n9115, n9116, n9117, n9120, n9121, n9122, n9123, n9124, 
      n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9135, n9136, 
      n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, 
      n9147, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, 
      n9159, n9160, n9161, n9162, n9165, n9166, n9167, n9168, n9169, n9170, 
      n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9180, n9181, n9182, 
      n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, 
      n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, 
      n9205, n9206, n9207, n9210, n9211, n9212, n9213, n9214, n9215, n9216, 
      n9217, n9218, n9219, n9220, n9221, n9222, n9225, n9226, n9227, n9228, 
      n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9240, 
      n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, 
      n9251, n9252, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, 
      n9263, n9264, n9265, n9266, n9267, n9270, n9271, n9272, n9273, n9274, 
      n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9285, n9286, 
      n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9923, n9924, 
      n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, 
      n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, 
      n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, 
      n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, 
      n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, 
      n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, 
      n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, 
      n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004
      , n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
      n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022, 
      n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031, 
      n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040, 
      n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, 
      n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058, 
      n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, 
      n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076, 
      n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085, 
      n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094, 
      n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103, 
      n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112, 
      n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121, 
      n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130, 
      n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139, 
      n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148, 
      n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157, 
      n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166, 
      n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175, 
      n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184, 
      n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193, 
      n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202, 
      n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211, 
      n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220, 
      n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229, 
      n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238, 
      n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247, 
      n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256, 
      n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265, 
      n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274, 
      n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283, 
      n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292, 
      n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301, 
      n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310, 
      n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319, 
      n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328, 
      n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337, 
      n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346, 
      n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355, 
      n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364, 
      n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373, 
      n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382, 
      n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391, 
      n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400, 
      n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409, 
      n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418, 
      n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427, 
      n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436, 
      n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445, 
      n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454, 
      n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463, 
      n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472, 
      n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481, 
      n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490, 
      n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499, 
      n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508, 
      n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517, 
      n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526, 
      n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535, 
      n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544, 
      n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553, 
      n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562, 
      n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571, 
      n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580, 
      n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589, 
      n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598, 
      n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607, 
      n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616, 
      n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625, 
      n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634, 
      n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643, 
      n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652, 
      n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661, 
      n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670, 
      n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679, 
      n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688, 
      n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697, 
      n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706, 
      n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715, 
      n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724, 
      n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733, 
      n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742, 
      n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751, 
      n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760, 
      n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769, 
      n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778, 
      n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787, 
      n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796, 
      n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805, 
      n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814, 
      n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823, 
      n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832, 
      n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841, 
      n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850, 
      n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859, 
      n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868, 
      n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877, 
      n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886, 
      n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895, 
      n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904, 
      n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913, 
      n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922, 
      n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931, 
      n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940, 
      n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949, 
      n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958, 
      n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967, 
      n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976, 
      n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985, 
      n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994, 
      n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003, 
      n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012, 
      n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021, 
      n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030, 
      n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039, 
      n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048, 
      n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057, 
      n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066, 
      n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075, 
      n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084, 
      n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093, 
      n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102, 
      n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111, 
      n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120, 
      n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129, 
      n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138, 
      n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147, 
      n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156, 
      n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165, 
      n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174, 
      n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183, 
      n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192, 
      n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201, 
      n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210, 
      n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219, 
      n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228, 
      n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237, 
      n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246, 
      n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255, 
      n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264, 
      n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273, 
      n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282, 
      n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291, 
      n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300, 
      n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309, 
      n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318, 
      n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327, 
      n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336, 
      n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345, 
      n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354, 
      n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363, 
      n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372, 
      n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381, 
      n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390, 
      n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399, 
      n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408, 
      n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417, 
      n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426, 
      n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435, 
      n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444, 
      n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453, 
      n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462, 
      n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471, 
      n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480, 
      n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489, 
      n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498, 
      n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507, 
      n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516, 
      n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525, 
      n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534, 
      n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543, 
      n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552, 
      n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561, 
      n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570, 
      n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579, 
      n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588, 
      n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597, 
      n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606, 
      n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615, 
      n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624, 
      n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633, 
      n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642, 
      n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651, 
      n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660, 
      n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669, 
      n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678, 
      n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687, 
      n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696, 
      n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705, 
      n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714, 
      n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723, 
      n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732, 
      n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741, 
      n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750, 
      n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759, 
      n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768, 
      n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777, 
      n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786, 
      n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795, 
      n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804, 
      n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813, 
      n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822, 
      n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831, 
      n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840, 
      n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849, 
      n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858, 
      n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867, 
      n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876, 
      n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885, 
      n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894, 
      n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903, 
      n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912, 
      n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921, 
      n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930, 
      n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939, 
      n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948, 
      n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957, 
      n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966, 
      n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975, 
      n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984, 
      n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993, 
      n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002, 
      n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011, 
      n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020, 
      n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029, 
      n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038, 
      n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047, 
      n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056, 
      n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065, 
      n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074, 
      n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083, 
      n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092, 
      n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101, 
      n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110, 
      n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119, 
      n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128, 
      n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137, 
      n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146, 
      n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155, 
      n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164, 
      n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173, 
      n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182, 
      n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191, 
      n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200, 
      n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209, 
      n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218, 
      n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227, 
      n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236, 
      n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245, 
      n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254, 
      n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263, 
      n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272, 
      n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281, 
      n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338, 
      n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12520, n12521, 
      n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530, 
      n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539, 
      n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548, 
      n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557, 
      n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566, 
      n12567, n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737, 
      n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746, 
      n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755, 
      n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764, 
      n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773, 
      n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782, 
      n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791, 
      n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800, 
      n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809, 
      n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818, 
      n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827, 
      n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836, 
      n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845, 
      n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854, 
      n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863, 
      n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872, 
      n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881, 
      n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890, 
      n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899, 
      n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908, 
      n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917, 
      n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926, 
      n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935, 
      n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944, 
      n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953, 
      n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962, 
      n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971, 
      n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980, 
      n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989, 
      n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998, 
      n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007, 
      n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016, 
      n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025, 
      n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034, 
      n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043, 
      n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052, 
      n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061, 
      n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070, 
      n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079, 
      n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088, 
      n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097, 
      n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106, 
      n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115, 
      n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124, 
      n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133, 
      n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142, 
      n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151, 
      n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160, 
      n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169, 
      n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178, 
      n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187, 
      n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196, 
      n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205, 
      n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214, 
      n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223, 
      n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232, 
      n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241, 
      n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250, 
      n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259, 
      n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268, 
      n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277, 
      n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286, 
      n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295, 
      n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304, 
      n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313, 
      n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322, 
      n13323, n13324, n_1000, n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, 
      n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, 
      n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, 
      n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, 
      n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, 
      n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, 
      n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, 
      n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, 
      n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, 
      n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, 
      n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, 
      n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, 
      n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, 
      n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, 
      n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, 
      n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, 
      n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, 
      n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, 
      n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, 
      n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, 
      n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, 
      n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, 
      n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, 
      n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, 
      n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, 
      n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, 
      n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, 
      n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, 
      n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, 
      n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, 
      n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, 
      n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, 
      n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, 
      n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, 
      n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, 
      n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, 
      n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, 
      n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, 
      n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, 
      n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, 
      n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, 
      n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, 
      n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, 
      n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, 
      n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, 
      n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, 
      n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, 
      n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, 
      n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, 
      n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1447 : 
      std_logic;

begin
   
   OUT2_reg_31_inst : DFF_X1 port map( D => n2589, CK => CLK, Q => OUT2(31), QN
                           => n8783);
   OUT2_reg_30_inst : DFF_X1 port map( D => n2588, CK => CLK, Q => OUT2(30), QN
                           => n8784);
   OUT2_reg_29_inst : DFF_X1 port map( D => n2587, CK => CLK, Q => OUT2(29), QN
                           => n8785);
   OUT2_reg_28_inst : DFF_X1 port map( D => n2586, CK => CLK, Q => OUT2(28), QN
                           => n8786);
   OUT2_reg_27_inst : DFF_X1 port map( D => n2585, CK => CLK, Q => OUT2(27), QN
                           => n8787);
   OUT2_reg_26_inst : DFF_X1 port map( D => n2584, CK => CLK, Q => OUT2(26), QN
                           => n8788);
   OUT2_reg_25_inst : DFF_X1 port map( D => n2583, CK => CLK, Q => OUT2(25), QN
                           => n8789);
   OUT2_reg_24_inst : DFF_X1 port map( D => n2582, CK => CLK, Q => OUT2(24), QN
                           => n8790);
   OUT2_reg_23_inst : DFF_X1 port map( D => n2581, CK => CLK, Q => OUT2(23), QN
                           => n8791);
   OUT2_reg_22_inst : DFF_X1 port map( D => n2580, CK => CLK, Q => OUT2(22), QN
                           => n8792);
   OUT2_reg_21_inst : DFF_X1 port map( D => n2579, CK => CLK, Q => OUT2(21), QN
                           => n8793);
   OUT2_reg_20_inst : DFF_X1 port map( D => n2578, CK => CLK, Q => OUT2(20), QN
                           => n8794);
   OUT2_reg_19_inst : DFF_X1 port map( D => n2577, CK => CLK, Q => OUT2(19), QN
                           => n8795);
   OUT2_reg_18_inst : DFF_X1 port map( D => n2576, CK => CLK, Q => OUT2(18), QN
                           => n8796);
   OUT2_reg_17_inst : DFF_X1 port map( D => n2575, CK => CLK, Q => OUT2(17), QN
                           => n8797);
   OUT2_reg_16_inst : DFF_X1 port map( D => n2574, CK => CLK, Q => OUT2(16), QN
                           => n8798);
   OUT2_reg_15_inst : DFF_X1 port map( D => n2573, CK => CLK, Q => OUT2(15), QN
                           => n8799);
   OUT2_reg_14_inst : DFF_X1 port map( D => n2572, CK => CLK, Q => OUT2(14), QN
                           => n8800);
   OUT2_reg_13_inst : DFF_X1 port map( D => n2571, CK => CLK, Q => OUT2(13), QN
                           => n8801);
   OUT2_reg_12_inst : DFF_X1 port map( D => n2570, CK => CLK, Q => OUT2(12), QN
                           => n8802);
   OUT2_reg_11_inst : DFF_X1 port map( D => n2569, CK => CLK, Q => OUT2(11), QN
                           => n8803);
   OUT2_reg_10_inst : DFF_X1 port map( D => n2568, CK => CLK, Q => OUT2(10), QN
                           => n8804);
   OUT2_reg_9_inst : DFF_X1 port map( D => n2567, CK => CLK, Q => OUT2(9), QN 
                           => n8805);
   OUT2_reg_8_inst : DFF_X1 port map( D => n2566, CK => CLK, Q => OUT2(8), QN 
                           => n8806);
   OUT2_reg_7_inst : DFF_X1 port map( D => n2565, CK => CLK, Q => OUT2(7), QN 
                           => n8807);
   OUT2_reg_6_inst : DFF_X1 port map( D => n2564, CK => CLK, Q => OUT2(6), QN 
                           => n8808);
   OUT2_reg_5_inst : DFF_X1 port map( D => n2563, CK => CLK, Q => OUT2(5), QN 
                           => n8809);
   OUT2_reg_4_inst : DFF_X1 port map( D => n2562, CK => CLK, Q => OUT2(4), QN 
                           => n8810);
   OUT2_reg_3_inst : DFF_X1 port map( D => n2561, CK => CLK, Q => OUT2(3), QN 
                           => n8811);
   OUT2_reg_2_inst : DFF_X1 port map( D => n2560, CK => CLK, Q => OUT2(2), QN 
                           => n8812);
   OUT2_reg_1_inst : DFF_X1 port map( D => n2559, CK => CLK, Q => OUT2(1), QN 
                           => n8813);
   OUT2_reg_0_inst : DFF_X1 port map( D => n2558, CK => CLK, Q => OUT2(0), QN 
                           => n8814);
   OUT1_reg_31_inst : DFF_X1 port map( D => n2557, CK => CLK, Q => OUT1(31), QN
                           => n8815);
   OUT1_reg_30_inst : DFF_X1 port map( D => n2556, CK => CLK, Q => OUT1(30), QN
                           => n8830);
   OUT1_reg_29_inst : DFF_X1 port map( D => n2555, CK => CLK, Q => OUT1(29), QN
                           => n8845);
   OUT1_reg_28_inst : DFF_X1 port map( D => n2554, CK => CLK, Q => OUT1(28), QN
                           => n8860);
   OUT1_reg_27_inst : DFF_X1 port map( D => n2553, CK => CLK, Q => OUT1(27), QN
                           => n8875);
   OUT1_reg_26_inst : DFF_X1 port map( D => n2552, CK => CLK, Q => OUT1(26), QN
                           => n8890);
   OUT1_reg_25_inst : DFF_X1 port map( D => n2551, CK => CLK, Q => OUT1(25), QN
                           => n8905);
   OUT1_reg_24_inst : DFF_X1 port map( D => n2550, CK => CLK, Q => OUT1(24), QN
                           => n8920);
   OUT1_reg_23_inst : DFF_X1 port map( D => n2549, CK => CLK, Q => OUT1(23), QN
                           => n8935);
   OUT1_reg_22_inst : DFF_X1 port map( D => n2548, CK => CLK, Q => OUT1(22), QN
                           => n8950);
   OUT1_reg_21_inst : DFF_X1 port map( D => n2547, CK => CLK, Q => OUT1(21), QN
                           => n8965);
   OUT1_reg_20_inst : DFF_X1 port map( D => n2546, CK => CLK, Q => OUT1(20), QN
                           => n8980);
   OUT1_reg_19_inst : DFF_X1 port map( D => n2545, CK => CLK, Q => OUT1(19), QN
                           => n8995);
   OUT1_reg_18_inst : DFF_X1 port map( D => n2544, CK => CLK, Q => OUT1(18), QN
                           => n9010);
   OUT1_reg_17_inst : DFF_X1 port map( D => n2543, CK => CLK, Q => OUT1(17), QN
                           => n9025);
   OUT1_reg_16_inst : DFF_X1 port map( D => n2542, CK => CLK, Q => OUT1(16), QN
                           => n9040);
   OUT1_reg_15_inst : DFF_X1 port map( D => n2541, CK => CLK, Q => OUT1(15), QN
                           => n9055);
   OUT1_reg_14_inst : DFF_X1 port map( D => n2540, CK => CLK, Q => OUT1(14), QN
                           => n9070);
   OUT1_reg_13_inst : DFF_X1 port map( D => n2539, CK => CLK, Q => OUT1(13), QN
                           => n9085);
   OUT1_reg_12_inst : DFF_X1 port map( D => n2538, CK => CLK, Q => OUT1(12), QN
                           => n9100);
   OUT1_reg_11_inst : DFF_X1 port map( D => n2537, CK => CLK, Q => OUT1(11), QN
                           => n9115);
   OUT1_reg_10_inst : DFF_X1 port map( D => n2536, CK => CLK, Q => OUT1(10), QN
                           => n9130);
   OUT1_reg_9_inst : DFF_X1 port map( D => n2535, CK => CLK, Q => OUT1(9), QN 
                           => n9145);
   OUT1_reg_8_inst : DFF_X1 port map( D => n2534, CK => CLK, Q => OUT1(8), QN 
                           => n9160);
   OUT1_reg_7_inst : DFF_X1 port map( D => n2533, CK => CLK, Q => OUT1(7), QN 
                           => n9175);
   OUT1_reg_6_inst : DFF_X1 port map( D => n2532, CK => CLK, Q => OUT1(6), QN 
                           => n9190);
   OUT1_reg_5_inst : DFF_X1 port map( D => n2531, CK => CLK, Q => OUT1(5), QN 
                           => n9205);
   OUT1_reg_4_inst : DFF_X1 port map( D => n2530, CK => CLK, Q => OUT1(4), QN 
                           => n9220);
   OUT1_reg_3_inst : DFF_X1 port map( D => n2529, CK => CLK, Q => OUT1(3), QN 
                           => n9235);
   OUT1_reg_2_inst : DFF_X1 port map( D => n2528, CK => CLK, Q => OUT1(2), QN 
                           => n9250);
   OUT1_reg_1_inst : DFF_X1 port map( D => n2527, CK => CLK, Q => OUT1(1), QN 
                           => n9265);
   OUT1_reg_0_inst : DFF_X1 port map( D => n2526, CK => CLK, Q => OUT1(0), QN 
                           => n9280);
   U9447 : NAND3_X1 port map( A1 => n9925, A2 => n9924, A3 => n10948, ZN => 
                           n10932);
   U9448 : NAND3_X1 port map( A1 => n10948, A2 => n9924, A3 => ADD_WR(3), ZN =>
                           n10950);
   U9449 : NAND3_X1 port map( A1 => n10948, A2 => n9925, A3 => ADD_WR(4), ZN =>
                           n10959);
   U9450 : NAND3_X1 port map( A1 => n9927, A2 => n9926, A3 => n9928, ZN => 
                           n10933);
   U9451 : NAND3_X1 port map( A1 => n9927, A2 => n9926, A3 => ADD_WR(0), ZN => 
                           n10935);
   U9452 : NAND3_X1 port map( A1 => n9928, A2 => n9926, A3 => ADD_WR(1), ZN => 
                           n10937);
   U9453 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n9926, A3 => ADD_WR(1), ZN
                           => n10939);
   U9454 : NAND3_X1 port map( A1 => n9928, A2 => n9927, A3 => ADD_WR(2), ZN => 
                           n10941);
   U9455 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n9927, A3 => ADD_WR(2), ZN
                           => n10943);
   U9456 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => n9928, A3 => ADD_WR(2), ZN
                           => n10945);
   U9457 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => n10948, A3 => ADD_WR(4), 
                           ZN => n10968);
   U9458 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), A3 => ADD_WR(2)
                           , ZN => n10947);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n2621, CK => CLK, Q => 
                           n10027, QN => n8828);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n2620, CK => CLK, Q => 
                           n10028, QN => n8843);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n2619, CK => CLK, Q => 
                           n10029, QN => n8858);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n2618, CK => CLK, Q => 
                           n10030, QN => n8873);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n2617, CK => CLK, Q => 
                           n10031, QN => n8888);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n2616, CK => CLK, Q => 
                           n10032, QN => n8903);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n2615, CK => CLK, Q => 
                           n10033, QN => n8918);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n2614, CK => CLK, Q => 
                           n10034, QN => n8933);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n2613, CK => CLK, Q => 
                           n10035, QN => n8948);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n2612, CK => CLK, Q => 
                           n10036, QN => n8963);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n2611, CK => CLK, Q => 
                           n10037, QN => n8978);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n2610, CK => CLK, Q => 
                           n10038, QN => n8993);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n2609, CK => CLK, Q => 
                           n10039, QN => n9008);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n2608, CK => CLK, Q => 
                           n10040, QN => n9023);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n2607, CK => CLK, Q => 
                           n10041, QN => n9038);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n2606, CK => CLK, Q => 
                           n10042, QN => n9053);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n2605, CK => CLK, Q => 
                           n10043, QN => n9068);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n2604, CK => CLK, Q => 
                           n10044, QN => n9083);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n2603, CK => CLK, Q => 
                           n10045, QN => n9098);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n2602, CK => CLK, Q => 
                           n10046, QN => n9113);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n2601, CK => CLK, Q => 
                           n10047, QN => n9128);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n2600, CK => CLK, Q => 
                           n10048, QN => n9143);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n2599, CK => CLK, Q => 
                           n10049, QN => n9158);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n2598, CK => CLK, Q => 
                           n10050, QN => n9173);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n2597, CK => CLK, Q => 
                           n10051, QN => n9188);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n2596, CK => CLK, Q => 
                           n10052, QN => n9203);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n2595, CK => CLK, Q => 
                           n10053, QN => n9218);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n2594, CK => CLK, Q => 
                           n10054, QN => n9233);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n2593, CK => CLK, Q => 
                           n10055, QN => n9248);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n2592, CK => CLK, Q => 
                           n10056, QN => n9263);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n2591, CK => CLK, Q => 
                           n10057, QN => n9278);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n2590, CK => CLK, Q => 
                           n10058, QN => n9293);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n2653, CK => CLK, Q => 
                           n10059, QN => n8829);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n2652, CK => CLK, Q => 
                           n10060, QN => n8844);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n2651, CK => CLK, Q => 
                           n10061, QN => n8859);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n2650, CK => CLK, Q => 
                           n10062, QN => n8874);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n2649, CK => CLK, Q => 
                           n10063, QN => n8889);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n2648, CK => CLK, Q => 
                           n10064, QN => n8904);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n2647, CK => CLK, Q => 
                           n10065, QN => n8919);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n2646, CK => CLK, Q => 
                           n10066, QN => n8934);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n2749, CK => CLK, Q => 
                           n10067, QN => n8826);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n2748, CK => CLK, Q => 
                           n10068, QN => n8841);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n2747, CK => CLK, Q => 
                           n10069, QN => n8856);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n2746, CK => CLK, Q => 
                           n10070, QN => n8871);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n2745, CK => CLK, Q => 
                           n10071, QN => n8886);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n2744, CK => CLK, Q => 
                           n10072, QN => n8901);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n2743, CK => CLK, Q => 
                           n10073, QN => n8916);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n2742, CK => CLK, Q => 
                           n10074, QN => n8931);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n2781, CK => CLK, Q => 
                           n10075, QN => n8827);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n2780, CK => CLK, Q => 
                           n10076, QN => n8842);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n2779, CK => CLK, Q => 
                           n10077, QN => n8857);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n2778, CK => CLK, Q => 
                           n10078, QN => n8872);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n2777, CK => CLK, Q => 
                           n10079, QN => n8887);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n2776, CK => CLK, Q => 
                           n10080, QN => n8902);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n2775, CK => CLK, Q => 
                           n10081, QN => n8917);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n2774, CK => CLK, Q => 
                           n10082, QN => n8932);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n2941, CK => CLK, Q => 
                           n10083, QN => n8824);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n2940, CK => CLK, Q => 
                           n10084, QN => n8839);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n2939, CK => CLK, Q => 
                           n10085, QN => n8854);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n2938, CK => CLK, Q => 
                           n10086, QN => n8869);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n2937, CK => CLK, Q => 
                           n10087, QN => n8884);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n2936, CK => CLK, Q => 
                           n10088, QN => n8899);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n2935, CK => CLK, Q => 
                           n10089, QN => n8914);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n2934, CK => CLK, Q => 
                           n10090, QN => n8929);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n2973, CK => CLK, Q => 
                           n10091, QN => n8825);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n2972, CK => CLK, Q => 
                           n10092, QN => n8840);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n2971, CK => CLK, Q => 
                           n10093, QN => n8855);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n2970, CK => CLK, Q => 
                           n10094, QN => n8870);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n2969, CK => CLK, Q => 
                           n10095, QN => n8885);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n2968, CK => CLK, Q => 
                           n10096, QN => n8900);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n2967, CK => CLK, Q => 
                           n10097, QN => n8915);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n2966, CK => CLK, Q => 
                           n10098, QN => n8930);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n3197, CK => CLK, Q => 
                           n10099, QN => n8820);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n3196, CK => CLK, Q => 
                           n10100, QN => n8835);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n3195, CK => CLK, Q => 
                           n10101, QN => n8850);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n3194, CK => CLK, Q => 
                           n10102, QN => n8865);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n3193, CK => CLK, Q => 
                           n10103, QN => n8880);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n3192, CK => CLK, Q => 
                           n10104, QN => n8895);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n3191, CK => CLK, Q => 
                           n10105, QN => n8910);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n3190, CK => CLK, Q => 
                           n10106, QN => n8925);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n3229, CK => CLK, Q => 
                           n10107, QN => n8821);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n3228, CK => CLK, Q => 
                           n10108, QN => n8836);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n3227, CK => CLK, Q => 
                           n10109, QN => n8851);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n3226, CK => CLK, Q => 
                           n10110, QN => n8866);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n3225, CK => CLK, Q => 
                           n10111, QN => n8881);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n3224, CK => CLK, Q => 
                           n10112, QN => n8896);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n3223, CK => CLK, Q => 
                           n10113, QN => n8911);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n3222, CK => CLK, Q => 
                           n10114, QN => n8926);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n3453, CK => CLK, Q => 
                           n10835, QN => n6600);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n3452, CK => CLK, Q => 
                           n10836, QN => n6601);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n3451, CK => CLK, Q => 
                           n10837, QN => n6602);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n3450, CK => CLK, Q => 
                           n10838, QN => n6603);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n3449, CK => CLK, Q => 
                           n10839, QN => n6604);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n3448, CK => CLK, Q => 
                           n10840, QN => n6605);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n3447, CK => CLK, Q => 
                           n10841, QN => n6606);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n3446, CK => CLK, Q => 
                           n10842, QN => n6607);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n3485, CK => CLK, Q => 
                           n10867, QN => n6568);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n3484, CK => CLK, Q => 
                           n10868, QN => n6569);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n3483, CK => CLK, Q => 
                           n10869, QN => n6570);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n3482, CK => CLK, Q => 
                           n10870, QN => n6571);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n3481, CK => CLK, Q => 
                           n10871, QN => n6572);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n3480, CK => CLK, Q => 
                           n10872, QN => n6573);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n3479, CK => CLK, Q => 
                           n10873, QN => n6574);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n3478, CK => CLK, Q => 
                           n10874, QN => n6575);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n3517, CK => CLK, Q => 
                           n10115, QN => n8817);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n3516, CK => CLK, Q => 
                           n10116, QN => n8832);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n3515, CK => CLK, Q => 
                           n10117, QN => n8847);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n3514, CK => CLK, Q => 
                           n10118, QN => n8862);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n3513, CK => CLK, Q => 
                           n10119, QN => n8877);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n3512, CK => CLK, Q => 
                           n10120, QN => n8892);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n3511, CK => CLK, Q => 
                           n10121, QN => n8907);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n3510, CK => CLK, Q => 
                           n10122, QN => n8922);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n3549, CK => CLK, Q => 
                           n10123, QN => n8816);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n3548, CK => CLK, Q => 
                           n10124, QN => n8831);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n3547, CK => CLK, Q => 
                           n10125, QN => n8846);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n3546, CK => CLK, Q => 
                           n10126, QN => n8861);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n3545, CK => CLK, Q => 
                           n10127, QN => n8876);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n3544, CK => CLK, Q => 
                           n10128, QN => n8891);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n3543, CK => CLK, Q => 
                           n10129, QN => n8906);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n3542, CK => CLK, Q => 
                           n10130, QN => n8921);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n2645, CK => CLK, Q => 
                           n10131, QN => n8949);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n2644, CK => CLK, Q => 
                           n10132, QN => n8964);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n2643, CK => CLK, Q => 
                           n10133, QN => n8979);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n2642, CK => CLK, Q => 
                           n10134, QN => n8994);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n2641, CK => CLK, Q => 
                           n10135, QN => n9009);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n2640, CK => CLK, Q => 
                           n10136, QN => n9024);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n2639, CK => CLK, Q => 
                           n10137, QN => n9039);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n2638, CK => CLK, Q => 
                           n10138, QN => n9054);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n2637, CK => CLK, Q => 
                           n10139, QN => n9069);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n2636, CK => CLK, Q => 
                           n10140, QN => n9084);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n2635, CK => CLK, Q => 
                           n10141, QN => n9099);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n2634, CK => CLK, Q => 
                           n10142, QN => n9114);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n2633, CK => CLK, Q => 
                           n10143, QN => n9129);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n2632, CK => CLK, Q => 
                           n10144, QN => n9144);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n2631, CK => CLK, Q => 
                           n10145, QN => n9159);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n2630, CK => CLK, Q => 
                           n10146, QN => n9174);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n2629, CK => CLK, Q => 
                           n10147, QN => n9189);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n2628, CK => CLK, Q => 
                           n10148, QN => n9204);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n2627, CK => CLK, Q => 
                           n10149, QN => n9219);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n2626, CK => CLK, Q => 
                           n10150, QN => n9234);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n2625, CK => CLK, Q => 
                           n10151, QN => n9249);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n2624, CK => CLK, Q => 
                           n10152, QN => n9264);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n2623, CK => CLK, Q => 
                           n10153, QN => n9279);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n2622, CK => CLK, Q => 
                           n10154, QN => n9294);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n2741, CK => CLK, Q => 
                           n10155, QN => n8946);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n2740, CK => CLK, Q => 
                           n10156, QN => n8961);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n2739, CK => CLK, Q => 
                           n10157, QN => n8976);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n2738, CK => CLK, Q => 
                           n10158, QN => n8991);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n2737, CK => CLK, Q => 
                           n10159, QN => n9006);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n2736, CK => CLK, Q => 
                           n10160, QN => n9021);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n2735, CK => CLK, Q => 
                           n10161, QN => n9036);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n2734, CK => CLK, Q => 
                           n10162, QN => n9051);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n2733, CK => CLK, Q => 
                           n10163, QN => n9066);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n2732, CK => CLK, Q => 
                           n10164, QN => n9081);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n2731, CK => CLK, Q => 
                           n10165, QN => n9096);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n2730, CK => CLK, Q => 
                           n10166, QN => n9111);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n2729, CK => CLK, Q => 
                           n10167, QN => n9126);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n2728, CK => CLK, Q => 
                           n10168, QN => n9141);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n2727, CK => CLK, Q => 
                           n10169, QN => n9156);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n2726, CK => CLK, Q => 
                           n10170, QN => n9171);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n2725, CK => CLK, Q => 
                           n10171, QN => n9186);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n2724, CK => CLK, Q => 
                           n10172, QN => n9201);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n2723, CK => CLK, Q => 
                           n10173, QN => n9216);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n2722, CK => CLK, Q => 
                           n10174, QN => n9231);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n2721, CK => CLK, Q => 
                           n10175, QN => n9246);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n2720, CK => CLK, Q => 
                           n10176, QN => n9261);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n2719, CK => CLK, Q => 
                           n10177, QN => n9276);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n2718, CK => CLK, Q => 
                           n10178, QN => n9291);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n2773, CK => CLK, Q => 
                           n10179, QN => n8947);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n2772, CK => CLK, Q => 
                           n10180, QN => n8962);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n2771, CK => CLK, Q => 
                           n10181, QN => n8977);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n2770, CK => CLK, Q => 
                           n10182, QN => n8992);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n2769, CK => CLK, Q => 
                           n10183, QN => n9007);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n2768, CK => CLK, Q => 
                           n10184, QN => n9022);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n2767, CK => CLK, Q => 
                           n10185, QN => n9037);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n2766, CK => CLK, Q => 
                           n10186, QN => n9052);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n2765, CK => CLK, Q => 
                           n10187, QN => n9067);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n2764, CK => CLK, Q => 
                           n10188, QN => n9082);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n2763, CK => CLK, Q => 
                           n10189, QN => n9097);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n2762, CK => CLK, Q => 
                           n10190, QN => n9112);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n2761, CK => CLK, Q => 
                           n10191, QN => n9127);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n2760, CK => CLK, Q => 
                           n10192, QN => n9142);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n2759, CK => CLK, Q => 
                           n10193, QN => n9157);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n2758, CK => CLK, Q => 
                           n10194, QN => n9172);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n2757, CK => CLK, Q => 
                           n10195, QN => n9187);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n2756, CK => CLK, Q => 
                           n10196, QN => n9202);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n2755, CK => CLK, Q => 
                           n10197, QN => n9217);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n2754, CK => CLK, Q => 
                           n10198, QN => n9232);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n2753, CK => CLK, Q => 
                           n10199, QN => n9247);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n2752, CK => CLK, Q => 
                           n10200, QN => n9262);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n2751, CK => CLK, Q => 
                           n10201, QN => n9277);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n2750, CK => CLK, Q => 
                           n10202, QN => n9292);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n2933, CK => CLK, Q => 
                           n10203, QN => n8944);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n2932, CK => CLK, Q => 
                           n10204, QN => n8959);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n2931, CK => CLK, Q => 
                           n10205, QN => n8974);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n2930, CK => CLK, Q => 
                           n10206, QN => n8989);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n2929, CK => CLK, Q => 
                           n10207, QN => n9004);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n2928, CK => CLK, Q => 
                           n10208, QN => n9019);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n2927, CK => CLK, Q => 
                           n10209, QN => n9034);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n2926, CK => CLK, Q => 
                           n10210, QN => n9049);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n2925, CK => CLK, Q => 
                           n10211, QN => n9064);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n2924, CK => CLK, Q => 
                           n10212, QN => n9079);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n2923, CK => CLK, Q => 
                           n10213, QN => n9094);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n2922, CK => CLK, Q => 
                           n10214, QN => n9109);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n2921, CK => CLK, Q => 
                           n10215, QN => n9124);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n2920, CK => CLK, Q => 
                           n10216, QN => n9139);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n2919, CK => CLK, Q => 
                           n10217, QN => n9154);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n2918, CK => CLK, Q => 
                           n10218, QN => n9169);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n2917, CK => CLK, Q => 
                           n10219, QN => n9184);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n2916, CK => CLK, Q => 
                           n10220, QN => n9199);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n2915, CK => CLK, Q => 
                           n10221, QN => n9214);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n2914, CK => CLK, Q => 
                           n10222, QN => n9229);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n2913, CK => CLK, Q => 
                           n10223, QN => n9244);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n2912, CK => CLK, Q => 
                           n10224, QN => n9259);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n2911, CK => CLK, Q => 
                           n10225, QN => n9274);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n2910, CK => CLK, Q => 
                           n10226, QN => n9289);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n2965, CK => CLK, Q => 
                           n10227, QN => n8945);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n2964, CK => CLK, Q => 
                           n10228, QN => n8960);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n2963, CK => CLK, Q => 
                           n10229, QN => n8975);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n2962, CK => CLK, Q => 
                           n10230, QN => n8990);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n2961, CK => CLK, Q => 
                           n10231, QN => n9005);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n2960, CK => CLK, Q => 
                           n10232, QN => n9020);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n2959, CK => CLK, Q => 
                           n10233, QN => n9035);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n2958, CK => CLK, Q => 
                           n10234, QN => n9050);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n2957, CK => CLK, Q => 
                           n10235, QN => n9065);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n2956, CK => CLK, Q => 
                           n10236, QN => n9080);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n2955, CK => CLK, Q => 
                           n10237, QN => n9095);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n2954, CK => CLK, Q => 
                           n10238, QN => n9110);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n2953, CK => CLK, Q => 
                           n10239, QN => n9125);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n2952, CK => CLK, Q => 
                           n10240, QN => n9140);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n2951, CK => CLK, Q => 
                           n10241, QN => n9155);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n2950, CK => CLK, Q => 
                           n10242, QN => n9170);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n2949, CK => CLK, Q => 
                           n10243, QN => n9185);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n2948, CK => CLK, Q => 
                           n10244, QN => n9200);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n2947, CK => CLK, Q => 
                           n10245, QN => n9215);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n2946, CK => CLK, Q => 
                           n10246, QN => n9230);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n2945, CK => CLK, Q => 
                           n10247, QN => n9245);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n2944, CK => CLK, Q => 
                           n10248, QN => n9260);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n2943, CK => CLK, Q => 
                           n10249, QN => n9275);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n2942, CK => CLK, Q => 
                           n10250, QN => n9290);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n3189, CK => CLK, Q => 
                           n10251, QN => n8940);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n3188, CK => CLK, Q => 
                           n10252, QN => n8955);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n3187, CK => CLK, Q => 
                           n10253, QN => n8970);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n3186, CK => CLK, Q => 
                           n10254, QN => n8985);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n3185, CK => CLK, Q => 
                           n10255, QN => n9000);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n3184, CK => CLK, Q => 
                           n10256, QN => n9015);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n3183, CK => CLK, Q => 
                           n10257, QN => n9030);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n3182, CK => CLK, Q => 
                           n10258, QN => n9045);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n3181, CK => CLK, Q => 
                           n10259, QN => n9060);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n3180, CK => CLK, Q => 
                           n10260, QN => n9075);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n3179, CK => CLK, Q => 
                           n10261, QN => n9090);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n3178, CK => CLK, Q => 
                           n10262, QN => n9105);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n3177, CK => CLK, Q => 
                           n10263, QN => n9120);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n3176, CK => CLK, Q => 
                           n10264, QN => n9135);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n3175, CK => CLK, Q => 
                           n10265, QN => n9150);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n3174, CK => CLK, Q => 
                           n10266, QN => n9165);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n3173, CK => CLK, Q => 
                           n10267, QN => n9180);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n3172, CK => CLK, Q => 
                           n10268, QN => n9195);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n3171, CK => CLK, Q => 
                           n10269, QN => n9210);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n3170, CK => CLK, Q => 
                           n10270, QN => n9225);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n3169, CK => CLK, Q => 
                           n10271, QN => n9240);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n3168, CK => CLK, Q => 
                           n10272, QN => n9255);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n3167, CK => CLK, Q => 
                           n10273, QN => n9270);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n3166, CK => CLK, Q => 
                           n10274, QN => n9285);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n3221, CK => CLK, Q => 
                           n10275, QN => n8941);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n3220, CK => CLK, Q => 
                           n10276, QN => n8956);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n3219, CK => CLK, Q => 
                           n10277, QN => n8971);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n3218, CK => CLK, Q => 
                           n10278, QN => n8986);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n3217, CK => CLK, Q => 
                           n10279, QN => n9001);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n3216, CK => CLK, Q => 
                           n10280, QN => n9016);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n3215, CK => CLK, Q => 
                           n10281, QN => n9031);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n3214, CK => CLK, Q => 
                           n10282, QN => n9046);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n3213, CK => CLK, Q => 
                           n10283, QN => n9061);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n3212, CK => CLK, Q => 
                           n10284, QN => n9076);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n3211, CK => CLK, Q => 
                           n10285, QN => n9091);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n3210, CK => CLK, Q => 
                           n10286, QN => n9106);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n3209, CK => CLK, Q => 
                           n10287, QN => n9121);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n3208, CK => CLK, Q => 
                           n10288, QN => n9136);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n3207, CK => CLK, Q => 
                           n10289, QN => n9151);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n3206, CK => CLK, Q => 
                           n10290, QN => n9166);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n3205, CK => CLK, Q => 
                           n10291, QN => n9181);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n3204, CK => CLK, Q => 
                           n10292, QN => n9196);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n3203, CK => CLK, Q => 
                           n10293, QN => n9211);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n3202, CK => CLK, Q => 
                           n10294, QN => n9226);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n3201, CK => CLK, Q => 
                           n10295, QN => n9241);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n3200, CK => CLK, Q => 
                           n10296, QN => n9256);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n3199, CK => CLK, Q => 
                           n10297, QN => n9271);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n3198, CK => CLK, Q => 
                           n10298, QN => n9286);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n3445, CK => CLK, Q => 
                           n10843, QN => n6608);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n3444, CK => CLK, Q => 
                           n10844, QN => n6609);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n3443, CK => CLK, Q => 
                           n10845, QN => n6610);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n3442, CK => CLK, Q => 
                           n10846, QN => n6611);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n3441, CK => CLK, Q => 
                           n10847, QN => n6612);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n3440, CK => CLK, Q => 
                           n10848, QN => n6613);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n3439, CK => CLK, Q => 
                           n10849, QN => n6614);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n3438, CK => CLK, Q => 
                           n10850, QN => n6615);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n3437, CK => CLK, Q => 
                           n10851, QN => n6616);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n3436, CK => CLK, Q => 
                           n10852, QN => n6617);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n3435, CK => CLK, Q => 
                           n10853, QN => n6618);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n3434, CK => CLK, Q => 
                           n10854, QN => n6619);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n3433, CK => CLK, Q => 
                           n10855, QN => n6620);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n3432, CK => CLK, Q => 
                           n10856, QN => n6621);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n3431, CK => CLK, Q => n10857
                           , QN => n6622);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n3430, CK => CLK, Q => n10858
                           , QN => n6623);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n3429, CK => CLK, Q => n10859
                           , QN => n6624);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n3428, CK => CLK, Q => n10860
                           , QN => n6625);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n3427, CK => CLK, Q => n10861
                           , QN => n6626);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n3426, CK => CLK, Q => n10862
                           , QN => n6627);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n3425, CK => CLK, Q => n10863
                           , QN => n6628);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n3424, CK => CLK, Q => n10864
                           , QN => n6629);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n3423, CK => CLK, Q => n10865
                           , QN => n6630);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n3422, CK => CLK, Q => n10866
                           , QN => n6631);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n3477, CK => CLK, Q => 
                           n10875, QN => n6576);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n3476, CK => CLK, Q => 
                           n10876, QN => n6577);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n3475, CK => CLK, Q => 
                           n10877, QN => n6578);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n3474, CK => CLK, Q => 
                           n10878, QN => n6579);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n3473, CK => CLK, Q => 
                           n10879, QN => n6580);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n3472, CK => CLK, Q => 
                           n10880, QN => n6581);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n3471, CK => CLK, Q => 
                           n10881, QN => n6582);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n3470, CK => CLK, Q => 
                           n10882, QN => n6583);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n3469, CK => CLK, Q => 
                           n10883, QN => n6584);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n3468, CK => CLK, Q => 
                           n10884, QN => n6585);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n3467, CK => CLK, Q => 
                           n10885, QN => n6586);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n3466, CK => CLK, Q => 
                           n10886, QN => n6587);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n3465, CK => CLK, Q => 
                           n10887, QN => n6588);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n3464, CK => CLK, Q => 
                           n10888, QN => n6589);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n3463, CK => CLK, Q => n10889
                           , QN => n6590);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n3462, CK => CLK, Q => n10890
                           , QN => n6591);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n3461, CK => CLK, Q => n10891
                           , QN => n6592);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n3460, CK => CLK, Q => n10892
                           , QN => n6593);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n3459, CK => CLK, Q => n10893
                           , QN => n6594);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n3458, CK => CLK, Q => n10894
                           , QN => n6595);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n3457, CK => CLK, Q => n10895
                           , QN => n6596);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n3456, CK => CLK, Q => n10896
                           , QN => n6597);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n3455, CK => CLK, Q => n10897
                           , QN => n6598);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n3454, CK => CLK, Q => n10898
                           , QN => n6599);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n3509, CK => CLK, Q => 
                           n10299, QN => n8937);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n3508, CK => CLK, Q => 
                           n10300, QN => n8952);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n3507, CK => CLK, Q => 
                           n10301, QN => n8967);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n3506, CK => CLK, Q => 
                           n10302, QN => n8982);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n3505, CK => CLK, Q => 
                           n10303, QN => n8997);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n3504, CK => CLK, Q => 
                           n10304, QN => n9012);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n3503, CK => CLK, Q => 
                           n10305, QN => n9027);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n3502, CK => CLK, Q => 
                           n10306, QN => n9042);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n3501, CK => CLK, Q => 
                           n10307, QN => n9057);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n3500, CK => CLK, Q => 
                           n10308, QN => n9072);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n3499, CK => CLK, Q => 
                           n10309, QN => n9087);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n3498, CK => CLK, Q => 
                           n10310, QN => n9102);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n3497, CK => CLK, Q => 
                           n10311, QN => n9117);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n3496, CK => CLK, Q => 
                           n10312, QN => n9132);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n3495, CK => CLK, Q => n10313
                           , QN => n9147);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n3494, CK => CLK, Q => n10314
                           , QN => n9162);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n3493, CK => CLK, Q => n10315
                           , QN => n9177);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n3492, CK => CLK, Q => n10316
                           , QN => n9192);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n3491, CK => CLK, Q => n10317
                           , QN => n9207);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n3490, CK => CLK, Q => n10318
                           , QN => n9222);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n3489, CK => CLK, Q => n10319
                           , QN => n9237);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n3488, CK => CLK, Q => n10320
                           , QN => n9252);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n3487, CK => CLK, Q => n10321
                           , QN => n9267);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n3486, CK => CLK, Q => n10322
                           , QN => n9282);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n3541, CK => CLK, Q => 
                           n10323, QN => n8936);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n3540, CK => CLK, Q => 
                           n10324, QN => n8951);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n3539, CK => CLK, Q => 
                           n10325, QN => n8966);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n3538, CK => CLK, Q => 
                           n10326, QN => n8981);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n3537, CK => CLK, Q => 
                           n10327, QN => n8996);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n3536, CK => CLK, Q => 
                           n10328, QN => n9011);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n3535, CK => CLK, Q => 
                           n10329, QN => n9026);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n3534, CK => CLK, Q => 
                           n10330, QN => n9041);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n3533, CK => CLK, Q => 
                           n10331, QN => n9056);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n3532, CK => CLK, Q => 
                           n10332, QN => n9071);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n3531, CK => CLK, Q => 
                           n10333, QN => n9086);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n3530, CK => CLK, Q => 
                           n10334, QN => n9101);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n3529, CK => CLK, Q => 
                           n10335, QN => n9116);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n3528, CK => CLK, Q => 
                           n10336, QN => n9131);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n3527, CK => CLK, Q => n10337
                           , QN => n9146);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n3526, CK => CLK, Q => n10338
                           , QN => n9161);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n3525, CK => CLK, Q => n10339
                           , QN => n9176);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n3524, CK => CLK, Q => n10340
                           , QN => n9191);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n3523, CK => CLK, Q => n10341
                           , QN => n9206);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n3522, CK => CLK, Q => n10342
                           , QN => n9221);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n3521, CK => CLK, Q => n10343
                           , QN => n9236);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n3520, CK => CLK, Q => n10344
                           , QN => n9251);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n3519, CK => CLK, Q => n10345
                           , QN => n9266);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n3518, CK => CLK, Q => n10346
                           , QN => n9281);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n3101, CK => CLK, Q => 
                           n_1000, QN => n8823);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n3100, CK => CLK, Q => 
                           n_1001, QN => n8838);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n3099, CK => CLK, Q => 
                           n_1002, QN => n8853);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n3098, CK => CLK, Q => 
                           n_1003, QN => n8868);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n3097, CK => CLK, Q => 
                           n_1004, QN => n8883);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n3096, CK => CLK, Q => 
                           n_1005, QN => n8898);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n3095, CK => CLK, Q => 
                           n_1006, QN => n8913);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n3094, CK => CLK, Q => 
                           n_1007, QN => n8928);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n3069, CK => CLK, Q => 
                           n_1008, QN => n8822);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n3068, CK => CLK, Q => 
                           n_1009, QN => n8837);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n3067, CK => CLK, Q => 
                           n_1010, QN => n8852);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n3066, CK => CLK, Q => 
                           n_1011, QN => n8867);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n3065, CK => CLK, Q => 
                           n_1012, QN => n8882);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n3064, CK => CLK, Q => 
                           n_1013, QN => n8897);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n3063, CK => CLK, Q => 
                           n_1014, QN => n8912);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n3062, CK => CLK, Q => 
                           n_1015, QN => n8927);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n3293, CK => CLK, Q => 
                           n10771, QN => n6696);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n3292, CK => CLK, Q => 
                           n10772, QN => n6697);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n3291, CK => CLK, Q => 
                           n10773, QN => n6698);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n3290, CK => CLK, Q => 
                           n10774, QN => n6699);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n3289, CK => CLK, Q => 
                           n10775, QN => n6700);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n3288, CK => CLK, Q => 
                           n10776, QN => n6701);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n3287, CK => CLK, Q => 
                           n10777, QN => n6702);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n3286, CK => CLK, Q => 
                           n10778, QN => n6703);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n3357, CK => CLK, Q => 
                           n10779, QN => n6632);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n3356, CK => CLK, Q => 
                           n10780, QN => n6633);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n3355, CK => CLK, Q => 
                           n10781, QN => n6634);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n3354, CK => CLK, Q => 
                           n10782, QN => n6635);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n3353, CK => CLK, Q => 
                           n10783, QN => n6636);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n3352, CK => CLK, Q => 
                           n10784, QN => n6637);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n3351, CK => CLK, Q => 
                           n10785, QN => n6638);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n3350, CK => CLK, Q => 
                           n10786, QN => n6639);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n3093, CK => CLK, Q => 
                           n_1016, QN => n8943);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n3092, CK => CLK, Q => 
                           n_1017, QN => n8958);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n3091, CK => CLK, Q => 
                           n_1018, QN => n8973);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n3090, CK => CLK, Q => 
                           n_1019, QN => n8988);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n3089, CK => CLK, Q => 
                           n_1020, QN => n9003);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n3088, CK => CLK, Q => 
                           n_1021, QN => n9018);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n3087, CK => CLK, Q => 
                           n_1022, QN => n9033);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n3086, CK => CLK, Q => 
                           n_1023, QN => n9048);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n3085, CK => CLK, Q => 
                           n_1024, QN => n9063);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n3084, CK => CLK, Q => 
                           n_1025, QN => n9078);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n3083, CK => CLK, Q => 
                           n_1026, QN => n9093);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n3082, CK => CLK, Q => 
                           n_1027, QN => n9108);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n3081, CK => CLK, Q => 
                           n_1028, QN => n9123);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n3080, CK => CLK, Q => 
                           n_1029, QN => n9138);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n3079, CK => CLK, Q => 
                           n_1030, QN => n9153);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n3078, CK => CLK, Q => 
                           n_1031, QN => n9168);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n3077, CK => CLK, Q => 
                           n_1032, QN => n9183);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n3076, CK => CLK, Q => 
                           n_1033, QN => n9198);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n3075, CK => CLK, Q => 
                           n_1034, QN => n9213);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n3074, CK => CLK, Q => 
                           n_1035, QN => n9228);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n3073, CK => CLK, Q => 
                           n_1036, QN => n9243);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n3072, CK => CLK, Q => 
                           n_1037, QN => n9258);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n3071, CK => CLK, Q => 
                           n_1038, QN => n9273);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n3070, CK => CLK, Q => 
                           n_1039, QN => n9288);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n3261, CK => CLK, Q => 
                           n10707, QN => n6728);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n3260, CK => CLK, Q => 
                           n10708, QN => n6729);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n3259, CK => CLK, Q => 
                           n10709, QN => n6730);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n3258, CK => CLK, Q => 
                           n10710, QN => n6731);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n3257, CK => CLK, Q => 
                           n10711, QN => n6732);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n3256, CK => CLK, Q => 
                           n10712, QN => n6733);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n3255, CK => CLK, Q => 
                           n10713, QN => n6734);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n3254, CK => CLK, Q => 
                           n10714, QN => n6735);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n3325, CK => CLK, Q => 
                           n10715, QN => n6664);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n3324, CK => CLK, Q => 
                           n10716, QN => n6665);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n3323, CK => CLK, Q => 
                           n10717, QN => n6666);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n3322, CK => CLK, Q => 
                           n10718, QN => n6667);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n3321, CK => CLK, Q => 
                           n10719, QN => n6668);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n3320, CK => CLK, Q => 
                           n10720, QN => n6669);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n3319, CK => CLK, Q => 
                           n10721, QN => n6670);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n3318, CK => CLK, Q => 
                           n10722, QN => n6671);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n3061, CK => CLK, Q => 
                           n_1040, QN => n8942);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n3060, CK => CLK, Q => 
                           n_1041, QN => n8957);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n3059, CK => CLK, Q => 
                           n_1042, QN => n8972);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n3058, CK => CLK, Q => 
                           n_1043, QN => n8987);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n3057, CK => CLK, Q => 
                           n_1044, QN => n9002);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n3056, CK => CLK, Q => 
                           n_1045, QN => n9017);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n3055, CK => CLK, Q => 
                           n_1046, QN => n9032);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n3054, CK => CLK, Q => 
                           n_1047, QN => n9047);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n3053, CK => CLK, Q => 
                           n_1048, QN => n9062);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n3052, CK => CLK, Q => 
                           n_1049, QN => n9077);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n3051, CK => CLK, Q => 
                           n_1050, QN => n9092);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n3050, CK => CLK, Q => 
                           n_1051, QN => n9107);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n3049, CK => CLK, Q => 
                           n_1052, QN => n9122);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n3048, CK => CLK, Q => 
                           n_1053, QN => n9137);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n3047, CK => CLK, Q => 
                           n_1054, QN => n9152);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n3046, CK => CLK, Q => 
                           n_1055, QN => n9167);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n3045, CK => CLK, Q => 
                           n_1056, QN => n9182);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n3044, CK => CLK, Q => 
                           n_1057, QN => n9197);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n3043, CK => CLK, Q => 
                           n_1058, QN => n9212);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n3042, CK => CLK, Q => 
                           n_1059, QN => n9227);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n3041, CK => CLK, Q => 
                           n_1060, QN => n9242);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n3040, CK => CLK, Q => 
                           n_1061, QN => n9257);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n3039, CK => CLK, Q => 
                           n_1062, QN => n9272);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n3038, CK => CLK, Q => 
                           n_1063, QN => n9287);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n3285, CK => CLK, Q => 
                           n10787, QN => n6704);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n3284, CK => CLK, Q => 
                           n10788, QN => n6705);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n3283, CK => CLK, Q => 
                           n10789, QN => n6706);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n3282, CK => CLK, Q => 
                           n10790, QN => n6707);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n3281, CK => CLK, Q => 
                           n10791, QN => n6708);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n3280, CK => CLK, Q => 
                           n10792, QN => n6709);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n3279, CK => CLK, Q => 
                           n10793, QN => n6710);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n3278, CK => CLK, Q => 
                           n10794, QN => n6711);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n3277, CK => CLK, Q => 
                           n10795, QN => n6712);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n3276, CK => CLK, Q => 
                           n10796, QN => n6713);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n3275, CK => CLK, Q => 
                           n10797, QN => n6714);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n3274, CK => CLK, Q => 
                           n10798, QN => n6715);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n3273, CK => CLK, Q => 
                           n10799, QN => n6716);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n3272, CK => CLK, Q => 
                           n10800, QN => n6717);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n3271, CK => CLK, Q => 
                           n10801, QN => n6718);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n3270, CK => CLK, Q => 
                           n10802, QN => n6719);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n3269, CK => CLK, Q => 
                           n10803, QN => n6720);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n3268, CK => CLK, Q => 
                           n10804, QN => n6721);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n3267, CK => CLK, Q => 
                           n10805, QN => n6722);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n3266, CK => CLK, Q => 
                           n10806, QN => n6723);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n3265, CK => CLK, Q => 
                           n10807, QN => n6724);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n3264, CK => CLK, Q => 
                           n10808, QN => n6725);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n3263, CK => CLK, Q => 
                           n10809, QN => n6726);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n3262, CK => CLK, Q => 
                           n10810, QN => n6727);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n3349, CK => CLK, Q => 
                           n10811, QN => n6640);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n3348, CK => CLK, Q => 
                           n10812, QN => n6641);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n3347, CK => CLK, Q => 
                           n10813, QN => n6642);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n3346, CK => CLK, Q => 
                           n10814, QN => n6643);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n3345, CK => CLK, Q => 
                           n10815, QN => n6644);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n3344, CK => CLK, Q => 
                           n10816, QN => n6645);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n3343, CK => CLK, Q => 
                           n10817, QN => n6646);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n3342, CK => CLK, Q => 
                           n10818, QN => n6647);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n3341, CK => CLK, Q => 
                           n10819, QN => n6648);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n3340, CK => CLK, Q => 
                           n10820, QN => n6649);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n3339, CK => CLK, Q => 
                           n10821, QN => n6650);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n3338, CK => CLK, Q => 
                           n10822, QN => n6651);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n3337, CK => CLK, Q => 
                           n10823, QN => n6652);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n3336, CK => CLK, Q => 
                           n10824, QN => n6653);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n3335, CK => CLK, Q => n10825
                           , QN => n6654);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n3334, CK => CLK, Q => n10826
                           , QN => n6655);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n3333, CK => CLK, Q => n10827
                           , QN => n6656);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n3332, CK => CLK, Q => n10828
                           , QN => n6657);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n3331, CK => CLK, Q => n10829
                           , QN => n6658);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n3330, CK => CLK, Q => n10830
                           , QN => n6659);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n3329, CK => CLK, Q => n10831
                           , QN => n6660);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n3328, CK => CLK, Q => n10832
                           , QN => n6661);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n3327, CK => CLK, Q => n10833
                           , QN => n6662);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n3326, CK => CLK, Q => n10834
                           , QN => n6663);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n3253, CK => CLK, Q => 
                           n10723, QN => n6736);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n3252, CK => CLK, Q => 
                           n10724, QN => n6737);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n3251, CK => CLK, Q => 
                           n10725, QN => n6738);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n3250, CK => CLK, Q => 
                           n10726, QN => n6739);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n3249, CK => CLK, Q => 
                           n10727, QN => n6740);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n3248, CK => CLK, Q => 
                           n10728, QN => n6741);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n3247, CK => CLK, Q => 
                           n10729, QN => n6742);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n3246, CK => CLK, Q => 
                           n10730, QN => n6743);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n3245, CK => CLK, Q => 
                           n10731, QN => n6744);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n3244, CK => CLK, Q => 
                           n10732, QN => n6745);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n3243, CK => CLK, Q => 
                           n10733, QN => n6746);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n3242, CK => CLK, Q => 
                           n10734, QN => n6747);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n3241, CK => CLK, Q => 
                           n10735, QN => n6748);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n3240, CK => CLK, Q => 
                           n10736, QN => n6749);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n3239, CK => CLK, Q => 
                           n10737, QN => n6750);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n3238, CK => CLK, Q => 
                           n10738, QN => n6751);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n3237, CK => CLK, Q => 
                           n10739, QN => n6752);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n3236, CK => CLK, Q => 
                           n10740, QN => n6753);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n3235, CK => CLK, Q => 
                           n10741, QN => n6754);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n3234, CK => CLK, Q => 
                           n10742, QN => n6755);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n3233, CK => CLK, Q => 
                           n10743, QN => n6756);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n3232, CK => CLK, Q => 
                           n10744, QN => n6757);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n3231, CK => CLK, Q => 
                           n10745, QN => n6758);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n3230, CK => CLK, Q => 
                           n10746, QN => n6759);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n3317, CK => CLK, Q => 
                           n10747, QN => n6672);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n3316, CK => CLK, Q => 
                           n10748, QN => n6673);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n3315, CK => CLK, Q => 
                           n10749, QN => n6674);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n3314, CK => CLK, Q => 
                           n10750, QN => n6675);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n3313, CK => CLK, Q => 
                           n10751, QN => n6676);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n3312, CK => CLK, Q => 
                           n10752, QN => n6677);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n3311, CK => CLK, Q => 
                           n10753, QN => n6678);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n3310, CK => CLK, Q => 
                           n10754, QN => n6679);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n3309, CK => CLK, Q => 
                           n10755, QN => n6680);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n3308, CK => CLK, Q => 
                           n10756, QN => n6681);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n3307, CK => CLK, Q => 
                           n10757, QN => n6682);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n3306, CK => CLK, Q => 
                           n10758, QN => n6683);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n3305, CK => CLK, Q => 
                           n10759, QN => n6684);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n3304, CK => CLK, Q => 
                           n10760, QN => n6685);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n3303, CK => CLK, Q => n10761
                           , QN => n6686);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n3302, CK => CLK, Q => n10762
                           , QN => n6687);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n3301, CK => CLK, Q => n10763
                           , QN => n6688);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n3300, CK => CLK, Q => n10764
                           , QN => n6689);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n3299, CK => CLK, Q => n10765
                           , QN => n6690);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n3298, CK => CLK, Q => n10766
                           , QN => n6691);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n3297, CK => CLK, Q => n10767
                           , QN => n6692);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n3296, CK => CLK, Q => n10768
                           , QN => n6693);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n3295, CK => CLK, Q => n10769
                           , QN => n6694);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n3294, CK => CLK, Q => n10770
                           , QN => n6695);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n2717, CK => CLK, Q => 
                           n_1064, QN => n10355);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n2716, CK => CLK, Q => 
                           n_1065, QN => n10356);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n2715, CK => CLK, Q => 
                           n_1066, QN => n10357);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n2714, CK => CLK, Q => 
                           n_1067, QN => n10358);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n2713, CK => CLK, Q => 
                           n_1068, QN => n10359);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n2712, CK => CLK, Q => 
                           n_1069, QN => n10360);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n2711, CK => CLK, Q => 
                           n_1070, QN => n10361);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n2710, CK => CLK, Q => 
                           n_1071, QN => n10362);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n2845, CK => CLK, Q => 
                           n_1072, QN => n10363);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n2844, CK => CLK, Q => 
                           n_1073, QN => n10364);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n2843, CK => CLK, Q => 
                           n_1074, QN => n10365);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n2842, CK => CLK, Q => 
                           n_1075, QN => n10366);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n2841, CK => CLK, Q => 
                           n_1076, QN => n10367);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n2840, CK => CLK, Q => 
                           n_1077, QN => n10368);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n2839, CK => CLK, Q => 
                           n_1078, QN => n10369);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n2838, CK => CLK, Q => 
                           n_1079, QN => n10370);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n2909, CK => CLK, Q => 
                           n_1080, QN => n10371);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n2908, CK => CLK, Q => 
                           n_1081, QN => n10372);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n2907, CK => CLK, Q => 
                           n_1082, QN => n10373);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n2906, CK => CLK, Q => 
                           n_1083, QN => n10374);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n2905, CK => CLK, Q => 
                           n_1084, QN => n10375);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n2904, CK => CLK, Q => 
                           n_1085, QN => n10376);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n2903, CK => CLK, Q => 
                           n_1086, QN => n10377);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n2902, CK => CLK, Q => 
                           n_1087, QN => n10378);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n3165, CK => CLK, Q => 
                           n_1088, QN => n10387);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n3164, CK => CLK, Q => 
                           n_1089, QN => n10388);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n3163, CK => CLK, Q => 
                           n_1090, QN => n10389);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n3162, CK => CLK, Q => 
                           n_1091, QN => n10390);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n3161, CK => CLK, Q => 
                           n_1092, QN => n10391);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n3160, CK => CLK, Q => 
                           n_1093, QN => n10392);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n3159, CK => CLK, Q => 
                           n_1094, QN => n10393);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n3158, CK => CLK, Q => 
                           n_1095, QN => n10394);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n3421, CK => CLK, Q => 
                           n_1096, QN => n10347);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n3420, CK => CLK, Q => 
                           n_1097, QN => n9964);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n3419, CK => CLK, Q => 
                           n_1098, QN => n9965);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n3418, CK => CLK, Q => 
                           n_1099, QN => n9966);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n3417, CK => CLK, Q => 
                           n_1100, QN => n9967);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n3416, CK => CLK, Q => 
                           n_1101, QN => n9968);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n3415, CK => CLK, Q => 
                           n_1102, QN => n9969);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n3414, CK => CLK, Q => 
                           n_1103, QN => n9970);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n3581, CK => CLK, Q => 
                           n_1104, QN => n10395);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n3580, CK => CLK, Q => 
                           n_1105, QN => n10396);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n3579, CK => CLK, Q => 
                           n_1106, QN => n10397);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n3578, CK => CLK, Q => 
                           n_1107, QN => n10398);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n3577, CK => CLK, Q => 
                           n_1108, QN => n10399);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n3576, CK => CLK, Q => 
                           n_1109, QN => n10400);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n3575, CK => CLK, Q => 
                           n_1110, QN => n10401);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n3574, CK => CLK, Q => 
                           n_1111, QN => n10402);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n2685, CK => CLK, Q => 
                           n_1112, QN => n10403);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n2684, CK => CLK, Q => 
                           n_1113, QN => n10404);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n2683, CK => CLK, Q => 
                           n_1114, QN => n10405);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n2682, CK => CLK, Q => 
                           n_1115, QN => n10406);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n2681, CK => CLK, Q => 
                           n_1116, QN => n10407);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n2680, CK => CLK, Q => 
                           n_1117, QN => n10408);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n2679, CK => CLK, Q => 
                           n_1118, QN => n10409);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n2678, CK => CLK, Q => 
                           n_1119, QN => n10410);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n2813, CK => CLK, Q => 
                           n_1120, QN => n10411);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n2812, CK => CLK, Q => 
                           n_1121, QN => n10412);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n2811, CK => CLK, Q => 
                           n_1122, QN => n10413);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n2810, CK => CLK, Q => 
                           n_1123, QN => n10414);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n2809, CK => CLK, Q => 
                           n_1124, QN => n10415);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n2808, CK => CLK, Q => 
                           n_1125, QN => n10416);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n2807, CK => CLK, Q => 
                           n_1126, QN => n10417);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n2806, CK => CLK, Q => 
                           n_1127, QN => n10418);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n2877, CK => CLK, Q => 
                           n_1128, QN => n10419);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n2876, CK => CLK, Q => 
                           n_1129, QN => n10420);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n2875, CK => CLK, Q => 
                           n_1130, QN => n10421);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n2874, CK => CLK, Q => 
                           n_1131, QN => n10422);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n2873, CK => CLK, Q => 
                           n_1132, QN => n10423);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n2872, CK => CLK, Q => 
                           n_1133, QN => n10424);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n2871, CK => CLK, Q => 
                           n_1134, QN => n10425);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n2870, CK => CLK, Q => 
                           n_1135, QN => n10426);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n3133, CK => CLK, Q => 
                           n_1136, QN => n10435);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n3132, CK => CLK, Q => 
                           n_1137, QN => n10436);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n3131, CK => CLK, Q => 
                           n_1138, QN => n10437);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n3130, CK => CLK, Q => 
                           n_1139, QN => n10438);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n3129, CK => CLK, Q => 
                           n_1140, QN => n10439);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n3128, CK => CLK, Q => 
                           n_1141, QN => n10440);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n3127, CK => CLK, Q => 
                           n_1142, QN => n10441);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n3126, CK => CLK, Q => 
                           n_1143, QN => n10442);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n3389, CK => CLK, Q => 
                           n_1144, QN => n9995);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n3388, CK => CLK, Q => 
                           n_1145, QN => n9996);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n3387, CK => CLK, Q => 
                           n_1146, QN => n9997);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n3386, CK => CLK, Q => 
                           n_1147, QN => n9998);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n3385, CK => CLK, Q => 
                           n_1148, QN => n9999);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n3384, CK => CLK, Q => 
                           n_1149, QN => n10000);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n3383, CK => CLK, Q => 
                           n_1150, QN => n10001);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n3382, CK => CLK, Q => 
                           n_1151, QN => n10002);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n3613, CK => CLK, Q => 
                           n_1152, QN => n10567);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n3612, CK => CLK, Q => 
                           n_1153, QN => n10568);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n3611, CK => CLK, Q => 
                           n_1154, QN => n10569);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n3610, CK => CLK, Q => 
                           n_1155, QN => n10570);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n3609, CK => CLK, Q => 
                           n_1156, QN => n9939);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n3608, CK => CLK, Q => 
                           n_1157, QN => n9940);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n3607, CK => CLK, Q => 
                           n_1158, QN => n9941);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n3606, CK => CLK, Q => 
                           n_1159, QN => n9942);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n2709, CK => CLK, Q => 
                           n_1160, QN => n10447);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n2708, CK => CLK, Q => 
                           n_1161, QN => n10448);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n2707, CK => CLK, Q => 
                           n_1162, QN => n10449);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n2706, CK => CLK, Q => 
                           n_1163, QN => n10450);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n2705, CK => CLK, Q => 
                           n_1164, QN => n10451);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n2704, CK => CLK, Q => 
                           n_1165, QN => n10452);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n2703, CK => CLK, Q => 
                           n_1166, QN => n10453);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n2702, CK => CLK, Q => 
                           n_1167, QN => n10454);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n2701, CK => CLK, Q => 
                           n_1168, QN => n10455);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n2700, CK => CLK, Q => 
                           n_1169, QN => n10456);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n2699, CK => CLK, Q => 
                           n_1170, QN => n10457);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n2698, CK => CLK, Q => 
                           n_1171, QN => n10458);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n2697, CK => CLK, Q => 
                           n_1172, QN => n10459);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n2696, CK => CLK, Q => 
                           n_1173, QN => n10460);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n2695, CK => CLK, Q => 
                           n_1174, QN => n10461);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n2694, CK => CLK, Q => 
                           n_1175, QN => n10462);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n2693, CK => CLK, Q => 
                           n_1176, QN => n10463);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n2692, CK => CLK, Q => 
                           n_1177, QN => n10464);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n2691, CK => CLK, Q => 
                           n_1178, QN => n10465);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n2690, CK => CLK, Q => 
                           n_1179, QN => n10466);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n2689, CK => CLK, Q => 
                           n_1180, QN => n10467);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n2688, CK => CLK, Q => 
                           n_1181, QN => n10468);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n2687, CK => CLK, Q => 
                           n_1182, QN => n10469);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n2686, CK => CLK, Q => 
                           n_1183, QN => n10470);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n2837, CK => CLK, Q => 
                           n_1184, QN => n10471);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n2836, CK => CLK, Q => 
                           n_1185, QN => n10472);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n2835, CK => CLK, Q => 
                           n_1186, QN => n10473);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n2834, CK => CLK, Q => 
                           n_1187, QN => n10474);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n2833, CK => CLK, Q => 
                           n_1188, QN => n10475);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n2832, CK => CLK, Q => 
                           n_1189, QN => n10476);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n2831, CK => CLK, Q => 
                           n_1190, QN => n10477);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n2830, CK => CLK, Q => 
                           n_1191, QN => n10478);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n2829, CK => CLK, Q => 
                           n_1192, QN => n10479);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n2828, CK => CLK, Q => 
                           n_1193, QN => n10480);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n2827, CK => CLK, Q => 
                           n_1194, QN => n10481);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n2826, CK => CLK, Q => 
                           n_1195, QN => n10482);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n2825, CK => CLK, Q => 
                           n_1196, QN => n10483);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n2824, CK => CLK, Q => 
                           n_1197, QN => n10484);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n2823, CK => CLK, Q => 
                           n_1198, QN => n10485);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n2822, CK => CLK, Q => 
                           n_1199, QN => n10486);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n2821, CK => CLK, Q => 
                           n_1200, QN => n10487);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n2820, CK => CLK, Q => 
                           n_1201, QN => n10488);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n2819, CK => CLK, Q => 
                           n_1202, QN => n10489);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n2818, CK => CLK, Q => 
                           n_1203, QN => n10490);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n2817, CK => CLK, Q => 
                           n_1204, QN => n10491);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n2816, CK => CLK, Q => 
                           n_1205, QN => n10492);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n2815, CK => CLK, Q => 
                           n_1206, QN => n10493);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n2814, CK => CLK, Q => 
                           n_1207, QN => n10494);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n2901, CK => CLK, Q => 
                           n_1208, QN => n10495);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n2900, CK => CLK, Q => 
                           n_1209, QN => n10496);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n2899, CK => CLK, Q => 
                           n_1210, QN => n10497);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n2898, CK => CLK, Q => 
                           n_1211, QN => n10498);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n2897, CK => CLK, Q => 
                           n_1212, QN => n10499);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n2896, CK => CLK, Q => 
                           n_1213, QN => n10500);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n2895, CK => CLK, Q => 
                           n_1214, QN => n10501);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n2894, CK => CLK, Q => 
                           n_1215, QN => n10502);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n2893, CK => CLK, Q => 
                           n_1216, QN => n10503);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n2892, CK => CLK, Q => 
                           n_1217, QN => n10504);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n2891, CK => CLK, Q => 
                           n_1218, QN => n10505);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n2890, CK => CLK, Q => 
                           n_1219, QN => n10506);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n2889, CK => CLK, Q => 
                           n_1220, QN => n10507);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n2888, CK => CLK, Q => 
                           n_1221, QN => n10508);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n2887, CK => CLK, Q => 
                           n_1222, QN => n10509);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n2886, CK => CLK, Q => 
                           n_1223, QN => n10510);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n2885, CK => CLK, Q => 
                           n_1224, QN => n10511);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n2884, CK => CLK, Q => 
                           n_1225, QN => n10512);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n2883, CK => CLK, Q => 
                           n_1226, QN => n10513);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n2882, CK => CLK, Q => 
                           n_1227, QN => n10514);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n2881, CK => CLK, Q => 
                           n_1228, QN => n10515);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n2880, CK => CLK, Q => 
                           n_1229, QN => n10516);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n2879, CK => CLK, Q => 
                           n_1230, QN => n10517);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n2878, CK => CLK, Q => 
                           n_1231, QN => n10518);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n3157, CK => CLK, Q => 
                           n_1232, QN => n10543);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n3156, CK => CLK, Q => 
                           n_1233, QN => n10544);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n3155, CK => CLK, Q => 
                           n_1234, QN => n10545);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n3154, CK => CLK, Q => 
                           n_1235, QN => n10546);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n3153, CK => CLK, Q => 
                           n_1236, QN => n10547);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n3152, CK => CLK, Q => 
                           n_1237, QN => n10548);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n3151, CK => CLK, Q => 
                           n_1238, QN => n10549);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n3150, CK => CLK, Q => 
                           n_1239, QN => n10550);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n3149, CK => CLK, Q => 
                           n_1240, QN => n10551);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n3148, CK => CLK, Q => 
                           n_1241, QN => n10552);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n3147, CK => CLK, Q => 
                           n_1242, QN => n10553);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n3146, CK => CLK, Q => 
                           n_1243, QN => n10554);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n3145, CK => CLK, Q => 
                           n_1244, QN => n10555);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n3144, CK => CLK, Q => 
                           n_1245, QN => n10556);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n3143, CK => CLK, Q => 
                           n_1246, QN => n10557);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n3142, CK => CLK, Q => 
                           n_1247, QN => n10558);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n3141, CK => CLK, Q => 
                           n_1248, QN => n10559);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n3140, CK => CLK, Q => 
                           n_1249, QN => n10560);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n3139, CK => CLK, Q => 
                           n_1250, QN => n10561);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n3138, CK => CLK, Q => 
                           n_1251, QN => n10562);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n3137, CK => CLK, Q => 
                           n_1252, QN => n10563);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n3136, CK => CLK, Q => 
                           n_1253, QN => n10564);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n3135, CK => CLK, Q => 
                           n_1254, QN => n10565);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n3134, CK => CLK, Q => 
                           n_1255, QN => n10566);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n3413, CK => CLK, Q => 
                           n_1256, QN => n9971);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n3412, CK => CLK, Q => 
                           n_1257, QN => n9972);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n3411, CK => CLK, Q => 
                           n_1258, QN => n9973);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n3410, CK => CLK, Q => 
                           n_1259, QN => n9974);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n3409, CK => CLK, Q => 
                           n_1260, QN => n9975);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n3408, CK => CLK, Q => 
                           n_1261, QN => n9976);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n3407, CK => CLK, Q => 
                           n_1262, QN => n9977);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n3406, CK => CLK, Q => 
                           n_1263, QN => n9978);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n3405, CK => CLK, Q => 
                           n_1264, QN => n9979);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n3404, CK => CLK, Q => 
                           n_1265, QN => n9980);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n3403, CK => CLK, Q => 
                           n_1266, QN => n9981);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n3402, CK => CLK, Q => 
                           n_1267, QN => n9982);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n3401, CK => CLK, Q => 
                           n_1268, QN => n9983);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n3400, CK => CLK, Q => 
                           n_1269, QN => n9984);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n3399, CK => CLK, Q => n_1270
                           , QN => n9985);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n3398, CK => CLK, Q => n_1271
                           , QN => n9986);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n3397, CK => CLK, Q => n_1272
                           , QN => n9987);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n3396, CK => CLK, Q => n_1273
                           , QN => n9988);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n3395, CK => CLK, Q => n_1274
                           , QN => n9989);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n3394, CK => CLK, Q => n_1275
                           , QN => n9990);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n3393, CK => CLK, Q => n_1276
                           , QN => n9991);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n3392, CK => CLK, Q => n_1277
                           , QN => n9992);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n3391, CK => CLK, Q => n_1278
                           , QN => n9993);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n3390, CK => CLK, Q => n_1279
                           , QN => n9994);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n3573, CK => CLK, Q => 
                           n_1280, QN => n10443);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n3572, CK => CLK, Q => 
                           n_1281, QN => n10444);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n3571, CK => CLK, Q => 
                           n_1282, QN => n10445);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n3570, CK => CLK, Q => 
                           n_1283, QN => n10446);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n3569, CK => CLK, Q => 
                           n_1284, QN => n9944);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n3568, CK => CLK, Q => 
                           n_1285, QN => n9945);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n3567, CK => CLK, Q => 
                           n_1286, QN => n9946);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n3566, CK => CLK, Q => 
                           n_1287, QN => n9947);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n3565, CK => CLK, Q => 
                           n_1288, QN => n9948);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n3564, CK => CLK, Q => 
                           n_1289, QN => n9949);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n3563, CK => CLK, Q => 
                           n_1290, QN => n9950);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n3562, CK => CLK, Q => 
                           n_1291, QN => n9951);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n3561, CK => CLK, Q => 
                           n_1292, QN => n9952);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n3560, CK => CLK, Q => 
                           n_1293, QN => n9953);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n3559, CK => CLK, Q => n_1294
                           , QN => n9954);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n3558, CK => CLK, Q => n_1295
                           , QN => n9955);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n3557, CK => CLK, Q => n_1296
                           , QN => n9956);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n3556, CK => CLK, Q => n_1297
                           , QN => n9957);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n3555, CK => CLK, Q => n_1298
                           , QN => n9958);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n3554, CK => CLK, Q => n_1299
                           , QN => n9959);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n3553, CK => CLK, Q => n_1300
                           , QN => n9960);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n3552, CK => CLK, Q => n_1301
                           , QN => n9961);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n3551, CK => CLK, Q => n_1302
                           , QN => n9962);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n3550, CK => CLK, Q => n_1303
                           , QN => n9963);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n2677, CK => CLK, Q => 
                           n_1304, QN => n10574);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n2676, CK => CLK, Q => 
                           n_1305, QN => n10575);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n2675, CK => CLK, Q => 
                           n_1306, QN => n10576);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n2674, CK => CLK, Q => 
                           n_1307, QN => n10577);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n2673, CK => CLK, Q => 
                           n_1308, QN => n10578);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n2672, CK => CLK, Q => 
                           n_1309, QN => n10579);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n2671, CK => CLK, Q => 
                           n_1310, QN => n10580);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n2670, CK => CLK, Q => 
                           n_1311, QN => n10581);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n2669, CK => CLK, Q => 
                           n_1312, QN => n10582);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n2668, CK => CLK, Q => 
                           n_1313, QN => n10583);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n2667, CK => CLK, Q => 
                           n_1314, QN => n10584);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n2666, CK => CLK, Q => 
                           n_1315, QN => n10585);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n2665, CK => CLK, Q => 
                           n_1316, QN => n10586);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n2664, CK => CLK, Q => 
                           n_1317, QN => n10587);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n2663, CK => CLK, Q => 
                           n_1318, QN => n10588);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n2662, CK => CLK, Q => 
                           n_1319, QN => n10589);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n2661, CK => CLK, Q => 
                           n_1320, QN => n10590);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n2660, CK => CLK, Q => 
                           n_1321, QN => n10591);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n2659, CK => CLK, Q => 
                           n_1322, QN => n10592);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n2658, CK => CLK, Q => 
                           n_1323, QN => n10593);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n2657, CK => CLK, Q => 
                           n_1324, QN => n10594);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n2656, CK => CLK, Q => 
                           n_1325, QN => n10595);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n2655, CK => CLK, Q => 
                           n_1326, QN => n10596);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n2654, CK => CLK, Q => 
                           n_1327, QN => n10597);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n2805, CK => CLK, Q => 
                           n_1328, QN => n10598);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n2804, CK => CLK, Q => 
                           n_1329, QN => n10599);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n2803, CK => CLK, Q => 
                           n_1330, QN => n10600);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n2802, CK => CLK, Q => 
                           n_1331, QN => n10601);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n2801, CK => CLK, Q => 
                           n_1332, QN => n10602);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n2800, CK => CLK, Q => 
                           n_1333, QN => n10603);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n2799, CK => CLK, Q => 
                           n_1334, QN => n10604);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n2798, CK => CLK, Q => 
                           n_1335, QN => n10605);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n2797, CK => CLK, Q => 
                           n_1336, QN => n10606);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n2796, CK => CLK, Q => 
                           n_1337, QN => n10607);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n2795, CK => CLK, Q => 
                           n_1338, QN => n10608);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n2794, CK => CLK, Q => 
                           n_1339, QN => n10609);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n2793, CK => CLK, Q => 
                           n_1340, QN => n10610);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n2792, CK => CLK, Q => 
                           n_1341, QN => n10611);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n2791, CK => CLK, Q => 
                           n_1342, QN => n10612);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n2790, CK => CLK, Q => 
                           n_1343, QN => n10613);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n2789, CK => CLK, Q => 
                           n_1344, QN => n10614);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n2788, CK => CLK, Q => 
                           n_1345, QN => n10615);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n2787, CK => CLK, Q => 
                           n_1346, QN => n10616);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n2786, CK => CLK, Q => 
                           n_1347, QN => n10617);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n2785, CK => CLK, Q => 
                           n_1348, QN => n10618);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n2784, CK => CLK, Q => 
                           n_1349, QN => n10619);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n2783, CK => CLK, Q => 
                           n_1350, QN => n10620);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n2782, CK => CLK, Q => 
                           n_1351, QN => n10621);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n2869, CK => CLK, Q => 
                           n_1352, QN => n10622);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n2868, CK => CLK, Q => 
                           n_1353, QN => n10623);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n2867, CK => CLK, Q => 
                           n_1354, QN => n10624);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n2866, CK => CLK, Q => 
                           n_1355, QN => n10625);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n2865, CK => CLK, Q => 
                           n_1356, QN => n10626);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n2864, CK => CLK, Q => 
                           n_1357, QN => n10627);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n2863, CK => CLK, Q => 
                           n_1358, QN => n10628);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n2862, CK => CLK, Q => 
                           n_1359, QN => n10629);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n2861, CK => CLK, Q => 
                           n_1360, QN => n10630);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n2860, CK => CLK, Q => 
                           n_1361, QN => n10631);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n2859, CK => CLK, Q => 
                           n_1362, QN => n10632);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n2858, CK => CLK, Q => 
                           n_1363, QN => n10633);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n2857, CK => CLK, Q => 
                           n_1364, QN => n10634);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n2856, CK => CLK, Q => 
                           n_1365, QN => n10635);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n2855, CK => CLK, Q => 
                           n_1366, QN => n10636);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n2854, CK => CLK, Q => 
                           n_1367, QN => n10637);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n2853, CK => CLK, Q => 
                           n_1368, QN => n10638);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n2852, CK => CLK, Q => 
                           n_1369, QN => n10639);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n2851, CK => CLK, Q => 
                           n_1370, QN => n10640);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n2850, CK => CLK, Q => 
                           n_1371, QN => n10641);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n2849, CK => CLK, Q => 
                           n_1372, QN => n10642);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n2848, CK => CLK, Q => 
                           n_1373, QN => n10643);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n2847, CK => CLK, Q => 
                           n_1374, QN => n10644);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n2846, CK => CLK, Q => 
                           n_1375, QN => n10645);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n3125, CK => CLK, Q => 
                           n_1376, QN => n10670);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n3124, CK => CLK, Q => 
                           n_1377, QN => n10671);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n3123, CK => CLK, Q => 
                           n_1378, QN => n10672);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n3122, CK => CLK, Q => 
                           n_1379, QN => n10673);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n3121, CK => CLK, Q => 
                           n_1380, QN => n10674);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n3120, CK => CLK, Q => 
                           n_1381, QN => n10675);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n3119, CK => CLK, Q => 
                           n_1382, QN => n10676);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n3118, CK => CLK, Q => 
                           n_1383, QN => n10677);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n3117, CK => CLK, Q => 
                           n_1384, QN => n10678);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n3116, CK => CLK, Q => 
                           n_1385, QN => n10679);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n3115, CK => CLK, Q => 
                           n_1386, QN => n10680);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n3114, CK => CLK, Q => 
                           n_1387, QN => n10681);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n3113, CK => CLK, Q => 
                           n_1388, QN => n10682);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n3112, CK => CLK, Q => 
                           n_1389, QN => n10683);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n3111, CK => CLK, Q => 
                           n_1390, QN => n10684);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n3110, CK => CLK, Q => 
                           n_1391, QN => n10685);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n3109, CK => CLK, Q => 
                           n_1392, QN => n10686);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n3108, CK => CLK, Q => 
                           n_1393, QN => n10687);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n3107, CK => CLK, Q => 
                           n_1394, QN => n10688);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n3106, CK => CLK, Q => 
                           n_1395, QN => n10689);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n3105, CK => CLK, Q => 
                           n_1396, QN => n10690);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n3104, CK => CLK, Q => 
                           n_1397, QN => n10691);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n3103, CK => CLK, Q => 
                           n_1398, QN => n10692);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n3102, CK => CLK, Q => 
                           n_1399, QN => n10693);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n3381, CK => CLK, Q => 
                           n_1400, QN => n10003);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n3380, CK => CLK, Q => 
                           n_1401, QN => n10004);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n3379, CK => CLK, Q => 
                           n_1402, QN => n10005);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n3378, CK => CLK, Q => 
                           n_1403, QN => n10006);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n3377, CK => CLK, Q => 
                           n_1404, QN => n10007);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n3376, CK => CLK, Q => 
                           n_1405, QN => n10008);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n3375, CK => CLK, Q => 
                           n_1406, QN => n10009);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n3374, CK => CLK, Q => 
                           n_1407, QN => n10010);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n3373, CK => CLK, Q => 
                           n_1408, QN => n10011);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n3372, CK => CLK, Q => 
                           n_1409, QN => n10012);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n3371, CK => CLK, Q => 
                           n_1410, QN => n10013);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n3370, CK => CLK, Q => 
                           n_1411, QN => n10014);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n3369, CK => CLK, Q => 
                           n_1412, QN => n10015);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n3368, CK => CLK, Q => 
                           n_1413, QN => n10016);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n3367, CK => CLK, Q => n_1414
                           , QN => n10017);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n3366, CK => CLK, Q => n_1415
                           , QN => n10018);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n3365, CK => CLK, Q => n_1416
                           , QN => n10019);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n3364, CK => CLK, Q => n_1417
                           , QN => n10020);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n3363, CK => CLK, Q => n_1418
                           , QN => n10021);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n3362, CK => CLK, Q => n_1419
                           , QN => n10022);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n3361, CK => CLK, Q => n_1420
                           , QN => n10023);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n3360, CK => CLK, Q => n_1421
                           , QN => n10024);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n3359, CK => CLK, Q => n_1422
                           , QN => n10025);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n3358, CK => CLK, Q => n_1423
                           , QN => n10026);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n3605, CK => CLK, Q => 
                           n_1424, QN => n9943);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n3604, CK => CLK, Q => 
                           n_1425, QN => n10571);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n3603, CK => CLK, Q => 
                           n_1426, QN => n10572);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n3602, CK => CLK, Q => 
                           n_1427, QN => n10573);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n3601, CK => CLK, Q => 
                           n_1428, QN => n10694);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n3600, CK => CLK, Q => 
                           n_1429, QN => n10695);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n3599, CK => CLK, Q => 
                           n_1430, QN => n10696);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n3598, CK => CLK, Q => 
                           n_1431, QN => n10697);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n3597, CK => CLK, Q => 
                           n_1432, QN => n10698);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n3596, CK => CLK, Q => 
                           n_1433, QN => n10699);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n3595, CK => CLK, Q => 
                           n_1434, QN => n10700);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n3594, CK => CLK, Q => 
                           n_1435, QN => n10701);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n3593, CK => CLK, Q => 
                           n_1436, QN => n10702);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n3592, CK => CLK, Q => 
                           n_1437, QN => n10703);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n3591, CK => CLK, Q => n_1438
                           , QN => n10704);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n3590, CK => CLK, Q => n_1439
                           , QN => n10705);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n3589, CK => CLK, Q => n_1440
                           , QN => n10348);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n3588, CK => CLK, Q => n_1441
                           , QN => n10349);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n3587, CK => CLK, Q => n_1442
                           , QN => n10350);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n3586, CK => CLK, Q => n_1443
                           , QN => n10351);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n3585, CK => CLK, Q => n_1444
                           , QN => n10352);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n3584, CK => CLK, Q => n_1445
                           , QN => n10353);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n3583, CK => CLK, Q => n_1446
                           , QN => n10354);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n3582, CK => CLK, Q => n_1447
                           , QN => n10706);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n3037, CK => CLK, Q => 
                           n12345, QN => n10379);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n3036, CK => CLK, Q => 
                           n12344, QN => n10380);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n3035, CK => CLK, Q => 
                           n12343, QN => n10381);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n3034, CK => CLK, Q => 
                           n12342, QN => n10382);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n3033, CK => CLK, Q => 
                           n12341, QN => n10383);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n3032, CK => CLK, Q => 
                           n12340, QN => n10384);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n3031, CK => CLK, Q => 
                           n12339, QN => n10385);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n3030, CK => CLK, Q => 
                           n12338, QN => n10386);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n3029, CK => CLK, Q => 
                           n12567, QN => n10519);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n3028, CK => CLK, Q => 
                           n12566, QN => n10520);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n3027, CK => CLK, Q => 
                           n12565, QN => n10521);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n3026, CK => CLK, Q => 
                           n12564, QN => n10522);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n3025, CK => CLK, Q => 
                           n12563, QN => n10523);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n3024, CK => CLK, Q => 
                           n12562, QN => n10524);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n3023, CK => CLK, Q => 
                           n12561, QN => n10525);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n3022, CK => CLK, Q => 
                           n12560, QN => n10526);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n3021, CK => CLK, Q => 
                           n12559, QN => n10527);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n3020, CK => CLK, Q => 
                           n12558, QN => n10528);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n3019, CK => CLK, Q => 
                           n12557, QN => n10529);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n3018, CK => CLK, Q => 
                           n12556, QN => n10530);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n3017, CK => CLK, Q => 
                           n12555, QN => n10531);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n3016, CK => CLK, Q => 
                           n12554, QN => n10532);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n3015, CK => CLK, Q => 
                           n12553, QN => n10533);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n3014, CK => CLK, Q => 
                           n12552, QN => n10534);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n3013, CK => CLK, Q => 
                           n12551, QN => n10535);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n3012, CK => CLK, Q => 
                           n12550, QN => n10536);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n3011, CK => CLK, Q => 
                           n12549, QN => n10537);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n3010, CK => CLK, Q => 
                           n12548, QN => n10538);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n3009, CK => CLK, Q => 
                           n12547, QN => n10539);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n3008, CK => CLK, Q => 
                           n12546, QN => n10540);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n3007, CK => CLK, Q => 
                           n12545, QN => n10541);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n3006, CK => CLK, Q => 
                           n12544, QN => n10542);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n3005, CK => CLK, Q => 
                           n12337, QN => n10427);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n3004, CK => CLK, Q => 
                           n12336, QN => n10428);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n3003, CK => CLK, Q => 
                           n12335, QN => n10429);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n3002, CK => CLK, Q => 
                           n12334, QN => n10430);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n3001, CK => CLK, Q => 
                           n12333, QN => n10431);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n3000, CK => CLK, Q => 
                           n12332, QN => n10432);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n2999, CK => CLK, Q => 
                           n12331, QN => n10433);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n2998, CK => CLK, Q => 
                           n12330, QN => n10434);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n2997, CK => CLK, Q => 
                           n12543, QN => n10646);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n2996, CK => CLK, Q => 
                           n12542, QN => n10647);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n2995, CK => CLK, Q => 
                           n12541, QN => n10648);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n2994, CK => CLK, Q => 
                           n12540, QN => n10649);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n2993, CK => CLK, Q => 
                           n12539, QN => n10650);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n2992, CK => CLK, Q => 
                           n12538, QN => n10651);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n2991, CK => CLK, Q => 
                           n12537, QN => n10652);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n2990, CK => CLK, Q => 
                           n12536, QN => n10653);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n2989, CK => CLK, Q => 
                           n12535, QN => n10654);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n2988, CK => CLK, Q => 
                           n12534, QN => n10655);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n2987, CK => CLK, Q => 
                           n12533, QN => n10656);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n2986, CK => CLK, Q => 
                           n12532, QN => n10657);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n2985, CK => CLK, Q => 
                           n12531, QN => n10658);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n2984, CK => CLK, Q => 
                           n12530, QN => n10659);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n2983, CK => CLK, Q => 
                           n12529, QN => n10660);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n2982, CK => CLK, Q => 
                           n12528, QN => n10661);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n2981, CK => CLK, Q => 
                           n12527, QN => n10662);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n2980, CK => CLK, Q => 
                           n12526, QN => n10663);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n2979, CK => CLK, Q => 
                           n12525, QN => n10664);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n2978, CK => CLK, Q => 
                           n12524, QN => n10665);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n2977, CK => CLK, Q => 
                           n12523, QN => n10666);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n2976, CK => CLK, Q => 
                           n12522, QN => n10667);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n2975, CK => CLK, Q => 
                           n12521, QN => n10668);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n2974, CK => CLK, Q => 
                           n12520, QN => n10669);
   U9459 : NOR2_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), ZN => n12260);
   U9460 : NOR2_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), ZN => n11607);
   U9461 : INV_X1 port map( A => n13314, ZN => n13307);
   U9462 : INV_X1 port map( A => n13185, ZN => n13178);
   U9463 : INV_X1 port map( A => n13176, ZN => n13169);
   U9464 : INV_X1 port map( A => n13149, ZN => n13142);
   U9465 : INV_X1 port map( A => n13131, ZN => n13124);
   U9466 : INV_X1 port map( A => n13140, ZN => n13133);
   U9467 : INV_X1 port map( A => n13122, ZN => n13115);
   U9468 : INV_X1 port map( A => n13203, ZN => n13196);
   U9469 : INV_X1 port map( A => n13194, ZN => n13187);
   U9470 : INV_X1 port map( A => n13113, ZN => n13106);
   U9471 : INV_X1 port map( A => n13104, ZN => n13097);
   U9472 : INV_X1 port map( A => n13077, ZN => n13070);
   U9473 : INV_X1 port map( A => n13068, ZN => n13061);
   U9474 : INV_X1 port map( A => n13041, ZN => n13034);
   U9475 : INV_X1 port map( A => n13032, ZN => n13025);
   U9476 : INV_X1 port map( A => n12987, ZN => n12980);
   U9477 : INV_X1 port map( A => n12978, ZN => n12971);
   U9478 : INV_X1 port map( A => n12951, ZN => n12944);
   U9479 : INV_X1 port map( A => n13086, ZN => n13079);
   U9480 : INV_X1 port map( A => n13050, ZN => n13043);
   U9481 : INV_X1 port map( A => n13014, ZN => n13007);
   U9482 : INV_X1 port map( A => n12996, ZN => n12989);
   U9483 : INV_X1 port map( A => n12960, ZN => n12953);
   U9484 : INV_X1 port map( A => n13095, ZN => n13088);
   U9485 : INV_X1 port map( A => n13059, ZN => n13052);
   U9486 : INV_X1 port map( A => n13023, ZN => n13016);
   U9487 : INV_X1 port map( A => n13005, ZN => n12998);
   U9488 : INV_X1 port map( A => n12969, ZN => n12962);
   U9489 : INV_X1 port map( A => n13158, ZN => n13151);
   U9490 : INV_X1 port map( A => n13167, ZN => n13160);
   U9491 : INV_X1 port map( A => n13212, ZN => n13205);
   U9492 : BUF_X1 port map( A => n11677, Z => n12736);
   U9493 : BUF_X1 port map( A => n11677, Z => n12737);
   U9494 : BUF_X1 port map( A => n11024, Z => n12838);
   U9495 : BUF_X1 port map( A => n11024, Z => n12839);
   U9496 : BUF_X1 port map( A => n11677, Z => n12738);
   U9497 : BUF_X1 port map( A => n11024, Z => n12840);
   U9498 : BUF_X1 port map( A => n13315, Z => n13310);
   U9499 : BUF_X1 port map( A => n13315, Z => n13311);
   U9500 : BUF_X1 port map( A => n13315, Z => n13308);
   U9501 : BUF_X1 port map( A => n13315, Z => n13309);
   U9502 : BUF_X1 port map( A => n13315, Z => n13312);
   U9503 : BUF_X1 port map( A => n13315, Z => n13313);
   U9504 : BUF_X1 port map( A => n13315, Z => n13314);
   U9505 : BUF_X1 port map( A => n12943, Z => n12935);
   U9506 : BUF_X1 port map( A => n12943, Z => n12936);
   U9507 : BUF_X1 port map( A => n12943, Z => n12937);
   U9508 : BUF_X1 port map( A => n12943, Z => n12938);
   U9509 : BUF_X1 port map( A => n12943, Z => n12939);
   U9510 : BUF_X1 port map( A => n12943, Z => n12940);
   U9511 : BUF_X1 port map( A => n12940, Z => n12941);
   U9512 : BUF_X1 port map( A => n12935, Z => n12942);
   U9513 : BUF_X1 port map( A => n11640, Z => n12817);
   U9514 : BUF_X1 port map( A => n11645, Z => n12805);
   U9515 : BUF_X1 port map( A => n11655, Z => n12781);
   U9516 : BUF_X1 port map( A => n11650, Z => n12793);
   U9517 : BUF_X1 port map( A => n11669, Z => n12757);
   U9518 : BUF_X1 port map( A => n11674, Z => n12745);
   U9519 : BUF_X1 port map( A => n11679, Z => n12733);
   U9520 : BUF_X1 port map( A => n11664, Z => n12769);
   U9521 : BUF_X1 port map( A => n11640, Z => n12818);
   U9522 : BUF_X1 port map( A => n11645, Z => n12806);
   U9523 : BUF_X1 port map( A => n11655, Z => n12782);
   U9524 : BUF_X1 port map( A => n11650, Z => n12794);
   U9525 : BUF_X1 port map( A => n11669, Z => n12758);
   U9526 : BUF_X1 port map( A => n11674, Z => n12746);
   U9527 : BUF_X1 port map( A => n11679, Z => n12734);
   U9528 : BUF_X1 port map( A => n11664, Z => n12770);
   U9529 : BUF_X1 port map( A => n10987, Z => n12919);
   U9530 : BUF_X1 port map( A => n10992, Z => n12907);
   U9531 : BUF_X1 port map( A => n11002, Z => n12883);
   U9532 : BUF_X1 port map( A => n10997, Z => n12895);
   U9533 : BUF_X1 port map( A => n11016, Z => n12859);
   U9534 : BUF_X1 port map( A => n11021, Z => n12847);
   U9535 : BUF_X1 port map( A => n11026, Z => n12835);
   U9536 : BUF_X1 port map( A => n11011, Z => n12871);
   U9537 : BUF_X1 port map( A => n10987, Z => n12920);
   U9538 : BUF_X1 port map( A => n10992, Z => n12908);
   U9539 : BUF_X1 port map( A => n11002, Z => n12884);
   U9540 : BUF_X1 port map( A => n10997, Z => n12896);
   U9541 : BUF_X1 port map( A => n11016, Z => n12860);
   U9542 : BUF_X1 port map( A => n11021, Z => n12848);
   U9543 : BUF_X1 port map( A => n11026, Z => n12836);
   U9544 : BUF_X1 port map( A => n11011, Z => n12872);
   U9545 : BUF_X1 port map( A => n11641, Z => n12814);
   U9546 : BUF_X1 port map( A => n11646, Z => n12802);
   U9547 : BUF_X1 port map( A => n11656, Z => n12778);
   U9548 : BUF_X1 port map( A => n11651, Z => n12790);
   U9549 : BUF_X1 port map( A => n11670, Z => n12754);
   U9550 : BUF_X1 port map( A => n11675, Z => n12742);
   U9551 : BUF_X1 port map( A => n11680, Z => n12730);
   U9552 : BUF_X1 port map( A => n11665, Z => n12766);
   U9553 : BUF_X1 port map( A => n11641, Z => n12815);
   U9554 : BUF_X1 port map( A => n11646, Z => n12803);
   U9555 : BUF_X1 port map( A => n11656, Z => n12779);
   U9556 : BUF_X1 port map( A => n11651, Z => n12791);
   U9557 : BUF_X1 port map( A => n11670, Z => n12755);
   U9558 : BUF_X1 port map( A => n11675, Z => n12743);
   U9559 : BUF_X1 port map( A => n11680, Z => n12731);
   U9560 : BUF_X1 port map( A => n11665, Z => n12767);
   U9561 : BUF_X1 port map( A => n10988, Z => n12916);
   U9562 : BUF_X1 port map( A => n10993, Z => n12904);
   U9563 : BUF_X1 port map( A => n11003, Z => n12880);
   U9564 : BUF_X1 port map( A => n10998, Z => n12892);
   U9565 : BUF_X1 port map( A => n11017, Z => n12856);
   U9566 : BUF_X1 port map( A => n11022, Z => n12844);
   U9567 : BUF_X1 port map( A => n11027, Z => n12832);
   U9568 : BUF_X1 port map( A => n11012, Z => n12868);
   U9569 : BUF_X1 port map( A => n10988, Z => n12917);
   U9570 : BUF_X1 port map( A => n10993, Z => n12905);
   U9571 : BUF_X1 port map( A => n11003, Z => n12881);
   U9572 : BUF_X1 port map( A => n10998, Z => n12893);
   U9573 : BUF_X1 port map( A => n11017, Z => n12857);
   U9574 : BUF_X1 port map( A => n11022, Z => n12845);
   U9575 : BUF_X1 port map( A => n11027, Z => n12833);
   U9576 : BUF_X1 port map( A => n11012, Z => n12869);
   U9577 : BUF_X1 port map( A => n11637, Z => n12823);
   U9578 : BUF_X1 port map( A => n11642, Z => n12811);
   U9579 : BUF_X1 port map( A => n11652, Z => n12787);
   U9580 : BUF_X1 port map( A => n11647, Z => n12799);
   U9581 : BUF_X1 port map( A => n11666, Z => n12763);
   U9582 : BUF_X1 port map( A => n11671, Z => n12751);
   U9583 : BUF_X1 port map( A => n11676, Z => n12739);
   U9584 : BUF_X1 port map( A => n11661, Z => n12775);
   U9585 : BUF_X1 port map( A => n11637, Z => n12824);
   U9586 : BUF_X1 port map( A => n11642, Z => n12812);
   U9587 : BUF_X1 port map( A => n11652, Z => n12788);
   U9588 : BUF_X1 port map( A => n11647, Z => n12800);
   U9589 : BUF_X1 port map( A => n11666, Z => n12764);
   U9590 : BUF_X1 port map( A => n11671, Z => n12752);
   U9591 : BUF_X1 port map( A => n11676, Z => n12740);
   U9592 : BUF_X1 port map( A => n11661, Z => n12776);
   U9593 : BUF_X1 port map( A => n10984, Z => n12925);
   U9594 : BUF_X1 port map( A => n10989, Z => n12913);
   U9595 : BUF_X1 port map( A => n10999, Z => n12889);
   U9596 : BUF_X1 port map( A => n10994, Z => n12901);
   U9597 : BUF_X1 port map( A => n11013, Z => n12865);
   U9598 : BUF_X1 port map( A => n11018, Z => n12853);
   U9599 : BUF_X1 port map( A => n11023, Z => n12841);
   U9600 : BUF_X1 port map( A => n11008, Z => n12877);
   U9601 : BUF_X1 port map( A => n10984, Z => n12926);
   U9602 : BUF_X1 port map( A => n10989, Z => n12914);
   U9603 : BUF_X1 port map( A => n10999, Z => n12890);
   U9604 : BUF_X1 port map( A => n10994, Z => n12902);
   U9605 : BUF_X1 port map( A => n11013, Z => n12866);
   U9606 : BUF_X1 port map( A => n11018, Z => n12854);
   U9607 : BUF_X1 port map( A => n11023, Z => n12842);
   U9608 : BUF_X1 port map( A => n11008, Z => n12878);
   U9609 : BUF_X1 port map( A => n11638, Z => n12820);
   U9610 : BUF_X1 port map( A => n11643, Z => n12808);
   U9611 : BUF_X1 port map( A => n11653, Z => n12784);
   U9612 : BUF_X1 port map( A => n11648, Z => n12796);
   U9613 : BUF_X1 port map( A => n11667, Z => n12760);
   U9614 : BUF_X1 port map( A => n11672, Z => n12748);
   U9615 : BUF_X1 port map( A => n11662, Z => n12772);
   U9616 : BUF_X1 port map( A => n11638, Z => n12821);
   U9617 : BUF_X1 port map( A => n11643, Z => n12809);
   U9618 : BUF_X1 port map( A => n11653, Z => n12785);
   U9619 : BUF_X1 port map( A => n11648, Z => n12797);
   U9620 : BUF_X1 port map( A => n11667, Z => n12761);
   U9621 : BUF_X1 port map( A => n11672, Z => n12749);
   U9622 : BUF_X1 port map( A => n11662, Z => n12773);
   U9623 : BUF_X1 port map( A => n10985, Z => n12922);
   U9624 : BUF_X1 port map( A => n10990, Z => n12910);
   U9625 : BUF_X1 port map( A => n11000, Z => n12886);
   U9626 : BUF_X1 port map( A => n10995, Z => n12898);
   U9627 : BUF_X1 port map( A => n11014, Z => n12862);
   U9628 : BUF_X1 port map( A => n11019, Z => n12850);
   U9629 : BUF_X1 port map( A => n11009, Z => n12874);
   U9630 : BUF_X1 port map( A => n10985, Z => n12923);
   U9631 : BUF_X1 port map( A => n10990, Z => n12911);
   U9632 : BUF_X1 port map( A => n11000, Z => n12887);
   U9633 : BUF_X1 port map( A => n10995, Z => n12899);
   U9634 : BUF_X1 port map( A => n11014, Z => n12863);
   U9635 : BUF_X1 port map( A => n11019, Z => n12851);
   U9636 : BUF_X1 port map( A => n11009, Z => n12875);
   U9637 : BUF_X1 port map( A => n11640, Z => n12819);
   U9638 : BUF_X1 port map( A => n11645, Z => n12807);
   U9639 : BUF_X1 port map( A => n11655, Z => n12783);
   U9640 : BUF_X1 port map( A => n11650, Z => n12795);
   U9641 : BUF_X1 port map( A => n11669, Z => n12759);
   U9642 : BUF_X1 port map( A => n11674, Z => n12747);
   U9643 : BUF_X1 port map( A => n11679, Z => n12735);
   U9644 : BUF_X1 port map( A => n11664, Z => n12771);
   U9645 : BUF_X1 port map( A => n10987, Z => n12921);
   U9646 : BUF_X1 port map( A => n10992, Z => n12909);
   U9647 : BUF_X1 port map( A => n11002, Z => n12885);
   U9648 : BUF_X1 port map( A => n10997, Z => n12897);
   U9649 : BUF_X1 port map( A => n11016, Z => n12861);
   U9650 : BUF_X1 port map( A => n11021, Z => n12849);
   U9651 : BUF_X1 port map( A => n11026, Z => n12837);
   U9652 : BUF_X1 port map( A => n11011, Z => n12873);
   U9653 : BUF_X1 port map( A => n11641, Z => n12816);
   U9654 : BUF_X1 port map( A => n11646, Z => n12804);
   U9655 : BUF_X1 port map( A => n11656, Z => n12780);
   U9656 : BUF_X1 port map( A => n11651, Z => n12792);
   U9657 : BUF_X1 port map( A => n11670, Z => n12756);
   U9658 : BUF_X1 port map( A => n11675, Z => n12744);
   U9659 : BUF_X1 port map( A => n11680, Z => n12732);
   U9660 : BUF_X1 port map( A => n11665, Z => n12768);
   U9661 : BUF_X1 port map( A => n10988, Z => n12918);
   U9662 : BUF_X1 port map( A => n10993, Z => n12906);
   U9663 : BUF_X1 port map( A => n11003, Z => n12882);
   U9664 : BUF_X1 port map( A => n10998, Z => n12894);
   U9665 : BUF_X1 port map( A => n11017, Z => n12858);
   U9666 : BUF_X1 port map( A => n11022, Z => n12846);
   U9667 : BUF_X1 port map( A => n11027, Z => n12834);
   U9668 : BUF_X1 port map( A => n11012, Z => n12870);
   U9669 : BUF_X1 port map( A => n11637, Z => n12825);
   U9670 : BUF_X1 port map( A => n11642, Z => n12813);
   U9671 : BUF_X1 port map( A => n11652, Z => n12789);
   U9672 : BUF_X1 port map( A => n11647, Z => n12801);
   U9673 : BUF_X1 port map( A => n11666, Z => n12765);
   U9674 : BUF_X1 port map( A => n11671, Z => n12753);
   U9675 : BUF_X1 port map( A => n11676, Z => n12741);
   U9676 : BUF_X1 port map( A => n11661, Z => n12777);
   U9677 : BUF_X1 port map( A => n10984, Z => n12927);
   U9678 : BUF_X1 port map( A => n10989, Z => n12915);
   U9679 : BUF_X1 port map( A => n10999, Z => n12891);
   U9680 : BUF_X1 port map( A => n10994, Z => n12903);
   U9681 : BUF_X1 port map( A => n11013, Z => n12867);
   U9682 : BUF_X1 port map( A => n11018, Z => n12855);
   U9683 : BUF_X1 port map( A => n11023, Z => n12843);
   U9684 : BUF_X1 port map( A => n11008, Z => n12879);
   U9685 : BUF_X1 port map( A => n11638, Z => n12822);
   U9686 : BUF_X1 port map( A => n11643, Z => n12810);
   U9687 : BUF_X1 port map( A => n11653, Z => n12786);
   U9688 : BUF_X1 port map( A => n11648, Z => n12798);
   U9689 : BUF_X1 port map( A => n11667, Z => n12762);
   U9690 : BUF_X1 port map( A => n11672, Z => n12750);
   U9691 : BUF_X1 port map( A => n11662, Z => n12774);
   U9692 : BUF_X1 port map( A => n10985, Z => n12924);
   U9693 : BUF_X1 port map( A => n10990, Z => n12912);
   U9694 : BUF_X1 port map( A => n11000, Z => n12888);
   U9695 : BUF_X1 port map( A => n10995, Z => n12900);
   U9696 : BUF_X1 port map( A => n11014, Z => n12864);
   U9697 : BUF_X1 port map( A => n11019, Z => n12852);
   U9698 : BUF_X1 port map( A => n11009, Z => n12876);
   U9699 : BUF_X1 port map( A => n13150, Z => n13143);
   U9700 : BUF_X1 port map( A => n13150, Z => n13144);
   U9701 : BUF_X1 port map( A => n13150, Z => n13145);
   U9702 : BUF_X1 port map( A => n13150, Z => n13146);
   U9703 : BUF_X1 port map( A => n13132, Z => n13125);
   U9704 : BUF_X1 port map( A => n13132, Z => n13126);
   U9705 : BUF_X1 port map( A => n13132, Z => n13127);
   U9706 : BUF_X1 port map( A => n13132, Z => n13128);
   U9707 : BUF_X1 port map( A => n13150, Z => n13147);
   U9708 : BUF_X1 port map( A => n13150, Z => n13148);
   U9709 : BUF_X1 port map( A => n13132, Z => n13129);
   U9710 : BUF_X1 port map( A => n13132, Z => n13130);
   U9711 : BUF_X1 port map( A => n13141, Z => n13134);
   U9712 : BUF_X1 port map( A => n13141, Z => n13135);
   U9713 : BUF_X1 port map( A => n13141, Z => n13136);
   U9714 : BUF_X1 port map( A => n13141, Z => n13137);
   U9715 : BUF_X1 port map( A => n13123, Z => n13116);
   U9716 : BUF_X1 port map( A => n13123, Z => n13117);
   U9717 : BUF_X1 port map( A => n13123, Z => n13118);
   U9718 : BUF_X1 port map( A => n13123, Z => n13119);
   U9719 : BUF_X1 port map( A => n13141, Z => n13138);
   U9720 : BUF_X1 port map( A => n13141, Z => n13139);
   U9721 : BUF_X1 port map( A => n13123, Z => n13120);
   U9722 : BUF_X1 port map( A => n13123, Z => n13121);
   U9723 : BUF_X1 port map( A => n13087, Z => n13080);
   U9724 : BUF_X1 port map( A => n13087, Z => n13081);
   U9725 : BUF_X1 port map( A => n13087, Z => n13082);
   U9726 : BUF_X1 port map( A => n13087, Z => n13083);
   U9727 : BUF_X1 port map( A => n13051, Z => n13044);
   U9728 : BUF_X1 port map( A => n13051, Z => n13045);
   U9729 : BUF_X1 port map( A => n13051, Z => n13046);
   U9730 : BUF_X1 port map( A => n13051, Z => n13047);
   U9731 : BUF_X1 port map( A => n13015, Z => n13008);
   U9732 : BUF_X1 port map( A => n13015, Z => n13009);
   U9733 : BUF_X1 port map( A => n13015, Z => n13010);
   U9734 : BUF_X1 port map( A => n13015, Z => n13011);
   U9735 : BUF_X1 port map( A => n12997, Z => n12990);
   U9736 : BUF_X1 port map( A => n12997, Z => n12991);
   U9737 : BUF_X1 port map( A => n12997, Z => n12992);
   U9738 : BUF_X1 port map( A => n12997, Z => n12993);
   U9739 : BUF_X1 port map( A => n12961, Z => n12954);
   U9740 : BUF_X1 port map( A => n12961, Z => n12955);
   U9741 : BUF_X1 port map( A => n12961, Z => n12956);
   U9742 : BUF_X1 port map( A => n12961, Z => n12957);
   U9743 : BUF_X1 port map( A => n13096, Z => n13089);
   U9744 : BUF_X1 port map( A => n13096, Z => n13090);
   U9745 : BUF_X1 port map( A => n13096, Z => n13091);
   U9746 : BUF_X1 port map( A => n13096, Z => n13092);
   U9747 : BUF_X1 port map( A => n13060, Z => n13053);
   U9748 : BUF_X1 port map( A => n13060, Z => n13054);
   U9749 : BUF_X1 port map( A => n13060, Z => n13055);
   U9750 : BUF_X1 port map( A => n13060, Z => n13056);
   U9751 : BUF_X1 port map( A => n13024, Z => n13017);
   U9752 : BUF_X1 port map( A => n13024, Z => n13018);
   U9753 : BUF_X1 port map( A => n13024, Z => n13019);
   U9754 : BUF_X1 port map( A => n13024, Z => n13020);
   U9755 : BUF_X1 port map( A => n13006, Z => n12999);
   U9756 : BUF_X1 port map( A => n13006, Z => n13000);
   U9757 : BUF_X1 port map( A => n13006, Z => n13001);
   U9758 : BUF_X1 port map( A => n13006, Z => n13002);
   U9759 : BUF_X1 port map( A => n12970, Z => n12963);
   U9760 : BUF_X1 port map( A => n12970, Z => n12964);
   U9761 : BUF_X1 port map( A => n12970, Z => n12965);
   U9762 : BUF_X1 port map( A => n12970, Z => n12966);
   U9763 : BUF_X1 port map( A => n13087, Z => n13084);
   U9764 : BUF_X1 port map( A => n13087, Z => n13085);
   U9765 : BUF_X1 port map( A => n13051, Z => n13048);
   U9766 : BUF_X1 port map( A => n13051, Z => n13049);
   U9767 : BUF_X1 port map( A => n13015, Z => n13012);
   U9768 : BUF_X1 port map( A => n13015, Z => n13013);
   U9769 : BUF_X1 port map( A => n12997, Z => n12994);
   U9770 : BUF_X1 port map( A => n12997, Z => n12995);
   U9771 : BUF_X1 port map( A => n12961, Z => n12958);
   U9772 : BUF_X1 port map( A => n12961, Z => n12959);
   U9773 : BUF_X1 port map( A => n13096, Z => n13093);
   U9774 : BUF_X1 port map( A => n13096, Z => n13094);
   U9775 : BUF_X1 port map( A => n13060, Z => n13057);
   U9776 : BUF_X1 port map( A => n13060, Z => n13058);
   U9777 : BUF_X1 port map( A => n13024, Z => n13021);
   U9778 : BUF_X1 port map( A => n13024, Z => n13022);
   U9779 : BUF_X1 port map( A => n13006, Z => n13003);
   U9780 : BUF_X1 port map( A => n13006, Z => n13004);
   U9781 : BUF_X1 port map( A => n12970, Z => n12967);
   U9782 : BUF_X1 port map( A => n12970, Z => n12968);
   U9783 : BUF_X1 port map( A => n13114, Z => n13107);
   U9784 : BUF_X1 port map( A => n13114, Z => n13108);
   U9785 : BUF_X1 port map( A => n13114, Z => n13109);
   U9786 : BUF_X1 port map( A => n13114, Z => n13110);
   U9787 : BUF_X1 port map( A => n13105, Z => n13098);
   U9788 : BUF_X1 port map( A => n13105, Z => n13099);
   U9789 : BUF_X1 port map( A => n13105, Z => n13100);
   U9790 : BUF_X1 port map( A => n13105, Z => n13101);
   U9791 : BUF_X1 port map( A => n13078, Z => n13071);
   U9792 : BUF_X1 port map( A => n13078, Z => n13072);
   U9793 : BUF_X1 port map( A => n13078, Z => n13073);
   U9794 : BUF_X1 port map( A => n13078, Z => n13074);
   U9795 : BUF_X1 port map( A => n13069, Z => n13062);
   U9796 : BUF_X1 port map( A => n13069, Z => n13063);
   U9797 : BUF_X1 port map( A => n13069, Z => n13064);
   U9798 : BUF_X1 port map( A => n13069, Z => n13065);
   U9799 : BUF_X1 port map( A => n13042, Z => n13035);
   U9800 : BUF_X1 port map( A => n13042, Z => n13036);
   U9801 : BUF_X1 port map( A => n13042, Z => n13037);
   U9802 : BUF_X1 port map( A => n13042, Z => n13038);
   U9803 : BUF_X1 port map( A => n13033, Z => n13026);
   U9804 : BUF_X1 port map( A => n13033, Z => n13027);
   U9805 : BUF_X1 port map( A => n13033, Z => n13028);
   U9806 : BUF_X1 port map( A => n13033, Z => n13029);
   U9807 : BUF_X1 port map( A => n12988, Z => n12981);
   U9808 : BUF_X1 port map( A => n12988, Z => n12982);
   U9809 : BUF_X1 port map( A => n12988, Z => n12983);
   U9810 : BUF_X1 port map( A => n12988, Z => n12984);
   U9811 : BUF_X1 port map( A => n12979, Z => n12972);
   U9812 : BUF_X1 port map( A => n12979, Z => n12973);
   U9813 : BUF_X1 port map( A => n12979, Z => n12974);
   U9814 : BUF_X1 port map( A => n12979, Z => n12975);
   U9815 : BUF_X1 port map( A => n12952, Z => n12945);
   U9816 : BUF_X1 port map( A => n12952, Z => n12946);
   U9817 : BUF_X1 port map( A => n12952, Z => n12947);
   U9818 : BUF_X1 port map( A => n12952, Z => n12948);
   U9819 : BUF_X1 port map( A => n13114, Z => n13111);
   U9820 : BUF_X1 port map( A => n13114, Z => n13112);
   U9821 : BUF_X1 port map( A => n13105, Z => n13102);
   U9822 : BUF_X1 port map( A => n13105, Z => n13103);
   U9823 : BUF_X1 port map( A => n13078, Z => n13075);
   U9824 : BUF_X1 port map( A => n13078, Z => n13076);
   U9825 : BUF_X1 port map( A => n13069, Z => n13066);
   U9826 : BUF_X1 port map( A => n13069, Z => n13067);
   U9827 : BUF_X1 port map( A => n13042, Z => n13039);
   U9828 : BUF_X1 port map( A => n13042, Z => n13040);
   U9829 : BUF_X1 port map( A => n13033, Z => n13030);
   U9830 : BUF_X1 port map( A => n13033, Z => n13031);
   U9831 : BUF_X1 port map( A => n12988, Z => n12985);
   U9832 : BUF_X1 port map( A => n12988, Z => n12986);
   U9833 : BUF_X1 port map( A => n12979, Z => n12976);
   U9834 : BUF_X1 port map( A => n12979, Z => n12977);
   U9835 : BUF_X1 port map( A => n12952, Z => n12949);
   U9836 : BUF_X1 port map( A => n12952, Z => n12950);
   U9837 : BUF_X1 port map( A => n13186, Z => n13179);
   U9838 : BUF_X1 port map( A => n13186, Z => n13180);
   U9839 : BUF_X1 port map( A => n13186, Z => n13181);
   U9840 : BUF_X1 port map( A => n13186, Z => n13182);
   U9841 : BUF_X1 port map( A => n13186, Z => n13183);
   U9842 : BUF_X1 port map( A => n13186, Z => n13184);
   U9843 : BUF_X1 port map( A => n13177, Z => n13170);
   U9844 : BUF_X1 port map( A => n13177, Z => n13171);
   U9845 : BUF_X1 port map( A => n13177, Z => n13172);
   U9846 : BUF_X1 port map( A => n13177, Z => n13173);
   U9847 : BUF_X1 port map( A => n13177, Z => n13174);
   U9848 : BUF_X1 port map( A => n13177, Z => n13175);
   U9849 : BUF_X1 port map( A => n13213, Z => n13210);
   U9850 : BUF_X1 port map( A => n13213, Z => n13211);
   U9851 : BUF_X1 port map( A => n13204, Z => n13197);
   U9852 : BUF_X1 port map( A => n13204, Z => n13198);
   U9853 : BUF_X1 port map( A => n13204, Z => n13199);
   U9854 : BUF_X1 port map( A => n13204, Z => n13200);
   U9855 : BUF_X1 port map( A => n13195, Z => n13188);
   U9856 : BUF_X1 port map( A => n13195, Z => n13189);
   U9857 : BUF_X1 port map( A => n13195, Z => n13190);
   U9858 : BUF_X1 port map( A => n13195, Z => n13191);
   U9859 : BUF_X1 port map( A => n13204, Z => n13201);
   U9860 : BUF_X1 port map( A => n13204, Z => n13202);
   U9861 : BUF_X1 port map( A => n13195, Z => n13192);
   U9862 : BUF_X1 port map( A => n13195, Z => n13193);
   U9863 : BUF_X1 port map( A => n13159, Z => n13152);
   U9864 : BUF_X1 port map( A => n13159, Z => n13153);
   U9865 : BUF_X1 port map( A => n13159, Z => n13154);
   U9866 : BUF_X1 port map( A => n13159, Z => n13155);
   U9867 : BUF_X1 port map( A => n13159, Z => n13156);
   U9868 : BUF_X1 port map( A => n13159, Z => n13157);
   U9869 : BUF_X1 port map( A => n13168, Z => n13161);
   U9870 : BUF_X1 port map( A => n13168, Z => n13162);
   U9871 : BUF_X1 port map( A => n13168, Z => n13163);
   U9872 : BUF_X1 port map( A => n13168, Z => n13164);
   U9873 : BUF_X1 port map( A => n13168, Z => n13165);
   U9874 : BUF_X1 port map( A => n13168, Z => n13166);
   U9875 : BUF_X1 port map( A => n13213, Z => n13206);
   U9876 : BUF_X1 port map( A => n13213, Z => n13207);
   U9877 : BUF_X1 port map( A => n13213, Z => n13208);
   U9878 : BUF_X1 port map( A => n13213, Z => n13209);
   U9879 : BUF_X1 port map( A => n13150, Z => n13149);
   U9880 : BUF_X1 port map( A => n13132, Z => n13131);
   U9881 : BUF_X1 port map( A => n13141, Z => n13140);
   U9882 : BUF_X1 port map( A => n13123, Z => n13122);
   U9883 : BUF_X1 port map( A => n13087, Z => n13086);
   U9884 : BUF_X1 port map( A => n13051, Z => n13050);
   U9885 : BUF_X1 port map( A => n13015, Z => n13014);
   U9886 : BUF_X1 port map( A => n12997, Z => n12996);
   U9887 : BUF_X1 port map( A => n12961, Z => n12960);
   U9888 : BUF_X1 port map( A => n13096, Z => n13095);
   U9889 : BUF_X1 port map( A => n13060, Z => n13059);
   U9890 : BUF_X1 port map( A => n13024, Z => n13023);
   U9891 : BUF_X1 port map( A => n13006, Z => n13005);
   U9892 : BUF_X1 port map( A => n12970, Z => n12969);
   U9893 : BUF_X1 port map( A => n13114, Z => n13113);
   U9894 : BUF_X1 port map( A => n13105, Z => n13104);
   U9895 : BUF_X1 port map( A => n13078, Z => n13077);
   U9896 : BUF_X1 port map( A => n13069, Z => n13068);
   U9897 : BUF_X1 port map( A => n13042, Z => n13041);
   U9898 : BUF_X1 port map( A => n13033, Z => n13032);
   U9899 : BUF_X1 port map( A => n12988, Z => n12987);
   U9900 : BUF_X1 port map( A => n12979, Z => n12978);
   U9901 : BUF_X1 port map( A => n12952, Z => n12951);
   U9902 : BUF_X1 port map( A => n13186, Z => n13185);
   U9903 : BUF_X1 port map( A => n13177, Z => n13176);
   U9904 : BUF_X1 port map( A => n13204, Z => n13203);
   U9905 : BUF_X1 port map( A => n13195, Z => n13194);
   U9906 : BUF_X1 port map( A => n13159, Z => n13158);
   U9907 : BUF_X1 port map( A => n13168, Z => n13167);
   U9908 : BUF_X1 port map( A => n13213, Z => n13212);
   U9909 : AND2_X1 port map( A1 => n12280, A2 => n12264, ZN => n11677);
   U9910 : AND2_X1 port map( A1 => n11627, A2 => n11611, ZN => n11024);
   U9911 : INV_X1 port map( A => n10900, ZN => n13315);
   U9912 : OAI21_X1 port map( B1 => n10932, B2 => n10933, A => n13321, ZN => 
                           n10900);
   U9913 : INV_X1 port map( A => n12934, ZN => n12943);
   U9914 : AOI221_X1 port map( B1 => n12823, B2 => n10322, C1 => n12820, C2 => 
                           n10346, A => n12258, ZN => n12257);
   U9915 : OAI22_X1 port map( A1 => n10706, A2 => n12817, B1 => n9963, B2 => 
                           n12814, ZN => n12258);
   U9916 : AOI221_X1 port map( B1 => n12823, B2 => n10321, C1 => n12820, C2 => 
                           n10345, A => n12239, ZN => n12238);
   U9917 : OAI22_X1 port map( A1 => n10354, A2 => n12817, B1 => n9962, B2 => 
                           n12814, ZN => n12239);
   U9918 : AOI221_X1 port map( B1 => n12823, B2 => n10320, C1 => n12820, C2 => 
                           n10344, A => n12220, ZN => n12219);
   U9919 : OAI22_X1 port map( A1 => n10353, A2 => n12817, B1 => n9961, B2 => 
                           n12814, ZN => n12220);
   U9920 : AOI221_X1 port map( B1 => n12823, B2 => n10319, C1 => n12820, C2 => 
                           n10343, A => n12201, ZN => n12200);
   U9921 : OAI22_X1 port map( A1 => n10352, A2 => n12817, B1 => n9960, B2 => 
                           n12814, ZN => n12201);
   U9922 : AOI221_X1 port map( B1 => n12823, B2 => n10318, C1 => n12820, C2 => 
                           n10342, A => n12182, ZN => n12181);
   U9923 : OAI22_X1 port map( A1 => n10351, A2 => n12817, B1 => n9959, B2 => 
                           n12814, ZN => n12182);
   U9924 : AOI221_X1 port map( B1 => n12823, B2 => n10317, C1 => n12820, C2 => 
                           n10341, A => n12163, ZN => n12162);
   U9925 : OAI22_X1 port map( A1 => n10350, A2 => n12817, B1 => n9958, B2 => 
                           n12814, ZN => n12163);
   U9926 : AOI221_X1 port map( B1 => n12823, B2 => n10316, C1 => n12820, C2 => 
                           n10340, A => n12144, ZN => n12143);
   U9927 : OAI22_X1 port map( A1 => n10349, A2 => n12817, B1 => n9957, B2 => 
                           n12814, ZN => n12144);
   U9928 : AOI221_X1 port map( B1 => n12823, B2 => n10315, C1 => n12820, C2 => 
                           n10339, A => n12125, ZN => n12124);
   U9929 : OAI22_X1 port map( A1 => n10348, A2 => n12817, B1 => n9956, B2 => 
                           n12814, ZN => n12125);
   U9930 : AOI221_X1 port map( B1 => n12823, B2 => n10314, C1 => n12820, C2 => 
                           n10338, A => n12106, ZN => n12105);
   U9931 : OAI22_X1 port map( A1 => n10705, A2 => n12817, B1 => n9955, B2 => 
                           n12814, ZN => n12106);
   U9932 : AOI221_X1 port map( B1 => n12823, B2 => n10313, C1 => n12820, C2 => 
                           n10337, A => n12087, ZN => n12086);
   U9933 : OAI22_X1 port map( A1 => n10704, A2 => n12817, B1 => n9954, B2 => 
                           n12814, ZN => n12087);
   U9934 : AOI221_X1 port map( B1 => n12823, B2 => n10312, C1 => n12820, C2 => 
                           n10336, A => n12068, ZN => n12067);
   U9935 : OAI22_X1 port map( A1 => n10703, A2 => n12817, B1 => n9953, B2 => 
                           n12814, ZN => n12068);
   U9936 : AOI221_X1 port map( B1 => n12823, B2 => n10311, C1 => n12820, C2 => 
                           n10335, A => n12049, ZN => n12048);
   U9937 : OAI22_X1 port map( A1 => n10702, A2 => n12817, B1 => n9952, B2 => 
                           n12814, ZN => n12049);
   U9938 : AOI221_X1 port map( B1 => n12824, B2 => n10310, C1 => n12821, C2 => 
                           n10334, A => n12030, ZN => n12029);
   U9939 : OAI22_X1 port map( A1 => n10701, A2 => n12818, B1 => n9951, B2 => 
                           n12815, ZN => n12030);
   U9940 : AOI221_X1 port map( B1 => n12824, B2 => n10309, C1 => n12821, C2 => 
                           n10333, A => n12011, ZN => n12010);
   U9941 : OAI22_X1 port map( A1 => n10700, A2 => n12818, B1 => n9950, B2 => 
                           n12815, ZN => n12011);
   U9942 : AOI221_X1 port map( B1 => n12824, B2 => n10308, C1 => n12821, C2 => 
                           n10332, A => n11992, ZN => n11991);
   U9943 : OAI22_X1 port map( A1 => n10699, A2 => n12818, B1 => n9949, B2 => 
                           n12815, ZN => n11992);
   U9944 : AOI221_X1 port map( B1 => n12824, B2 => n10307, C1 => n12821, C2 => 
                           n10331, A => n11973, ZN => n11972);
   U9945 : OAI22_X1 port map( A1 => n10698, A2 => n12818, B1 => n9948, B2 => 
                           n12815, ZN => n11973);
   U9946 : AOI221_X1 port map( B1 => n12824, B2 => n10306, C1 => n12821, C2 => 
                           n10330, A => n11954, ZN => n11953);
   U9947 : OAI22_X1 port map( A1 => n10697, A2 => n12818, B1 => n9947, B2 => 
                           n12815, ZN => n11954);
   U9948 : AOI221_X1 port map( B1 => n12824, B2 => n10305, C1 => n12821, C2 => 
                           n10329, A => n11935, ZN => n11934);
   U9949 : OAI22_X1 port map( A1 => n10696, A2 => n12818, B1 => n9946, B2 => 
                           n12815, ZN => n11935);
   U9950 : AOI221_X1 port map( B1 => n12824, B2 => n10304, C1 => n12821, C2 => 
                           n10328, A => n11916, ZN => n11915);
   U9951 : OAI22_X1 port map( A1 => n10695, A2 => n12818, B1 => n9945, B2 => 
                           n12815, ZN => n11916);
   U9952 : AOI221_X1 port map( B1 => n12824, B2 => n10303, C1 => n12821, C2 => 
                           n10327, A => n11897, ZN => n11896);
   U9953 : OAI22_X1 port map( A1 => n10694, A2 => n12818, B1 => n9944, B2 => 
                           n12815, ZN => n11897);
   U9954 : AOI221_X1 port map( B1 => n12824, B2 => n10302, C1 => n12821, C2 => 
                           n10326, A => n11878, ZN => n11877);
   U9955 : OAI22_X1 port map( A1 => n10573, A2 => n12818, B1 => n10446, B2 => 
                           n12815, ZN => n11878);
   U9956 : AOI221_X1 port map( B1 => n12824, B2 => n10301, C1 => n12821, C2 => 
                           n10325, A => n11859, ZN => n11858);
   U9957 : OAI22_X1 port map( A1 => n10572, A2 => n12818, B1 => n10445, B2 => 
                           n12815, ZN => n11859);
   U9958 : AOI221_X1 port map( B1 => n12824, B2 => n10300, C1 => n12821, C2 => 
                           n10324, A => n11840, ZN => n11839);
   U9959 : OAI22_X1 port map( A1 => n10571, A2 => n12818, B1 => n10444, B2 => 
                           n12815, ZN => n11840);
   U9960 : AOI221_X1 port map( B1 => n12824, B2 => n10299, C1 => n12821, C2 => 
                           n10323, A => n11821, ZN => n11820);
   U9961 : OAI22_X1 port map( A1 => n9943, A2 => n12818, B1 => n10443, B2 => 
                           n12815, ZN => n11821);
   U9962 : AOI221_X1 port map( B1 => n12925, B2 => n10322, C1 => n12922, C2 => 
                           n10346, A => n11605, ZN => n11604);
   U9963 : OAI22_X1 port map( A1 => n10706, A2 => n12919, B1 => n9963, B2 => 
                           n12916, ZN => n11605);
   U9964 : AOI221_X1 port map( B1 => n12925, B2 => n10321, C1 => n12922, C2 => 
                           n10345, A => n11586, ZN => n11585);
   U9965 : OAI22_X1 port map( A1 => n10354, A2 => n12919, B1 => n9962, B2 => 
                           n12916, ZN => n11586);
   U9966 : AOI221_X1 port map( B1 => n12925, B2 => n10320, C1 => n12922, C2 => 
                           n10344, A => n11567, ZN => n11566);
   U9967 : OAI22_X1 port map( A1 => n10353, A2 => n12919, B1 => n9961, B2 => 
                           n12916, ZN => n11567);
   U9968 : AOI221_X1 port map( B1 => n12925, B2 => n10319, C1 => n12922, C2 => 
                           n10343, A => n11548, ZN => n11547);
   U9969 : OAI22_X1 port map( A1 => n10352, A2 => n12919, B1 => n9960, B2 => 
                           n12916, ZN => n11548);
   U9970 : AOI221_X1 port map( B1 => n12925, B2 => n10318, C1 => n12922, C2 => 
                           n10342, A => n11529, ZN => n11528);
   U9971 : OAI22_X1 port map( A1 => n10351, A2 => n12919, B1 => n9959, B2 => 
                           n12916, ZN => n11529);
   U9972 : AOI221_X1 port map( B1 => n12925, B2 => n10317, C1 => n12922, C2 => 
                           n10341, A => n11510, ZN => n11509);
   U9973 : OAI22_X1 port map( A1 => n10350, A2 => n12919, B1 => n9958, B2 => 
                           n12916, ZN => n11510);
   U9974 : AOI221_X1 port map( B1 => n12925, B2 => n10316, C1 => n12922, C2 => 
                           n10340, A => n11491, ZN => n11490);
   U9975 : OAI22_X1 port map( A1 => n10349, A2 => n12919, B1 => n9957, B2 => 
                           n12916, ZN => n11491);
   U9976 : AOI221_X1 port map( B1 => n12925, B2 => n10315, C1 => n12922, C2 => 
                           n10339, A => n11472, ZN => n11471);
   U9977 : OAI22_X1 port map( A1 => n10348, A2 => n12919, B1 => n9956, B2 => 
                           n12916, ZN => n11472);
   U9978 : AOI221_X1 port map( B1 => n12925, B2 => n10314, C1 => n12922, C2 => 
                           n10338, A => n11453, ZN => n11452);
   U9979 : OAI22_X1 port map( A1 => n10705, A2 => n12919, B1 => n9955, B2 => 
                           n12916, ZN => n11453);
   U9980 : AOI221_X1 port map( B1 => n12925, B2 => n10313, C1 => n12922, C2 => 
                           n10337, A => n11434, ZN => n11433);
   U9981 : OAI22_X1 port map( A1 => n10704, A2 => n12919, B1 => n9954, B2 => 
                           n12916, ZN => n11434);
   U9982 : AOI221_X1 port map( B1 => n12925, B2 => n10312, C1 => n12922, C2 => 
                           n10336, A => n11415, ZN => n11414);
   U9983 : OAI22_X1 port map( A1 => n10703, A2 => n12919, B1 => n9953, B2 => 
                           n12916, ZN => n11415);
   U9984 : AOI221_X1 port map( B1 => n12925, B2 => n10311, C1 => n12922, C2 => 
                           n10335, A => n11396, ZN => n11395);
   U9985 : OAI22_X1 port map( A1 => n10702, A2 => n12919, B1 => n9952, B2 => 
                           n12916, ZN => n11396);
   U9986 : AOI221_X1 port map( B1 => n12926, B2 => n10310, C1 => n12923, C2 => 
                           n10334, A => n11377, ZN => n11376);
   U9987 : OAI22_X1 port map( A1 => n10701, A2 => n12920, B1 => n9951, B2 => 
                           n12917, ZN => n11377);
   U9988 : AOI221_X1 port map( B1 => n12926, B2 => n10309, C1 => n12923, C2 => 
                           n10333, A => n11358, ZN => n11357);
   U9989 : OAI22_X1 port map( A1 => n10700, A2 => n12920, B1 => n9950, B2 => 
                           n12917, ZN => n11358);
   U9990 : AOI221_X1 port map( B1 => n12926, B2 => n10308, C1 => n12923, C2 => 
                           n10332, A => n11339, ZN => n11338);
   U9991 : OAI22_X1 port map( A1 => n10699, A2 => n12920, B1 => n9949, B2 => 
                           n12917, ZN => n11339);
   U9992 : AOI221_X1 port map( B1 => n12926, B2 => n10307, C1 => n12923, C2 => 
                           n10331, A => n11320, ZN => n11319);
   U9993 : OAI22_X1 port map( A1 => n10698, A2 => n12920, B1 => n9948, B2 => 
                           n12917, ZN => n11320);
   U9994 : AOI221_X1 port map( B1 => n12926, B2 => n10306, C1 => n12923, C2 => 
                           n10330, A => n11301, ZN => n11300);
   U9995 : OAI22_X1 port map( A1 => n10697, A2 => n12920, B1 => n9947, B2 => 
                           n12917, ZN => n11301);
   U9996 : AOI221_X1 port map( B1 => n12926, B2 => n10305, C1 => n12923, C2 => 
                           n10329, A => n11282, ZN => n11281);
   U9997 : OAI22_X1 port map( A1 => n10696, A2 => n12920, B1 => n9946, B2 => 
                           n12917, ZN => n11282);
   U9998 : AOI221_X1 port map( B1 => n12926, B2 => n10304, C1 => n12923, C2 => 
                           n10328, A => n11263, ZN => n11262);
   U9999 : OAI22_X1 port map( A1 => n10695, A2 => n12920, B1 => n9945, B2 => 
                           n12917, ZN => n11263);
   U10000 : AOI221_X1 port map( B1 => n12926, B2 => n10303, C1 => n12923, C2 =>
                           n10327, A => n11244, ZN => n11243);
   U10001 : OAI22_X1 port map( A1 => n10694, A2 => n12920, B1 => n9944, B2 => 
                           n12917, ZN => n11244);
   U10002 : AOI221_X1 port map( B1 => n12926, B2 => n10302, C1 => n12923, C2 =>
                           n10326, A => n11225, ZN => n11224);
   U10003 : OAI22_X1 port map( A1 => n10573, A2 => n12920, B1 => n10446, B2 => 
                           n12917, ZN => n11225);
   U10004 : AOI221_X1 port map( B1 => n12926, B2 => n10301, C1 => n12923, C2 =>
                           n10325, A => n11206, ZN => n11205);
   U10005 : OAI22_X1 port map( A1 => n10572, A2 => n12920, B1 => n10445, B2 => 
                           n12917, ZN => n11206);
   U10006 : AOI221_X1 port map( B1 => n12926, B2 => n10300, C1 => n12923, C2 =>
                           n10324, A => n11187, ZN => n11186);
   U10007 : OAI22_X1 port map( A1 => n10571, A2 => n12920, B1 => n10444, B2 => 
                           n12917, ZN => n11187);
   U10008 : AOI221_X1 port map( B1 => n12926, B2 => n10299, C1 => n12923, C2 =>
                           n10323, A => n11168, ZN => n11167);
   U10009 : OAI22_X1 port map( A1 => n9943, A2 => n12920, B1 => n10443, B2 => 
                           n12917, ZN => n11168);
   U10010 : AOI221_X1 port map( B1 => n12927, B2 => n10122, C1 => n12924, C2 =>
                           n10130, A => n11149, ZN => n11148);
   U10011 : OAI22_X1 port map( A1 => n9942, A2 => n12921, B1 => n10402, B2 => 
                           n12918, ZN => n11149);
   U10012 : AOI221_X1 port map( B1 => n12927, B2 => n10121, C1 => n12924, C2 =>
                           n10129, A => n11130, ZN => n11129);
   U10013 : OAI22_X1 port map( A1 => n9941, A2 => n12921, B1 => n10401, B2 => 
                           n12918, ZN => n11130);
   U10014 : AOI221_X1 port map( B1 => n12927, B2 => n10120, C1 => n12924, C2 =>
                           n10128, A => n11111, ZN => n11110);
   U10015 : OAI22_X1 port map( A1 => n9940, A2 => n12921, B1 => n10400, B2 => 
                           n12918, ZN => n11111);
   U10016 : AOI221_X1 port map( B1 => n12927, B2 => n10119, C1 => n12924, C2 =>
                           n10127, A => n11092, ZN => n11091);
   U10017 : OAI22_X1 port map( A1 => n9939, A2 => n12921, B1 => n10399, B2 => 
                           n12918, ZN => n11092);
   U10018 : AOI221_X1 port map( B1 => n12927, B2 => n10118, C1 => n12924, C2 =>
                           n10126, A => n11073, ZN => n11072);
   U10019 : OAI22_X1 port map( A1 => n10570, A2 => n12921, B1 => n10398, B2 => 
                           n12918, ZN => n11073);
   U10020 : AOI221_X1 port map( B1 => n12927, B2 => n10117, C1 => n12924, C2 =>
                           n10125, A => n11054, ZN => n11053);
   U10021 : OAI22_X1 port map( A1 => n10569, A2 => n12921, B1 => n10397, B2 => 
                           n12918, ZN => n11054);
   U10022 : AOI221_X1 port map( B1 => n12927, B2 => n10116, C1 => n12924, C2 =>
                           n10124, A => n11035, ZN => n11034);
   U10023 : OAI22_X1 port map( A1 => n10568, A2 => n12921, B1 => n10396, B2 => 
                           n12918, ZN => n11035);
   U10024 : AOI221_X1 port map( B1 => n12927, B2 => n10115, C1 => n12924, C2 =>
                           n10123, A => n10986, ZN => n10983);
   U10025 : OAI22_X1 port map( A1 => n10567, A2 => n12921, B1 => n10395, B2 => 
                           n12918, ZN => n10986);
   U10026 : AOI221_X1 port map( B1 => n12811, B2 => n10898, C1 => n12808, C2 =>
                           n10866, A => n12263, ZN => n12256);
   U10027 : OAI22_X1 port map( A1 => n10026, A2 => n12805, B1 => n9994, B2 => 
                           n12802, ZN => n12263);
   U10028 : AOI221_X1 port map( B1 => n12763, B2 => n10250, C1 => n12760, C2 =>
                           n10226, A => n12277, ZN => n12272);
   U10029 : OAI22_X1 port map( A1 => n10645, A2 => n12757, B1 => n10518, B2 => 
                           n12754, ZN => n12277);
   U10030 : AOI221_X1 port map( B1 => n12811, B2 => n10897, C1 => n12808, C2 =>
                           n10865, A => n12240, ZN => n12237);
   U10031 : OAI22_X1 port map( A1 => n10025, A2 => n12805, B1 => n9993, B2 => 
                           n12802, ZN => n12240);
   U10032 : AOI221_X1 port map( B1 => n12763, B2 => n10249, C1 => n12760, C2 =>
                           n10225, A => n12248, ZN => n12245);
   U10033 : OAI22_X1 port map( A1 => n10644, A2 => n12757, B1 => n10517, B2 => 
                           n12754, ZN => n12248);
   U10034 : AOI221_X1 port map( B1 => n12811, B2 => n10896, C1 => n12808, C2 =>
                           n10864, A => n12221, ZN => n12218);
   U10035 : OAI22_X1 port map( A1 => n10024, A2 => n12805, B1 => n9992, B2 => 
                           n12802, ZN => n12221);
   U10036 : AOI221_X1 port map( B1 => n12763, B2 => n10248, C1 => n12760, C2 =>
                           n10224, A => n12229, ZN => n12226);
   U10037 : OAI22_X1 port map( A1 => n10643, A2 => n12757, B1 => n10516, B2 => 
                           n12754, ZN => n12229);
   U10038 : AOI221_X1 port map( B1 => n12811, B2 => n10895, C1 => n12808, C2 =>
                           n10863, A => n12202, ZN => n12199);
   U10039 : OAI22_X1 port map( A1 => n10023, A2 => n12805, B1 => n9991, B2 => 
                           n12802, ZN => n12202);
   U10040 : AOI221_X1 port map( B1 => n12763, B2 => n10247, C1 => n12760, C2 =>
                           n10223, A => n12210, ZN => n12207);
   U10041 : OAI22_X1 port map( A1 => n10642, A2 => n12757, B1 => n10515, B2 => 
                           n12754, ZN => n12210);
   U10042 : AOI221_X1 port map( B1 => n12811, B2 => n10894, C1 => n12808, C2 =>
                           n10862, A => n12183, ZN => n12180);
   U10043 : OAI22_X1 port map( A1 => n10022, A2 => n12805, B1 => n9990, B2 => 
                           n12802, ZN => n12183);
   U10044 : AOI221_X1 port map( B1 => n12763, B2 => n10246, C1 => n12760, C2 =>
                           n10222, A => n12191, ZN => n12188);
   U10045 : OAI22_X1 port map( A1 => n10641, A2 => n12757, B1 => n10514, B2 => 
                           n12754, ZN => n12191);
   U10046 : AOI221_X1 port map( B1 => n12811, B2 => n10893, C1 => n12808, C2 =>
                           n10861, A => n12164, ZN => n12161);
   U10047 : OAI22_X1 port map( A1 => n10021, A2 => n12805, B1 => n9989, B2 => 
                           n12802, ZN => n12164);
   U10048 : AOI221_X1 port map( B1 => n12763, B2 => n10245, C1 => n12760, C2 =>
                           n10221, A => n12172, ZN => n12169);
   U10049 : OAI22_X1 port map( A1 => n10640, A2 => n12757, B1 => n10513, B2 => 
                           n12754, ZN => n12172);
   U10050 : AOI221_X1 port map( B1 => n12811, B2 => n10892, C1 => n12808, C2 =>
                           n10860, A => n12145, ZN => n12142);
   U10051 : OAI22_X1 port map( A1 => n10020, A2 => n12805, B1 => n9988, B2 => 
                           n12802, ZN => n12145);
   U10052 : AOI221_X1 port map( B1 => n12763, B2 => n10244, C1 => n12760, C2 =>
                           n10220, A => n12153, ZN => n12150);
   U10053 : OAI22_X1 port map( A1 => n10639, A2 => n12757, B1 => n10512, B2 => 
                           n12754, ZN => n12153);
   U10054 : AOI221_X1 port map( B1 => n12811, B2 => n10891, C1 => n12808, C2 =>
                           n10859, A => n12126, ZN => n12123);
   U10055 : OAI22_X1 port map( A1 => n10019, A2 => n12805, B1 => n9987, B2 => 
                           n12802, ZN => n12126);
   U10056 : AOI221_X1 port map( B1 => n12763, B2 => n10243, C1 => n12760, C2 =>
                           n10219, A => n12134, ZN => n12131);
   U10057 : OAI22_X1 port map( A1 => n10638, A2 => n12757, B1 => n10511, B2 => 
                           n12754, ZN => n12134);
   U10058 : AOI221_X1 port map( B1 => n12811, B2 => n10890, C1 => n12808, C2 =>
                           n10858, A => n12107, ZN => n12104);
   U10059 : OAI22_X1 port map( A1 => n10018, A2 => n12805, B1 => n9986, B2 => 
                           n12802, ZN => n12107);
   U10060 : AOI221_X1 port map( B1 => n12763, B2 => n10242, C1 => n12760, C2 =>
                           n10218, A => n12115, ZN => n12112);
   U10061 : OAI22_X1 port map( A1 => n10637, A2 => n12757, B1 => n10510, B2 => 
                           n12754, ZN => n12115);
   U10062 : AOI221_X1 port map( B1 => n12811, B2 => n10889, C1 => n12808, C2 =>
                           n10857, A => n12088, ZN => n12085);
   U10063 : OAI22_X1 port map( A1 => n10017, A2 => n12805, B1 => n9985, B2 => 
                           n12802, ZN => n12088);
   U10064 : AOI221_X1 port map( B1 => n12763, B2 => n10241, C1 => n12760, C2 =>
                           n10217, A => n12096, ZN => n12093);
   U10065 : OAI22_X1 port map( A1 => n10636, A2 => n12757, B1 => n10509, B2 => 
                           n12754, ZN => n12096);
   U10066 : AOI221_X1 port map( B1 => n12811, B2 => n10888, C1 => n12808, C2 =>
                           n10856, A => n12069, ZN => n12066);
   U10067 : OAI22_X1 port map( A1 => n10016, A2 => n12805, B1 => n9984, B2 => 
                           n12802, ZN => n12069);
   U10068 : AOI221_X1 port map( B1 => n12763, B2 => n10240, C1 => n12760, C2 =>
                           n10216, A => n12077, ZN => n12074);
   U10069 : OAI22_X1 port map( A1 => n10635, A2 => n12757, B1 => n10508, B2 => 
                           n12754, ZN => n12077);
   U10070 : AOI221_X1 port map( B1 => n12811, B2 => n10887, C1 => n12808, C2 =>
                           n10855, A => n12050, ZN => n12047);
   U10071 : OAI22_X1 port map( A1 => n10015, A2 => n12805, B1 => n9983, B2 => 
                           n12802, ZN => n12050);
   U10072 : AOI221_X1 port map( B1 => n12763, B2 => n10239, C1 => n12760, C2 =>
                           n10215, A => n12058, ZN => n12055);
   U10073 : OAI22_X1 port map( A1 => n10634, A2 => n12757, B1 => n10507, B2 => 
                           n12754, ZN => n12058);
   U10074 : AOI221_X1 port map( B1 => n12812, B2 => n10886, C1 => n12809, C2 =>
                           n10854, A => n12031, ZN => n12028);
   U10075 : OAI22_X1 port map( A1 => n10014, A2 => n12806, B1 => n9982, B2 => 
                           n12803, ZN => n12031);
   U10076 : AOI221_X1 port map( B1 => n12764, B2 => n10238, C1 => n12761, C2 =>
                           n10214, A => n12039, ZN => n12036);
   U10077 : OAI22_X1 port map( A1 => n10633, A2 => n12758, B1 => n10506, B2 => 
                           n12755, ZN => n12039);
   U10078 : AOI221_X1 port map( B1 => n12812, B2 => n10885, C1 => n12809, C2 =>
                           n10853, A => n12012, ZN => n12009);
   U10079 : OAI22_X1 port map( A1 => n10013, A2 => n12806, B1 => n9981, B2 => 
                           n12803, ZN => n12012);
   U10080 : AOI221_X1 port map( B1 => n12764, B2 => n10237, C1 => n12761, C2 =>
                           n10213, A => n12020, ZN => n12017);
   U10081 : OAI22_X1 port map( A1 => n10632, A2 => n12758, B1 => n10505, B2 => 
                           n12755, ZN => n12020);
   U10082 : AOI221_X1 port map( B1 => n12812, B2 => n10884, C1 => n12809, C2 =>
                           n10852, A => n11993, ZN => n11990);
   U10083 : OAI22_X1 port map( A1 => n10012, A2 => n12806, B1 => n9980, B2 => 
                           n12803, ZN => n11993);
   U10084 : AOI221_X1 port map( B1 => n12764, B2 => n10236, C1 => n12761, C2 =>
                           n10212, A => n12001, ZN => n11998);
   U10085 : OAI22_X1 port map( A1 => n10631, A2 => n12758, B1 => n10504, B2 => 
                           n12755, ZN => n12001);
   U10086 : AOI221_X1 port map( B1 => n12812, B2 => n10883, C1 => n12809, C2 =>
                           n10851, A => n11974, ZN => n11971);
   U10087 : OAI22_X1 port map( A1 => n10011, A2 => n12806, B1 => n9979, B2 => 
                           n12803, ZN => n11974);
   U10088 : AOI221_X1 port map( B1 => n12764, B2 => n10235, C1 => n12761, C2 =>
                           n10211, A => n11982, ZN => n11979);
   U10089 : OAI22_X1 port map( A1 => n10630, A2 => n12758, B1 => n10503, B2 => 
                           n12755, ZN => n11982);
   U10090 : AOI221_X1 port map( B1 => n12812, B2 => n10882, C1 => n12809, C2 =>
                           n10850, A => n11955, ZN => n11952);
   U10091 : OAI22_X1 port map( A1 => n10010, A2 => n12806, B1 => n9978, B2 => 
                           n12803, ZN => n11955);
   U10092 : AOI221_X1 port map( B1 => n12764, B2 => n10234, C1 => n12761, C2 =>
                           n10210, A => n11963, ZN => n11960);
   U10093 : OAI22_X1 port map( A1 => n10629, A2 => n12758, B1 => n10502, B2 => 
                           n12755, ZN => n11963);
   U10094 : AOI221_X1 port map( B1 => n12812, B2 => n10881, C1 => n12809, C2 =>
                           n10849, A => n11936, ZN => n11933);
   U10095 : OAI22_X1 port map( A1 => n10009, A2 => n12806, B1 => n9977, B2 => 
                           n12803, ZN => n11936);
   U10096 : AOI221_X1 port map( B1 => n12764, B2 => n10233, C1 => n12761, C2 =>
                           n10209, A => n11944, ZN => n11941);
   U10097 : OAI22_X1 port map( A1 => n10628, A2 => n12758, B1 => n10501, B2 => 
                           n12755, ZN => n11944);
   U10098 : AOI221_X1 port map( B1 => n12812, B2 => n10880, C1 => n12809, C2 =>
                           n10848, A => n11917, ZN => n11914);
   U10099 : OAI22_X1 port map( A1 => n10008, A2 => n12806, B1 => n9976, B2 => 
                           n12803, ZN => n11917);
   U10100 : AOI221_X1 port map( B1 => n12764, B2 => n10232, C1 => n12761, C2 =>
                           n10208, A => n11925, ZN => n11922);
   U10101 : OAI22_X1 port map( A1 => n10627, A2 => n12758, B1 => n10500, B2 => 
                           n12755, ZN => n11925);
   U10102 : AOI221_X1 port map( B1 => n12812, B2 => n10879, C1 => n12809, C2 =>
                           n10847, A => n11898, ZN => n11895);
   U10103 : OAI22_X1 port map( A1 => n10007, A2 => n12806, B1 => n9975, B2 => 
                           n12803, ZN => n11898);
   U10104 : AOI221_X1 port map( B1 => n12764, B2 => n10231, C1 => n12761, C2 =>
                           n10207, A => n11906, ZN => n11903);
   U10105 : OAI22_X1 port map( A1 => n10626, A2 => n12758, B1 => n10499, B2 => 
                           n12755, ZN => n11906);
   U10106 : AOI221_X1 port map( B1 => n12812, B2 => n10878, C1 => n12809, C2 =>
                           n10846, A => n11879, ZN => n11876);
   U10107 : OAI22_X1 port map( A1 => n10006, A2 => n12806, B1 => n9974, B2 => 
                           n12803, ZN => n11879);
   U10108 : AOI221_X1 port map( B1 => n12764, B2 => n10230, C1 => n12761, C2 =>
                           n10206, A => n11887, ZN => n11884);
   U10109 : OAI22_X1 port map( A1 => n10625, A2 => n12758, B1 => n10498, B2 => 
                           n12755, ZN => n11887);
   U10110 : AOI221_X1 port map( B1 => n12812, B2 => n10877, C1 => n12809, C2 =>
                           n10845, A => n11860, ZN => n11857);
   U10111 : OAI22_X1 port map( A1 => n10005, A2 => n12806, B1 => n9973, B2 => 
                           n12803, ZN => n11860);
   U10112 : AOI221_X1 port map( B1 => n12764, B2 => n10229, C1 => n12761, C2 =>
                           n10205, A => n11868, ZN => n11865);
   U10113 : OAI22_X1 port map( A1 => n10624, A2 => n12758, B1 => n10497, B2 => 
                           n12755, ZN => n11868);
   U10114 : AOI221_X1 port map( B1 => n12812, B2 => n10876, C1 => n12809, C2 =>
                           n10844, A => n11841, ZN => n11838);
   U10115 : OAI22_X1 port map( A1 => n10004, A2 => n12806, B1 => n9972, B2 => 
                           n12803, ZN => n11841);
   U10116 : AOI221_X1 port map( B1 => n12764, B2 => n10228, C1 => n12761, C2 =>
                           n10204, A => n11849, ZN => n11846);
   U10117 : OAI22_X1 port map( A1 => n10623, A2 => n12758, B1 => n10496, B2 => 
                           n12755, ZN => n11849);
   U10118 : AOI221_X1 port map( B1 => n12812, B2 => n10875, C1 => n12809, C2 =>
                           n10843, A => n11822, ZN => n11819);
   U10119 : OAI22_X1 port map( A1 => n10003, A2 => n12806, B1 => n9971, B2 => 
                           n12803, ZN => n11822);
   U10120 : AOI221_X1 port map( B1 => n12764, B2 => n10227, C1 => n12761, C2 =>
                           n10203, A => n11830, ZN => n11827);
   U10121 : OAI22_X1 port map( A1 => n10622, A2 => n12758, B1 => n10495, B2 => 
                           n12755, ZN => n11830);
   U10122 : AOI221_X1 port map( B1 => n12765, B2 => n10098, C1 => n12762, C2 =>
                           n10090, A => n11811, ZN => n11808);
   U10123 : OAI22_X1 port map( A1 => n10426, A2 => n12759, B1 => n10378, B2 => 
                           n12756, ZN => n11811);
   U10124 : AOI221_X1 port map( B1 => n12765, B2 => n10097, C1 => n12762, C2 =>
                           n10089, A => n11792, ZN => n11789);
   U10125 : OAI22_X1 port map( A1 => n10425, A2 => n12759, B1 => n10377, B2 => 
                           n12756, ZN => n11792);
   U10126 : AOI221_X1 port map( B1 => n12765, B2 => n10096, C1 => n12762, C2 =>
                           n10088, A => n11773, ZN => n11770);
   U10127 : OAI22_X1 port map( A1 => n10424, A2 => n12759, B1 => n10376, B2 => 
                           n12756, ZN => n11773);
   U10128 : AOI221_X1 port map( B1 => n12765, B2 => n10095, C1 => n12762, C2 =>
                           n10087, A => n11754, ZN => n11751);
   U10129 : OAI22_X1 port map( A1 => n10423, A2 => n12759, B1 => n10375, B2 => 
                           n12756, ZN => n11754);
   U10130 : AOI221_X1 port map( B1 => n12765, B2 => n10094, C1 => n12762, C2 =>
                           n10086, A => n11735, ZN => n11732);
   U10131 : OAI22_X1 port map( A1 => n10422, A2 => n12759, B1 => n10374, B2 => 
                           n12756, ZN => n11735);
   U10132 : AOI221_X1 port map( B1 => n12765, B2 => n10093, C1 => n12762, C2 =>
                           n10085, A => n11716, ZN => n11713);
   U10133 : OAI22_X1 port map( A1 => n10421, A2 => n12759, B1 => n10373, B2 => 
                           n12756, ZN => n11716);
   U10134 : AOI221_X1 port map( B1 => n12765, B2 => n10092, C1 => n12762, C2 =>
                           n10084, A => n11697, ZN => n11694);
   U10135 : OAI22_X1 port map( A1 => n10420, A2 => n12759, B1 => n10372, B2 => 
                           n12756, ZN => n11697);
   U10136 : AOI221_X1 port map( B1 => n12765, B2 => n10091, C1 => n12762, C2 =>
                           n10083, A => n11668, ZN => n11659);
   U10137 : OAI22_X1 port map( A1 => n10419, A2 => n12759, B1 => n10371, B2 => 
                           n12756, ZN => n11668);
   U10138 : AOI221_X1 port map( B1 => n12913, B2 => n10898, C1 => n12910, C2 =>
                           n10866, A => n11610, ZN => n11603);
   U10139 : OAI22_X1 port map( A1 => n10026, A2 => n12907, B1 => n9994, B2 => 
                           n12904, ZN => n11610);
   U10140 : AOI221_X1 port map( B1 => n12865, B2 => n10250, C1 => n12862, C2 =>
                           n10226, A => n11624, ZN => n11619);
   U10141 : OAI22_X1 port map( A1 => n10645, A2 => n12859, B1 => n10518, B2 => 
                           n12856, ZN => n11624);
   U10142 : AOI221_X1 port map( B1 => n12913, B2 => n10897, C1 => n12910, C2 =>
                           n10865, A => n11587, ZN => n11584);
   U10143 : OAI22_X1 port map( A1 => n10025, A2 => n12907, B1 => n9993, B2 => 
                           n12904, ZN => n11587);
   U10144 : AOI221_X1 port map( B1 => n12865, B2 => n10249, C1 => n12862, C2 =>
                           n10225, A => n11595, ZN => n11592);
   U10145 : OAI22_X1 port map( A1 => n10644, A2 => n12859, B1 => n10517, B2 => 
                           n12856, ZN => n11595);
   U10146 : AOI221_X1 port map( B1 => n12913, B2 => n10896, C1 => n12910, C2 =>
                           n10864, A => n11568, ZN => n11565);
   U10147 : OAI22_X1 port map( A1 => n10024, A2 => n12907, B1 => n9992, B2 => 
                           n12904, ZN => n11568);
   U10148 : AOI221_X1 port map( B1 => n12865, B2 => n10248, C1 => n12862, C2 =>
                           n10224, A => n11576, ZN => n11573);
   U10149 : OAI22_X1 port map( A1 => n10643, A2 => n12859, B1 => n10516, B2 => 
                           n12856, ZN => n11576);
   U10150 : AOI221_X1 port map( B1 => n12913, B2 => n10895, C1 => n12910, C2 =>
                           n10863, A => n11549, ZN => n11546);
   U10151 : OAI22_X1 port map( A1 => n10023, A2 => n12907, B1 => n9991, B2 => 
                           n12904, ZN => n11549);
   U10152 : AOI221_X1 port map( B1 => n12865, B2 => n10247, C1 => n12862, C2 =>
                           n10223, A => n11557, ZN => n11554);
   U10153 : OAI22_X1 port map( A1 => n10642, A2 => n12859, B1 => n10515, B2 => 
                           n12856, ZN => n11557);
   U10154 : AOI221_X1 port map( B1 => n12913, B2 => n10894, C1 => n12910, C2 =>
                           n10862, A => n11530, ZN => n11527);
   U10155 : OAI22_X1 port map( A1 => n10022, A2 => n12907, B1 => n9990, B2 => 
                           n12904, ZN => n11530);
   U10156 : AOI221_X1 port map( B1 => n12865, B2 => n10246, C1 => n12862, C2 =>
                           n10222, A => n11538, ZN => n11535);
   U10157 : OAI22_X1 port map( A1 => n10641, A2 => n12859, B1 => n10514, B2 => 
                           n12856, ZN => n11538);
   U10158 : AOI221_X1 port map( B1 => n12913, B2 => n10893, C1 => n12910, C2 =>
                           n10861, A => n11511, ZN => n11508);
   U10159 : OAI22_X1 port map( A1 => n10021, A2 => n12907, B1 => n9989, B2 => 
                           n12904, ZN => n11511);
   U10160 : AOI221_X1 port map( B1 => n12865, B2 => n10245, C1 => n12862, C2 =>
                           n10221, A => n11519, ZN => n11516);
   U10161 : OAI22_X1 port map( A1 => n10640, A2 => n12859, B1 => n10513, B2 => 
                           n12856, ZN => n11519);
   U10162 : AOI221_X1 port map( B1 => n12913, B2 => n10892, C1 => n12910, C2 =>
                           n10860, A => n11492, ZN => n11489);
   U10163 : OAI22_X1 port map( A1 => n10020, A2 => n12907, B1 => n9988, B2 => 
                           n12904, ZN => n11492);
   U10164 : AOI221_X1 port map( B1 => n12865, B2 => n10244, C1 => n12862, C2 =>
                           n10220, A => n11500, ZN => n11497);
   U10165 : OAI22_X1 port map( A1 => n10639, A2 => n12859, B1 => n10512, B2 => 
                           n12856, ZN => n11500);
   U10166 : AOI221_X1 port map( B1 => n12913, B2 => n10891, C1 => n12910, C2 =>
                           n10859, A => n11473, ZN => n11470);
   U10167 : OAI22_X1 port map( A1 => n10019, A2 => n12907, B1 => n9987, B2 => 
                           n12904, ZN => n11473);
   U10168 : AOI221_X1 port map( B1 => n12865, B2 => n10243, C1 => n12862, C2 =>
                           n10219, A => n11481, ZN => n11478);
   U10169 : OAI22_X1 port map( A1 => n10638, A2 => n12859, B1 => n10511, B2 => 
                           n12856, ZN => n11481);
   U10170 : AOI221_X1 port map( B1 => n12913, B2 => n10890, C1 => n12910, C2 =>
                           n10858, A => n11454, ZN => n11451);
   U10171 : OAI22_X1 port map( A1 => n10018, A2 => n12907, B1 => n9986, B2 => 
                           n12904, ZN => n11454);
   U10172 : AOI221_X1 port map( B1 => n12865, B2 => n10242, C1 => n12862, C2 =>
                           n10218, A => n11462, ZN => n11459);
   U10173 : OAI22_X1 port map( A1 => n10637, A2 => n12859, B1 => n10510, B2 => 
                           n12856, ZN => n11462);
   U10174 : AOI221_X1 port map( B1 => n12913, B2 => n10889, C1 => n12910, C2 =>
                           n10857, A => n11435, ZN => n11432);
   U10175 : OAI22_X1 port map( A1 => n10017, A2 => n12907, B1 => n9985, B2 => 
                           n12904, ZN => n11435);
   U10176 : AOI221_X1 port map( B1 => n12865, B2 => n10241, C1 => n12862, C2 =>
                           n10217, A => n11443, ZN => n11440);
   U10177 : OAI22_X1 port map( A1 => n10636, A2 => n12859, B1 => n10509, B2 => 
                           n12856, ZN => n11443);
   U10178 : AOI221_X1 port map( B1 => n12913, B2 => n10888, C1 => n12910, C2 =>
                           n10856, A => n11416, ZN => n11413);
   U10179 : OAI22_X1 port map( A1 => n10016, A2 => n12907, B1 => n9984, B2 => 
                           n12904, ZN => n11416);
   U10180 : AOI221_X1 port map( B1 => n12865, B2 => n10240, C1 => n12862, C2 =>
                           n10216, A => n11424, ZN => n11421);
   U10181 : OAI22_X1 port map( A1 => n10635, A2 => n12859, B1 => n10508, B2 => 
                           n12856, ZN => n11424);
   U10182 : AOI221_X1 port map( B1 => n12913, B2 => n10887, C1 => n12910, C2 =>
                           n10855, A => n11397, ZN => n11394);
   U10183 : OAI22_X1 port map( A1 => n10015, A2 => n12907, B1 => n9983, B2 => 
                           n12904, ZN => n11397);
   U10184 : AOI221_X1 port map( B1 => n12865, B2 => n10239, C1 => n12862, C2 =>
                           n10215, A => n11405, ZN => n11402);
   U10185 : OAI22_X1 port map( A1 => n10634, A2 => n12859, B1 => n10507, B2 => 
                           n12856, ZN => n11405);
   U10186 : AOI221_X1 port map( B1 => n12914, B2 => n10886, C1 => n12911, C2 =>
                           n10854, A => n11378, ZN => n11375);
   U10187 : OAI22_X1 port map( A1 => n10014, A2 => n12908, B1 => n9982, B2 => 
                           n12905, ZN => n11378);
   U10188 : AOI221_X1 port map( B1 => n12866, B2 => n10238, C1 => n12863, C2 =>
                           n10214, A => n11386, ZN => n11383);
   U10189 : OAI22_X1 port map( A1 => n10633, A2 => n12860, B1 => n10506, B2 => 
                           n12857, ZN => n11386);
   U10190 : AOI221_X1 port map( B1 => n12914, B2 => n10885, C1 => n12911, C2 =>
                           n10853, A => n11359, ZN => n11356);
   U10191 : OAI22_X1 port map( A1 => n10013, A2 => n12908, B1 => n9981, B2 => 
                           n12905, ZN => n11359);
   U10192 : AOI221_X1 port map( B1 => n12866, B2 => n10237, C1 => n12863, C2 =>
                           n10213, A => n11367, ZN => n11364);
   U10193 : OAI22_X1 port map( A1 => n10632, A2 => n12860, B1 => n10505, B2 => 
                           n12857, ZN => n11367);
   U10194 : AOI221_X1 port map( B1 => n12914, B2 => n10884, C1 => n12911, C2 =>
                           n10852, A => n11340, ZN => n11337);
   U10195 : OAI22_X1 port map( A1 => n10012, A2 => n12908, B1 => n9980, B2 => 
                           n12905, ZN => n11340);
   U10196 : AOI221_X1 port map( B1 => n12866, B2 => n10236, C1 => n12863, C2 =>
                           n10212, A => n11348, ZN => n11345);
   U10197 : OAI22_X1 port map( A1 => n10631, A2 => n12860, B1 => n10504, B2 => 
                           n12857, ZN => n11348);
   U10198 : AOI221_X1 port map( B1 => n12914, B2 => n10883, C1 => n12911, C2 =>
                           n10851, A => n11321, ZN => n11318);
   U10199 : OAI22_X1 port map( A1 => n10011, A2 => n12908, B1 => n9979, B2 => 
                           n12905, ZN => n11321);
   U10200 : AOI221_X1 port map( B1 => n12866, B2 => n10235, C1 => n12863, C2 =>
                           n10211, A => n11329, ZN => n11326);
   U10201 : OAI22_X1 port map( A1 => n10630, A2 => n12860, B1 => n10503, B2 => 
                           n12857, ZN => n11329);
   U10202 : AOI221_X1 port map( B1 => n12914, B2 => n10882, C1 => n12911, C2 =>
                           n10850, A => n11302, ZN => n11299);
   U10203 : OAI22_X1 port map( A1 => n10010, A2 => n12908, B1 => n9978, B2 => 
                           n12905, ZN => n11302);
   U10204 : AOI221_X1 port map( B1 => n12866, B2 => n10234, C1 => n12863, C2 =>
                           n10210, A => n11310, ZN => n11307);
   U10205 : OAI22_X1 port map( A1 => n10629, A2 => n12860, B1 => n10502, B2 => 
                           n12857, ZN => n11310);
   U10206 : AOI221_X1 port map( B1 => n12914, B2 => n10881, C1 => n12911, C2 =>
                           n10849, A => n11283, ZN => n11280);
   U10207 : OAI22_X1 port map( A1 => n10009, A2 => n12908, B1 => n9977, B2 => 
                           n12905, ZN => n11283);
   U10208 : AOI221_X1 port map( B1 => n12866, B2 => n10233, C1 => n12863, C2 =>
                           n10209, A => n11291, ZN => n11288);
   U10209 : OAI22_X1 port map( A1 => n10628, A2 => n12860, B1 => n10501, B2 => 
                           n12857, ZN => n11291);
   U10210 : AOI221_X1 port map( B1 => n12914, B2 => n10880, C1 => n12911, C2 =>
                           n10848, A => n11264, ZN => n11261);
   U10211 : OAI22_X1 port map( A1 => n10008, A2 => n12908, B1 => n9976, B2 => 
                           n12905, ZN => n11264);
   U10212 : AOI221_X1 port map( B1 => n12866, B2 => n10232, C1 => n12863, C2 =>
                           n10208, A => n11272, ZN => n11269);
   U10213 : OAI22_X1 port map( A1 => n10627, A2 => n12860, B1 => n10500, B2 => 
                           n12857, ZN => n11272);
   U10214 : AOI221_X1 port map( B1 => n12914, B2 => n10879, C1 => n12911, C2 =>
                           n10847, A => n11245, ZN => n11242);
   U10215 : OAI22_X1 port map( A1 => n10007, A2 => n12908, B1 => n9975, B2 => 
                           n12905, ZN => n11245);
   U10216 : AOI221_X1 port map( B1 => n12866, B2 => n10231, C1 => n12863, C2 =>
                           n10207, A => n11253, ZN => n11250);
   U10217 : OAI22_X1 port map( A1 => n10626, A2 => n12860, B1 => n10499, B2 => 
                           n12857, ZN => n11253);
   U10218 : AOI221_X1 port map( B1 => n12914, B2 => n10878, C1 => n12911, C2 =>
                           n10846, A => n11226, ZN => n11223);
   U10219 : OAI22_X1 port map( A1 => n10006, A2 => n12908, B1 => n9974, B2 => 
                           n12905, ZN => n11226);
   U10220 : AOI221_X1 port map( B1 => n12866, B2 => n10230, C1 => n12863, C2 =>
                           n10206, A => n11234, ZN => n11231);
   U10221 : OAI22_X1 port map( A1 => n10625, A2 => n12860, B1 => n10498, B2 => 
                           n12857, ZN => n11234);
   U10222 : AOI221_X1 port map( B1 => n12914, B2 => n10877, C1 => n12911, C2 =>
                           n10845, A => n11207, ZN => n11204);
   U10223 : OAI22_X1 port map( A1 => n10005, A2 => n12908, B1 => n9973, B2 => 
                           n12905, ZN => n11207);
   U10224 : AOI221_X1 port map( B1 => n12866, B2 => n10229, C1 => n12863, C2 =>
                           n10205, A => n11215, ZN => n11212);
   U10225 : OAI22_X1 port map( A1 => n10624, A2 => n12860, B1 => n10497, B2 => 
                           n12857, ZN => n11215);
   U10226 : AOI221_X1 port map( B1 => n12914, B2 => n10876, C1 => n12911, C2 =>
                           n10844, A => n11188, ZN => n11185);
   U10227 : OAI22_X1 port map( A1 => n10004, A2 => n12908, B1 => n9972, B2 => 
                           n12905, ZN => n11188);
   U10228 : AOI221_X1 port map( B1 => n12866, B2 => n10228, C1 => n12863, C2 =>
                           n10204, A => n11196, ZN => n11193);
   U10229 : OAI22_X1 port map( A1 => n10623, A2 => n12860, B1 => n10496, B2 => 
                           n12857, ZN => n11196);
   U10230 : AOI221_X1 port map( B1 => n12914, B2 => n10875, C1 => n12911, C2 =>
                           n10843, A => n11169, ZN => n11166);
   U10231 : OAI22_X1 port map( A1 => n10003, A2 => n12908, B1 => n9971, B2 => 
                           n12905, ZN => n11169);
   U10232 : AOI221_X1 port map( B1 => n12866, B2 => n10227, C1 => n12863, C2 =>
                           n10203, A => n11177, ZN => n11174);
   U10233 : OAI22_X1 port map( A1 => n10622, A2 => n12860, B1 => n10495, B2 => 
                           n12857, ZN => n11177);
   U10234 : AOI221_X1 port map( B1 => n12867, B2 => n10098, C1 => n12864, C2 =>
                           n10090, A => n11158, ZN => n11155);
   U10235 : OAI22_X1 port map( A1 => n10426, A2 => n12861, B1 => n10378, B2 => 
                           n12858, ZN => n11158);
   U10236 : AOI221_X1 port map( B1 => n12867, B2 => n10097, C1 => n12864, C2 =>
                           n10089, A => n11139, ZN => n11136);
   U10237 : OAI22_X1 port map( A1 => n10425, A2 => n12861, B1 => n10377, B2 => 
                           n12858, ZN => n11139);
   U10238 : AOI221_X1 port map( B1 => n12867, B2 => n10096, C1 => n12864, C2 =>
                           n10088, A => n11120, ZN => n11117);
   U10239 : OAI22_X1 port map( A1 => n10424, A2 => n12861, B1 => n10376, B2 => 
                           n12858, ZN => n11120);
   U10240 : AOI221_X1 port map( B1 => n12867, B2 => n10095, C1 => n12864, C2 =>
                           n10087, A => n11101, ZN => n11098);
   U10241 : OAI22_X1 port map( A1 => n10423, A2 => n12861, B1 => n10375, B2 => 
                           n12858, ZN => n11101);
   U10242 : AOI221_X1 port map( B1 => n12867, B2 => n10094, C1 => n12864, C2 =>
                           n10086, A => n11082, ZN => n11079);
   U10243 : OAI22_X1 port map( A1 => n10422, A2 => n12861, B1 => n10374, B2 => 
                           n12858, ZN => n11082);
   U10244 : AOI221_X1 port map( B1 => n12867, B2 => n10093, C1 => n12864, C2 =>
                           n10085, A => n11063, ZN => n11060);
   U10245 : OAI22_X1 port map( A1 => n10421, A2 => n12861, B1 => n10373, B2 => 
                           n12858, ZN => n11063);
   U10246 : AOI221_X1 port map( B1 => n12867, B2 => n10092, C1 => n12864, C2 =>
                           n10084, A => n11044, ZN => n11041);
   U10247 : OAI22_X1 port map( A1 => n10420, A2 => n12861, B1 => n10372, B2 => 
                           n12858, ZN => n11044);
   U10248 : AOI221_X1 port map( B1 => n12867, B2 => n10091, C1 => n12864, C2 =>
                           n10083, A => n11015, ZN => n11006);
   U10249 : OAI22_X1 port map( A1 => n10419, A2 => n12861, B1 => n10371, B2 => 
                           n12858, ZN => n11015);
   U10250 : AOI221_X1 port map( B1 => n12751, B2 => n10202, C1 => n12748, C2 =>
                           n10178, A => n12278, ZN => n12271);
   U10251 : OAI22_X1 port map( A1 => n10621, A2 => n12745, B1 => n10494, B2 => 
                           n12742, ZN => n12278);
   U10252 : AOI221_X1 port map( B1 => n12751, B2 => n10201, C1 => n12748, C2 =>
                           n10177, A => n12249, ZN => n12244);
   U10253 : OAI22_X1 port map( A1 => n10620, A2 => n12745, B1 => n10493, B2 => 
                           n12742, ZN => n12249);
   U10254 : AOI221_X1 port map( B1 => n12751, B2 => n10200, C1 => n12748, C2 =>
                           n10176, A => n12230, ZN => n12225);
   U10255 : OAI22_X1 port map( A1 => n10619, A2 => n12745, B1 => n10492, B2 => 
                           n12742, ZN => n12230);
   U10256 : AOI221_X1 port map( B1 => n12751, B2 => n10199, C1 => n12748, C2 =>
                           n10175, A => n12211, ZN => n12206);
   U10257 : OAI22_X1 port map( A1 => n10618, A2 => n12745, B1 => n10491, B2 => 
                           n12742, ZN => n12211);
   U10258 : AOI221_X1 port map( B1 => n12751, B2 => n10198, C1 => n12748, C2 =>
                           n10174, A => n12192, ZN => n12187);
   U10259 : OAI22_X1 port map( A1 => n10617, A2 => n12745, B1 => n10490, B2 => 
                           n12742, ZN => n12192);
   U10260 : AOI221_X1 port map( B1 => n12751, B2 => n10197, C1 => n12748, C2 =>
                           n10173, A => n12173, ZN => n12168);
   U10261 : OAI22_X1 port map( A1 => n10616, A2 => n12745, B1 => n10489, B2 => 
                           n12742, ZN => n12173);
   U10262 : AOI221_X1 port map( B1 => n12751, B2 => n10196, C1 => n12748, C2 =>
                           n10172, A => n12154, ZN => n12149);
   U10263 : OAI22_X1 port map( A1 => n10615, A2 => n12745, B1 => n10488, B2 => 
                           n12742, ZN => n12154);
   U10264 : AOI221_X1 port map( B1 => n12751, B2 => n10195, C1 => n12748, C2 =>
                           n10171, A => n12135, ZN => n12130);
   U10265 : OAI22_X1 port map( A1 => n10614, A2 => n12745, B1 => n10487, B2 => 
                           n12742, ZN => n12135);
   U10266 : AOI221_X1 port map( B1 => n12751, B2 => n10194, C1 => n12748, C2 =>
                           n10170, A => n12116, ZN => n12111);
   U10267 : OAI22_X1 port map( A1 => n10613, A2 => n12745, B1 => n10486, B2 => 
                           n12742, ZN => n12116);
   U10268 : AOI221_X1 port map( B1 => n12751, B2 => n10193, C1 => n12748, C2 =>
                           n10169, A => n12097, ZN => n12092);
   U10269 : OAI22_X1 port map( A1 => n10612, A2 => n12745, B1 => n10485, B2 => 
                           n12742, ZN => n12097);
   U10270 : AOI221_X1 port map( B1 => n12751, B2 => n10192, C1 => n12748, C2 =>
                           n10168, A => n12078, ZN => n12073);
   U10271 : OAI22_X1 port map( A1 => n10611, A2 => n12745, B1 => n10484, B2 => 
                           n12742, ZN => n12078);
   U10272 : AOI221_X1 port map( B1 => n12751, B2 => n10191, C1 => n12748, C2 =>
                           n10167, A => n12059, ZN => n12054);
   U10273 : OAI22_X1 port map( A1 => n10610, A2 => n12745, B1 => n10483, B2 => 
                           n12742, ZN => n12059);
   U10274 : AOI221_X1 port map( B1 => n12752, B2 => n10190, C1 => n12749, C2 =>
                           n10166, A => n12040, ZN => n12035);
   U10275 : OAI22_X1 port map( A1 => n10609, A2 => n12746, B1 => n10482, B2 => 
                           n12743, ZN => n12040);
   U10276 : AOI221_X1 port map( B1 => n12752, B2 => n10189, C1 => n12749, C2 =>
                           n10165, A => n12021, ZN => n12016);
   U10277 : OAI22_X1 port map( A1 => n10608, A2 => n12746, B1 => n10481, B2 => 
                           n12743, ZN => n12021);
   U10278 : AOI221_X1 port map( B1 => n12752, B2 => n10188, C1 => n12749, C2 =>
                           n10164, A => n12002, ZN => n11997);
   U10279 : OAI22_X1 port map( A1 => n10607, A2 => n12746, B1 => n10480, B2 => 
                           n12743, ZN => n12002);
   U10280 : AOI221_X1 port map( B1 => n12752, B2 => n10187, C1 => n12749, C2 =>
                           n10163, A => n11983, ZN => n11978);
   U10281 : OAI22_X1 port map( A1 => n10606, A2 => n12746, B1 => n10479, B2 => 
                           n12743, ZN => n11983);
   U10282 : AOI221_X1 port map( B1 => n12752, B2 => n10186, C1 => n12749, C2 =>
                           n10162, A => n11964, ZN => n11959);
   U10283 : OAI22_X1 port map( A1 => n10605, A2 => n12746, B1 => n10478, B2 => 
                           n12743, ZN => n11964);
   U10284 : AOI221_X1 port map( B1 => n12752, B2 => n10185, C1 => n12749, C2 =>
                           n10161, A => n11945, ZN => n11940);
   U10285 : OAI22_X1 port map( A1 => n10604, A2 => n12746, B1 => n10477, B2 => 
                           n12743, ZN => n11945);
   U10286 : AOI221_X1 port map( B1 => n12752, B2 => n10184, C1 => n12749, C2 =>
                           n10160, A => n11926, ZN => n11921);
   U10287 : OAI22_X1 port map( A1 => n10603, A2 => n12746, B1 => n10476, B2 => 
                           n12743, ZN => n11926);
   U10288 : AOI221_X1 port map( B1 => n12752, B2 => n10183, C1 => n12749, C2 =>
                           n10159, A => n11907, ZN => n11902);
   U10289 : OAI22_X1 port map( A1 => n10602, A2 => n12746, B1 => n10475, B2 => 
                           n12743, ZN => n11907);
   U10290 : AOI221_X1 port map( B1 => n12752, B2 => n10182, C1 => n12749, C2 =>
                           n10158, A => n11888, ZN => n11883);
   U10291 : OAI22_X1 port map( A1 => n10601, A2 => n12746, B1 => n10474, B2 => 
                           n12743, ZN => n11888);
   U10292 : AOI221_X1 port map( B1 => n12752, B2 => n10181, C1 => n12749, C2 =>
                           n10157, A => n11869, ZN => n11864);
   U10293 : OAI22_X1 port map( A1 => n10600, A2 => n12746, B1 => n10473, B2 => 
                           n12743, ZN => n11869);
   U10294 : AOI221_X1 port map( B1 => n12752, B2 => n10180, C1 => n12749, C2 =>
                           n10156, A => n11850, ZN => n11845);
   U10295 : OAI22_X1 port map( A1 => n10599, A2 => n12746, B1 => n10472, B2 => 
                           n12743, ZN => n11850);
   U10296 : AOI221_X1 port map( B1 => n12752, B2 => n10179, C1 => n12749, C2 =>
                           n10155, A => n11831, ZN => n11826);
   U10297 : OAI22_X1 port map( A1 => n10598, A2 => n12746, B1 => n10471, B2 => 
                           n12743, ZN => n11831);
   U10298 : AOI221_X1 port map( B1 => n12853, B2 => n10202, C1 => n12850, C2 =>
                           n10178, A => n11625, ZN => n11618);
   U10299 : OAI22_X1 port map( A1 => n10621, A2 => n12847, B1 => n10494, B2 => 
                           n12844, ZN => n11625);
   U10300 : AOI221_X1 port map( B1 => n12853, B2 => n10201, C1 => n12850, C2 =>
                           n10177, A => n11596, ZN => n11591);
   U10301 : OAI22_X1 port map( A1 => n10620, A2 => n12847, B1 => n10493, B2 => 
                           n12844, ZN => n11596);
   U10302 : AOI221_X1 port map( B1 => n12853, B2 => n10200, C1 => n12850, C2 =>
                           n10176, A => n11577, ZN => n11572);
   U10303 : OAI22_X1 port map( A1 => n10619, A2 => n12847, B1 => n10492, B2 => 
                           n12844, ZN => n11577);
   U10304 : AOI221_X1 port map( B1 => n12853, B2 => n10199, C1 => n12850, C2 =>
                           n10175, A => n11558, ZN => n11553);
   U10305 : OAI22_X1 port map( A1 => n10618, A2 => n12847, B1 => n10491, B2 => 
                           n12844, ZN => n11558);
   U10306 : AOI221_X1 port map( B1 => n12853, B2 => n10198, C1 => n12850, C2 =>
                           n10174, A => n11539, ZN => n11534);
   U10307 : OAI22_X1 port map( A1 => n10617, A2 => n12847, B1 => n10490, B2 => 
                           n12844, ZN => n11539);
   U10308 : AOI221_X1 port map( B1 => n12853, B2 => n10197, C1 => n12850, C2 =>
                           n10173, A => n11520, ZN => n11515);
   U10309 : OAI22_X1 port map( A1 => n10616, A2 => n12847, B1 => n10489, B2 => 
                           n12844, ZN => n11520);
   U10310 : AOI221_X1 port map( B1 => n12853, B2 => n10196, C1 => n12850, C2 =>
                           n10172, A => n11501, ZN => n11496);
   U10311 : OAI22_X1 port map( A1 => n10615, A2 => n12847, B1 => n10488, B2 => 
                           n12844, ZN => n11501);
   U10312 : AOI221_X1 port map( B1 => n12853, B2 => n10195, C1 => n12850, C2 =>
                           n10171, A => n11482, ZN => n11477);
   U10313 : OAI22_X1 port map( A1 => n10614, A2 => n12847, B1 => n10487, B2 => 
                           n12844, ZN => n11482);
   U10314 : AOI221_X1 port map( B1 => n12853, B2 => n10194, C1 => n12850, C2 =>
                           n10170, A => n11463, ZN => n11458);
   U10315 : OAI22_X1 port map( A1 => n10613, A2 => n12847, B1 => n10486, B2 => 
                           n12844, ZN => n11463);
   U10316 : AOI221_X1 port map( B1 => n12853, B2 => n10193, C1 => n12850, C2 =>
                           n10169, A => n11444, ZN => n11439);
   U10317 : OAI22_X1 port map( A1 => n10612, A2 => n12847, B1 => n10485, B2 => 
                           n12844, ZN => n11444);
   U10318 : AOI221_X1 port map( B1 => n12853, B2 => n10192, C1 => n12850, C2 =>
                           n10168, A => n11425, ZN => n11420);
   U10319 : OAI22_X1 port map( A1 => n10611, A2 => n12847, B1 => n10484, B2 => 
                           n12844, ZN => n11425);
   U10320 : AOI221_X1 port map( B1 => n12853, B2 => n10191, C1 => n12850, C2 =>
                           n10167, A => n11406, ZN => n11401);
   U10321 : OAI22_X1 port map( A1 => n10610, A2 => n12847, B1 => n10483, B2 => 
                           n12844, ZN => n11406);
   U10322 : AOI221_X1 port map( B1 => n12854, B2 => n10190, C1 => n12851, C2 =>
                           n10166, A => n11387, ZN => n11382);
   U10323 : OAI22_X1 port map( A1 => n10609, A2 => n12848, B1 => n10482, B2 => 
                           n12845, ZN => n11387);
   U10324 : AOI221_X1 port map( B1 => n12854, B2 => n10189, C1 => n12851, C2 =>
                           n10165, A => n11368, ZN => n11363);
   U10325 : OAI22_X1 port map( A1 => n10608, A2 => n12848, B1 => n10481, B2 => 
                           n12845, ZN => n11368);
   U10326 : AOI221_X1 port map( B1 => n12854, B2 => n10188, C1 => n12851, C2 =>
                           n10164, A => n11349, ZN => n11344);
   U10327 : OAI22_X1 port map( A1 => n10607, A2 => n12848, B1 => n10480, B2 => 
                           n12845, ZN => n11349);
   U10328 : AOI221_X1 port map( B1 => n12854, B2 => n10187, C1 => n12851, C2 =>
                           n10163, A => n11330, ZN => n11325);
   U10329 : OAI22_X1 port map( A1 => n10606, A2 => n12848, B1 => n10479, B2 => 
                           n12845, ZN => n11330);
   U10330 : AOI221_X1 port map( B1 => n12854, B2 => n10186, C1 => n12851, C2 =>
                           n10162, A => n11311, ZN => n11306);
   U10331 : OAI22_X1 port map( A1 => n10605, A2 => n12848, B1 => n10478, B2 => 
                           n12845, ZN => n11311);
   U10332 : AOI221_X1 port map( B1 => n12854, B2 => n10185, C1 => n12851, C2 =>
                           n10161, A => n11292, ZN => n11287);
   U10333 : OAI22_X1 port map( A1 => n10604, A2 => n12848, B1 => n10477, B2 => 
                           n12845, ZN => n11292);
   U10334 : AOI221_X1 port map( B1 => n12854, B2 => n10184, C1 => n12851, C2 =>
                           n10160, A => n11273, ZN => n11268);
   U10335 : OAI22_X1 port map( A1 => n10603, A2 => n12848, B1 => n10476, B2 => 
                           n12845, ZN => n11273);
   U10336 : AOI221_X1 port map( B1 => n12854, B2 => n10183, C1 => n12851, C2 =>
                           n10159, A => n11254, ZN => n11249);
   U10337 : OAI22_X1 port map( A1 => n10602, A2 => n12848, B1 => n10475, B2 => 
                           n12845, ZN => n11254);
   U10338 : AOI221_X1 port map( B1 => n12854, B2 => n10182, C1 => n12851, C2 =>
                           n10158, A => n11235, ZN => n11230);
   U10339 : OAI22_X1 port map( A1 => n10601, A2 => n12848, B1 => n10474, B2 => 
                           n12845, ZN => n11235);
   U10340 : AOI221_X1 port map( B1 => n12854, B2 => n10181, C1 => n12851, C2 =>
                           n10157, A => n11216, ZN => n11211);
   U10341 : OAI22_X1 port map( A1 => n10600, A2 => n12848, B1 => n10473, B2 => 
                           n12845, ZN => n11216);
   U10342 : AOI221_X1 port map( B1 => n12854, B2 => n10180, C1 => n12851, C2 =>
                           n10156, A => n11197, ZN => n11192);
   U10343 : OAI22_X1 port map( A1 => n10599, A2 => n12848, B1 => n10472, B2 => 
                           n12845, ZN => n11197);
   U10344 : AOI221_X1 port map( B1 => n12854, B2 => n10179, C1 => n12851, C2 =>
                           n10155, A => n11178, ZN => n11173);
   U10345 : OAI22_X1 port map( A1 => n10598, A2 => n12848, B1 => n10471, B2 => 
                           n12845, ZN => n11178);
   U10346 : AOI221_X1 port map( B1 => n12855, B2 => n10082, C1 => n12852, C2 =>
                           n10074, A => n11159, ZN => n11154);
   U10347 : OAI22_X1 port map( A1 => n10418, A2 => n12849, B1 => n10370, B2 => 
                           n12846, ZN => n11159);
   U10348 : AOI221_X1 port map( B1 => n12855, B2 => n10081, C1 => n12852, C2 =>
                           n10073, A => n11140, ZN => n11135);
   U10349 : OAI22_X1 port map( A1 => n10417, A2 => n12849, B1 => n10369, B2 => 
                           n12846, ZN => n11140);
   U10350 : AOI221_X1 port map( B1 => n12855, B2 => n10080, C1 => n12852, C2 =>
                           n10072, A => n11121, ZN => n11116);
   U10351 : OAI22_X1 port map( A1 => n10416, A2 => n12849, B1 => n10368, B2 => 
                           n12846, ZN => n11121);
   U10352 : AOI221_X1 port map( B1 => n12855, B2 => n10079, C1 => n12852, C2 =>
                           n10071, A => n11102, ZN => n11097);
   U10353 : OAI22_X1 port map( A1 => n10415, A2 => n12849, B1 => n10367, B2 => 
                           n12846, ZN => n11102);
   U10354 : AOI221_X1 port map( B1 => n12855, B2 => n10078, C1 => n12852, C2 =>
                           n10070, A => n11083, ZN => n11078);
   U10355 : OAI22_X1 port map( A1 => n10414, A2 => n12849, B1 => n10366, B2 => 
                           n12846, ZN => n11083);
   U10356 : AOI221_X1 port map( B1 => n12855, B2 => n10077, C1 => n12852, C2 =>
                           n10069, A => n11064, ZN => n11059);
   U10357 : OAI22_X1 port map( A1 => n10413, A2 => n12849, B1 => n10365, B2 => 
                           n12846, ZN => n11064);
   U10358 : AOI221_X1 port map( B1 => n12855, B2 => n10076, C1 => n12852, C2 =>
                           n10068, A => n11045, ZN => n11040);
   U10359 : OAI22_X1 port map( A1 => n10412, A2 => n12849, B1 => n10364, B2 => 
                           n12846, ZN => n11045);
   U10360 : AOI221_X1 port map( B1 => n12855, B2 => n10075, C1 => n12852, C2 =>
                           n10067, A => n11020, ZN => n11005);
   U10361 : OAI22_X1 port map( A1 => n10411, A2 => n12849, B1 => n10363, B2 => 
                           n12846, ZN => n11020);
   U10362 : AOI221_X1 port map( B1 => n12787, B2 => n10298, C1 => n12784, C2 =>
                           n10274, A => n12269, ZN => n12254);
   U10363 : OAI22_X1 port map( A1 => n10693, A2 => n12781, B1 => n10566, B2 => 
                           n12778, ZN => n12269);
   U10364 : AOI221_X1 port map( B1 => n12739, B2 => n10154, C1 => n12736, C2 =>
                           n10058, A => n12281, ZN => n12270);
   U10365 : OAI22_X1 port map( A1 => n10597, A2 => n12733, B1 => n10470, B2 => 
                           n12730, ZN => n12281);
   U10366 : AOI221_X1 port map( B1 => n12787, B2 => n10297, C1 => n12784, C2 =>
                           n10273, A => n12242, ZN => n12235);
   U10367 : OAI22_X1 port map( A1 => n10692, A2 => n12781, B1 => n10565, B2 => 
                           n12778, ZN => n12242);
   U10368 : AOI221_X1 port map( B1 => n12739, B2 => n10153, C1 => n12736, C2 =>
                           n10057, A => n12250, ZN => n12243);
   U10369 : OAI22_X1 port map( A1 => n10596, A2 => n12733, B1 => n10469, B2 => 
                           n12730, ZN => n12250);
   U10370 : AOI221_X1 port map( B1 => n12787, B2 => n10296, C1 => n12784, C2 =>
                           n10272, A => n12223, ZN => n12216);
   U10371 : OAI22_X1 port map( A1 => n10691, A2 => n12781, B1 => n10564, B2 => 
                           n12778, ZN => n12223);
   U10372 : AOI221_X1 port map( B1 => n12739, B2 => n10152, C1 => n12736, C2 =>
                           n10056, A => n12231, ZN => n12224);
   U10373 : OAI22_X1 port map( A1 => n10595, A2 => n12733, B1 => n10468, B2 => 
                           n12730, ZN => n12231);
   U10374 : AOI221_X1 port map( B1 => n12787, B2 => n10295, C1 => n12784, C2 =>
                           n10271, A => n12204, ZN => n12197);
   U10375 : OAI22_X1 port map( A1 => n10690, A2 => n12781, B1 => n10563, B2 => 
                           n12778, ZN => n12204);
   U10376 : AOI221_X1 port map( B1 => n12739, B2 => n10151, C1 => n12736, C2 =>
                           n10055, A => n12212, ZN => n12205);
   U10377 : OAI22_X1 port map( A1 => n10594, A2 => n12733, B1 => n10467, B2 => 
                           n12730, ZN => n12212);
   U10378 : AOI221_X1 port map( B1 => n12787, B2 => n10294, C1 => n12784, C2 =>
                           n10270, A => n12185, ZN => n12178);
   U10379 : OAI22_X1 port map( A1 => n10689, A2 => n12781, B1 => n10562, B2 => 
                           n12778, ZN => n12185);
   U10380 : AOI221_X1 port map( B1 => n12739, B2 => n10150, C1 => n12736, C2 =>
                           n10054, A => n12193, ZN => n12186);
   U10381 : OAI22_X1 port map( A1 => n10593, A2 => n12733, B1 => n10466, B2 => 
                           n12730, ZN => n12193);
   U10382 : AOI221_X1 port map( B1 => n12787, B2 => n10293, C1 => n12784, C2 =>
                           n10269, A => n12166, ZN => n12159);
   U10383 : OAI22_X1 port map( A1 => n10688, A2 => n12781, B1 => n10561, B2 => 
                           n12778, ZN => n12166);
   U10384 : AOI221_X1 port map( B1 => n12739, B2 => n10149, C1 => n12736, C2 =>
                           n10053, A => n12174, ZN => n12167);
   U10385 : OAI22_X1 port map( A1 => n10592, A2 => n12733, B1 => n10465, B2 => 
                           n12730, ZN => n12174);
   U10386 : AOI221_X1 port map( B1 => n12787, B2 => n10292, C1 => n12784, C2 =>
                           n10268, A => n12147, ZN => n12140);
   U10387 : OAI22_X1 port map( A1 => n10687, A2 => n12781, B1 => n10560, B2 => 
                           n12778, ZN => n12147);
   U10388 : AOI221_X1 port map( B1 => n12739, B2 => n10148, C1 => n12736, C2 =>
                           n10052, A => n12155, ZN => n12148);
   U10389 : OAI22_X1 port map( A1 => n10591, A2 => n12733, B1 => n10464, B2 => 
                           n12730, ZN => n12155);
   U10390 : AOI221_X1 port map( B1 => n12787, B2 => n10291, C1 => n12784, C2 =>
                           n10267, A => n12128, ZN => n12121);
   U10391 : OAI22_X1 port map( A1 => n10686, A2 => n12781, B1 => n10559, B2 => 
                           n12778, ZN => n12128);
   U10392 : AOI221_X1 port map( B1 => n12739, B2 => n10147, C1 => n12736, C2 =>
                           n10051, A => n12136, ZN => n12129);
   U10393 : OAI22_X1 port map( A1 => n10590, A2 => n12733, B1 => n10463, B2 => 
                           n12730, ZN => n12136);
   U10394 : AOI221_X1 port map( B1 => n12787, B2 => n10290, C1 => n12784, C2 =>
                           n10266, A => n12109, ZN => n12102);
   U10395 : OAI22_X1 port map( A1 => n10685, A2 => n12781, B1 => n10558, B2 => 
                           n12778, ZN => n12109);
   U10396 : AOI221_X1 port map( B1 => n12739, B2 => n10146, C1 => n12736, C2 =>
                           n10050, A => n12117, ZN => n12110);
   U10397 : OAI22_X1 port map( A1 => n10589, A2 => n12733, B1 => n10462, B2 => 
                           n12730, ZN => n12117);
   U10398 : AOI221_X1 port map( B1 => n12787, B2 => n10289, C1 => n12784, C2 =>
                           n10265, A => n12090, ZN => n12083);
   U10399 : OAI22_X1 port map( A1 => n10684, A2 => n12781, B1 => n10557, B2 => 
                           n12778, ZN => n12090);
   U10400 : AOI221_X1 port map( B1 => n12739, B2 => n10145, C1 => n12736, C2 =>
                           n10049, A => n12098, ZN => n12091);
   U10401 : OAI22_X1 port map( A1 => n10588, A2 => n12733, B1 => n10461, B2 => 
                           n12730, ZN => n12098);
   U10402 : AOI221_X1 port map( B1 => n12787, B2 => n10288, C1 => n12784, C2 =>
                           n10264, A => n12071, ZN => n12064);
   U10403 : OAI22_X1 port map( A1 => n10683, A2 => n12781, B1 => n10556, B2 => 
                           n12778, ZN => n12071);
   U10404 : AOI221_X1 port map( B1 => n12739, B2 => n10144, C1 => n12736, C2 =>
                           n10048, A => n12079, ZN => n12072);
   U10405 : OAI22_X1 port map( A1 => n10587, A2 => n12733, B1 => n10460, B2 => 
                           n12730, ZN => n12079);
   U10406 : AOI221_X1 port map( B1 => n12787, B2 => n10287, C1 => n12784, C2 =>
                           n10263, A => n12052, ZN => n12045);
   U10407 : OAI22_X1 port map( A1 => n10682, A2 => n12781, B1 => n10555, B2 => 
                           n12778, ZN => n12052);
   U10408 : AOI221_X1 port map( B1 => n12739, B2 => n10143, C1 => n12736, C2 =>
                           n10047, A => n12060, ZN => n12053);
   U10409 : OAI22_X1 port map( A1 => n10586, A2 => n12733, B1 => n10459, B2 => 
                           n12730, ZN => n12060);
   U10410 : AOI221_X1 port map( B1 => n12788, B2 => n10286, C1 => n12785, C2 =>
                           n10262, A => n12033, ZN => n12026);
   U10411 : OAI22_X1 port map( A1 => n10681, A2 => n12782, B1 => n10554, B2 => 
                           n12779, ZN => n12033);
   U10412 : AOI221_X1 port map( B1 => n12740, B2 => n10142, C1 => n12737, C2 =>
                           n10046, A => n12041, ZN => n12034);
   U10413 : OAI22_X1 port map( A1 => n10585, A2 => n12734, B1 => n10458, B2 => 
                           n12731, ZN => n12041);
   U10414 : AOI221_X1 port map( B1 => n12788, B2 => n10285, C1 => n12785, C2 =>
                           n10261, A => n12014, ZN => n12007);
   U10415 : OAI22_X1 port map( A1 => n10680, A2 => n12782, B1 => n10553, B2 => 
                           n12779, ZN => n12014);
   U10416 : AOI221_X1 port map( B1 => n12740, B2 => n10141, C1 => n12737, C2 =>
                           n10045, A => n12022, ZN => n12015);
   U10417 : OAI22_X1 port map( A1 => n10584, A2 => n12734, B1 => n10457, B2 => 
                           n12731, ZN => n12022);
   U10418 : AOI221_X1 port map( B1 => n12788, B2 => n10284, C1 => n12785, C2 =>
                           n10260, A => n11995, ZN => n11988);
   U10419 : OAI22_X1 port map( A1 => n10679, A2 => n12782, B1 => n10552, B2 => 
                           n12779, ZN => n11995);
   U10420 : AOI221_X1 port map( B1 => n12740, B2 => n10140, C1 => n12737, C2 =>
                           n10044, A => n12003, ZN => n11996);
   U10421 : OAI22_X1 port map( A1 => n10583, A2 => n12734, B1 => n10456, B2 => 
                           n12731, ZN => n12003);
   U10422 : AOI221_X1 port map( B1 => n12788, B2 => n10283, C1 => n12785, C2 =>
                           n10259, A => n11976, ZN => n11969);
   U10423 : OAI22_X1 port map( A1 => n10678, A2 => n12782, B1 => n10551, B2 => 
                           n12779, ZN => n11976);
   U10424 : AOI221_X1 port map( B1 => n12740, B2 => n10139, C1 => n12737, C2 =>
                           n10043, A => n11984, ZN => n11977);
   U10425 : OAI22_X1 port map( A1 => n10582, A2 => n12734, B1 => n10455, B2 => 
                           n12731, ZN => n11984);
   U10426 : AOI221_X1 port map( B1 => n12788, B2 => n10282, C1 => n12785, C2 =>
                           n10258, A => n11957, ZN => n11950);
   U10427 : OAI22_X1 port map( A1 => n10677, A2 => n12782, B1 => n10550, B2 => 
                           n12779, ZN => n11957);
   U10428 : AOI221_X1 port map( B1 => n12740, B2 => n10138, C1 => n12737, C2 =>
                           n10042, A => n11965, ZN => n11958);
   U10429 : OAI22_X1 port map( A1 => n10581, A2 => n12734, B1 => n10454, B2 => 
                           n12731, ZN => n11965);
   U10430 : AOI221_X1 port map( B1 => n12788, B2 => n10281, C1 => n12785, C2 =>
                           n10257, A => n11938, ZN => n11931);
   U10431 : OAI22_X1 port map( A1 => n10676, A2 => n12782, B1 => n10549, B2 => 
                           n12779, ZN => n11938);
   U10432 : AOI221_X1 port map( B1 => n12740, B2 => n10137, C1 => n12737, C2 =>
                           n10041, A => n11946, ZN => n11939);
   U10433 : OAI22_X1 port map( A1 => n10580, A2 => n12734, B1 => n10453, B2 => 
                           n12731, ZN => n11946);
   U10434 : AOI221_X1 port map( B1 => n12788, B2 => n10280, C1 => n12785, C2 =>
                           n10256, A => n11919, ZN => n11912);
   U10435 : OAI22_X1 port map( A1 => n10675, A2 => n12782, B1 => n10548, B2 => 
                           n12779, ZN => n11919);
   U10436 : AOI221_X1 port map( B1 => n12740, B2 => n10136, C1 => n12737, C2 =>
                           n10040, A => n11927, ZN => n11920);
   U10437 : OAI22_X1 port map( A1 => n10579, A2 => n12734, B1 => n10452, B2 => 
                           n12731, ZN => n11927);
   U10438 : AOI221_X1 port map( B1 => n12788, B2 => n10279, C1 => n12785, C2 =>
                           n10255, A => n11900, ZN => n11893);
   U10439 : OAI22_X1 port map( A1 => n10674, A2 => n12782, B1 => n10547, B2 => 
                           n12779, ZN => n11900);
   U10440 : AOI221_X1 port map( B1 => n12740, B2 => n10135, C1 => n12737, C2 =>
                           n10039, A => n11908, ZN => n11901);
   U10441 : OAI22_X1 port map( A1 => n10578, A2 => n12734, B1 => n10451, B2 => 
                           n12731, ZN => n11908);
   U10442 : AOI221_X1 port map( B1 => n12788, B2 => n10278, C1 => n12785, C2 =>
                           n10254, A => n11881, ZN => n11874);
   U10443 : OAI22_X1 port map( A1 => n10673, A2 => n12782, B1 => n10546, B2 => 
                           n12779, ZN => n11881);
   U10444 : AOI221_X1 port map( B1 => n12740, B2 => n10134, C1 => n12737, C2 =>
                           n10038, A => n11889, ZN => n11882);
   U10445 : OAI22_X1 port map( A1 => n10577, A2 => n12734, B1 => n10450, B2 => 
                           n12731, ZN => n11889);
   U10446 : AOI221_X1 port map( B1 => n12788, B2 => n10277, C1 => n12785, C2 =>
                           n10253, A => n11862, ZN => n11855);
   U10447 : OAI22_X1 port map( A1 => n10672, A2 => n12782, B1 => n10545, B2 => 
                           n12779, ZN => n11862);
   U10448 : AOI221_X1 port map( B1 => n12740, B2 => n10133, C1 => n12737, C2 =>
                           n10037, A => n11870, ZN => n11863);
   U10449 : OAI22_X1 port map( A1 => n10576, A2 => n12734, B1 => n10449, B2 => 
                           n12731, ZN => n11870);
   U10450 : AOI221_X1 port map( B1 => n12788, B2 => n10276, C1 => n12785, C2 =>
                           n10252, A => n11843, ZN => n11836);
   U10451 : OAI22_X1 port map( A1 => n10671, A2 => n12782, B1 => n10544, B2 => 
                           n12779, ZN => n11843);
   U10452 : AOI221_X1 port map( B1 => n12740, B2 => n10132, C1 => n12737, C2 =>
                           n10036, A => n11851, ZN => n11844);
   U10453 : OAI22_X1 port map( A1 => n10575, A2 => n12734, B1 => n10448, B2 => 
                           n12731, ZN => n11851);
   U10454 : AOI221_X1 port map( B1 => n12788, B2 => n10275, C1 => n12785, C2 =>
                           n10251, A => n11824, ZN => n11817);
   U10455 : OAI22_X1 port map( A1 => n10670, A2 => n12782, B1 => n10543, B2 => 
                           n12779, ZN => n11824);
   U10456 : AOI221_X1 port map( B1 => n12740, B2 => n10131, C1 => n12737, C2 =>
                           n10035, A => n11832, ZN => n11825);
   U10457 : OAI22_X1 port map( A1 => n10574, A2 => n12734, B1 => n10447, B2 => 
                           n12731, ZN => n11832);
   U10458 : AOI221_X1 port map( B1 => n12789, B2 => n10114, C1 => n12786, C2 =>
                           n10106, A => n11805, ZN => n11798);
   U10459 : OAI22_X1 port map( A1 => n10442, A2 => n12783, B1 => n10394, B2 => 
                           n12780, ZN => n11805);
   U10460 : AOI221_X1 port map( B1 => n12741, B2 => n10066, C1 => n12738, C2 =>
                           n10034, A => n11813, ZN => n11806);
   U10461 : OAI22_X1 port map( A1 => n10410, A2 => n12735, B1 => n10362, B2 => 
                           n12732, ZN => n11813);
   U10462 : AOI221_X1 port map( B1 => n12789, B2 => n10113, C1 => n12786, C2 =>
                           n10105, A => n11786, ZN => n11779);
   U10463 : OAI22_X1 port map( A1 => n10441, A2 => n12783, B1 => n10393, B2 => 
                           n12780, ZN => n11786);
   U10464 : AOI221_X1 port map( B1 => n12741, B2 => n10065, C1 => n12738, C2 =>
                           n10033, A => n11794, ZN => n11787);
   U10465 : OAI22_X1 port map( A1 => n10409, A2 => n12735, B1 => n10361, B2 => 
                           n12732, ZN => n11794);
   U10466 : AOI221_X1 port map( B1 => n12789, B2 => n10112, C1 => n12786, C2 =>
                           n10104, A => n11767, ZN => n11760);
   U10467 : OAI22_X1 port map( A1 => n10440, A2 => n12783, B1 => n10392, B2 => 
                           n12780, ZN => n11767);
   U10468 : AOI221_X1 port map( B1 => n12741, B2 => n10064, C1 => n12738, C2 =>
                           n10032, A => n11775, ZN => n11768);
   U10469 : OAI22_X1 port map( A1 => n10408, A2 => n12735, B1 => n10360, B2 => 
                           n12732, ZN => n11775);
   U10470 : AOI221_X1 port map( B1 => n12789, B2 => n10111, C1 => n12786, C2 =>
                           n10103, A => n11748, ZN => n11741);
   U10471 : OAI22_X1 port map( A1 => n10439, A2 => n12783, B1 => n10391, B2 => 
                           n12780, ZN => n11748);
   U10472 : AOI221_X1 port map( B1 => n12741, B2 => n10063, C1 => n12738, C2 =>
                           n10031, A => n11756, ZN => n11749);
   U10473 : OAI22_X1 port map( A1 => n10407, A2 => n12735, B1 => n10359, B2 => 
                           n12732, ZN => n11756);
   U10474 : AOI221_X1 port map( B1 => n12789, B2 => n10110, C1 => n12786, C2 =>
                           n10102, A => n11729, ZN => n11722);
   U10475 : OAI22_X1 port map( A1 => n10438, A2 => n12783, B1 => n10390, B2 => 
                           n12780, ZN => n11729);
   U10476 : AOI221_X1 port map( B1 => n12741, B2 => n10062, C1 => n12738, C2 =>
                           n10030, A => n11737, ZN => n11730);
   U10477 : OAI22_X1 port map( A1 => n10406, A2 => n12735, B1 => n10358, B2 => 
                           n12732, ZN => n11737);
   U10478 : AOI221_X1 port map( B1 => n12789, B2 => n10109, C1 => n12786, C2 =>
                           n10101, A => n11710, ZN => n11703);
   U10479 : OAI22_X1 port map( A1 => n10437, A2 => n12783, B1 => n10389, B2 => 
                           n12780, ZN => n11710);
   U10480 : AOI221_X1 port map( B1 => n12741, B2 => n10061, C1 => n12738, C2 =>
                           n10029, A => n11718, ZN => n11711);
   U10481 : OAI22_X1 port map( A1 => n10405, A2 => n12735, B1 => n10357, B2 => 
                           n12732, ZN => n11718);
   U10482 : AOI221_X1 port map( B1 => n12789, B2 => n10108, C1 => n12786, C2 =>
                           n10100, A => n11691, ZN => n11684);
   U10483 : OAI22_X1 port map( A1 => n10436, A2 => n12783, B1 => n10388, B2 => 
                           n12780, ZN => n11691);
   U10484 : AOI221_X1 port map( B1 => n12741, B2 => n10060, C1 => n12738, C2 =>
                           n10028, A => n11699, ZN => n11692);
   U10485 : OAI22_X1 port map( A1 => n10404, A2 => n12735, B1 => n10356, B2 => 
                           n12732, ZN => n11699);
   U10486 : AOI221_X1 port map( B1 => n12789, B2 => n10107, C1 => n12786, C2 =>
                           n10099, A => n11654, ZN => n11633);
   U10487 : OAI22_X1 port map( A1 => n10435, A2 => n12783, B1 => n10387, B2 => 
                           n12780, ZN => n11654);
   U10488 : AOI221_X1 port map( B1 => n12741, B2 => n10059, C1 => n12738, C2 =>
                           n10027, A => n11678, ZN => n11657);
   U10489 : OAI22_X1 port map( A1 => n10403, A2 => n12735, B1 => n10355, B2 => 
                           n12732, ZN => n11678);
   U10490 : AOI221_X1 port map( B1 => n12889, B2 => n10298, C1 => n12886, C2 =>
                           n10274, A => n11616, ZN => n11601);
   U10491 : OAI22_X1 port map( A1 => n10693, A2 => n12883, B1 => n10566, B2 => 
                           n12880, ZN => n11616);
   U10492 : AOI221_X1 port map( B1 => n12841, B2 => n10154, C1 => n12838, C2 =>
                           n10058, A => n11628, ZN => n11617);
   U10493 : OAI22_X1 port map( A1 => n10597, A2 => n12835, B1 => n10470, B2 => 
                           n12832, ZN => n11628);
   U10494 : AOI221_X1 port map( B1 => n12889, B2 => n10297, C1 => n12886, C2 =>
                           n10273, A => n11589, ZN => n11582);
   U10495 : OAI22_X1 port map( A1 => n10692, A2 => n12883, B1 => n10565, B2 => 
                           n12880, ZN => n11589);
   U10496 : AOI221_X1 port map( B1 => n12841, B2 => n10153, C1 => n12838, C2 =>
                           n10057, A => n11597, ZN => n11590);
   U10497 : OAI22_X1 port map( A1 => n10596, A2 => n12835, B1 => n10469, B2 => 
                           n12832, ZN => n11597);
   U10498 : AOI221_X1 port map( B1 => n12889, B2 => n10296, C1 => n12886, C2 =>
                           n10272, A => n11570, ZN => n11563);
   U10499 : OAI22_X1 port map( A1 => n10691, A2 => n12883, B1 => n10564, B2 => 
                           n12880, ZN => n11570);
   U10500 : AOI221_X1 port map( B1 => n12841, B2 => n10152, C1 => n12838, C2 =>
                           n10056, A => n11578, ZN => n11571);
   U10501 : OAI22_X1 port map( A1 => n10595, A2 => n12835, B1 => n10468, B2 => 
                           n12832, ZN => n11578);
   U10502 : AOI221_X1 port map( B1 => n12889, B2 => n10295, C1 => n12886, C2 =>
                           n10271, A => n11551, ZN => n11544);
   U10503 : OAI22_X1 port map( A1 => n10690, A2 => n12883, B1 => n10563, B2 => 
                           n12880, ZN => n11551);
   U10504 : AOI221_X1 port map( B1 => n12841, B2 => n10151, C1 => n12838, C2 =>
                           n10055, A => n11559, ZN => n11552);
   U10505 : OAI22_X1 port map( A1 => n10594, A2 => n12835, B1 => n10467, B2 => 
                           n12832, ZN => n11559);
   U10506 : AOI221_X1 port map( B1 => n12889, B2 => n10294, C1 => n12886, C2 =>
                           n10270, A => n11532, ZN => n11525);
   U10507 : OAI22_X1 port map( A1 => n10689, A2 => n12883, B1 => n10562, B2 => 
                           n12880, ZN => n11532);
   U10508 : AOI221_X1 port map( B1 => n12841, B2 => n10150, C1 => n12838, C2 =>
                           n10054, A => n11540, ZN => n11533);
   U10509 : OAI22_X1 port map( A1 => n10593, A2 => n12835, B1 => n10466, B2 => 
                           n12832, ZN => n11540);
   U10510 : AOI221_X1 port map( B1 => n12889, B2 => n10293, C1 => n12886, C2 =>
                           n10269, A => n11513, ZN => n11506);
   U10511 : OAI22_X1 port map( A1 => n10688, A2 => n12883, B1 => n10561, B2 => 
                           n12880, ZN => n11513);
   U10512 : AOI221_X1 port map( B1 => n12841, B2 => n10149, C1 => n12838, C2 =>
                           n10053, A => n11521, ZN => n11514);
   U10513 : OAI22_X1 port map( A1 => n10592, A2 => n12835, B1 => n10465, B2 => 
                           n12832, ZN => n11521);
   U10514 : AOI221_X1 port map( B1 => n12889, B2 => n10292, C1 => n12886, C2 =>
                           n10268, A => n11494, ZN => n11487);
   U10515 : OAI22_X1 port map( A1 => n10687, A2 => n12883, B1 => n10560, B2 => 
                           n12880, ZN => n11494);
   U10516 : AOI221_X1 port map( B1 => n12841, B2 => n10148, C1 => n12838, C2 =>
                           n10052, A => n11502, ZN => n11495);
   U10517 : OAI22_X1 port map( A1 => n10591, A2 => n12835, B1 => n10464, B2 => 
                           n12832, ZN => n11502);
   U10518 : AOI221_X1 port map( B1 => n12889, B2 => n10291, C1 => n12886, C2 =>
                           n10267, A => n11475, ZN => n11468);
   U10519 : OAI22_X1 port map( A1 => n10686, A2 => n12883, B1 => n10559, B2 => 
                           n12880, ZN => n11475);
   U10520 : AOI221_X1 port map( B1 => n12841, B2 => n10147, C1 => n12838, C2 =>
                           n10051, A => n11483, ZN => n11476);
   U10521 : OAI22_X1 port map( A1 => n10590, A2 => n12835, B1 => n10463, B2 => 
                           n12832, ZN => n11483);
   U10522 : AOI221_X1 port map( B1 => n12889, B2 => n10290, C1 => n12886, C2 =>
                           n10266, A => n11456, ZN => n11449);
   U10523 : OAI22_X1 port map( A1 => n10685, A2 => n12883, B1 => n10558, B2 => 
                           n12880, ZN => n11456);
   U10524 : AOI221_X1 port map( B1 => n12841, B2 => n10146, C1 => n12838, C2 =>
                           n10050, A => n11464, ZN => n11457);
   U10525 : OAI22_X1 port map( A1 => n10589, A2 => n12835, B1 => n10462, B2 => 
                           n12832, ZN => n11464);
   U10526 : AOI221_X1 port map( B1 => n12889, B2 => n10289, C1 => n12886, C2 =>
                           n10265, A => n11437, ZN => n11430);
   U10527 : OAI22_X1 port map( A1 => n10684, A2 => n12883, B1 => n10557, B2 => 
                           n12880, ZN => n11437);
   U10528 : AOI221_X1 port map( B1 => n12841, B2 => n10145, C1 => n12838, C2 =>
                           n10049, A => n11445, ZN => n11438);
   U10529 : OAI22_X1 port map( A1 => n10588, A2 => n12835, B1 => n10461, B2 => 
                           n12832, ZN => n11445);
   U10530 : AOI221_X1 port map( B1 => n12889, B2 => n10288, C1 => n12886, C2 =>
                           n10264, A => n11418, ZN => n11411);
   U10531 : OAI22_X1 port map( A1 => n10683, A2 => n12883, B1 => n10556, B2 => 
                           n12880, ZN => n11418);
   U10532 : AOI221_X1 port map( B1 => n12841, B2 => n10144, C1 => n12838, C2 =>
                           n10048, A => n11426, ZN => n11419);
   U10533 : OAI22_X1 port map( A1 => n10587, A2 => n12835, B1 => n10460, B2 => 
                           n12832, ZN => n11426);
   U10534 : AOI221_X1 port map( B1 => n12889, B2 => n10287, C1 => n12886, C2 =>
                           n10263, A => n11399, ZN => n11392);
   U10535 : OAI22_X1 port map( A1 => n10682, A2 => n12883, B1 => n10555, B2 => 
                           n12880, ZN => n11399);
   U10536 : AOI221_X1 port map( B1 => n12841, B2 => n10143, C1 => n12838, C2 =>
                           n10047, A => n11407, ZN => n11400);
   U10537 : OAI22_X1 port map( A1 => n10586, A2 => n12835, B1 => n10459, B2 => 
                           n12832, ZN => n11407);
   U10538 : AOI221_X1 port map( B1 => n12890, B2 => n10286, C1 => n12887, C2 =>
                           n10262, A => n11380, ZN => n11373);
   U10539 : OAI22_X1 port map( A1 => n10681, A2 => n12884, B1 => n10554, B2 => 
                           n12881, ZN => n11380);
   U10540 : AOI221_X1 port map( B1 => n12842, B2 => n10142, C1 => n12839, C2 =>
                           n10046, A => n11388, ZN => n11381);
   U10541 : OAI22_X1 port map( A1 => n10585, A2 => n12836, B1 => n10458, B2 => 
                           n12833, ZN => n11388);
   U10542 : AOI221_X1 port map( B1 => n12890, B2 => n10285, C1 => n12887, C2 =>
                           n10261, A => n11361, ZN => n11354);
   U10543 : OAI22_X1 port map( A1 => n10680, A2 => n12884, B1 => n10553, B2 => 
                           n12881, ZN => n11361);
   U10544 : AOI221_X1 port map( B1 => n12842, B2 => n10141, C1 => n12839, C2 =>
                           n10045, A => n11369, ZN => n11362);
   U10545 : OAI22_X1 port map( A1 => n10584, A2 => n12836, B1 => n10457, B2 => 
                           n12833, ZN => n11369);
   U10546 : AOI221_X1 port map( B1 => n12890, B2 => n10284, C1 => n12887, C2 =>
                           n10260, A => n11342, ZN => n11335);
   U10547 : OAI22_X1 port map( A1 => n10679, A2 => n12884, B1 => n10552, B2 => 
                           n12881, ZN => n11342);
   U10548 : AOI221_X1 port map( B1 => n12842, B2 => n10140, C1 => n12839, C2 =>
                           n10044, A => n11350, ZN => n11343);
   U10549 : OAI22_X1 port map( A1 => n10583, A2 => n12836, B1 => n10456, B2 => 
                           n12833, ZN => n11350);
   U10550 : AOI221_X1 port map( B1 => n12890, B2 => n10283, C1 => n12887, C2 =>
                           n10259, A => n11323, ZN => n11316);
   U10551 : OAI22_X1 port map( A1 => n10678, A2 => n12884, B1 => n10551, B2 => 
                           n12881, ZN => n11323);
   U10552 : AOI221_X1 port map( B1 => n12842, B2 => n10139, C1 => n12839, C2 =>
                           n10043, A => n11331, ZN => n11324);
   U10553 : OAI22_X1 port map( A1 => n10582, A2 => n12836, B1 => n10455, B2 => 
                           n12833, ZN => n11331);
   U10554 : AOI221_X1 port map( B1 => n12890, B2 => n10282, C1 => n12887, C2 =>
                           n10258, A => n11304, ZN => n11297);
   U10555 : OAI22_X1 port map( A1 => n10677, A2 => n12884, B1 => n10550, B2 => 
                           n12881, ZN => n11304);
   U10556 : AOI221_X1 port map( B1 => n12842, B2 => n10138, C1 => n12839, C2 =>
                           n10042, A => n11312, ZN => n11305);
   U10557 : OAI22_X1 port map( A1 => n10581, A2 => n12836, B1 => n10454, B2 => 
                           n12833, ZN => n11312);
   U10558 : AOI221_X1 port map( B1 => n12890, B2 => n10281, C1 => n12887, C2 =>
                           n10257, A => n11285, ZN => n11278);
   U10559 : OAI22_X1 port map( A1 => n10676, A2 => n12884, B1 => n10549, B2 => 
                           n12881, ZN => n11285);
   U10560 : AOI221_X1 port map( B1 => n12842, B2 => n10137, C1 => n12839, C2 =>
                           n10041, A => n11293, ZN => n11286);
   U10561 : OAI22_X1 port map( A1 => n10580, A2 => n12836, B1 => n10453, B2 => 
                           n12833, ZN => n11293);
   U10562 : AOI221_X1 port map( B1 => n12890, B2 => n10280, C1 => n12887, C2 =>
                           n10256, A => n11266, ZN => n11259);
   U10563 : OAI22_X1 port map( A1 => n10675, A2 => n12884, B1 => n10548, B2 => 
                           n12881, ZN => n11266);
   U10564 : AOI221_X1 port map( B1 => n12842, B2 => n10136, C1 => n12839, C2 =>
                           n10040, A => n11274, ZN => n11267);
   U10565 : OAI22_X1 port map( A1 => n10579, A2 => n12836, B1 => n10452, B2 => 
                           n12833, ZN => n11274);
   U10566 : AOI221_X1 port map( B1 => n12890, B2 => n10279, C1 => n12887, C2 =>
                           n10255, A => n11247, ZN => n11240);
   U10567 : OAI22_X1 port map( A1 => n10674, A2 => n12884, B1 => n10547, B2 => 
                           n12881, ZN => n11247);
   U10568 : AOI221_X1 port map( B1 => n12842, B2 => n10135, C1 => n12839, C2 =>
                           n10039, A => n11255, ZN => n11248);
   U10569 : OAI22_X1 port map( A1 => n10578, A2 => n12836, B1 => n10451, B2 => 
                           n12833, ZN => n11255);
   U10570 : AOI221_X1 port map( B1 => n12890, B2 => n10278, C1 => n12887, C2 =>
                           n10254, A => n11228, ZN => n11221);
   U10571 : OAI22_X1 port map( A1 => n10673, A2 => n12884, B1 => n10546, B2 => 
                           n12881, ZN => n11228);
   U10572 : AOI221_X1 port map( B1 => n12842, B2 => n10134, C1 => n12839, C2 =>
                           n10038, A => n11236, ZN => n11229);
   U10573 : OAI22_X1 port map( A1 => n10577, A2 => n12836, B1 => n10450, B2 => 
                           n12833, ZN => n11236);
   U10574 : AOI221_X1 port map( B1 => n12890, B2 => n10277, C1 => n12887, C2 =>
                           n10253, A => n11209, ZN => n11202);
   U10575 : OAI22_X1 port map( A1 => n10672, A2 => n12884, B1 => n10545, B2 => 
                           n12881, ZN => n11209);
   U10576 : AOI221_X1 port map( B1 => n12842, B2 => n10133, C1 => n12839, C2 =>
                           n10037, A => n11217, ZN => n11210);
   U10577 : OAI22_X1 port map( A1 => n10576, A2 => n12836, B1 => n10449, B2 => 
                           n12833, ZN => n11217);
   U10578 : AOI221_X1 port map( B1 => n12890, B2 => n10276, C1 => n12887, C2 =>
                           n10252, A => n11190, ZN => n11183);
   U10579 : OAI22_X1 port map( A1 => n10671, A2 => n12884, B1 => n10544, B2 => 
                           n12881, ZN => n11190);
   U10580 : AOI221_X1 port map( B1 => n12842, B2 => n10132, C1 => n12839, C2 =>
                           n10036, A => n11198, ZN => n11191);
   U10581 : OAI22_X1 port map( A1 => n10575, A2 => n12836, B1 => n10448, B2 => 
                           n12833, ZN => n11198);
   U10582 : AOI221_X1 port map( B1 => n12890, B2 => n10275, C1 => n12887, C2 =>
                           n10251, A => n11171, ZN => n11164);
   U10583 : OAI22_X1 port map( A1 => n10670, A2 => n12884, B1 => n10543, B2 => 
                           n12881, ZN => n11171);
   U10584 : AOI221_X1 port map( B1 => n12842, B2 => n10131, C1 => n12839, C2 =>
                           n10035, A => n11179, ZN => n11172);
   U10585 : OAI22_X1 port map( A1 => n10574, A2 => n12836, B1 => n10447, B2 => 
                           n12833, ZN => n11179);
   U10586 : AOI221_X1 port map( B1 => n12891, B2 => n10114, C1 => n12888, C2 =>
                           n10106, A => n11152, ZN => n11145);
   U10587 : OAI22_X1 port map( A1 => n10442, A2 => n12885, B1 => n10394, B2 => 
                           n12882, ZN => n11152);
   U10588 : AOI221_X1 port map( B1 => n12843, B2 => n10066, C1 => n12840, C2 =>
                           n10034, A => n11160, ZN => n11153);
   U10589 : OAI22_X1 port map( A1 => n10410, A2 => n12837, B1 => n10362, B2 => 
                           n12834, ZN => n11160);
   U10590 : AOI221_X1 port map( B1 => n12891, B2 => n10113, C1 => n12888, C2 =>
                           n10105, A => n11133, ZN => n11126);
   U10591 : OAI22_X1 port map( A1 => n10441, A2 => n12885, B1 => n10393, B2 => 
                           n12882, ZN => n11133);
   U10592 : AOI221_X1 port map( B1 => n12843, B2 => n10065, C1 => n12840, C2 =>
                           n10033, A => n11141, ZN => n11134);
   U10593 : OAI22_X1 port map( A1 => n10409, A2 => n12837, B1 => n10361, B2 => 
                           n12834, ZN => n11141);
   U10594 : AOI221_X1 port map( B1 => n12891, B2 => n10112, C1 => n12888, C2 =>
                           n10104, A => n11114, ZN => n11107);
   U10595 : OAI22_X1 port map( A1 => n10440, A2 => n12885, B1 => n10392, B2 => 
                           n12882, ZN => n11114);
   U10596 : AOI221_X1 port map( B1 => n12843, B2 => n10064, C1 => n12840, C2 =>
                           n10032, A => n11122, ZN => n11115);
   U10597 : OAI22_X1 port map( A1 => n10408, A2 => n12837, B1 => n10360, B2 => 
                           n12834, ZN => n11122);
   U10598 : AOI221_X1 port map( B1 => n12891, B2 => n10111, C1 => n12888, C2 =>
                           n10103, A => n11095, ZN => n11088);
   U10599 : OAI22_X1 port map( A1 => n10439, A2 => n12885, B1 => n10391, B2 => 
                           n12882, ZN => n11095);
   U10600 : AOI221_X1 port map( B1 => n12843, B2 => n10063, C1 => n12840, C2 =>
                           n10031, A => n11103, ZN => n11096);
   U10601 : OAI22_X1 port map( A1 => n10407, A2 => n12837, B1 => n10359, B2 => 
                           n12834, ZN => n11103);
   U10602 : AOI221_X1 port map( B1 => n12891, B2 => n10110, C1 => n12888, C2 =>
                           n10102, A => n11076, ZN => n11069);
   U10603 : OAI22_X1 port map( A1 => n10438, A2 => n12885, B1 => n10390, B2 => 
                           n12882, ZN => n11076);
   U10604 : AOI221_X1 port map( B1 => n12843, B2 => n10062, C1 => n12840, C2 =>
                           n10030, A => n11084, ZN => n11077);
   U10605 : OAI22_X1 port map( A1 => n10406, A2 => n12837, B1 => n10358, B2 => 
                           n12834, ZN => n11084);
   U10606 : AOI221_X1 port map( B1 => n12891, B2 => n10109, C1 => n12888, C2 =>
                           n10101, A => n11057, ZN => n11050);
   U10607 : OAI22_X1 port map( A1 => n10437, A2 => n12885, B1 => n10389, B2 => 
                           n12882, ZN => n11057);
   U10608 : AOI221_X1 port map( B1 => n12843, B2 => n10061, C1 => n12840, C2 =>
                           n10029, A => n11065, ZN => n11058);
   U10609 : OAI22_X1 port map( A1 => n10405, A2 => n12837, B1 => n10357, B2 => 
                           n12834, ZN => n11065);
   U10610 : AOI221_X1 port map( B1 => n12891, B2 => n10108, C1 => n12888, C2 =>
                           n10100, A => n11038, ZN => n11031);
   U10611 : OAI22_X1 port map( A1 => n10436, A2 => n12885, B1 => n10388, B2 => 
                           n12882, ZN => n11038);
   U10612 : AOI221_X1 port map( B1 => n12843, B2 => n10060, C1 => n12840, C2 =>
                           n10028, A => n11046, ZN => n11039);
   U10613 : OAI22_X1 port map( A1 => n10404, A2 => n12837, B1 => n10356, B2 => 
                           n12834, ZN => n11046);
   U10614 : AOI221_X1 port map( B1 => n12891, B2 => n10107, C1 => n12888, C2 =>
                           n10099, A => n11001, ZN => n10980);
   U10615 : OAI22_X1 port map( A1 => n10435, A2 => n12885, B1 => n10387, B2 => 
                           n12882, ZN => n11001);
   U10616 : AOI221_X1 port map( B1 => n12843, B2 => n10059, C1 => n12840, C2 =>
                           n10027, A => n11025, ZN => n11004);
   U10617 : OAI22_X1 port map( A1 => n10403, A2 => n12837, B1 => n10355, B2 => 
                           n12834, ZN => n11025);
   U10618 : AOI221_X1 port map( B1 => n12825, B2 => n10122, C1 => n12822, C2 =>
                           n10130, A => n11802, ZN => n11801);
   U10619 : OAI22_X1 port map( A1 => n9942, A2 => n12819, B1 => n10402, B2 => 
                           n12816, ZN => n11802);
   U10620 : AOI221_X1 port map( B1 => n12813, B2 => n10874, C1 => n12810, C2 =>
                           n10842, A => n11803, ZN => n11800);
   U10621 : OAI22_X1 port map( A1 => n10002, A2 => n12807, B1 => n9970, B2 => 
                           n12804, ZN => n11803);
   U10622 : AOI221_X1 port map( B1 => n12753, B2 => n10082, C1 => n12750, C2 =>
                           n10074, A => n11812, ZN => n11807);
   U10623 : OAI22_X1 port map( A1 => n10418, A2 => n12747, B1 => n10370, B2 => 
                           n12744, ZN => n11812);
   U10624 : AOI221_X1 port map( B1 => n12825, B2 => n10121, C1 => n12822, C2 =>
                           n10129, A => n11783, ZN => n11782);
   U10625 : OAI22_X1 port map( A1 => n9941, A2 => n12819, B1 => n10401, B2 => 
                           n12816, ZN => n11783);
   U10626 : AOI221_X1 port map( B1 => n12813, B2 => n10873, C1 => n12810, C2 =>
                           n10841, A => n11784, ZN => n11781);
   U10627 : OAI22_X1 port map( A1 => n10001, A2 => n12807, B1 => n9969, B2 => 
                           n12804, ZN => n11784);
   U10628 : AOI221_X1 port map( B1 => n12753, B2 => n10081, C1 => n12750, C2 =>
                           n10073, A => n11793, ZN => n11788);
   U10629 : OAI22_X1 port map( A1 => n10417, A2 => n12747, B1 => n10369, B2 => 
                           n12744, ZN => n11793);
   U10630 : AOI221_X1 port map( B1 => n12825, B2 => n10120, C1 => n12822, C2 =>
                           n10128, A => n11764, ZN => n11763);
   U10631 : OAI22_X1 port map( A1 => n9940, A2 => n12819, B1 => n10400, B2 => 
                           n12816, ZN => n11764);
   U10632 : AOI221_X1 port map( B1 => n12813, B2 => n10872, C1 => n12810, C2 =>
                           n10840, A => n11765, ZN => n11762);
   U10633 : OAI22_X1 port map( A1 => n10000, A2 => n12807, B1 => n9968, B2 => 
                           n12804, ZN => n11765);
   U10634 : AOI221_X1 port map( B1 => n12753, B2 => n10080, C1 => n12750, C2 =>
                           n10072, A => n11774, ZN => n11769);
   U10635 : OAI22_X1 port map( A1 => n10416, A2 => n12747, B1 => n10368, B2 => 
                           n12744, ZN => n11774);
   U10636 : AOI221_X1 port map( B1 => n12825, B2 => n10119, C1 => n12822, C2 =>
                           n10127, A => n11745, ZN => n11744);
   U10637 : OAI22_X1 port map( A1 => n9939, A2 => n12819, B1 => n10399, B2 => 
                           n12816, ZN => n11745);
   U10638 : AOI221_X1 port map( B1 => n12813, B2 => n10871, C1 => n12810, C2 =>
                           n10839, A => n11746, ZN => n11743);
   U10639 : OAI22_X1 port map( A1 => n9999, A2 => n12807, B1 => n9967, B2 => 
                           n12804, ZN => n11746);
   U10640 : AOI221_X1 port map( B1 => n12753, B2 => n10079, C1 => n12750, C2 =>
                           n10071, A => n11755, ZN => n11750);
   U10641 : OAI22_X1 port map( A1 => n10415, A2 => n12747, B1 => n10367, B2 => 
                           n12744, ZN => n11755);
   U10642 : AOI221_X1 port map( B1 => n12825, B2 => n10118, C1 => n12822, C2 =>
                           n10126, A => n11726, ZN => n11725);
   U10643 : OAI22_X1 port map( A1 => n10570, A2 => n12819, B1 => n10398, B2 => 
                           n12816, ZN => n11726);
   U10644 : AOI221_X1 port map( B1 => n12813, B2 => n10870, C1 => n12810, C2 =>
                           n10838, A => n11727, ZN => n11724);
   U10645 : OAI22_X1 port map( A1 => n9998, A2 => n12807, B1 => n9966, B2 => 
                           n12804, ZN => n11727);
   U10646 : AOI221_X1 port map( B1 => n12753, B2 => n10078, C1 => n12750, C2 =>
                           n10070, A => n11736, ZN => n11731);
   U10647 : OAI22_X1 port map( A1 => n10414, A2 => n12747, B1 => n10366, B2 => 
                           n12744, ZN => n11736);
   U10648 : AOI221_X1 port map( B1 => n12825, B2 => n10117, C1 => n12822, C2 =>
                           n10125, A => n11707, ZN => n11706);
   U10649 : OAI22_X1 port map( A1 => n10569, A2 => n12819, B1 => n10397, B2 => 
                           n12816, ZN => n11707);
   U10650 : AOI221_X1 port map( B1 => n12813, B2 => n10869, C1 => n12810, C2 =>
                           n10837, A => n11708, ZN => n11705);
   U10651 : OAI22_X1 port map( A1 => n9997, A2 => n12807, B1 => n9965, B2 => 
                           n12804, ZN => n11708);
   U10652 : AOI221_X1 port map( B1 => n12753, B2 => n10077, C1 => n12750, C2 =>
                           n10069, A => n11717, ZN => n11712);
   U10653 : OAI22_X1 port map( A1 => n10413, A2 => n12747, B1 => n10365, B2 => 
                           n12744, ZN => n11717);
   U10654 : AOI221_X1 port map( B1 => n12825, B2 => n10116, C1 => n12822, C2 =>
                           n10124, A => n11688, ZN => n11687);
   U10655 : OAI22_X1 port map( A1 => n10568, A2 => n12819, B1 => n10396, B2 => 
                           n12816, ZN => n11688);
   U10656 : AOI221_X1 port map( B1 => n12813, B2 => n10868, C1 => n12810, C2 =>
                           n10836, A => n11689, ZN => n11686);
   U10657 : OAI22_X1 port map( A1 => n9996, A2 => n12807, B1 => n9964, B2 => 
                           n12804, ZN => n11689);
   U10658 : AOI221_X1 port map( B1 => n12753, B2 => n10076, C1 => n12750, C2 =>
                           n10068, A => n11698, ZN => n11693);
   U10659 : OAI22_X1 port map( A1 => n10412, A2 => n12747, B1 => n10364, B2 => 
                           n12744, ZN => n11698);
   U10660 : AOI221_X1 port map( B1 => n12825, B2 => n10115, C1 => n12822, C2 =>
                           n10123, A => n11639, ZN => n11636);
   U10661 : OAI22_X1 port map( A1 => n10567, A2 => n12819, B1 => n10395, B2 => 
                           n12816, ZN => n11639);
   U10662 : AOI221_X1 port map( B1 => n12813, B2 => n10867, C1 => n12810, C2 =>
                           n10835, A => n11644, ZN => n11635);
   U10663 : OAI22_X1 port map( A1 => n9995, A2 => n12807, B1 => n10347, B2 => 
                           n12804, ZN => n11644);
   U10664 : AOI221_X1 port map( B1 => n12753, B2 => n10075, C1 => n12750, C2 =>
                           n10067, A => n11673, ZN => n11658);
   U10665 : OAI22_X1 port map( A1 => n10411, A2 => n12747, B1 => n10363, B2 => 
                           n12744, ZN => n11673);
   U10666 : AOI221_X1 port map( B1 => n12915, B2 => n10874, C1 => n12912, C2 =>
                           n10842, A => n11150, ZN => n11147);
   U10667 : OAI22_X1 port map( A1 => n10002, A2 => n12909, B1 => n9970, B2 => 
                           n12906, ZN => n11150);
   U10668 : AOI221_X1 port map( B1 => n12915, B2 => n10873, C1 => n12912, C2 =>
                           n10841, A => n11131, ZN => n11128);
   U10669 : OAI22_X1 port map( A1 => n10001, A2 => n12909, B1 => n9969, B2 => 
                           n12906, ZN => n11131);
   U10670 : AOI221_X1 port map( B1 => n12915, B2 => n10872, C1 => n12912, C2 =>
                           n10840, A => n11112, ZN => n11109);
   U10671 : OAI22_X1 port map( A1 => n10000, A2 => n12909, B1 => n9968, B2 => 
                           n12906, ZN => n11112);
   U10672 : AOI221_X1 port map( B1 => n12915, B2 => n10871, C1 => n12912, C2 =>
                           n10839, A => n11093, ZN => n11090);
   U10673 : OAI22_X1 port map( A1 => n9999, A2 => n12909, B1 => n9967, B2 => 
                           n12906, ZN => n11093);
   U10674 : AOI221_X1 port map( B1 => n12915, B2 => n10870, C1 => n12912, C2 =>
                           n10838, A => n11074, ZN => n11071);
   U10675 : OAI22_X1 port map( A1 => n9998, A2 => n12909, B1 => n9966, B2 => 
                           n12906, ZN => n11074);
   U10676 : AOI221_X1 port map( B1 => n12915, B2 => n10869, C1 => n12912, C2 =>
                           n10837, A => n11055, ZN => n11052);
   U10677 : OAI22_X1 port map( A1 => n9997, A2 => n12909, B1 => n9965, B2 => 
                           n12906, ZN => n11055);
   U10678 : AOI221_X1 port map( B1 => n12915, B2 => n10868, C1 => n12912, C2 =>
                           n10836, A => n11036, ZN => n11033);
   U10679 : OAI22_X1 port map( A1 => n9996, A2 => n12909, B1 => n9964, B2 => 
                           n12906, ZN => n11036);
   U10680 : AOI221_X1 port map( B1 => n12915, B2 => n10867, C1 => n12912, C2 =>
                           n10835, A => n10991, ZN => n10982);
   U10681 : OAI22_X1 port map( A1 => n9995, A2 => n12909, B1 => n10347, B2 => 
                           n12906, ZN => n10991);
   U10682 : OAI22_X1 port map( A1 => n13313, A2 => n13298, B1 => n10900, B2 => 
                           n10570, ZN => n3610);
   U10683 : OAI22_X1 port map( A1 => n13313, A2 => n13301, B1 => n10900, B2 => 
                           n10569, ZN => n3611);
   U10684 : OAI22_X1 port map( A1 => n13314, A2 => n13304, B1 => n10900, B2 => 
                           n10568, ZN => n3612);
   U10685 : OAI22_X1 port map( A1 => n13314, A2 => n13316, B1 => n10900, B2 => 
                           n10567, ZN => n3613);
   U10686 : OAI22_X1 port map( A1 => n13084, A2 => n13287, B1 => n10957, B2 => 
                           n10442, ZN => n3126);
   U10687 : OAI22_X1 port map( A1 => n13085, A2 => n13290, B1 => n10957, B2 => 
                           n10441, ZN => n3127);
   U10688 : OAI22_X1 port map( A1 => n13085, A2 => n13293, B1 => n10957, B2 => 
                           n10440, ZN => n3128);
   U10689 : OAI22_X1 port map( A1 => n13085, A2 => n13296, B1 => n10957, B2 => 
                           n10439, ZN => n3129);
   U10690 : OAI22_X1 port map( A1 => n13085, A2 => n13299, B1 => n10957, B2 => 
                           n10438, ZN => n3130);
   U10691 : OAI22_X1 port map( A1 => n13085, A2 => n13302, B1 => n10957, B2 => 
                           n10437, ZN => n3131);
   U10692 : OAI22_X1 port map( A1 => n13086, A2 => n13305, B1 => n10957, B2 => 
                           n10436, ZN => n3132);
   U10693 : OAI22_X1 port map( A1 => n13086, A2 => n13317, B1 => n10957, B2 => 
                           n10435, ZN => n3133);
   U10694 : OAI22_X1 port map( A1 => n13012, A2 => n13287, B1 => n10966, B2 => 
                           n10426, ZN => n2870);
   U10695 : OAI22_X1 port map( A1 => n13013, A2 => n13290, B1 => n10966, B2 => 
                           n10425, ZN => n2871);
   U10696 : OAI22_X1 port map( A1 => n13013, A2 => n13293, B1 => n10966, B2 => 
                           n10424, ZN => n2872);
   U10697 : OAI22_X1 port map( A1 => n13013, A2 => n13296, B1 => n10966, B2 => 
                           n10423, ZN => n2873);
   U10698 : OAI22_X1 port map( A1 => n13013, A2 => n13299, B1 => n10966, B2 => 
                           n10422, ZN => n2874);
   U10699 : OAI22_X1 port map( A1 => n13013, A2 => n13302, B1 => n10966, B2 => 
                           n10421, ZN => n2875);
   U10700 : OAI22_X1 port map( A1 => n13014, A2 => n13305, B1 => n10966, B2 => 
                           n10420, ZN => n2876);
   U10701 : OAI22_X1 port map( A1 => n13014, A2 => n13317, B1 => n10966, B2 => 
                           n10419, ZN => n2877);
   U10702 : OAI22_X1 port map( A1 => n12994, A2 => n13288, B1 => n10969, B2 => 
                           n10418, ZN => n2806);
   U10703 : OAI22_X1 port map( A1 => n12995, A2 => n13291, B1 => n10969, B2 => 
                           n10417, ZN => n2807);
   U10704 : OAI22_X1 port map( A1 => n12995, A2 => n13294, B1 => n10969, B2 => 
                           n10416, ZN => n2808);
   U10705 : OAI22_X1 port map( A1 => n12995, A2 => n13297, B1 => n10969, B2 => 
                           n10415, ZN => n2809);
   U10706 : OAI22_X1 port map( A1 => n12995, A2 => n13300, B1 => n10969, B2 => 
                           n10414, ZN => n2810);
   U10707 : OAI22_X1 port map( A1 => n12995, A2 => n13303, B1 => n10969, B2 => 
                           n10413, ZN => n2811);
   U10708 : OAI22_X1 port map( A1 => n12996, A2 => n13306, B1 => n10969, B2 => 
                           n10412, ZN => n2812);
   U10709 : OAI22_X1 port map( A1 => n12996, A2 => n13318, B1 => n10969, B2 => 
                           n10411, ZN => n2813);
   U10710 : OAI22_X1 port map( A1 => n12958, A2 => n13288, B1 => n10973, B2 => 
                           n10410, ZN => n2678);
   U10711 : OAI22_X1 port map( A1 => n12959, A2 => n13291, B1 => n10973, B2 => 
                           n10409, ZN => n2679);
   U10712 : OAI22_X1 port map( A1 => n12959, A2 => n13294, B1 => n10973, B2 => 
                           n10408, ZN => n2680);
   U10713 : OAI22_X1 port map( A1 => n12959, A2 => n13297, B1 => n10973, B2 => 
                           n10407, ZN => n2681);
   U10714 : OAI22_X1 port map( A1 => n12959, A2 => n13300, B1 => n10973, B2 => 
                           n10406, ZN => n2682);
   U10715 : OAI22_X1 port map( A1 => n12959, A2 => n13303, B1 => n10973, B2 => 
                           n10405, ZN => n2683);
   U10716 : OAI22_X1 port map( A1 => n12960, A2 => n13306, B1 => n10973, B2 => 
                           n10404, ZN => n2684);
   U10717 : OAI22_X1 port map( A1 => n12960, A2 => n13318, B1 => n10973, B2 => 
                           n10403, ZN => n2685);
   U10718 : OAI22_X1 port map( A1 => n13210, A2 => n13286, B1 => n10934, B2 => 
                           n10402, ZN => n3574);
   U10719 : OAI22_X1 port map( A1 => n13211, A2 => n13289, B1 => n10934, B2 => 
                           n10401, ZN => n3575);
   U10720 : OAI22_X1 port map( A1 => n13211, A2 => n13292, B1 => n10934, B2 => 
                           n10400, ZN => n3576);
   U10721 : OAI22_X1 port map( A1 => n13211, A2 => n13295, B1 => n10934, B2 => 
                           n10399, ZN => n3577);
   U10722 : OAI22_X1 port map( A1 => n13211, A2 => n13298, B1 => n10934, B2 => 
                           n10398, ZN => n3578);
   U10723 : OAI22_X1 port map( A1 => n13211, A2 => n13301, B1 => n10934, B2 => 
                           n10397, ZN => n3579);
   U10724 : OAI22_X1 port map( A1 => n13212, A2 => n13304, B1 => n10934, B2 => 
                           n10396, ZN => n3580);
   U10725 : OAI22_X1 port map( A1 => n13212, A2 => n13316, B1 => n10934, B2 => 
                           n10395, ZN => n3581);
   U10726 : OAI22_X1 port map( A1 => n13093, A2 => n13287, B1 => n10956, B2 => 
                           n10394, ZN => n3158);
   U10727 : OAI22_X1 port map( A1 => n13094, A2 => n13290, B1 => n10956, B2 => 
                           n10393, ZN => n3159);
   U10728 : OAI22_X1 port map( A1 => n13094, A2 => n13293, B1 => n10956, B2 => 
                           n10392, ZN => n3160);
   U10729 : OAI22_X1 port map( A1 => n13094, A2 => n13296, B1 => n10956, B2 => 
                           n10391, ZN => n3161);
   U10730 : OAI22_X1 port map( A1 => n13094, A2 => n13299, B1 => n10956, B2 => 
                           n10390, ZN => n3162);
   U10731 : OAI22_X1 port map( A1 => n13094, A2 => n13302, B1 => n10956, B2 => 
                           n10389, ZN => n3163);
   U10732 : OAI22_X1 port map( A1 => n13095, A2 => n13305, B1 => n10956, B2 => 
                           n10388, ZN => n3164);
   U10733 : OAI22_X1 port map( A1 => n13095, A2 => n13317, B1 => n10956, B2 => 
                           n10387, ZN => n3165);
   U10734 : OAI22_X1 port map( A1 => n13021, A2 => n13287, B1 => n10965, B2 => 
                           n10378, ZN => n2902);
   U10735 : OAI22_X1 port map( A1 => n13022, A2 => n13290, B1 => n10965, B2 => 
                           n10377, ZN => n2903);
   U10736 : OAI22_X1 port map( A1 => n13022, A2 => n13293, B1 => n10965, B2 => 
                           n10376, ZN => n2904);
   U10737 : OAI22_X1 port map( A1 => n13022, A2 => n13296, B1 => n10965, B2 => 
                           n10375, ZN => n2905);
   U10738 : OAI22_X1 port map( A1 => n13022, A2 => n13299, B1 => n10965, B2 => 
                           n10374, ZN => n2906);
   U10739 : OAI22_X1 port map( A1 => n13022, A2 => n13302, B1 => n10965, B2 => 
                           n10373, ZN => n2907);
   U10740 : OAI22_X1 port map( A1 => n13023, A2 => n13305, B1 => n10965, B2 => 
                           n10372, ZN => n2908);
   U10741 : OAI22_X1 port map( A1 => n13023, A2 => n13317, B1 => n10965, B2 => 
                           n10371, ZN => n2909);
   U10742 : OAI22_X1 port map( A1 => n13003, A2 => n13288, B1 => n10967, B2 => 
                           n10370, ZN => n2838);
   U10743 : OAI22_X1 port map( A1 => n13004, A2 => n13291, B1 => n10967, B2 => 
                           n10369, ZN => n2839);
   U10744 : OAI22_X1 port map( A1 => n13004, A2 => n13294, B1 => n10967, B2 => 
                           n10368, ZN => n2840);
   U10745 : OAI22_X1 port map( A1 => n13004, A2 => n13297, B1 => n10967, B2 => 
                           n10367, ZN => n2841);
   U10746 : OAI22_X1 port map( A1 => n13004, A2 => n13300, B1 => n10967, B2 => 
                           n10366, ZN => n2842);
   U10747 : OAI22_X1 port map( A1 => n13004, A2 => n13303, B1 => n10967, B2 => 
                           n10365, ZN => n2843);
   U10748 : OAI22_X1 port map( A1 => n13005, A2 => n13306, B1 => n10967, B2 => 
                           n10364, ZN => n2844);
   U10749 : OAI22_X1 port map( A1 => n13005, A2 => n13318, B1 => n10967, B2 => 
                           n10363, ZN => n2845);
   U10750 : OAI22_X1 port map( A1 => n12967, A2 => n13288, B1 => n10972, B2 => 
                           n10362, ZN => n2710);
   U10751 : OAI22_X1 port map( A1 => n12968, A2 => n13291, B1 => n10972, B2 => 
                           n10361, ZN => n2711);
   U10752 : OAI22_X1 port map( A1 => n12968, A2 => n13294, B1 => n10972, B2 => 
                           n10360, ZN => n2712);
   U10753 : OAI22_X1 port map( A1 => n12968, A2 => n13297, B1 => n10972, B2 => 
                           n10359, ZN => n2713);
   U10754 : OAI22_X1 port map( A1 => n12968, A2 => n13300, B1 => n10972, B2 => 
                           n10358, ZN => n2714);
   U10755 : OAI22_X1 port map( A1 => n12968, A2 => n13303, B1 => n10972, B2 => 
                           n10357, ZN => n2715);
   U10756 : OAI22_X1 port map( A1 => n12969, A2 => n13306, B1 => n10972, B2 => 
                           n10356, ZN => n2716);
   U10757 : OAI22_X1 port map( A1 => n12969, A2 => n13318, B1 => n10972, B2 => 
                           n10355, ZN => n2717);
   U10758 : OAI22_X1 port map( A1 => n13167, A2 => n13316, B1 => n10944, B2 => 
                           n10347, ZN => n3421);
   U10759 : OAI22_X1 port map( A1 => n13156, A2 => n13286, B1 => n10946, B2 => 
                           n10002, ZN => n3382);
   U10760 : OAI22_X1 port map( A1 => n13157, A2 => n13289, B1 => n10946, B2 => 
                           n10001, ZN => n3383);
   U10761 : OAI22_X1 port map( A1 => n13157, A2 => n13292, B1 => n10946, B2 => 
                           n10000, ZN => n3384);
   U10762 : OAI22_X1 port map( A1 => n13157, A2 => n13295, B1 => n10946, B2 => 
                           n9999, ZN => n3385);
   U10763 : OAI22_X1 port map( A1 => n13157, A2 => n13298, B1 => n10946, B2 => 
                           n9998, ZN => n3386);
   U10764 : OAI22_X1 port map( A1 => n13157, A2 => n13301, B1 => n10946, B2 => 
                           n9997, ZN => n3387);
   U10765 : OAI22_X1 port map( A1 => n13158, A2 => n13304, B1 => n10946, B2 => 
                           n9996, ZN => n3388);
   U10766 : OAI22_X1 port map( A1 => n13158, A2 => n13316, B1 => n10946, B2 => 
                           n9995, ZN => n3389);
   U10767 : OAI22_X1 port map( A1 => n13165, A2 => n13286, B1 => n10944, B2 => 
                           n9970, ZN => n3414);
   U10768 : OAI22_X1 port map( A1 => n13166, A2 => n13289, B1 => n10944, B2 => 
                           n9969, ZN => n3415);
   U10769 : OAI22_X1 port map( A1 => n13166, A2 => n13292, B1 => n10944, B2 => 
                           n9968, ZN => n3416);
   U10770 : OAI22_X1 port map( A1 => n13166, A2 => n13295, B1 => n10944, B2 => 
                           n9967, ZN => n3417);
   U10771 : OAI22_X1 port map( A1 => n13166, A2 => n13298, B1 => n10944, B2 => 
                           n9966, ZN => n3418);
   U10772 : OAI22_X1 port map( A1 => n13166, A2 => n13301, B1 => n10944, B2 => 
                           n9965, ZN => n3419);
   U10773 : OAI22_X1 port map( A1 => n13167, A2 => n13304, B1 => n10944, B2 => 
                           n9964, ZN => n3420);
   U10774 : OAI22_X1 port map( A1 => n13312, A2 => n13286, B1 => n10900, B2 => 
                           n9942, ZN => n3606);
   U10775 : OAI22_X1 port map( A1 => n13313, A2 => n13289, B1 => n10900, B2 => 
                           n9941, ZN => n3607);
   U10776 : OAI22_X1 port map( A1 => n13313, A2 => n13292, B1 => n10900, B2 => 
                           n9940, ZN => n3608);
   U10777 : OAI22_X1 port map( A1 => n13313, A2 => n13295, B1 => n10900, B2 => 
                           n9939, ZN => n3609);
   U10778 : OAI22_X1 port map( A1 => n13308, A2 => n13214, B1 => n13307, B2 => 
                           n10706, ZN => n3582);
   U10779 : OAI22_X1 port map( A1 => n13309, A2 => n13238, B1 => n13307, B2 => 
                           n10705, ZN => n3590);
   U10780 : OAI22_X1 port map( A1 => n13309, A2 => n13241, B1 => n13307, B2 => 
                           n10704, ZN => n3591);
   U10781 : OAI22_X1 port map( A1 => n13310, A2 => n13244, B1 => n13307, B2 => 
                           n10703, ZN => n3592);
   U10782 : OAI22_X1 port map( A1 => n13310, A2 => n13247, B1 => n13307, B2 => 
                           n10702, ZN => n3593);
   U10783 : OAI22_X1 port map( A1 => n13310, A2 => n13250, B1 => n10900, B2 => 
                           n10701, ZN => n3594);
   U10784 : OAI22_X1 port map( A1 => n13310, A2 => n13253, B1 => n10900, B2 => 
                           n10700, ZN => n3595);
   U10785 : OAI22_X1 port map( A1 => n13310, A2 => n13256, B1 => n10900, B2 => 
                           n10699, ZN => n3596);
   U10786 : OAI22_X1 port map( A1 => n13311, A2 => n13259, B1 => n13307, B2 => 
                           n10698, ZN => n3597);
   U10787 : OAI22_X1 port map( A1 => n13311, A2 => n13262, B1 => n13307, B2 => 
                           n10697, ZN => n3598);
   U10788 : OAI22_X1 port map( A1 => n13311, A2 => n13265, B1 => n13307, B2 => 
                           n10696, ZN => n3599);
   U10789 : OAI22_X1 port map( A1 => n13311, A2 => n13268, B1 => n13307, B2 => 
                           n10695, ZN => n3600);
   U10790 : OAI22_X1 port map( A1 => n13311, A2 => n13271, B1 => n13307, B2 => 
                           n10694, ZN => n3601);
   U10791 : OAI22_X1 port map( A1 => n13080, A2 => n13215, B1 => n13079, B2 => 
                           n10693, ZN => n3102);
   U10792 : OAI22_X1 port map( A1 => n13080, A2 => n13218, B1 => n13079, B2 => 
                           n10692, ZN => n3103);
   U10793 : OAI22_X1 port map( A1 => n13080, A2 => n13221, B1 => n13079, B2 => 
                           n10691, ZN => n3104);
   U10794 : OAI22_X1 port map( A1 => n13080, A2 => n13224, B1 => n13079, B2 => 
                           n10690, ZN => n3105);
   U10795 : OAI22_X1 port map( A1 => n13080, A2 => n13227, B1 => n13079, B2 => 
                           n10689, ZN => n3106);
   U10796 : OAI22_X1 port map( A1 => n13081, A2 => n13230, B1 => n13079, B2 => 
                           n10688, ZN => n3107);
   U10797 : OAI22_X1 port map( A1 => n13081, A2 => n13233, B1 => n13079, B2 => 
                           n10687, ZN => n3108);
   U10798 : OAI22_X1 port map( A1 => n13081, A2 => n13236, B1 => n13079, B2 => 
                           n10686, ZN => n3109);
   U10799 : OAI22_X1 port map( A1 => n13081, A2 => n13239, B1 => n13079, B2 => 
                           n10685, ZN => n3110);
   U10800 : OAI22_X1 port map( A1 => n13081, A2 => n13242, B1 => n13079, B2 => 
                           n10684, ZN => n3111);
   U10801 : OAI22_X1 port map( A1 => n13082, A2 => n13245, B1 => n13079, B2 => 
                           n10683, ZN => n3112);
   U10802 : OAI22_X1 port map( A1 => n13082, A2 => n13248, B1 => n13079, B2 => 
                           n10682, ZN => n3113);
   U10803 : OAI22_X1 port map( A1 => n13082, A2 => n13251, B1 => n10957, B2 => 
                           n10681, ZN => n3114);
   U10804 : OAI22_X1 port map( A1 => n13082, A2 => n13254, B1 => n10957, B2 => 
                           n10680, ZN => n3115);
   U10805 : OAI22_X1 port map( A1 => n13082, A2 => n13257, B1 => n10957, B2 => 
                           n10679, ZN => n3116);
   U10806 : OAI22_X1 port map( A1 => n13083, A2 => n13260, B1 => n13079, B2 => 
                           n10678, ZN => n3117);
   U10807 : OAI22_X1 port map( A1 => n13083, A2 => n13263, B1 => n13079, B2 => 
                           n10677, ZN => n3118);
   U10808 : OAI22_X1 port map( A1 => n13083, A2 => n13266, B1 => n13079, B2 => 
                           n10676, ZN => n3119);
   U10809 : OAI22_X1 port map( A1 => n13083, A2 => n13269, B1 => n13079, B2 => 
                           n10675, ZN => n3120);
   U10810 : OAI22_X1 port map( A1 => n13083, A2 => n13272, B1 => n13079, B2 => 
                           n10674, ZN => n3121);
   U10811 : OAI22_X1 port map( A1 => n13084, A2 => n13275, B1 => n13079, B2 => 
                           n10673, ZN => n3122);
   U10812 : OAI22_X1 port map( A1 => n13084, A2 => n13278, B1 => n13079, B2 => 
                           n10672, ZN => n3123);
   U10813 : OAI22_X1 port map( A1 => n13084, A2 => n13281, B1 => n13079, B2 => 
                           n10671, ZN => n3124);
   U10814 : OAI22_X1 port map( A1 => n13084, A2 => n13284, B1 => n13079, B2 => 
                           n10670, ZN => n3125);
   U10815 : OAI22_X1 port map( A1 => n13008, A2 => n13215, B1 => n13007, B2 => 
                           n10645, ZN => n2846);
   U10816 : OAI22_X1 port map( A1 => n13008, A2 => n13218, B1 => n13007, B2 => 
                           n10644, ZN => n2847);
   U10817 : OAI22_X1 port map( A1 => n13008, A2 => n13221, B1 => n13007, B2 => 
                           n10643, ZN => n2848);
   U10818 : OAI22_X1 port map( A1 => n13008, A2 => n13224, B1 => n13007, B2 => 
                           n10642, ZN => n2849);
   U10819 : OAI22_X1 port map( A1 => n13008, A2 => n13227, B1 => n13007, B2 => 
                           n10641, ZN => n2850);
   U10820 : OAI22_X1 port map( A1 => n13009, A2 => n13230, B1 => n13007, B2 => 
                           n10640, ZN => n2851);
   U10821 : OAI22_X1 port map( A1 => n13009, A2 => n13233, B1 => n13007, B2 => 
                           n10639, ZN => n2852);
   U10822 : OAI22_X1 port map( A1 => n13009, A2 => n13236, B1 => n13007, B2 => 
                           n10638, ZN => n2853);
   U10823 : OAI22_X1 port map( A1 => n13009, A2 => n13239, B1 => n13007, B2 => 
                           n10637, ZN => n2854);
   U10824 : OAI22_X1 port map( A1 => n13009, A2 => n13242, B1 => n13007, B2 => 
                           n10636, ZN => n2855);
   U10825 : OAI22_X1 port map( A1 => n13010, A2 => n13245, B1 => n13007, B2 => 
                           n10635, ZN => n2856);
   U10826 : OAI22_X1 port map( A1 => n13010, A2 => n13248, B1 => n13007, B2 => 
                           n10634, ZN => n2857);
   U10827 : OAI22_X1 port map( A1 => n13010, A2 => n13251, B1 => n10966, B2 => 
                           n10633, ZN => n2858);
   U10828 : OAI22_X1 port map( A1 => n13010, A2 => n13254, B1 => n10966, B2 => 
                           n10632, ZN => n2859);
   U10829 : OAI22_X1 port map( A1 => n13010, A2 => n13257, B1 => n10966, B2 => 
                           n10631, ZN => n2860);
   U10830 : OAI22_X1 port map( A1 => n13011, A2 => n13260, B1 => n13007, B2 => 
                           n10630, ZN => n2861);
   U10831 : OAI22_X1 port map( A1 => n13011, A2 => n13263, B1 => n13007, B2 => 
                           n10629, ZN => n2862);
   U10832 : OAI22_X1 port map( A1 => n13011, A2 => n13266, B1 => n13007, B2 => 
                           n10628, ZN => n2863);
   U10833 : OAI22_X1 port map( A1 => n13011, A2 => n13269, B1 => n13007, B2 => 
                           n10627, ZN => n2864);
   U10834 : OAI22_X1 port map( A1 => n13011, A2 => n13272, B1 => n13007, B2 => 
                           n10626, ZN => n2865);
   U10835 : OAI22_X1 port map( A1 => n13012, A2 => n13275, B1 => n13007, B2 => 
                           n10625, ZN => n2866);
   U10836 : OAI22_X1 port map( A1 => n13012, A2 => n13278, B1 => n13007, B2 => 
                           n10624, ZN => n2867);
   U10837 : OAI22_X1 port map( A1 => n13012, A2 => n13281, B1 => n13007, B2 => 
                           n10623, ZN => n2868);
   U10838 : OAI22_X1 port map( A1 => n13012, A2 => n13284, B1 => n13007, B2 => 
                           n10622, ZN => n2869);
   U10839 : OAI22_X1 port map( A1 => n12990, A2 => n13216, B1 => n12989, B2 => 
                           n10621, ZN => n2782);
   U10840 : OAI22_X1 port map( A1 => n12990, A2 => n13219, B1 => n12989, B2 => 
                           n10620, ZN => n2783);
   U10841 : OAI22_X1 port map( A1 => n12990, A2 => n13222, B1 => n12989, B2 => 
                           n10619, ZN => n2784);
   U10842 : OAI22_X1 port map( A1 => n12990, A2 => n13225, B1 => n12989, B2 => 
                           n10618, ZN => n2785);
   U10843 : OAI22_X1 port map( A1 => n12990, A2 => n13228, B1 => n12989, B2 => 
                           n10617, ZN => n2786);
   U10844 : OAI22_X1 port map( A1 => n12991, A2 => n13231, B1 => n12989, B2 => 
                           n10616, ZN => n2787);
   U10845 : OAI22_X1 port map( A1 => n12991, A2 => n13234, B1 => n12989, B2 => 
                           n10615, ZN => n2788);
   U10846 : OAI22_X1 port map( A1 => n12991, A2 => n13237, B1 => n12989, B2 => 
                           n10614, ZN => n2789);
   U10847 : OAI22_X1 port map( A1 => n12991, A2 => n13240, B1 => n12989, B2 => 
                           n10613, ZN => n2790);
   U10848 : OAI22_X1 port map( A1 => n12991, A2 => n13243, B1 => n12989, B2 => 
                           n10612, ZN => n2791);
   U10849 : OAI22_X1 port map( A1 => n12992, A2 => n13246, B1 => n12989, B2 => 
                           n10611, ZN => n2792);
   U10850 : OAI22_X1 port map( A1 => n12992, A2 => n13249, B1 => n12989, B2 => 
                           n10610, ZN => n2793);
   U10851 : OAI22_X1 port map( A1 => n12992, A2 => n13252, B1 => n10969, B2 => 
                           n10609, ZN => n2794);
   U10852 : OAI22_X1 port map( A1 => n12992, A2 => n13255, B1 => n10969, B2 => 
                           n10608, ZN => n2795);
   U10853 : OAI22_X1 port map( A1 => n12992, A2 => n13258, B1 => n10969, B2 => 
                           n10607, ZN => n2796);
   U10854 : OAI22_X1 port map( A1 => n12993, A2 => n13261, B1 => n12989, B2 => 
                           n10606, ZN => n2797);
   U10855 : OAI22_X1 port map( A1 => n12993, A2 => n13264, B1 => n12989, B2 => 
                           n10605, ZN => n2798);
   U10856 : OAI22_X1 port map( A1 => n12993, A2 => n13267, B1 => n12989, B2 => 
                           n10604, ZN => n2799);
   U10857 : OAI22_X1 port map( A1 => n12993, A2 => n13270, B1 => n12989, B2 => 
                           n10603, ZN => n2800);
   U10858 : OAI22_X1 port map( A1 => n12993, A2 => n13273, B1 => n12989, B2 => 
                           n10602, ZN => n2801);
   U10859 : OAI22_X1 port map( A1 => n12994, A2 => n13276, B1 => n12989, B2 => 
                           n10601, ZN => n2802);
   U10860 : OAI22_X1 port map( A1 => n12994, A2 => n13279, B1 => n12989, B2 => 
                           n10600, ZN => n2803);
   U10861 : OAI22_X1 port map( A1 => n12994, A2 => n13282, B1 => n12989, B2 => 
                           n10599, ZN => n2804);
   U10862 : OAI22_X1 port map( A1 => n12994, A2 => n13285, B1 => n12989, B2 => 
                           n10598, ZN => n2805);
   U10863 : OAI22_X1 port map( A1 => n12954, A2 => n13216, B1 => n12953, B2 => 
                           n10597, ZN => n2654);
   U10864 : OAI22_X1 port map( A1 => n12954, A2 => n13219, B1 => n12953, B2 => 
                           n10596, ZN => n2655);
   U10865 : OAI22_X1 port map( A1 => n12954, A2 => n13222, B1 => n12953, B2 => 
                           n10595, ZN => n2656);
   U10866 : OAI22_X1 port map( A1 => n12954, A2 => n13225, B1 => n12953, B2 => 
                           n10594, ZN => n2657);
   U10867 : OAI22_X1 port map( A1 => n12954, A2 => n13228, B1 => n12953, B2 => 
                           n10593, ZN => n2658);
   U10868 : OAI22_X1 port map( A1 => n12955, A2 => n13231, B1 => n12953, B2 => 
                           n10592, ZN => n2659);
   U10869 : OAI22_X1 port map( A1 => n12955, A2 => n13234, B1 => n12953, B2 => 
                           n10591, ZN => n2660);
   U10870 : OAI22_X1 port map( A1 => n12955, A2 => n13237, B1 => n12953, B2 => 
                           n10590, ZN => n2661);
   U10871 : OAI22_X1 port map( A1 => n12955, A2 => n13240, B1 => n12953, B2 => 
                           n10589, ZN => n2662);
   U10872 : OAI22_X1 port map( A1 => n12955, A2 => n13243, B1 => n12953, B2 => 
                           n10588, ZN => n2663);
   U10873 : OAI22_X1 port map( A1 => n12956, A2 => n13246, B1 => n12953, B2 => 
                           n10587, ZN => n2664);
   U10874 : OAI22_X1 port map( A1 => n12956, A2 => n13249, B1 => n12953, B2 => 
                           n10586, ZN => n2665);
   U10875 : OAI22_X1 port map( A1 => n12956, A2 => n13252, B1 => n10973, B2 => 
                           n10585, ZN => n2666);
   U10876 : OAI22_X1 port map( A1 => n12956, A2 => n13255, B1 => n10973, B2 => 
                           n10584, ZN => n2667);
   U10877 : OAI22_X1 port map( A1 => n12956, A2 => n13258, B1 => n10973, B2 => 
                           n10583, ZN => n2668);
   U10878 : OAI22_X1 port map( A1 => n12957, A2 => n13261, B1 => n12953, B2 => 
                           n10582, ZN => n2669);
   U10879 : OAI22_X1 port map( A1 => n12957, A2 => n13264, B1 => n12953, B2 => 
                           n10581, ZN => n2670);
   U10880 : OAI22_X1 port map( A1 => n12957, A2 => n13267, B1 => n12953, B2 => 
                           n10580, ZN => n2671);
   U10881 : OAI22_X1 port map( A1 => n12957, A2 => n13270, B1 => n12953, B2 => 
                           n10579, ZN => n2672);
   U10882 : OAI22_X1 port map( A1 => n12957, A2 => n13273, B1 => n12953, B2 => 
                           n10578, ZN => n2673);
   U10883 : OAI22_X1 port map( A1 => n12958, A2 => n13276, B1 => n12953, B2 => 
                           n10577, ZN => n2674);
   U10884 : OAI22_X1 port map( A1 => n12958, A2 => n13279, B1 => n12953, B2 => 
                           n10576, ZN => n2675);
   U10885 : OAI22_X1 port map( A1 => n12958, A2 => n13282, B1 => n12953, B2 => 
                           n10575, ZN => n2676);
   U10886 : OAI22_X1 port map( A1 => n12958, A2 => n13285, B1 => n12953, B2 => 
                           n10574, ZN => n2677);
   U10887 : OAI22_X1 port map( A1 => n13312, A2 => n13274, B1 => n13307, B2 => 
                           n10573, ZN => n3602);
   U10888 : OAI22_X1 port map( A1 => n13312, A2 => n13277, B1 => n13307, B2 => 
                           n10572, ZN => n3603);
   U10889 : OAI22_X1 port map( A1 => n13312, A2 => n13280, B1 => n13307, B2 => 
                           n10571, ZN => n3604);
   U10890 : OAI22_X1 port map( A1 => n13089, A2 => n13215, B1 => n13088, B2 => 
                           n10566, ZN => n3134);
   U10891 : OAI22_X1 port map( A1 => n13089, A2 => n13218, B1 => n13088, B2 => 
                           n10565, ZN => n3135);
   U10892 : OAI22_X1 port map( A1 => n13089, A2 => n13221, B1 => n13088, B2 => 
                           n10564, ZN => n3136);
   U10893 : OAI22_X1 port map( A1 => n13089, A2 => n13224, B1 => n13088, B2 => 
                           n10563, ZN => n3137);
   U10894 : OAI22_X1 port map( A1 => n13089, A2 => n13227, B1 => n13088, B2 => 
                           n10562, ZN => n3138);
   U10895 : OAI22_X1 port map( A1 => n13090, A2 => n13230, B1 => n13088, B2 => 
                           n10561, ZN => n3139);
   U10896 : OAI22_X1 port map( A1 => n13090, A2 => n13233, B1 => n13088, B2 => 
                           n10560, ZN => n3140);
   U10897 : OAI22_X1 port map( A1 => n13090, A2 => n13236, B1 => n13088, B2 => 
                           n10559, ZN => n3141);
   U10898 : OAI22_X1 port map( A1 => n13090, A2 => n13239, B1 => n13088, B2 => 
                           n10558, ZN => n3142);
   U10899 : OAI22_X1 port map( A1 => n13090, A2 => n13242, B1 => n13088, B2 => 
                           n10557, ZN => n3143);
   U10900 : OAI22_X1 port map( A1 => n13091, A2 => n13245, B1 => n13088, B2 => 
                           n10556, ZN => n3144);
   U10901 : OAI22_X1 port map( A1 => n13091, A2 => n13248, B1 => n13088, B2 => 
                           n10555, ZN => n3145);
   U10902 : OAI22_X1 port map( A1 => n13091, A2 => n13251, B1 => n10956, B2 => 
                           n10554, ZN => n3146);
   U10903 : OAI22_X1 port map( A1 => n13091, A2 => n13254, B1 => n10956, B2 => 
                           n10553, ZN => n3147);
   U10904 : OAI22_X1 port map( A1 => n13091, A2 => n13257, B1 => n10956, B2 => 
                           n10552, ZN => n3148);
   U10905 : OAI22_X1 port map( A1 => n13092, A2 => n13260, B1 => n13088, B2 => 
                           n10551, ZN => n3149);
   U10906 : OAI22_X1 port map( A1 => n13092, A2 => n13263, B1 => n13088, B2 => 
                           n10550, ZN => n3150);
   U10907 : OAI22_X1 port map( A1 => n13092, A2 => n13266, B1 => n13088, B2 => 
                           n10549, ZN => n3151);
   U10908 : OAI22_X1 port map( A1 => n13092, A2 => n13269, B1 => n13088, B2 => 
                           n10548, ZN => n3152);
   U10909 : OAI22_X1 port map( A1 => n13092, A2 => n13272, B1 => n13088, B2 => 
                           n10547, ZN => n3153);
   U10910 : OAI22_X1 port map( A1 => n13093, A2 => n13275, B1 => n13088, B2 => 
                           n10546, ZN => n3154);
   U10911 : OAI22_X1 port map( A1 => n13093, A2 => n13278, B1 => n13088, B2 => 
                           n10545, ZN => n3155);
   U10912 : OAI22_X1 port map( A1 => n13093, A2 => n13281, B1 => n13088, B2 => 
                           n10544, ZN => n3156);
   U10913 : OAI22_X1 port map( A1 => n13093, A2 => n13284, B1 => n13088, B2 => 
                           n10543, ZN => n3157);
   U10914 : OAI22_X1 port map( A1 => n13017, A2 => n13215, B1 => n13016, B2 => 
                           n10518, ZN => n2878);
   U10915 : OAI22_X1 port map( A1 => n13017, A2 => n13218, B1 => n13016, B2 => 
                           n10517, ZN => n2879);
   U10916 : OAI22_X1 port map( A1 => n13017, A2 => n13221, B1 => n13016, B2 => 
                           n10516, ZN => n2880);
   U10917 : OAI22_X1 port map( A1 => n13017, A2 => n13224, B1 => n13016, B2 => 
                           n10515, ZN => n2881);
   U10918 : OAI22_X1 port map( A1 => n13017, A2 => n13227, B1 => n13016, B2 => 
                           n10514, ZN => n2882);
   U10919 : OAI22_X1 port map( A1 => n13018, A2 => n13230, B1 => n13016, B2 => 
                           n10513, ZN => n2883);
   U10920 : OAI22_X1 port map( A1 => n13018, A2 => n13233, B1 => n13016, B2 => 
                           n10512, ZN => n2884);
   U10921 : OAI22_X1 port map( A1 => n13018, A2 => n13236, B1 => n13016, B2 => 
                           n10511, ZN => n2885);
   U10922 : OAI22_X1 port map( A1 => n13018, A2 => n13239, B1 => n13016, B2 => 
                           n10510, ZN => n2886);
   U10923 : OAI22_X1 port map( A1 => n13018, A2 => n13242, B1 => n13016, B2 => 
                           n10509, ZN => n2887);
   U10924 : OAI22_X1 port map( A1 => n13019, A2 => n13245, B1 => n13016, B2 => 
                           n10508, ZN => n2888);
   U10925 : OAI22_X1 port map( A1 => n13019, A2 => n13248, B1 => n13016, B2 => 
                           n10507, ZN => n2889);
   U10926 : OAI22_X1 port map( A1 => n13019, A2 => n13251, B1 => n10965, B2 => 
                           n10506, ZN => n2890);
   U10927 : OAI22_X1 port map( A1 => n13019, A2 => n13254, B1 => n10965, B2 => 
                           n10505, ZN => n2891);
   U10928 : OAI22_X1 port map( A1 => n13019, A2 => n13257, B1 => n10965, B2 => 
                           n10504, ZN => n2892);
   U10929 : OAI22_X1 port map( A1 => n13020, A2 => n13260, B1 => n13016, B2 => 
                           n10503, ZN => n2893);
   U10930 : OAI22_X1 port map( A1 => n13020, A2 => n13263, B1 => n13016, B2 => 
                           n10502, ZN => n2894);
   U10931 : OAI22_X1 port map( A1 => n13020, A2 => n13266, B1 => n13016, B2 => 
                           n10501, ZN => n2895);
   U10932 : OAI22_X1 port map( A1 => n13020, A2 => n13269, B1 => n13016, B2 => 
                           n10500, ZN => n2896);
   U10933 : OAI22_X1 port map( A1 => n13020, A2 => n13272, B1 => n13016, B2 => 
                           n10499, ZN => n2897);
   U10934 : OAI22_X1 port map( A1 => n13021, A2 => n13275, B1 => n13016, B2 => 
                           n10498, ZN => n2898);
   U10935 : OAI22_X1 port map( A1 => n13021, A2 => n13278, B1 => n13016, B2 => 
                           n10497, ZN => n2899);
   U10936 : OAI22_X1 port map( A1 => n13021, A2 => n13281, B1 => n13016, B2 => 
                           n10496, ZN => n2900);
   U10937 : OAI22_X1 port map( A1 => n13021, A2 => n13284, B1 => n13016, B2 => 
                           n10495, ZN => n2901);
   U10938 : OAI22_X1 port map( A1 => n12999, A2 => n13216, B1 => n12998, B2 => 
                           n10494, ZN => n2814);
   U10939 : OAI22_X1 port map( A1 => n12999, A2 => n13219, B1 => n12998, B2 => 
                           n10493, ZN => n2815);
   U10940 : OAI22_X1 port map( A1 => n12999, A2 => n13222, B1 => n12998, B2 => 
                           n10492, ZN => n2816);
   U10941 : OAI22_X1 port map( A1 => n12999, A2 => n13225, B1 => n12998, B2 => 
                           n10491, ZN => n2817);
   U10942 : OAI22_X1 port map( A1 => n12999, A2 => n13228, B1 => n12998, B2 => 
                           n10490, ZN => n2818);
   U10943 : OAI22_X1 port map( A1 => n13000, A2 => n13231, B1 => n12998, B2 => 
                           n10489, ZN => n2819);
   U10944 : OAI22_X1 port map( A1 => n13000, A2 => n13234, B1 => n12998, B2 => 
                           n10488, ZN => n2820);
   U10945 : OAI22_X1 port map( A1 => n13000, A2 => n13237, B1 => n12998, B2 => 
                           n10487, ZN => n2821);
   U10946 : OAI22_X1 port map( A1 => n13000, A2 => n13240, B1 => n12998, B2 => 
                           n10486, ZN => n2822);
   U10947 : OAI22_X1 port map( A1 => n13000, A2 => n13243, B1 => n12998, B2 => 
                           n10485, ZN => n2823);
   U10948 : OAI22_X1 port map( A1 => n13001, A2 => n13246, B1 => n12998, B2 => 
                           n10484, ZN => n2824);
   U10949 : OAI22_X1 port map( A1 => n13001, A2 => n13249, B1 => n12998, B2 => 
                           n10483, ZN => n2825);
   U10950 : OAI22_X1 port map( A1 => n13001, A2 => n13252, B1 => n10967, B2 => 
                           n10482, ZN => n2826);
   U10951 : OAI22_X1 port map( A1 => n13001, A2 => n13255, B1 => n10967, B2 => 
                           n10481, ZN => n2827);
   U10952 : OAI22_X1 port map( A1 => n13001, A2 => n13258, B1 => n10967, B2 => 
                           n10480, ZN => n2828);
   U10953 : OAI22_X1 port map( A1 => n13002, A2 => n13261, B1 => n12998, B2 => 
                           n10479, ZN => n2829);
   U10954 : OAI22_X1 port map( A1 => n13002, A2 => n13264, B1 => n12998, B2 => 
                           n10478, ZN => n2830);
   U10955 : OAI22_X1 port map( A1 => n13002, A2 => n13267, B1 => n12998, B2 => 
                           n10477, ZN => n2831);
   U10956 : OAI22_X1 port map( A1 => n13002, A2 => n13270, B1 => n12998, B2 => 
                           n10476, ZN => n2832);
   U10957 : OAI22_X1 port map( A1 => n13002, A2 => n13273, B1 => n12998, B2 => 
                           n10475, ZN => n2833);
   U10958 : OAI22_X1 port map( A1 => n13003, A2 => n13276, B1 => n12998, B2 => 
                           n10474, ZN => n2834);
   U10959 : OAI22_X1 port map( A1 => n13003, A2 => n13279, B1 => n12998, B2 => 
                           n10473, ZN => n2835);
   U10960 : OAI22_X1 port map( A1 => n13003, A2 => n13282, B1 => n12998, B2 => 
                           n10472, ZN => n2836);
   U10961 : OAI22_X1 port map( A1 => n13003, A2 => n13285, B1 => n12998, B2 => 
                           n10471, ZN => n2837);
   U10962 : OAI22_X1 port map( A1 => n12963, A2 => n13216, B1 => n12962, B2 => 
                           n10470, ZN => n2686);
   U10963 : OAI22_X1 port map( A1 => n12963, A2 => n13219, B1 => n12962, B2 => 
                           n10469, ZN => n2687);
   U10964 : OAI22_X1 port map( A1 => n12963, A2 => n13222, B1 => n12962, B2 => 
                           n10468, ZN => n2688);
   U10965 : OAI22_X1 port map( A1 => n12963, A2 => n13225, B1 => n12962, B2 => 
                           n10467, ZN => n2689);
   U10966 : OAI22_X1 port map( A1 => n12963, A2 => n13228, B1 => n12962, B2 => 
                           n10466, ZN => n2690);
   U10967 : OAI22_X1 port map( A1 => n12964, A2 => n13231, B1 => n12962, B2 => 
                           n10465, ZN => n2691);
   U10968 : OAI22_X1 port map( A1 => n12964, A2 => n13234, B1 => n12962, B2 => 
                           n10464, ZN => n2692);
   U10969 : OAI22_X1 port map( A1 => n12964, A2 => n13237, B1 => n12962, B2 => 
                           n10463, ZN => n2693);
   U10970 : OAI22_X1 port map( A1 => n12964, A2 => n13240, B1 => n12962, B2 => 
                           n10462, ZN => n2694);
   U10971 : OAI22_X1 port map( A1 => n12964, A2 => n13243, B1 => n12962, B2 => 
                           n10461, ZN => n2695);
   U10972 : OAI22_X1 port map( A1 => n12965, A2 => n13246, B1 => n12962, B2 => 
                           n10460, ZN => n2696);
   U10973 : OAI22_X1 port map( A1 => n12965, A2 => n13249, B1 => n12962, B2 => 
                           n10459, ZN => n2697);
   U10974 : OAI22_X1 port map( A1 => n12965, A2 => n13252, B1 => n10972, B2 => 
                           n10458, ZN => n2698);
   U10975 : OAI22_X1 port map( A1 => n12965, A2 => n13255, B1 => n10972, B2 => 
                           n10457, ZN => n2699);
   U10976 : OAI22_X1 port map( A1 => n12965, A2 => n13258, B1 => n10972, B2 => 
                           n10456, ZN => n2700);
   U10977 : OAI22_X1 port map( A1 => n12966, A2 => n13261, B1 => n12962, B2 => 
                           n10455, ZN => n2701);
   U10978 : OAI22_X1 port map( A1 => n12966, A2 => n13264, B1 => n12962, B2 => 
                           n10454, ZN => n2702);
   U10979 : OAI22_X1 port map( A1 => n12966, A2 => n13267, B1 => n12962, B2 => 
                           n10453, ZN => n2703);
   U10980 : OAI22_X1 port map( A1 => n12966, A2 => n13270, B1 => n12962, B2 => 
                           n10452, ZN => n2704);
   U10981 : OAI22_X1 port map( A1 => n12966, A2 => n13273, B1 => n12962, B2 => 
                           n10451, ZN => n2705);
   U10982 : OAI22_X1 port map( A1 => n12967, A2 => n13276, B1 => n12962, B2 => 
                           n10450, ZN => n2706);
   U10983 : OAI22_X1 port map( A1 => n12967, A2 => n13279, B1 => n12962, B2 => 
                           n10449, ZN => n2707);
   U10984 : OAI22_X1 port map( A1 => n12967, A2 => n13282, B1 => n12962, B2 => 
                           n10448, ZN => n2708);
   U10985 : OAI22_X1 port map( A1 => n12967, A2 => n13285, B1 => n12962, B2 => 
                           n10447, ZN => n2709);
   U10986 : OAI22_X1 port map( A1 => n13210, A2 => n13274, B1 => n10934, B2 => 
                           n10446, ZN => n3570);
   U10987 : OAI22_X1 port map( A1 => n13210, A2 => n13277, B1 => n10934, B2 => 
                           n10445, ZN => n3571);
   U10988 : OAI22_X1 port map( A1 => n13210, A2 => n13280, B1 => n10934, B2 => 
                           n10444, ZN => n3572);
   U10989 : OAI22_X1 port map( A1 => n13210, A2 => n13283, B1 => n13205, B2 => 
                           n10443, ZN => n3573);
   U10990 : OAI22_X1 port map( A1 => n13308, A2 => n13217, B1 => n13307, B2 => 
                           n10354, ZN => n3583);
   U10991 : OAI22_X1 port map( A1 => n13308, A2 => n13220, B1 => n13307, B2 => 
                           n10353, ZN => n3584);
   U10992 : OAI22_X1 port map( A1 => n13308, A2 => n13223, B1 => n13307, B2 => 
                           n10352, ZN => n3585);
   U10993 : OAI22_X1 port map( A1 => n13308, A2 => n13226, B1 => n13307, B2 => 
                           n10351, ZN => n3586);
   U10994 : OAI22_X1 port map( A1 => n13309, A2 => n13229, B1 => n13307, B2 => 
                           n10350, ZN => n3587);
   U10995 : OAI22_X1 port map( A1 => n13309, A2 => n13232, B1 => n13307, B2 => 
                           n10349, ZN => n3588);
   U10996 : OAI22_X1 port map( A1 => n13309, A2 => n13235, B1 => n13307, B2 => 
                           n10348, ZN => n3589);
   U10997 : OAI22_X1 port map( A1 => n13152, A2 => n13214, B1 => n13151, B2 => 
                           n10026, ZN => n3358);
   U10998 : OAI22_X1 port map( A1 => n13152, A2 => n13217, B1 => n13151, B2 => 
                           n10025, ZN => n3359);
   U10999 : OAI22_X1 port map( A1 => n13152, A2 => n13220, B1 => n13151, B2 => 
                           n10024, ZN => n3360);
   U11000 : OAI22_X1 port map( A1 => n13152, A2 => n13223, B1 => n13151, B2 => 
                           n10023, ZN => n3361);
   U11001 : OAI22_X1 port map( A1 => n13152, A2 => n13226, B1 => n13151, B2 => 
                           n10022, ZN => n3362);
   U11002 : OAI22_X1 port map( A1 => n13153, A2 => n13229, B1 => n13151, B2 => 
                           n10021, ZN => n3363);
   U11003 : OAI22_X1 port map( A1 => n13153, A2 => n13232, B1 => n13151, B2 => 
                           n10020, ZN => n3364);
   U11004 : OAI22_X1 port map( A1 => n13153, A2 => n13235, B1 => n13151, B2 => 
                           n10019, ZN => n3365);
   U11005 : OAI22_X1 port map( A1 => n13153, A2 => n13238, B1 => n13151, B2 => 
                           n10018, ZN => n3366);
   U11006 : OAI22_X1 port map( A1 => n13153, A2 => n13241, B1 => n13151, B2 => 
                           n10017, ZN => n3367);
   U11007 : OAI22_X1 port map( A1 => n13154, A2 => n13244, B1 => n13151, B2 => 
                           n10016, ZN => n3368);
   U11008 : OAI22_X1 port map( A1 => n13154, A2 => n13247, B1 => n13151, B2 => 
                           n10015, ZN => n3369);
   U11009 : OAI22_X1 port map( A1 => n13154, A2 => n13250, B1 => n10946, B2 => 
                           n10014, ZN => n3370);
   U11010 : OAI22_X1 port map( A1 => n13154, A2 => n13253, B1 => n10946, B2 => 
                           n10013, ZN => n3371);
   U11011 : OAI22_X1 port map( A1 => n13154, A2 => n13256, B1 => n10946, B2 => 
                           n10012, ZN => n3372);
   U11012 : OAI22_X1 port map( A1 => n13155, A2 => n13259, B1 => n13151, B2 => 
                           n10011, ZN => n3373);
   U11013 : OAI22_X1 port map( A1 => n13155, A2 => n13262, B1 => n13151, B2 => 
                           n10010, ZN => n3374);
   U11014 : OAI22_X1 port map( A1 => n13155, A2 => n13265, B1 => n13151, B2 => 
                           n10009, ZN => n3375);
   U11015 : OAI22_X1 port map( A1 => n13155, A2 => n13268, B1 => n13151, B2 => 
                           n10008, ZN => n3376);
   U11016 : OAI22_X1 port map( A1 => n13155, A2 => n13271, B1 => n13151, B2 => 
                           n10007, ZN => n3377);
   U11017 : OAI22_X1 port map( A1 => n13156, A2 => n13274, B1 => n13151, B2 => 
                           n10006, ZN => n3378);
   U11018 : OAI22_X1 port map( A1 => n13156, A2 => n13277, B1 => n13151, B2 => 
                           n10005, ZN => n3379);
   U11019 : OAI22_X1 port map( A1 => n13156, A2 => n13280, B1 => n13151, B2 => 
                           n10004, ZN => n3380);
   U11020 : OAI22_X1 port map( A1 => n13156, A2 => n13283, B1 => n13151, B2 => 
                           n10003, ZN => n3381);
   U11021 : OAI22_X1 port map( A1 => n13161, A2 => n13214, B1 => n13160, B2 => 
                           n9994, ZN => n3390);
   U11022 : OAI22_X1 port map( A1 => n13161, A2 => n13217, B1 => n13160, B2 => 
                           n9993, ZN => n3391);
   U11023 : OAI22_X1 port map( A1 => n13161, A2 => n13220, B1 => n13160, B2 => 
                           n9992, ZN => n3392);
   U11024 : OAI22_X1 port map( A1 => n13161, A2 => n13223, B1 => n13160, B2 => 
                           n9991, ZN => n3393);
   U11025 : OAI22_X1 port map( A1 => n13161, A2 => n13226, B1 => n13160, B2 => 
                           n9990, ZN => n3394);
   U11026 : OAI22_X1 port map( A1 => n13162, A2 => n13229, B1 => n13160, B2 => 
                           n9989, ZN => n3395);
   U11027 : OAI22_X1 port map( A1 => n13162, A2 => n13232, B1 => n13160, B2 => 
                           n9988, ZN => n3396);
   U11028 : OAI22_X1 port map( A1 => n13162, A2 => n13235, B1 => n13160, B2 => 
                           n9987, ZN => n3397);
   U11029 : OAI22_X1 port map( A1 => n13162, A2 => n13238, B1 => n13160, B2 => 
                           n9986, ZN => n3398);
   U11030 : OAI22_X1 port map( A1 => n13162, A2 => n13241, B1 => n13160, B2 => 
                           n9985, ZN => n3399);
   U11031 : OAI22_X1 port map( A1 => n13163, A2 => n13244, B1 => n13160, B2 => 
                           n9984, ZN => n3400);
   U11032 : OAI22_X1 port map( A1 => n13163, A2 => n13247, B1 => n13160, B2 => 
                           n9983, ZN => n3401);
   U11033 : OAI22_X1 port map( A1 => n13163, A2 => n13250, B1 => n10944, B2 => 
                           n9982, ZN => n3402);
   U11034 : OAI22_X1 port map( A1 => n13163, A2 => n13253, B1 => n10944, B2 => 
                           n9981, ZN => n3403);
   U11035 : OAI22_X1 port map( A1 => n13163, A2 => n13256, B1 => n10944, B2 => 
                           n9980, ZN => n3404);
   U11036 : OAI22_X1 port map( A1 => n13164, A2 => n13259, B1 => n13160, B2 => 
                           n9979, ZN => n3405);
   U11037 : OAI22_X1 port map( A1 => n13164, A2 => n13262, B1 => n13160, B2 => 
                           n9978, ZN => n3406);
   U11038 : OAI22_X1 port map( A1 => n13164, A2 => n13265, B1 => n13160, B2 => 
                           n9977, ZN => n3407);
   U11039 : OAI22_X1 port map( A1 => n13164, A2 => n13268, B1 => n13160, B2 => 
                           n9976, ZN => n3408);
   U11040 : OAI22_X1 port map( A1 => n13164, A2 => n13271, B1 => n13160, B2 => 
                           n9975, ZN => n3409);
   U11041 : OAI22_X1 port map( A1 => n13165, A2 => n13274, B1 => n13160, B2 => 
                           n9974, ZN => n3410);
   U11042 : OAI22_X1 port map( A1 => n13165, A2 => n13277, B1 => n13160, B2 => 
                           n9973, ZN => n3411);
   U11043 : OAI22_X1 port map( A1 => n13165, A2 => n13280, B1 => n13160, B2 => 
                           n9972, ZN => n3412);
   U11044 : OAI22_X1 port map( A1 => n13165, A2 => n13283, B1 => n13160, B2 => 
                           n9971, ZN => n3413);
   U11045 : OAI22_X1 port map( A1 => n13206, A2 => n13214, B1 => n13205, B2 => 
                           n9963, ZN => n3550);
   U11046 : OAI22_X1 port map( A1 => n13206, A2 => n13217, B1 => n13205, B2 => 
                           n9962, ZN => n3551);
   U11047 : OAI22_X1 port map( A1 => n13206, A2 => n13220, B1 => n13205, B2 => 
                           n9961, ZN => n3552);
   U11048 : OAI22_X1 port map( A1 => n13206, A2 => n13223, B1 => n13205, B2 => 
                           n9960, ZN => n3553);
   U11049 : OAI22_X1 port map( A1 => n13206, A2 => n13226, B1 => n13205, B2 => 
                           n9959, ZN => n3554);
   U11050 : OAI22_X1 port map( A1 => n13207, A2 => n13229, B1 => n13205, B2 => 
                           n9958, ZN => n3555);
   U11051 : OAI22_X1 port map( A1 => n13207, A2 => n13232, B1 => n13205, B2 => 
                           n9957, ZN => n3556);
   U11052 : OAI22_X1 port map( A1 => n13207, A2 => n13235, B1 => n13205, B2 => 
                           n9956, ZN => n3557);
   U11053 : OAI22_X1 port map( A1 => n13207, A2 => n13238, B1 => n13205, B2 => 
                           n9955, ZN => n3558);
   U11054 : OAI22_X1 port map( A1 => n13207, A2 => n13241, B1 => n13205, B2 => 
                           n9954, ZN => n3559);
   U11055 : OAI22_X1 port map( A1 => n13208, A2 => n13244, B1 => n13205, B2 => 
                           n9953, ZN => n3560);
   U11056 : OAI22_X1 port map( A1 => n13208, A2 => n13247, B1 => n13205, B2 => 
                           n9952, ZN => n3561);
   U11057 : OAI22_X1 port map( A1 => n13208, A2 => n13250, B1 => n13205, B2 => 
                           n9951, ZN => n3562);
   U11058 : OAI22_X1 port map( A1 => n13208, A2 => n13253, B1 => n13205, B2 => 
                           n9950, ZN => n3563);
   U11059 : OAI22_X1 port map( A1 => n13208, A2 => n13256, B1 => n13205, B2 => 
                           n9949, ZN => n3564);
   U11060 : OAI22_X1 port map( A1 => n13209, A2 => n13259, B1 => n13205, B2 => 
                           n9948, ZN => n3565);
   U11061 : OAI22_X1 port map( A1 => n13209, A2 => n13262, B1 => n13205, B2 => 
                           n9947, ZN => n3566);
   U11062 : OAI22_X1 port map( A1 => n13209, A2 => n13265, B1 => n13205, B2 => 
                           n9946, ZN => n3567);
   U11063 : OAI22_X1 port map( A1 => n13209, A2 => n13268, B1 => n13205, B2 => 
                           n9945, ZN => n3568);
   U11064 : OAI22_X1 port map( A1 => n13209, A2 => n13271, B1 => n13205, B2 => 
                           n9944, ZN => n3569);
   U11065 : OAI22_X1 port map( A1 => n13312, A2 => n13283, B1 => n13307, B2 => 
                           n9943, ZN => n3605);
   U11066 : NOR2_X1 port map( A1 => n9931, A2 => n9932, ZN => n12264);
   U11067 : NOR2_X1 port map( A1 => n9936, A2 => n9937, ZN => n11611);
   U11068 : NOR3_X1 port map( A1 => n9933, A2 => n9929, A3 => n9930, ZN => 
                           n12280);
   U11069 : NOR3_X1 port map( A1 => n9938, A2 => n9934, A3 => n9935, ZN => 
                           n11627);
   U11070 : BUF_X1 port map( A => n11629, Z => n12828);
   U11071 : BUF_X1 port map( A => n10976, Z => n12930);
   U11072 : BUF_X1 port map( A => n11629, Z => n12829);
   U11073 : BUF_X1 port map( A => n11629, Z => n12830);
   U11074 : BUF_X1 port map( A => n10976, Z => n12931);
   U11075 : BUF_X1 port map( A => n10976, Z => n12932);
   U11076 : BUF_X1 port map( A => n9923, Z => n13322);
   U11077 : BUF_X1 port map( A => n9923, Z => n13323);
   U11078 : BUF_X1 port map( A => n9923, Z => n13320);
   U11079 : BUF_X1 port map( A => n9923, Z => n13319);
   U11080 : BUF_X1 port map( A => n10931, Z => n13215);
   U11081 : BUF_X1 port map( A => n10930, Z => n13218);
   U11082 : BUF_X1 port map( A => n10929, Z => n13221);
   U11083 : BUF_X1 port map( A => n10928, Z => n13224);
   U11084 : BUF_X1 port map( A => n10927, Z => n13227);
   U11085 : BUF_X1 port map( A => n10926, Z => n13230);
   U11086 : BUF_X1 port map( A => n10925, Z => n13233);
   U11087 : BUF_X1 port map( A => n10924, Z => n13236);
   U11088 : BUF_X1 port map( A => n10923, Z => n13239);
   U11089 : BUF_X1 port map( A => n10922, Z => n13242);
   U11090 : BUF_X1 port map( A => n10921, Z => n13245);
   U11091 : BUF_X1 port map( A => n10920, Z => n13248);
   U11092 : BUF_X1 port map( A => n10919, Z => n13251);
   U11093 : BUF_X1 port map( A => n10918, Z => n13254);
   U11094 : BUF_X1 port map( A => n10917, Z => n13257);
   U11095 : BUF_X1 port map( A => n10916, Z => n13260);
   U11096 : BUF_X1 port map( A => n10915, Z => n13263);
   U11097 : BUF_X1 port map( A => n10914, Z => n13266);
   U11098 : BUF_X1 port map( A => n10913, Z => n13269);
   U11099 : BUF_X1 port map( A => n10912, Z => n13272);
   U11100 : BUF_X1 port map( A => n10911, Z => n13275);
   U11101 : BUF_X1 port map( A => n10910, Z => n13278);
   U11102 : BUF_X1 port map( A => n10909, Z => n13281);
   U11103 : BUF_X1 port map( A => n10908, Z => n13284);
   U11104 : BUF_X1 port map( A => n10907, Z => n13287);
   U11105 : BUF_X1 port map( A => n10906, Z => n13290);
   U11106 : BUF_X1 port map( A => n10905, Z => n13293);
   U11107 : BUF_X1 port map( A => n10904, Z => n13296);
   U11108 : BUF_X1 port map( A => n10903, Z => n13299);
   U11109 : BUF_X1 port map( A => n10902, Z => n13302);
   U11110 : BUF_X1 port map( A => n10901, Z => n13305);
   U11111 : BUF_X1 port map( A => n10899, Z => n13317);
   U11112 : BUF_X1 port map( A => n10899, Z => n13316);
   U11113 : BUF_X1 port map( A => n10911, Z => n13274);
   U11114 : BUF_X1 port map( A => n10910, Z => n13277);
   U11115 : BUF_X1 port map( A => n10909, Z => n13280);
   U11116 : BUF_X1 port map( A => n10903, Z => n13298);
   U11117 : BUF_X1 port map( A => n10902, Z => n13301);
   U11118 : BUF_X1 port map( A => n10901, Z => n13304);
   U11119 : BUF_X1 port map( A => n10931, Z => n13214);
   U11120 : BUF_X1 port map( A => n10930, Z => n13217);
   U11121 : BUF_X1 port map( A => n10929, Z => n13220);
   U11122 : BUF_X1 port map( A => n10928, Z => n13223);
   U11123 : BUF_X1 port map( A => n10927, Z => n13226);
   U11124 : BUF_X1 port map( A => n10926, Z => n13229);
   U11125 : BUF_X1 port map( A => n10925, Z => n13232);
   U11126 : BUF_X1 port map( A => n10924, Z => n13235);
   U11127 : BUF_X1 port map( A => n10923, Z => n13238);
   U11128 : BUF_X1 port map( A => n10922, Z => n13241);
   U11129 : BUF_X1 port map( A => n10921, Z => n13244);
   U11130 : BUF_X1 port map( A => n10920, Z => n13247);
   U11131 : BUF_X1 port map( A => n10919, Z => n13250);
   U11132 : BUF_X1 port map( A => n10918, Z => n13253);
   U11133 : BUF_X1 port map( A => n10917, Z => n13256);
   U11134 : BUF_X1 port map( A => n10916, Z => n13259);
   U11135 : BUF_X1 port map( A => n10915, Z => n13262);
   U11136 : BUF_X1 port map( A => n10914, Z => n13265);
   U11137 : BUF_X1 port map( A => n10913, Z => n13268);
   U11138 : BUF_X1 port map( A => n10912, Z => n13271);
   U11139 : BUF_X1 port map( A => n10908, Z => n13283);
   U11140 : BUF_X1 port map( A => n10907, Z => n13286);
   U11141 : BUF_X1 port map( A => n10906, Z => n13289);
   U11142 : BUF_X1 port map( A => n10905, Z => n13292);
   U11143 : BUF_X1 port map( A => n10904, Z => n13295);
   U11144 : BUF_X1 port map( A => n9923, Z => n13321);
   U11145 : BUF_X1 port map( A => n11629, Z => n12826);
   U11146 : BUF_X1 port map( A => n11629, Z => n12827);
   U11147 : BUF_X1 port map( A => n10976, Z => n12928);
   U11148 : BUF_X1 port map( A => n10976, Z => n12929);
   U11149 : BUF_X1 port map( A => n10931, Z => n13216);
   U11150 : BUF_X1 port map( A => n10930, Z => n13219);
   U11151 : BUF_X1 port map( A => n10929, Z => n13222);
   U11152 : BUF_X1 port map( A => n10928, Z => n13225);
   U11153 : BUF_X1 port map( A => n10927, Z => n13228);
   U11154 : BUF_X1 port map( A => n10926, Z => n13231);
   U11155 : BUF_X1 port map( A => n10925, Z => n13234);
   U11156 : BUF_X1 port map( A => n10924, Z => n13237);
   U11157 : BUF_X1 port map( A => n10923, Z => n13240);
   U11158 : BUF_X1 port map( A => n10922, Z => n13243);
   U11159 : BUF_X1 port map( A => n10921, Z => n13246);
   U11160 : BUF_X1 port map( A => n10920, Z => n13249);
   U11161 : BUF_X1 port map( A => n10919, Z => n13252);
   U11162 : BUF_X1 port map( A => n10918, Z => n13255);
   U11163 : BUF_X1 port map( A => n10917, Z => n13258);
   U11164 : BUF_X1 port map( A => n10916, Z => n13261);
   U11165 : BUF_X1 port map( A => n10915, Z => n13264);
   U11166 : BUF_X1 port map( A => n10914, Z => n13267);
   U11167 : BUF_X1 port map( A => n10913, Z => n13270);
   U11168 : BUF_X1 port map( A => n10912, Z => n13273);
   U11169 : BUF_X1 port map( A => n10911, Z => n13276);
   U11170 : BUF_X1 port map( A => n10910, Z => n13279);
   U11171 : BUF_X1 port map( A => n10909, Z => n13282);
   U11172 : BUF_X1 port map( A => n10908, Z => n13285);
   U11173 : BUF_X1 port map( A => n10907, Z => n13288);
   U11174 : BUF_X1 port map( A => n10906, Z => n13291);
   U11175 : BUF_X1 port map( A => n10905, Z => n13294);
   U11176 : BUF_X1 port map( A => n10904, Z => n13297);
   U11177 : BUF_X1 port map( A => n10903, Z => n13300);
   U11178 : BUF_X1 port map( A => n10902, Z => n13303);
   U11179 : BUF_X1 port map( A => n10901, Z => n13306);
   U11180 : BUF_X1 port map( A => n10899, Z => n13318);
   U11181 : NAND2_X1 port map( A1 => n12260, A2 => n12276, ZN => n11664);
   U11182 : NAND2_X1 port map( A1 => n12260, A2 => n12275, ZN => n11665);
   U11183 : NAND2_X1 port map( A1 => n11607, A2 => n11623, ZN => n11011);
   U11184 : NAND2_X1 port map( A1 => n11607, A2 => n11622, ZN => n11012);
   U11185 : NAND2_X1 port map( A1 => n12264, A2 => n12276, ZN => n11669);
   U11186 : NAND2_X1 port map( A1 => n12264, A2 => n12275, ZN => n11670);
   U11187 : NAND2_X1 port map( A1 => n11611, A2 => n11623, ZN => n11016);
   U11188 : NAND2_X1 port map( A1 => n11611, A2 => n11622, ZN => n11017);
   U11189 : NAND2_X1 port map( A1 => n12261, A2 => n12260, ZN => n11640);
   U11190 : NAND2_X1 port map( A1 => n12261, A2 => n12264, ZN => n11646);
   U11191 : NAND2_X1 port map( A1 => n12280, A2 => n12260, ZN => n11674);
   U11192 : NAND2_X1 port map( A1 => n12280, A2 => n12265, ZN => n11679);
   U11193 : NAND2_X1 port map( A1 => n11608, A2 => n11607, ZN => n10987);
   U11194 : NAND2_X1 port map( A1 => n11608, A2 => n11611, ZN => n10993);
   U11195 : NAND2_X1 port map( A1 => n11627, A2 => n11607, ZN => n11021);
   U11196 : NAND2_X1 port map( A1 => n11627, A2 => n11612, ZN => n11026);
   U11197 : NAND2_X1 port map( A1 => n12259, A2 => n12260, ZN => n11641);
   U11198 : NAND2_X1 port map( A1 => n12259, A2 => n12264, ZN => n11645);
   U11199 : NAND2_X1 port map( A1 => n12268, A2 => n12264, ZN => n11655);
   U11200 : NAND2_X1 port map( A1 => n12267, A2 => n12264, ZN => n11656);
   U11201 : NAND2_X1 port map( A1 => n12268, A2 => n12260, ZN => n11650);
   U11202 : NAND2_X1 port map( A1 => n12267, A2 => n12260, ZN => n11651);
   U11203 : NAND2_X1 port map( A1 => n12279, A2 => n12260, ZN => n11675);
   U11204 : NAND2_X1 port map( A1 => n12279, A2 => n12265, ZN => n11680);
   U11205 : NAND2_X1 port map( A1 => n11606, A2 => n11607, ZN => n10988);
   U11206 : NAND2_X1 port map( A1 => n11606, A2 => n11611, ZN => n10992);
   U11207 : NAND2_X1 port map( A1 => n11615, A2 => n11611, ZN => n11002);
   U11208 : NAND2_X1 port map( A1 => n11614, A2 => n11611, ZN => n11003);
   U11209 : NAND2_X1 port map( A1 => n11615, A2 => n11609, ZN => n10997);
   U11210 : NAND2_X1 port map( A1 => n11614, A2 => n11609, ZN => n10998);
   U11211 : NAND2_X1 port map( A1 => n11626, A2 => n11607, ZN => n11022);
   U11212 : NAND2_X1 port map( A1 => n11626, A2 => n11612, ZN => n11027);
   U11213 : AND2_X1 port map( A1 => n12276, A2 => n12262, ZN => n11662);
   U11214 : AND2_X1 port map( A1 => n11623, A2 => n11609, ZN => n11009);
   U11215 : AND2_X1 port map( A1 => n11609, A2 => n11622, ZN => n11008);
   U11216 : AND2_X1 port map( A1 => n12265, A2 => n12275, ZN => n11666);
   U11217 : AND2_X1 port map( A1 => n12265, A2 => n12276, ZN => n11667);
   U11218 : AND2_X1 port map( A1 => n11612, A2 => n11622, ZN => n11013);
   U11219 : AND2_X1 port map( A1 => n11612, A2 => n11623, ZN => n11014);
   U11220 : AND2_X1 port map( A1 => n12279, A2 => n12264, ZN => n11676);
   U11221 : AND2_X1 port map( A1 => n11614, A2 => n11607, ZN => n10994);
   U11222 : AND2_X1 port map( A1 => n11615, A2 => n11607, ZN => n10995);
   U11223 : AND2_X1 port map( A1 => n11626, A2 => n11611, ZN => n11023);
   U11224 : AND2_X1 port map( A1 => n12259, A2 => n12262, ZN => n11637);
   U11225 : AND2_X1 port map( A1 => n12261, A2 => n12262, ZN => n11638);
   U11226 : AND2_X1 port map( A1 => n12261, A2 => n12265, ZN => n11642);
   U11227 : AND2_X1 port map( A1 => n12259, A2 => n12265, ZN => n11643);
   U11228 : AND2_X1 port map( A1 => n12267, A2 => n12265, ZN => n11652);
   U11229 : AND2_X1 port map( A1 => n12268, A2 => n12265, ZN => n11653);
   U11230 : AND2_X1 port map( A1 => n12267, A2 => n12262, ZN => n11647);
   U11231 : AND2_X1 port map( A1 => n12268, A2 => n12262, ZN => n11648);
   U11232 : AND2_X1 port map( A1 => n12279, A2 => n12262, ZN => n11671);
   U11233 : AND2_X1 port map( A1 => n12280, A2 => n12262, ZN => n11672);
   U11234 : AND2_X1 port map( A1 => n11606, A2 => n11609, ZN => n10984);
   U11235 : AND2_X1 port map( A1 => n11608, A2 => n11609, ZN => n10985);
   U11236 : AND2_X1 port map( A1 => n11608, A2 => n11612, ZN => n10989);
   U11237 : AND2_X1 port map( A1 => n11606, A2 => n11612, ZN => n10990);
   U11238 : AND2_X1 port map( A1 => n11614, A2 => n11612, ZN => n10999);
   U11239 : AND2_X1 port map( A1 => n11615, A2 => n11612, ZN => n11000);
   U11240 : AND2_X1 port map( A1 => n11626, A2 => n11609, ZN => n11018);
   U11241 : AND2_X1 port map( A1 => n11627, A2 => n11609, ZN => n11019);
   U11242 : AND2_X1 port map( A1 => n12262, A2 => n12275, ZN => n11661);
   U11243 : BUF_X1 port map( A => n10975, Z => n12934);
   U11244 : OAI21_X1 port map( B1 => n10947, B2 => n10968, A => n13321, ZN => 
                           n10975);
   U11245 : INV_X1 port map( A => n10949, ZN => n13150);
   U11246 : OAI21_X1 port map( B1 => n10933, B2 => n10950, A => n13323, ZN => 
                           n10949);
   U11247 : INV_X1 port map( A => n10952, ZN => n13132);
   U11248 : OAI21_X1 port map( B1 => n10937, B2 => n10950, A => n13323, ZN => 
                           n10952);
   U11249 : INV_X1 port map( A => n10951, ZN => n13141);
   U11250 : OAI21_X1 port map( B1 => n10935, B2 => n10950, A => n13323, ZN => 
                           n10951);
   U11251 : INV_X1 port map( A => n10953, ZN => n13123);
   U11252 : OAI21_X1 port map( B1 => n10939, B2 => n10950, A => n13323, ZN => 
                           n10953);
   U11253 : INV_X1 port map( A => n10957, ZN => n13087);
   U11254 : OAI21_X1 port map( B1 => n10947, B2 => n10950, A => n13323, ZN => 
                           n10957);
   U11255 : INV_X1 port map( A => n10962, ZN => n13051);
   U11256 : OAI21_X1 port map( B1 => n10939, B2 => n10959, A => n13322, ZN => 
                           n10962);
   U11257 : INV_X1 port map( A => n10966, ZN => n13015);
   U11258 : OAI21_X1 port map( B1 => n10947, B2 => n10959, A => n13322, ZN => 
                           n10966);
   U11259 : INV_X1 port map( A => n10969, ZN => n12997);
   U11260 : OAI21_X1 port map( B1 => n10935, B2 => n10968, A => n13322, ZN => 
                           n10969);
   U11261 : INV_X1 port map( A => n10973, ZN => n12961);
   U11262 : OAI21_X1 port map( B1 => n10943, B2 => n10968, A => n13321, ZN => 
                           n10973);
   U11263 : INV_X1 port map( A => n10956, ZN => n13096);
   U11264 : OAI21_X1 port map( B1 => n10945, B2 => n10950, A => n13323, ZN => 
                           n10956);
   U11265 : INV_X1 port map( A => n10961, ZN => n13060);
   U11266 : OAI21_X1 port map( B1 => n10937, B2 => n10959, A => n13322, ZN => 
                           n10961);
   U11267 : INV_X1 port map( A => n10965, ZN => n13024);
   U11268 : OAI21_X1 port map( B1 => n10945, B2 => n10959, A => n13322, ZN => 
                           n10965);
   U11269 : INV_X1 port map( A => n10967, ZN => n13006);
   U11270 : OAI21_X1 port map( B1 => n10933, B2 => n10968, A => n13322, ZN => 
                           n10967);
   U11271 : INV_X1 port map( A => n10972, ZN => n12970);
   U11272 : OAI21_X1 port map( B1 => n10941, B2 => n10968, A => n13322, ZN => 
                           n10972);
   U11273 : INV_X1 port map( A => n10954, ZN => n13114);
   U11274 : OAI21_X1 port map( B1 => n10941, B2 => n10950, A => n13323, ZN => 
                           n10954);
   U11275 : INV_X1 port map( A => n10955, ZN => n13105);
   U11276 : OAI21_X1 port map( B1 => n10943, B2 => n10950, A => n13323, ZN => 
                           n10955);
   U11277 : INV_X1 port map( A => n10958, ZN => n13078);
   U11278 : OAI21_X1 port map( B1 => n10933, B2 => n10959, A => n13322, ZN => 
                           n10958);
   U11279 : INV_X1 port map( A => n10960, ZN => n13069);
   U11280 : OAI21_X1 port map( B1 => n10935, B2 => n10959, A => n13322, ZN => 
                           n10960);
   U11281 : INV_X1 port map( A => n10963, ZN => n13042);
   U11282 : OAI21_X1 port map( B1 => n10941, B2 => n10959, A => n13322, ZN => 
                           n10963);
   U11283 : INV_X1 port map( A => n10964, ZN => n13033);
   U11284 : OAI21_X1 port map( B1 => n10943, B2 => n10959, A => n13322, ZN => 
                           n10964);
   U11285 : INV_X1 port map( A => n10970, ZN => n12988);
   U11286 : OAI21_X1 port map( B1 => n10937, B2 => n10968, A => n13322, ZN => 
                           n10970);
   U11287 : INV_X1 port map( A => n10971, ZN => n12979);
   U11288 : OAI21_X1 port map( B1 => n10939, B2 => n10968, A => n13322, ZN => 
                           n10971);
   U11289 : INV_X1 port map( A => n10974, ZN => n12952);
   U11290 : OAI21_X1 port map( B1 => n10945, B2 => n10968, A => n13321, ZN => 
                           n10974);
   U11291 : INV_X1 port map( A => n10940, ZN => n13186);
   U11292 : OAI21_X1 port map( B1 => n10932, B2 => n10941, A => n13323, ZN => 
                           n10940);
   U11293 : INV_X1 port map( A => n10942, ZN => n13177);
   U11294 : OAI21_X1 port map( B1 => n10932, B2 => n10943, A => n13323, ZN => 
                           n10942);
   U11295 : INV_X1 port map( A => n10936, ZN => n13204);
   U11296 : OAI21_X1 port map( B1 => n10932, B2 => n10937, A => n13324, ZN => 
                           n10936);
   U11297 : INV_X1 port map( A => n10938, ZN => n13195);
   U11298 : OAI21_X1 port map( B1 => n10932, B2 => n10939, A => n13323, ZN => 
                           n10938);
   U11299 : INV_X1 port map( A => n10946, ZN => n13159);
   U11300 : OAI21_X1 port map( B1 => n10932, B2 => n10947, A => n13323, ZN => 
                           n10946);
   U11301 : INV_X1 port map( A => n10944, ZN => n13168);
   U11302 : OAI21_X1 port map( B1 => n10932, B2 => n10945, A => n13323, ZN => 
                           n10944);
   U11303 : INV_X1 port map( A => n10934, ZN => n13213);
   U11304 : OAI21_X1 port map( B1 => n10932, B2 => n10935, A => n13324, ZN => 
                           n10934);
   U11305 : AOI221_X1 port map( B1 => n12775, B2 => n12544, C1 => n12772, C2 =>
                           n12520, A => n12274, ZN => n12273);
   U11306 : OAI22_X1 port map( A1 => n9287, A2 => n12769, B1 => n9288, B2 => 
                           n12766, ZN => n12274);
   U11307 : AOI221_X1 port map( B1 => n12775, B2 => n12545, C1 => n12772, C2 =>
                           n12521, A => n12247, ZN => n12246);
   U11308 : OAI22_X1 port map( A1 => n9272, A2 => n12769, B1 => n9273, B2 => 
                           n12766, ZN => n12247);
   U11309 : AOI221_X1 port map( B1 => n12775, B2 => n12546, C1 => n12772, C2 =>
                           n12522, A => n12228, ZN => n12227);
   U11310 : OAI22_X1 port map( A1 => n9257, A2 => n12769, B1 => n9258, B2 => 
                           n12766, ZN => n12228);
   U11311 : AOI221_X1 port map( B1 => n12775, B2 => n12547, C1 => n12772, C2 =>
                           n12523, A => n12209, ZN => n12208);
   U11312 : OAI22_X1 port map( A1 => n9242, A2 => n12769, B1 => n9243, B2 => 
                           n12766, ZN => n12209);
   U11313 : AOI221_X1 port map( B1 => n12775, B2 => n12548, C1 => n12772, C2 =>
                           n12524, A => n12190, ZN => n12189);
   U11314 : OAI22_X1 port map( A1 => n9227, A2 => n12769, B1 => n9228, B2 => 
                           n12766, ZN => n12190);
   U11315 : AOI221_X1 port map( B1 => n12775, B2 => n12549, C1 => n12772, C2 =>
                           n12525, A => n12171, ZN => n12170);
   U11316 : OAI22_X1 port map( A1 => n9212, A2 => n12769, B1 => n9213, B2 => 
                           n12766, ZN => n12171);
   U11317 : AOI221_X1 port map( B1 => n12775, B2 => n12550, C1 => n12772, C2 =>
                           n12526, A => n12152, ZN => n12151);
   U11318 : OAI22_X1 port map( A1 => n9197, A2 => n12769, B1 => n9198, B2 => 
                           n12766, ZN => n12152);
   U11319 : AOI221_X1 port map( B1 => n12775, B2 => n12551, C1 => n12772, C2 =>
                           n12527, A => n12133, ZN => n12132);
   U11320 : OAI22_X1 port map( A1 => n9182, A2 => n12769, B1 => n9183, B2 => 
                           n12766, ZN => n12133);
   U11321 : AOI221_X1 port map( B1 => n12775, B2 => n12552, C1 => n12772, C2 =>
                           n12528, A => n12114, ZN => n12113);
   U11322 : OAI22_X1 port map( A1 => n9167, A2 => n12769, B1 => n9168, B2 => 
                           n12766, ZN => n12114);
   U11323 : AOI221_X1 port map( B1 => n12775, B2 => n12553, C1 => n12772, C2 =>
                           n12529, A => n12095, ZN => n12094);
   U11324 : OAI22_X1 port map( A1 => n9152, A2 => n12769, B1 => n9153, B2 => 
                           n12766, ZN => n12095);
   U11325 : AOI221_X1 port map( B1 => n12775, B2 => n12554, C1 => n12772, C2 =>
                           n12530, A => n12076, ZN => n12075);
   U11326 : OAI22_X1 port map( A1 => n9137, A2 => n12769, B1 => n9138, B2 => 
                           n12766, ZN => n12076);
   U11327 : AOI221_X1 port map( B1 => n12775, B2 => n12555, C1 => n12772, C2 =>
                           n12531, A => n12057, ZN => n12056);
   U11328 : OAI22_X1 port map( A1 => n9122, A2 => n12769, B1 => n9123, B2 => 
                           n12766, ZN => n12057);
   U11329 : AOI221_X1 port map( B1 => n12776, B2 => n12556, C1 => n12773, C2 =>
                           n12532, A => n12038, ZN => n12037);
   U11330 : OAI22_X1 port map( A1 => n9107, A2 => n12770, B1 => n9108, B2 => 
                           n12767, ZN => n12038);
   U11331 : AOI221_X1 port map( B1 => n12776, B2 => n12557, C1 => n12773, C2 =>
                           n12533, A => n12019, ZN => n12018);
   U11332 : OAI22_X1 port map( A1 => n9092, A2 => n12770, B1 => n9093, B2 => 
                           n12767, ZN => n12019);
   U11333 : AOI221_X1 port map( B1 => n12776, B2 => n12558, C1 => n12773, C2 =>
                           n12534, A => n12000, ZN => n11999);
   U11334 : OAI22_X1 port map( A1 => n9077, A2 => n12770, B1 => n9078, B2 => 
                           n12767, ZN => n12000);
   U11335 : AOI221_X1 port map( B1 => n12776, B2 => n12559, C1 => n12773, C2 =>
                           n12535, A => n11981, ZN => n11980);
   U11336 : OAI22_X1 port map( A1 => n9062, A2 => n12770, B1 => n9063, B2 => 
                           n12767, ZN => n11981);
   U11337 : AOI221_X1 port map( B1 => n12776, B2 => n12560, C1 => n12773, C2 =>
                           n12536, A => n11962, ZN => n11961);
   U11338 : OAI22_X1 port map( A1 => n9047, A2 => n12770, B1 => n9048, B2 => 
                           n12767, ZN => n11962);
   U11339 : AOI221_X1 port map( B1 => n12776, B2 => n12561, C1 => n12773, C2 =>
                           n12537, A => n11943, ZN => n11942);
   U11340 : OAI22_X1 port map( A1 => n9032, A2 => n12770, B1 => n9033, B2 => 
                           n12767, ZN => n11943);
   U11341 : AOI221_X1 port map( B1 => n12776, B2 => n12562, C1 => n12773, C2 =>
                           n12538, A => n11924, ZN => n11923);
   U11342 : OAI22_X1 port map( A1 => n9017, A2 => n12770, B1 => n9018, B2 => 
                           n12767, ZN => n11924);
   U11343 : AOI221_X1 port map( B1 => n12776, B2 => n12563, C1 => n12773, C2 =>
                           n12539, A => n11905, ZN => n11904);
   U11344 : OAI22_X1 port map( A1 => n9002, A2 => n12770, B1 => n9003, B2 => 
                           n12767, ZN => n11905);
   U11345 : AOI221_X1 port map( B1 => n12776, B2 => n12564, C1 => n12773, C2 =>
                           n12540, A => n11886, ZN => n11885);
   U11346 : OAI22_X1 port map( A1 => n8987, A2 => n12770, B1 => n8988, B2 => 
                           n12767, ZN => n11886);
   U11347 : AOI221_X1 port map( B1 => n12776, B2 => n12565, C1 => n12773, C2 =>
                           n12541, A => n11867, ZN => n11866);
   U11348 : OAI22_X1 port map( A1 => n8972, A2 => n12770, B1 => n8973, B2 => 
                           n12767, ZN => n11867);
   U11349 : AOI221_X1 port map( B1 => n12776, B2 => n12566, C1 => n12773, C2 =>
                           n12542, A => n11848, ZN => n11847);
   U11350 : OAI22_X1 port map( A1 => n8957, A2 => n12770, B1 => n8958, B2 => 
                           n12767, ZN => n11848);
   U11351 : AOI221_X1 port map( B1 => n12776, B2 => n12567, C1 => n12773, C2 =>
                           n12543, A => n11829, ZN => n11828);
   U11352 : OAI22_X1 port map( A1 => n8942, A2 => n12770, B1 => n8943, B2 => 
                           n12767, ZN => n11829);
   U11353 : AOI221_X1 port map( B1 => n12777, B2 => n12338, C1 => n12774, C2 =>
                           n12330, A => n11810, ZN => n11809);
   U11354 : OAI22_X1 port map( A1 => n8927, A2 => n12771, B1 => n8928, B2 => 
                           n12768, ZN => n11810);
   U11355 : AOI221_X1 port map( B1 => n12777, B2 => n12339, C1 => n12774, C2 =>
                           n12331, A => n11791, ZN => n11790);
   U11356 : OAI22_X1 port map( A1 => n8912, A2 => n12771, B1 => n8913, B2 => 
                           n12768, ZN => n11791);
   U11357 : AOI221_X1 port map( B1 => n12777, B2 => n12340, C1 => n12774, C2 =>
                           n12332, A => n11772, ZN => n11771);
   U11358 : OAI22_X1 port map( A1 => n8897, A2 => n12771, B1 => n8898, B2 => 
                           n12768, ZN => n11772);
   U11359 : AOI221_X1 port map( B1 => n12777, B2 => n12341, C1 => n12774, C2 =>
                           n12333, A => n11753, ZN => n11752);
   U11360 : OAI22_X1 port map( A1 => n8882, A2 => n12771, B1 => n8883, B2 => 
                           n12768, ZN => n11753);
   U11361 : AOI221_X1 port map( B1 => n12777, B2 => n12342, C1 => n12774, C2 =>
                           n12334, A => n11734, ZN => n11733);
   U11362 : OAI22_X1 port map( A1 => n8867, A2 => n12771, B1 => n8868, B2 => 
                           n12768, ZN => n11734);
   U11363 : AOI221_X1 port map( B1 => n12777, B2 => n12343, C1 => n12774, C2 =>
                           n12335, A => n11715, ZN => n11714);
   U11364 : OAI22_X1 port map( A1 => n8852, A2 => n12771, B1 => n8853, B2 => 
                           n12768, ZN => n11715);
   U11365 : AOI221_X1 port map( B1 => n12777, B2 => n12344, C1 => n12774, C2 =>
                           n12336, A => n11696, ZN => n11695);
   U11366 : OAI22_X1 port map( A1 => n8837, A2 => n12771, B1 => n8838, B2 => 
                           n12768, ZN => n11696);
   U11367 : AOI221_X1 port map( B1 => n12777, B2 => n12345, C1 => n12774, C2 =>
                           n12337, A => n11663, ZN => n11660);
   U11368 : OAI22_X1 port map( A1 => n8822, A2 => n12771, B1 => n8823, B2 => 
                           n12768, ZN => n11663);
   U11369 : AOI221_X1 port map( B1 => n12877, B2 => n12544, C1 => n12874, C2 =>
                           n12520, A => n11621, ZN => n11620);
   U11370 : OAI22_X1 port map( A1 => n9287, A2 => n12871, B1 => n9288, B2 => 
                           n12868, ZN => n11621);
   U11371 : AOI221_X1 port map( B1 => n12877, B2 => n12545, C1 => n12874, C2 =>
                           n12521, A => n11594, ZN => n11593);
   U11372 : OAI22_X1 port map( A1 => n9272, A2 => n12871, B1 => n9273, B2 => 
                           n12868, ZN => n11594);
   U11373 : AOI221_X1 port map( B1 => n12877, B2 => n12546, C1 => n12874, C2 =>
                           n12522, A => n11575, ZN => n11574);
   U11374 : OAI22_X1 port map( A1 => n9257, A2 => n12871, B1 => n9258, B2 => 
                           n12868, ZN => n11575);
   U11375 : AOI221_X1 port map( B1 => n12877, B2 => n12547, C1 => n12874, C2 =>
                           n12523, A => n11556, ZN => n11555);
   U11376 : OAI22_X1 port map( A1 => n9242, A2 => n12871, B1 => n9243, B2 => 
                           n12868, ZN => n11556);
   U11377 : AOI221_X1 port map( B1 => n12877, B2 => n12548, C1 => n12874, C2 =>
                           n12524, A => n11537, ZN => n11536);
   U11378 : OAI22_X1 port map( A1 => n9227, A2 => n12871, B1 => n9228, B2 => 
                           n12868, ZN => n11537);
   U11379 : AOI221_X1 port map( B1 => n12877, B2 => n12549, C1 => n12874, C2 =>
                           n12525, A => n11518, ZN => n11517);
   U11380 : OAI22_X1 port map( A1 => n9212, A2 => n12871, B1 => n9213, B2 => 
                           n12868, ZN => n11518);
   U11381 : AOI221_X1 port map( B1 => n12877, B2 => n12550, C1 => n12874, C2 =>
                           n12526, A => n11499, ZN => n11498);
   U11382 : OAI22_X1 port map( A1 => n9197, A2 => n12871, B1 => n9198, B2 => 
                           n12868, ZN => n11499);
   U11383 : AOI221_X1 port map( B1 => n12877, B2 => n12551, C1 => n12874, C2 =>
                           n12527, A => n11480, ZN => n11479);
   U11384 : OAI22_X1 port map( A1 => n9182, A2 => n12871, B1 => n9183, B2 => 
                           n12868, ZN => n11480);
   U11385 : AOI221_X1 port map( B1 => n12877, B2 => n12552, C1 => n12874, C2 =>
                           n12528, A => n11461, ZN => n11460);
   U11386 : OAI22_X1 port map( A1 => n9167, A2 => n12871, B1 => n9168, B2 => 
                           n12868, ZN => n11461);
   U11387 : AOI221_X1 port map( B1 => n12877, B2 => n12553, C1 => n12874, C2 =>
                           n12529, A => n11442, ZN => n11441);
   U11388 : OAI22_X1 port map( A1 => n9152, A2 => n12871, B1 => n9153, B2 => 
                           n12868, ZN => n11442);
   U11389 : AOI221_X1 port map( B1 => n12877, B2 => n12554, C1 => n12874, C2 =>
                           n12530, A => n11423, ZN => n11422);
   U11390 : OAI22_X1 port map( A1 => n9137, A2 => n12871, B1 => n9138, B2 => 
                           n12868, ZN => n11423);
   U11391 : AOI221_X1 port map( B1 => n12877, B2 => n12555, C1 => n12874, C2 =>
                           n12531, A => n11404, ZN => n11403);
   U11392 : OAI22_X1 port map( A1 => n9122, A2 => n12871, B1 => n9123, B2 => 
                           n12868, ZN => n11404);
   U11393 : AOI221_X1 port map( B1 => n12878, B2 => n12556, C1 => n12875, C2 =>
                           n12532, A => n11385, ZN => n11384);
   U11394 : OAI22_X1 port map( A1 => n9107, A2 => n12872, B1 => n9108, B2 => 
                           n12869, ZN => n11385);
   U11395 : AOI221_X1 port map( B1 => n12878, B2 => n12557, C1 => n12875, C2 =>
                           n12533, A => n11366, ZN => n11365);
   U11396 : OAI22_X1 port map( A1 => n9092, A2 => n12872, B1 => n9093, B2 => 
                           n12869, ZN => n11366);
   U11397 : AOI221_X1 port map( B1 => n12878, B2 => n12558, C1 => n12875, C2 =>
                           n12534, A => n11347, ZN => n11346);
   U11398 : OAI22_X1 port map( A1 => n9077, A2 => n12872, B1 => n9078, B2 => 
                           n12869, ZN => n11347);
   U11399 : AOI221_X1 port map( B1 => n12878, B2 => n12559, C1 => n12875, C2 =>
                           n12535, A => n11328, ZN => n11327);
   U11400 : OAI22_X1 port map( A1 => n9062, A2 => n12872, B1 => n9063, B2 => 
                           n12869, ZN => n11328);
   U11401 : AOI221_X1 port map( B1 => n12878, B2 => n12560, C1 => n12875, C2 =>
                           n12536, A => n11309, ZN => n11308);
   U11402 : OAI22_X1 port map( A1 => n9047, A2 => n12872, B1 => n9048, B2 => 
                           n12869, ZN => n11309);
   U11403 : AOI221_X1 port map( B1 => n12878, B2 => n12561, C1 => n12875, C2 =>
                           n12537, A => n11290, ZN => n11289);
   U11404 : OAI22_X1 port map( A1 => n9032, A2 => n12872, B1 => n9033, B2 => 
                           n12869, ZN => n11290);
   U11405 : AOI221_X1 port map( B1 => n12878, B2 => n12562, C1 => n12875, C2 =>
                           n12538, A => n11271, ZN => n11270);
   U11406 : OAI22_X1 port map( A1 => n9017, A2 => n12872, B1 => n9018, B2 => 
                           n12869, ZN => n11271);
   U11407 : AOI221_X1 port map( B1 => n12878, B2 => n12563, C1 => n12875, C2 =>
                           n12539, A => n11252, ZN => n11251);
   U11408 : OAI22_X1 port map( A1 => n9002, A2 => n12872, B1 => n9003, B2 => 
                           n12869, ZN => n11252);
   U11409 : AOI221_X1 port map( B1 => n12878, B2 => n12564, C1 => n12875, C2 =>
                           n12540, A => n11233, ZN => n11232);
   U11410 : OAI22_X1 port map( A1 => n8987, A2 => n12872, B1 => n8988, B2 => 
                           n12869, ZN => n11233);
   U11411 : AOI221_X1 port map( B1 => n12878, B2 => n12565, C1 => n12875, C2 =>
                           n12541, A => n11214, ZN => n11213);
   U11412 : OAI22_X1 port map( A1 => n8972, A2 => n12872, B1 => n8973, B2 => 
                           n12869, ZN => n11214);
   U11413 : AOI221_X1 port map( B1 => n12878, B2 => n12566, C1 => n12875, C2 =>
                           n12542, A => n11195, ZN => n11194);
   U11414 : OAI22_X1 port map( A1 => n8957, A2 => n12872, B1 => n8958, B2 => 
                           n12869, ZN => n11195);
   U11415 : AOI221_X1 port map( B1 => n12878, B2 => n12567, C1 => n12875, C2 =>
                           n12543, A => n11176, ZN => n11175);
   U11416 : OAI22_X1 port map( A1 => n8942, A2 => n12872, B1 => n8943, B2 => 
                           n12869, ZN => n11176);
   U11417 : AOI221_X1 port map( B1 => n12879, B2 => n12338, C1 => n12876, C2 =>
                           n12330, A => n11157, ZN => n11156);
   U11418 : OAI22_X1 port map( A1 => n8927, A2 => n12873, B1 => n8928, B2 => 
                           n12870, ZN => n11157);
   U11419 : AOI221_X1 port map( B1 => n12879, B2 => n12339, C1 => n12876, C2 =>
                           n12331, A => n11138, ZN => n11137);
   U11420 : OAI22_X1 port map( A1 => n8912, A2 => n12873, B1 => n8913, B2 => 
                           n12870, ZN => n11138);
   U11421 : AOI221_X1 port map( B1 => n12879, B2 => n12340, C1 => n12876, C2 =>
                           n12332, A => n11119, ZN => n11118);
   U11422 : OAI22_X1 port map( A1 => n8897, A2 => n12873, B1 => n8898, B2 => 
                           n12870, ZN => n11119);
   U11423 : AOI221_X1 port map( B1 => n12879, B2 => n12341, C1 => n12876, C2 =>
                           n12333, A => n11100, ZN => n11099);
   U11424 : OAI22_X1 port map( A1 => n8882, A2 => n12873, B1 => n8883, B2 => 
                           n12870, ZN => n11100);
   U11425 : AOI221_X1 port map( B1 => n12879, B2 => n12342, C1 => n12876, C2 =>
                           n12334, A => n11081, ZN => n11080);
   U11426 : OAI22_X1 port map( A1 => n8867, A2 => n12873, B1 => n8868, B2 => 
                           n12870, ZN => n11081);
   U11427 : AOI221_X1 port map( B1 => n12879, B2 => n12343, C1 => n12876, C2 =>
                           n12335, A => n11062, ZN => n11061);
   U11428 : OAI22_X1 port map( A1 => n8852, A2 => n12873, B1 => n8853, B2 => 
                           n12870, ZN => n11062);
   U11429 : AOI221_X1 port map( B1 => n12879, B2 => n12344, C1 => n12876, C2 =>
                           n12336, A => n11043, ZN => n11042);
   U11430 : OAI22_X1 port map( A1 => n8837, A2 => n12873, B1 => n8838, B2 => 
                           n12870, ZN => n11043);
   U11431 : AOI221_X1 port map( B1 => n12879, B2 => n12345, C1 => n12876, C2 =>
                           n12337, A => n11010, ZN => n11007);
   U11432 : OAI22_X1 port map( A1 => n8822, A2 => n12873, B1 => n8823, B2 => 
                           n12870, ZN => n11010);
   U11433 : AOI221_X1 port map( B1 => n12799, B2 => n10810, C1 => n12796, C2 =>
                           n10746, A => n12266, ZN => n12255);
   U11434 : OAI22_X1 port map( A1 => n6695, A2 => n12793, B1 => n6663, B2 => 
                           n12790, ZN => n12266);
   U11435 : AOI221_X1 port map( B1 => n12799, B2 => n10809, C1 => n12796, C2 =>
                           n10745, A => n12241, ZN => n12236);
   U11436 : OAI22_X1 port map( A1 => n6694, A2 => n12793, B1 => n6662, B2 => 
                           n12790, ZN => n12241);
   U11437 : AOI221_X1 port map( B1 => n12799, B2 => n10808, C1 => n12796, C2 =>
                           n10744, A => n12222, ZN => n12217);
   U11438 : OAI22_X1 port map( A1 => n6693, A2 => n12793, B1 => n6661, B2 => 
                           n12790, ZN => n12222);
   U11439 : AOI221_X1 port map( B1 => n12799, B2 => n10807, C1 => n12796, C2 =>
                           n10743, A => n12203, ZN => n12198);
   U11440 : OAI22_X1 port map( A1 => n6692, A2 => n12793, B1 => n6660, B2 => 
                           n12790, ZN => n12203);
   U11441 : AOI221_X1 port map( B1 => n12799, B2 => n10806, C1 => n12796, C2 =>
                           n10742, A => n12184, ZN => n12179);
   U11442 : OAI22_X1 port map( A1 => n6691, A2 => n12793, B1 => n6659, B2 => 
                           n12790, ZN => n12184);
   U11443 : AOI221_X1 port map( B1 => n12799, B2 => n10805, C1 => n12796, C2 =>
                           n10741, A => n12165, ZN => n12160);
   U11444 : OAI22_X1 port map( A1 => n6690, A2 => n12793, B1 => n6658, B2 => 
                           n12790, ZN => n12165);
   U11445 : AOI221_X1 port map( B1 => n12799, B2 => n10804, C1 => n12796, C2 =>
                           n10740, A => n12146, ZN => n12141);
   U11446 : OAI22_X1 port map( A1 => n6689, A2 => n12793, B1 => n6657, B2 => 
                           n12790, ZN => n12146);
   U11447 : AOI221_X1 port map( B1 => n12799, B2 => n10803, C1 => n12796, C2 =>
                           n10739, A => n12127, ZN => n12122);
   U11448 : OAI22_X1 port map( A1 => n6688, A2 => n12793, B1 => n6656, B2 => 
                           n12790, ZN => n12127);
   U11449 : AOI221_X1 port map( B1 => n12799, B2 => n10802, C1 => n12796, C2 =>
                           n10738, A => n12108, ZN => n12103);
   U11450 : OAI22_X1 port map( A1 => n6687, A2 => n12793, B1 => n6655, B2 => 
                           n12790, ZN => n12108);
   U11451 : AOI221_X1 port map( B1 => n12799, B2 => n10801, C1 => n12796, C2 =>
                           n10737, A => n12089, ZN => n12084);
   U11452 : OAI22_X1 port map( A1 => n6686, A2 => n12793, B1 => n6654, B2 => 
                           n12790, ZN => n12089);
   U11453 : AOI221_X1 port map( B1 => n12799, B2 => n10800, C1 => n12796, C2 =>
                           n10736, A => n12070, ZN => n12065);
   U11454 : OAI22_X1 port map( A1 => n6685, A2 => n12793, B1 => n6653, B2 => 
                           n12790, ZN => n12070);
   U11455 : AOI221_X1 port map( B1 => n12799, B2 => n10799, C1 => n12796, C2 =>
                           n10735, A => n12051, ZN => n12046);
   U11456 : OAI22_X1 port map( A1 => n6684, A2 => n12793, B1 => n6652, B2 => 
                           n12790, ZN => n12051);
   U11457 : AOI221_X1 port map( B1 => n12800, B2 => n10798, C1 => n12797, C2 =>
                           n10734, A => n12032, ZN => n12027);
   U11458 : OAI22_X1 port map( A1 => n6683, A2 => n12794, B1 => n6651, B2 => 
                           n12791, ZN => n12032);
   U11459 : AOI221_X1 port map( B1 => n12800, B2 => n10797, C1 => n12797, C2 =>
                           n10733, A => n12013, ZN => n12008);
   U11460 : OAI22_X1 port map( A1 => n6682, A2 => n12794, B1 => n6650, B2 => 
                           n12791, ZN => n12013);
   U11461 : AOI221_X1 port map( B1 => n12800, B2 => n10796, C1 => n12797, C2 =>
                           n10732, A => n11994, ZN => n11989);
   U11462 : OAI22_X1 port map( A1 => n6681, A2 => n12794, B1 => n6649, B2 => 
                           n12791, ZN => n11994);
   U11463 : AOI221_X1 port map( B1 => n12800, B2 => n10795, C1 => n12797, C2 =>
                           n10731, A => n11975, ZN => n11970);
   U11464 : OAI22_X1 port map( A1 => n6680, A2 => n12794, B1 => n6648, B2 => 
                           n12791, ZN => n11975);
   U11465 : AOI221_X1 port map( B1 => n12800, B2 => n10794, C1 => n12797, C2 =>
                           n10730, A => n11956, ZN => n11951);
   U11466 : OAI22_X1 port map( A1 => n6679, A2 => n12794, B1 => n6647, B2 => 
                           n12791, ZN => n11956);
   U11467 : AOI221_X1 port map( B1 => n12800, B2 => n10793, C1 => n12797, C2 =>
                           n10729, A => n11937, ZN => n11932);
   U11468 : OAI22_X1 port map( A1 => n6678, A2 => n12794, B1 => n6646, B2 => 
                           n12791, ZN => n11937);
   U11469 : AOI221_X1 port map( B1 => n12800, B2 => n10792, C1 => n12797, C2 =>
                           n10728, A => n11918, ZN => n11913);
   U11470 : OAI22_X1 port map( A1 => n6677, A2 => n12794, B1 => n6645, B2 => 
                           n12791, ZN => n11918);
   U11471 : AOI221_X1 port map( B1 => n12800, B2 => n10791, C1 => n12797, C2 =>
                           n10727, A => n11899, ZN => n11894);
   U11472 : OAI22_X1 port map( A1 => n6676, A2 => n12794, B1 => n6644, B2 => 
                           n12791, ZN => n11899);
   U11473 : AOI221_X1 port map( B1 => n12800, B2 => n10790, C1 => n12797, C2 =>
                           n10726, A => n11880, ZN => n11875);
   U11474 : OAI22_X1 port map( A1 => n6675, A2 => n12794, B1 => n6643, B2 => 
                           n12791, ZN => n11880);
   U11475 : AOI221_X1 port map( B1 => n12800, B2 => n10789, C1 => n12797, C2 =>
                           n10725, A => n11861, ZN => n11856);
   U11476 : OAI22_X1 port map( A1 => n6674, A2 => n12794, B1 => n6642, B2 => 
                           n12791, ZN => n11861);
   U11477 : AOI221_X1 port map( B1 => n12800, B2 => n10788, C1 => n12797, C2 =>
                           n10724, A => n11842, ZN => n11837);
   U11478 : OAI22_X1 port map( A1 => n6673, A2 => n12794, B1 => n6641, B2 => 
                           n12791, ZN => n11842);
   U11479 : AOI221_X1 port map( B1 => n12800, B2 => n10787, C1 => n12797, C2 =>
                           n10723, A => n11823, ZN => n11818);
   U11480 : OAI22_X1 port map( A1 => n6672, A2 => n12794, B1 => n6640, B2 => 
                           n12791, ZN => n11823);
   U11481 : AOI221_X1 port map( B1 => n12801, B2 => n10778, C1 => n12798, C2 =>
                           n10714, A => n11804, ZN => n11799);
   U11482 : OAI22_X1 port map( A1 => n6671, A2 => n12795, B1 => n6639, B2 => 
                           n12792, ZN => n11804);
   U11483 : AOI221_X1 port map( B1 => n12801, B2 => n10777, C1 => n12798, C2 =>
                           n10713, A => n11785, ZN => n11780);
   U11484 : OAI22_X1 port map( A1 => n6670, A2 => n12795, B1 => n6638, B2 => 
                           n12792, ZN => n11785);
   U11485 : AOI221_X1 port map( B1 => n12801, B2 => n10776, C1 => n12798, C2 =>
                           n10712, A => n11766, ZN => n11761);
   U11486 : OAI22_X1 port map( A1 => n6669, A2 => n12795, B1 => n6637, B2 => 
                           n12792, ZN => n11766);
   U11487 : AOI221_X1 port map( B1 => n12801, B2 => n10775, C1 => n12798, C2 =>
                           n10711, A => n11747, ZN => n11742);
   U11488 : OAI22_X1 port map( A1 => n6668, A2 => n12795, B1 => n6636, B2 => 
                           n12792, ZN => n11747);
   U11489 : AOI221_X1 port map( B1 => n12801, B2 => n10774, C1 => n12798, C2 =>
                           n10710, A => n11728, ZN => n11723);
   U11490 : OAI22_X1 port map( A1 => n6667, A2 => n12795, B1 => n6635, B2 => 
                           n12792, ZN => n11728);
   U11491 : AOI221_X1 port map( B1 => n12801, B2 => n10773, C1 => n12798, C2 =>
                           n10709, A => n11709, ZN => n11704);
   U11492 : OAI22_X1 port map( A1 => n6666, A2 => n12795, B1 => n6634, B2 => 
                           n12792, ZN => n11709);
   U11493 : AOI221_X1 port map( B1 => n12801, B2 => n10772, C1 => n12798, C2 =>
                           n10708, A => n11690, ZN => n11685);
   U11494 : OAI22_X1 port map( A1 => n6665, A2 => n12795, B1 => n6633, B2 => 
                           n12792, ZN => n11690);
   U11495 : AOI221_X1 port map( B1 => n12801, B2 => n10771, C1 => n12798, C2 =>
                           n10707, A => n11649, ZN => n11634);
   U11496 : OAI22_X1 port map( A1 => n6664, A2 => n12795, B1 => n6632, B2 => 
                           n12792, ZN => n11649);
   U11497 : AOI221_X1 port map( B1 => n12901, B2 => n10834, C1 => n12898, C2 =>
                           n10770, A => n11613, ZN => n11602);
   U11498 : OAI22_X1 port map( A1 => n6759, A2 => n12895, B1 => n6727, B2 => 
                           n12892, ZN => n11613);
   U11499 : AOI221_X1 port map( B1 => n12901, B2 => n10833, C1 => n12898, C2 =>
                           n10769, A => n11588, ZN => n11583);
   U11500 : OAI22_X1 port map( A1 => n6758, A2 => n12895, B1 => n6726, B2 => 
                           n12892, ZN => n11588);
   U11501 : AOI221_X1 port map( B1 => n12901, B2 => n10832, C1 => n12898, C2 =>
                           n10768, A => n11569, ZN => n11564);
   U11502 : OAI22_X1 port map( A1 => n6757, A2 => n12895, B1 => n6725, B2 => 
                           n12892, ZN => n11569);
   U11503 : AOI221_X1 port map( B1 => n12901, B2 => n10831, C1 => n12898, C2 =>
                           n10767, A => n11550, ZN => n11545);
   U11504 : OAI22_X1 port map( A1 => n6756, A2 => n12895, B1 => n6724, B2 => 
                           n12892, ZN => n11550);
   U11505 : AOI221_X1 port map( B1 => n12901, B2 => n10830, C1 => n12898, C2 =>
                           n10766, A => n11531, ZN => n11526);
   U11506 : OAI22_X1 port map( A1 => n6755, A2 => n12895, B1 => n6723, B2 => 
                           n12892, ZN => n11531);
   U11507 : AOI221_X1 port map( B1 => n12901, B2 => n10829, C1 => n12898, C2 =>
                           n10765, A => n11512, ZN => n11507);
   U11508 : OAI22_X1 port map( A1 => n6754, A2 => n12895, B1 => n6722, B2 => 
                           n12892, ZN => n11512);
   U11509 : AOI221_X1 port map( B1 => n12901, B2 => n10828, C1 => n12898, C2 =>
                           n10764, A => n11493, ZN => n11488);
   U11510 : OAI22_X1 port map( A1 => n6753, A2 => n12895, B1 => n6721, B2 => 
                           n12892, ZN => n11493);
   U11511 : AOI221_X1 port map( B1 => n12901, B2 => n10827, C1 => n12898, C2 =>
                           n10763, A => n11474, ZN => n11469);
   U11512 : OAI22_X1 port map( A1 => n6752, A2 => n12895, B1 => n6720, B2 => 
                           n12892, ZN => n11474);
   U11513 : AOI221_X1 port map( B1 => n12901, B2 => n10826, C1 => n12898, C2 =>
                           n10762, A => n11455, ZN => n11450);
   U11514 : OAI22_X1 port map( A1 => n6751, A2 => n12895, B1 => n6719, B2 => 
                           n12892, ZN => n11455);
   U11515 : AOI221_X1 port map( B1 => n12901, B2 => n10825, C1 => n12898, C2 =>
                           n10761, A => n11436, ZN => n11431);
   U11516 : OAI22_X1 port map( A1 => n6750, A2 => n12895, B1 => n6718, B2 => 
                           n12892, ZN => n11436);
   U11517 : AOI221_X1 port map( B1 => n12901, B2 => n10824, C1 => n12898, C2 =>
                           n10760, A => n11417, ZN => n11412);
   U11518 : OAI22_X1 port map( A1 => n6749, A2 => n12895, B1 => n6717, B2 => 
                           n12892, ZN => n11417);
   U11519 : AOI221_X1 port map( B1 => n12901, B2 => n10823, C1 => n12898, C2 =>
                           n10759, A => n11398, ZN => n11393);
   U11520 : OAI22_X1 port map( A1 => n6748, A2 => n12895, B1 => n6716, B2 => 
                           n12892, ZN => n11398);
   U11521 : AOI221_X1 port map( B1 => n12902, B2 => n10822, C1 => n12899, C2 =>
                           n10758, A => n11379, ZN => n11374);
   U11522 : OAI22_X1 port map( A1 => n6747, A2 => n12896, B1 => n6715, B2 => 
                           n12893, ZN => n11379);
   U11523 : AOI221_X1 port map( B1 => n12902, B2 => n10821, C1 => n12899, C2 =>
                           n10757, A => n11360, ZN => n11355);
   U11524 : OAI22_X1 port map( A1 => n6746, A2 => n12896, B1 => n6714, B2 => 
                           n12893, ZN => n11360);
   U11525 : AOI221_X1 port map( B1 => n12902, B2 => n10820, C1 => n12899, C2 =>
                           n10756, A => n11341, ZN => n11336);
   U11526 : OAI22_X1 port map( A1 => n6745, A2 => n12896, B1 => n6713, B2 => 
                           n12893, ZN => n11341);
   U11527 : AOI221_X1 port map( B1 => n12902, B2 => n10819, C1 => n12899, C2 =>
                           n10755, A => n11322, ZN => n11317);
   U11528 : OAI22_X1 port map( A1 => n6744, A2 => n12896, B1 => n6712, B2 => 
                           n12893, ZN => n11322);
   U11529 : AOI221_X1 port map( B1 => n12902, B2 => n10818, C1 => n12899, C2 =>
                           n10754, A => n11303, ZN => n11298);
   U11530 : OAI22_X1 port map( A1 => n6743, A2 => n12896, B1 => n6711, B2 => 
                           n12893, ZN => n11303);
   U11531 : AOI221_X1 port map( B1 => n12902, B2 => n10817, C1 => n12899, C2 =>
                           n10753, A => n11284, ZN => n11279);
   U11532 : OAI22_X1 port map( A1 => n6742, A2 => n12896, B1 => n6710, B2 => 
                           n12893, ZN => n11284);
   U11533 : AOI221_X1 port map( B1 => n12902, B2 => n10816, C1 => n12899, C2 =>
                           n10752, A => n11265, ZN => n11260);
   U11534 : OAI22_X1 port map( A1 => n6741, A2 => n12896, B1 => n6709, B2 => 
                           n12893, ZN => n11265);
   U11535 : AOI221_X1 port map( B1 => n12902, B2 => n10815, C1 => n12899, C2 =>
                           n10751, A => n11246, ZN => n11241);
   U11536 : OAI22_X1 port map( A1 => n6740, A2 => n12896, B1 => n6708, B2 => 
                           n12893, ZN => n11246);
   U11537 : AOI221_X1 port map( B1 => n12902, B2 => n10814, C1 => n12899, C2 =>
                           n10750, A => n11227, ZN => n11222);
   U11538 : OAI22_X1 port map( A1 => n6739, A2 => n12896, B1 => n6707, B2 => 
                           n12893, ZN => n11227);
   U11539 : AOI221_X1 port map( B1 => n12902, B2 => n10813, C1 => n12899, C2 =>
                           n10749, A => n11208, ZN => n11203);
   U11540 : OAI22_X1 port map( A1 => n6738, A2 => n12896, B1 => n6706, B2 => 
                           n12893, ZN => n11208);
   U11541 : AOI221_X1 port map( B1 => n12902, B2 => n10812, C1 => n12899, C2 =>
                           n10748, A => n11189, ZN => n11184);
   U11542 : OAI22_X1 port map( A1 => n6737, A2 => n12896, B1 => n6705, B2 => 
                           n12893, ZN => n11189);
   U11543 : AOI221_X1 port map( B1 => n12902, B2 => n10811, C1 => n12899, C2 =>
                           n10747, A => n11170, ZN => n11165);
   U11544 : OAI22_X1 port map( A1 => n6736, A2 => n12896, B1 => n6704, B2 => 
                           n12893, ZN => n11170);
   U11545 : AOI221_X1 port map( B1 => n12903, B2 => n10786, C1 => n12900, C2 =>
                           n10722, A => n11151, ZN => n11146);
   U11546 : OAI22_X1 port map( A1 => n6735, A2 => n12897, B1 => n6703, B2 => 
                           n12894, ZN => n11151);
   U11547 : AOI221_X1 port map( B1 => n12903, B2 => n10785, C1 => n12900, C2 =>
                           n10721, A => n11132, ZN => n11127);
   U11548 : OAI22_X1 port map( A1 => n6734, A2 => n12897, B1 => n6702, B2 => 
                           n12894, ZN => n11132);
   U11549 : AOI221_X1 port map( B1 => n12903, B2 => n10784, C1 => n12900, C2 =>
                           n10720, A => n11113, ZN => n11108);
   U11550 : OAI22_X1 port map( A1 => n6733, A2 => n12897, B1 => n6701, B2 => 
                           n12894, ZN => n11113);
   U11551 : AOI221_X1 port map( B1 => n12903, B2 => n10783, C1 => n12900, C2 =>
                           n10719, A => n11094, ZN => n11089);
   U11552 : OAI22_X1 port map( A1 => n6732, A2 => n12897, B1 => n6700, B2 => 
                           n12894, ZN => n11094);
   U11553 : AOI221_X1 port map( B1 => n12903, B2 => n10782, C1 => n12900, C2 =>
                           n10718, A => n11075, ZN => n11070);
   U11554 : OAI22_X1 port map( A1 => n6731, A2 => n12897, B1 => n6699, B2 => 
                           n12894, ZN => n11075);
   U11555 : AOI221_X1 port map( B1 => n12903, B2 => n10781, C1 => n12900, C2 =>
                           n10717, A => n11056, ZN => n11051);
   U11556 : OAI22_X1 port map( A1 => n6730, A2 => n12897, B1 => n6698, B2 => 
                           n12894, ZN => n11056);
   U11557 : AOI221_X1 port map( B1 => n12903, B2 => n10780, C1 => n12900, C2 =>
                           n10716, A => n11037, ZN => n11032);
   U11558 : OAI22_X1 port map( A1 => n6729, A2 => n12897, B1 => n6697, B2 => 
                           n12894, ZN => n11037);
   U11559 : AOI221_X1 port map( B1 => n12903, B2 => n10779, C1 => n12900, C2 =>
                           n10715, A => n10996, ZN => n10981);
   U11560 : OAI22_X1 port map( A1 => n6728, A2 => n12897, B1 => n6696, B2 => 
                           n12894, ZN => n10996);
   U11561 : OAI22_X1 port map( A1 => n13048, A2 => n13287, B1 => n10962, B2 => 
                           n10434, ZN => n2998);
   U11562 : OAI22_X1 port map( A1 => n13049, A2 => n13290, B1 => n10962, B2 => 
                           n10433, ZN => n2999);
   U11563 : OAI22_X1 port map( A1 => n13049, A2 => n13293, B1 => n10962, B2 => 
                           n10432, ZN => n3000);
   U11564 : OAI22_X1 port map( A1 => n13049, A2 => n13296, B1 => n10962, B2 => 
                           n10431, ZN => n3001);
   U11565 : OAI22_X1 port map( A1 => n13049, A2 => n13299, B1 => n10962, B2 => 
                           n10430, ZN => n3002);
   U11566 : OAI22_X1 port map( A1 => n13049, A2 => n13302, B1 => n10962, B2 => 
                           n10429, ZN => n3003);
   U11567 : OAI22_X1 port map( A1 => n13050, A2 => n13305, B1 => n10962, B2 => 
                           n10428, ZN => n3004);
   U11568 : OAI22_X1 port map( A1 => n13050, A2 => n13317, B1 => n10962, B2 => 
                           n10427, ZN => n3005);
   U11569 : OAI22_X1 port map( A1 => n13183, A2 => n13286, B1 => n6575, B2 => 
                           n10940, ZN => n3478);
   U11570 : OAI22_X1 port map( A1 => n13184, A2 => n13289, B1 => n6574, B2 => 
                           n10940, ZN => n3479);
   U11571 : OAI22_X1 port map( A1 => n13184, A2 => n13292, B1 => n6573, B2 => 
                           n10940, ZN => n3480);
   U11572 : OAI22_X1 port map( A1 => n13184, A2 => n13295, B1 => n6572, B2 => 
                           n10940, ZN => n3481);
   U11573 : OAI22_X1 port map( A1 => n13184, A2 => n13298, B1 => n6571, B2 => 
                           n10940, ZN => n3482);
   U11574 : OAI22_X1 port map( A1 => n13184, A2 => n13301, B1 => n6570, B2 => 
                           n10940, ZN => n3483);
   U11575 : OAI22_X1 port map( A1 => n13185, A2 => n13304, B1 => n6569, B2 => 
                           n10940, ZN => n3484);
   U11576 : OAI22_X1 port map( A1 => n13185, A2 => n13316, B1 => n6568, B2 => 
                           n10940, ZN => n3485);
   U11577 : OAI22_X1 port map( A1 => n13174, A2 => n13286, B1 => n6607, B2 => 
                           n10942, ZN => n3446);
   U11578 : OAI22_X1 port map( A1 => n13175, A2 => n13289, B1 => n6606, B2 => 
                           n10942, ZN => n3447);
   U11579 : OAI22_X1 port map( A1 => n13175, A2 => n13292, B1 => n6605, B2 => 
                           n10942, ZN => n3448);
   U11580 : OAI22_X1 port map( A1 => n13175, A2 => n13295, B1 => n6604, B2 => 
                           n10942, ZN => n3449);
   U11581 : OAI22_X1 port map( A1 => n13175, A2 => n13298, B1 => n6603, B2 => 
                           n10942, ZN => n3450);
   U11582 : OAI22_X1 port map( A1 => n13175, A2 => n13301, B1 => n6602, B2 => 
                           n10942, ZN => n3451);
   U11583 : OAI22_X1 port map( A1 => n13176, A2 => n13304, B1 => n6601, B2 => 
                           n10942, ZN => n3452);
   U11584 : OAI22_X1 port map( A1 => n13176, A2 => n13316, B1 => n6600, B2 => 
                           n10942, ZN => n3453);
   U11585 : OAI22_X1 port map( A1 => n13147, A2 => n13286, B1 => n6639, B2 => 
                           n10949, ZN => n3350);
   U11586 : OAI22_X1 port map( A1 => n13148, A2 => n13289, B1 => n6638, B2 => 
                           n10949, ZN => n3351);
   U11587 : OAI22_X1 port map( A1 => n13148, A2 => n13292, B1 => n6637, B2 => 
                           n10949, ZN => n3352);
   U11588 : OAI22_X1 port map( A1 => n13148, A2 => n13295, B1 => n6636, B2 => 
                           n10949, ZN => n3353);
   U11589 : OAI22_X1 port map( A1 => n13148, A2 => n13298, B1 => n6635, B2 => 
                           n10949, ZN => n3354);
   U11590 : OAI22_X1 port map( A1 => n13148, A2 => n13301, B1 => n6634, B2 => 
                           n10949, ZN => n3355);
   U11591 : OAI22_X1 port map( A1 => n13149, A2 => n13304, B1 => n6633, B2 => 
                           n10949, ZN => n3356);
   U11592 : OAI22_X1 port map( A1 => n13149, A2 => n13316, B1 => n6632, B2 => 
                           n10949, ZN => n3357);
   U11593 : OAI22_X1 port map( A1 => n13129, A2 => n13286, B1 => n6703, B2 => 
                           n10952, ZN => n3286);
   U11594 : OAI22_X1 port map( A1 => n13130, A2 => n13289, B1 => n6702, B2 => 
                           n10952, ZN => n3287);
   U11595 : OAI22_X1 port map( A1 => n13130, A2 => n13292, B1 => n6701, B2 => 
                           n10952, ZN => n3288);
   U11596 : OAI22_X1 port map( A1 => n13130, A2 => n13295, B1 => n6700, B2 => 
                           n10952, ZN => n3289);
   U11597 : OAI22_X1 port map( A1 => n13130, A2 => n13298, B1 => n6699, B2 => 
                           n10952, ZN => n3290);
   U11598 : OAI22_X1 port map( A1 => n13130, A2 => n13301, B1 => n6698, B2 => 
                           n10952, ZN => n3291);
   U11599 : OAI22_X1 port map( A1 => n13131, A2 => n13304, B1 => n6697, B2 => 
                           n10952, ZN => n3292);
   U11600 : OAI22_X1 port map( A1 => n13131, A2 => n13316, B1 => n6696, B2 => 
                           n10952, ZN => n3293);
   U11601 : OAI22_X1 port map( A1 => n13138, A2 => n13286, B1 => n6671, B2 => 
                           n10951, ZN => n3318);
   U11602 : OAI22_X1 port map( A1 => n13139, A2 => n13289, B1 => n6670, B2 => 
                           n10951, ZN => n3319);
   U11603 : OAI22_X1 port map( A1 => n13139, A2 => n13292, B1 => n6669, B2 => 
                           n10951, ZN => n3320);
   U11604 : OAI22_X1 port map( A1 => n13139, A2 => n13295, B1 => n6668, B2 => 
                           n10951, ZN => n3321);
   U11605 : OAI22_X1 port map( A1 => n13139, A2 => n13298, B1 => n6667, B2 => 
                           n10951, ZN => n3322);
   U11606 : OAI22_X1 port map( A1 => n13139, A2 => n13301, B1 => n6666, B2 => 
                           n10951, ZN => n3323);
   U11607 : OAI22_X1 port map( A1 => n13140, A2 => n13304, B1 => n6665, B2 => 
                           n10951, ZN => n3324);
   U11608 : OAI22_X1 port map( A1 => n13140, A2 => n13316, B1 => n6664, B2 => 
                           n10951, ZN => n3325);
   U11609 : OAI22_X1 port map( A1 => n13120, A2 => n13286, B1 => n6735, B2 => 
                           n10953, ZN => n3254);
   U11610 : OAI22_X1 port map( A1 => n13121, A2 => n13289, B1 => n6734, B2 => 
                           n10953, ZN => n3255);
   U11611 : OAI22_X1 port map( A1 => n13121, A2 => n13292, B1 => n6733, B2 => 
                           n10953, ZN => n3256);
   U11612 : OAI22_X1 port map( A1 => n13121, A2 => n13295, B1 => n6732, B2 => 
                           n10953, ZN => n3257);
   U11613 : OAI22_X1 port map( A1 => n13121, A2 => n13298, B1 => n6731, B2 => 
                           n10953, ZN => n3258);
   U11614 : OAI22_X1 port map( A1 => n13121, A2 => n13301, B1 => n6730, B2 => 
                           n10953, ZN => n3259);
   U11615 : OAI22_X1 port map( A1 => n13122, A2 => n13304, B1 => n6729, B2 => 
                           n10953, ZN => n3260);
   U11616 : OAI22_X1 port map( A1 => n13122, A2 => n13316, B1 => n6728, B2 => 
                           n10953, ZN => n3261);
   U11617 : OAI22_X1 port map( A1 => n13201, A2 => n13286, B1 => n8921, B2 => 
                           n10936, ZN => n3542);
   U11618 : OAI22_X1 port map( A1 => n13202, A2 => n13289, B1 => n8906, B2 => 
                           n10936, ZN => n3543);
   U11619 : OAI22_X1 port map( A1 => n13202, A2 => n13292, B1 => n8891, B2 => 
                           n10936, ZN => n3544);
   U11620 : OAI22_X1 port map( A1 => n13202, A2 => n13295, B1 => n8876, B2 => 
                           n10936, ZN => n3545);
   U11621 : OAI22_X1 port map( A1 => n13202, A2 => n13298, B1 => n8861, B2 => 
                           n10936, ZN => n3546);
   U11622 : OAI22_X1 port map( A1 => n13202, A2 => n13301, B1 => n8846, B2 => 
                           n10936, ZN => n3547);
   U11623 : OAI22_X1 port map( A1 => n13203, A2 => n13304, B1 => n8831, B2 => 
                           n10936, ZN => n3548);
   U11624 : OAI22_X1 port map( A1 => n13203, A2 => n13316, B1 => n8816, B2 => 
                           n10936, ZN => n3549);
   U11625 : OAI22_X1 port map( A1 => n13192, A2 => n13286, B1 => n8922, B2 => 
                           n10938, ZN => n3510);
   U11626 : OAI22_X1 port map( A1 => n13193, A2 => n13289, B1 => n8907, B2 => 
                           n10938, ZN => n3511);
   U11627 : OAI22_X1 port map( A1 => n13193, A2 => n13292, B1 => n8892, B2 => 
                           n10938, ZN => n3512);
   U11628 : OAI22_X1 port map( A1 => n13193, A2 => n13295, B1 => n8877, B2 => 
                           n10938, ZN => n3513);
   U11629 : OAI22_X1 port map( A1 => n13193, A2 => n13298, B1 => n8862, B2 => 
                           n10938, ZN => n3514);
   U11630 : OAI22_X1 port map( A1 => n13193, A2 => n13301, B1 => n8847, B2 => 
                           n10938, ZN => n3515);
   U11631 : OAI22_X1 port map( A1 => n13194, A2 => n13304, B1 => n8832, B2 => 
                           n10938, ZN => n3516);
   U11632 : OAI22_X1 port map( A1 => n13194, A2 => n13316, B1 => n8817, B2 => 
                           n10938, ZN => n3517);
   U11633 : OAI22_X1 port map( A1 => n13111, A2 => n13287, B1 => n8926, B2 => 
                           n10954, ZN => n3222);
   U11634 : OAI22_X1 port map( A1 => n13112, A2 => n13290, B1 => n8911, B2 => 
                           n10954, ZN => n3223);
   U11635 : OAI22_X1 port map( A1 => n13112, A2 => n13293, B1 => n8896, B2 => 
                           n10954, ZN => n3224);
   U11636 : OAI22_X1 port map( A1 => n13112, A2 => n13296, B1 => n8881, B2 => 
                           n10954, ZN => n3225);
   U11637 : OAI22_X1 port map( A1 => n13112, A2 => n13299, B1 => n8866, B2 => 
                           n10954, ZN => n3226);
   U11638 : OAI22_X1 port map( A1 => n13112, A2 => n13302, B1 => n8851, B2 => 
                           n10954, ZN => n3227);
   U11639 : OAI22_X1 port map( A1 => n13113, A2 => n13305, B1 => n8836, B2 => 
                           n10954, ZN => n3228);
   U11640 : OAI22_X1 port map( A1 => n13113, A2 => n13317, B1 => n8821, B2 => 
                           n10954, ZN => n3229);
   U11641 : OAI22_X1 port map( A1 => n13102, A2 => n13287, B1 => n8925, B2 => 
                           n10955, ZN => n3190);
   U11642 : OAI22_X1 port map( A1 => n13103, A2 => n13290, B1 => n8910, B2 => 
                           n10955, ZN => n3191);
   U11643 : OAI22_X1 port map( A1 => n13103, A2 => n13293, B1 => n8895, B2 => 
                           n10955, ZN => n3192);
   U11644 : OAI22_X1 port map( A1 => n13103, A2 => n13296, B1 => n8880, B2 => 
                           n10955, ZN => n3193);
   U11645 : OAI22_X1 port map( A1 => n13103, A2 => n13299, B1 => n8865, B2 => 
                           n10955, ZN => n3194);
   U11646 : OAI22_X1 port map( A1 => n13103, A2 => n13302, B1 => n8850, B2 => 
                           n10955, ZN => n3195);
   U11647 : OAI22_X1 port map( A1 => n13104, A2 => n13305, B1 => n8835, B2 => 
                           n10955, ZN => n3196);
   U11648 : OAI22_X1 port map( A1 => n13104, A2 => n13317, B1 => n8820, B2 => 
                           n10955, ZN => n3197);
   U11649 : OAI22_X1 port map( A1 => n13075, A2 => n13287, B1 => n8928, B2 => 
                           n10958, ZN => n3094);
   U11650 : OAI22_X1 port map( A1 => n13076, A2 => n13290, B1 => n8913, B2 => 
                           n10958, ZN => n3095);
   U11651 : OAI22_X1 port map( A1 => n13076, A2 => n13293, B1 => n8898, B2 => 
                           n10958, ZN => n3096);
   U11652 : OAI22_X1 port map( A1 => n13076, A2 => n13296, B1 => n8883, B2 => 
                           n10958, ZN => n3097);
   U11653 : OAI22_X1 port map( A1 => n13076, A2 => n13299, B1 => n8868, B2 => 
                           n10958, ZN => n3098);
   U11654 : OAI22_X1 port map( A1 => n13076, A2 => n13302, B1 => n8853, B2 => 
                           n10958, ZN => n3099);
   U11655 : OAI22_X1 port map( A1 => n13077, A2 => n13305, B1 => n8838, B2 => 
                           n10958, ZN => n3100);
   U11656 : OAI22_X1 port map( A1 => n13077, A2 => n13317, B1 => n8823, B2 => 
                           n10958, ZN => n3101);
   U11657 : OAI22_X1 port map( A1 => n13066, A2 => n13287, B1 => n8927, B2 => 
                           n10960, ZN => n3062);
   U11658 : OAI22_X1 port map( A1 => n13067, A2 => n13290, B1 => n8912, B2 => 
                           n10960, ZN => n3063);
   U11659 : OAI22_X1 port map( A1 => n13067, A2 => n13293, B1 => n8897, B2 => 
                           n10960, ZN => n3064);
   U11660 : OAI22_X1 port map( A1 => n13067, A2 => n13296, B1 => n8882, B2 => 
                           n10960, ZN => n3065);
   U11661 : OAI22_X1 port map( A1 => n13067, A2 => n13299, B1 => n8867, B2 => 
                           n10960, ZN => n3066);
   U11662 : OAI22_X1 port map( A1 => n13067, A2 => n13302, B1 => n8852, B2 => 
                           n10960, ZN => n3067);
   U11663 : OAI22_X1 port map( A1 => n13068, A2 => n13305, B1 => n8837, B2 => 
                           n10960, ZN => n3068);
   U11664 : OAI22_X1 port map( A1 => n13068, A2 => n13317, B1 => n8822, B2 => 
                           n10960, ZN => n3069);
   U11665 : OAI22_X1 port map( A1 => n13039, A2 => n13287, B1 => n8930, B2 => 
                           n10963, ZN => n2966);
   U11666 : OAI22_X1 port map( A1 => n13040, A2 => n13290, B1 => n8915, B2 => 
                           n10963, ZN => n2967);
   U11667 : OAI22_X1 port map( A1 => n13040, A2 => n13293, B1 => n8900, B2 => 
                           n10963, ZN => n2968);
   U11668 : OAI22_X1 port map( A1 => n13040, A2 => n13296, B1 => n8885, B2 => 
                           n10963, ZN => n2969);
   U11669 : OAI22_X1 port map( A1 => n13040, A2 => n13299, B1 => n8870, B2 => 
                           n10963, ZN => n2970);
   U11670 : OAI22_X1 port map( A1 => n13040, A2 => n13302, B1 => n8855, B2 => 
                           n10963, ZN => n2971);
   U11671 : OAI22_X1 port map( A1 => n13041, A2 => n13305, B1 => n8840, B2 => 
                           n10963, ZN => n2972);
   U11672 : OAI22_X1 port map( A1 => n13041, A2 => n13317, B1 => n8825, B2 => 
                           n10963, ZN => n2973);
   U11673 : OAI22_X1 port map( A1 => n13030, A2 => n13287, B1 => n8929, B2 => 
                           n10964, ZN => n2934);
   U11674 : OAI22_X1 port map( A1 => n13031, A2 => n13290, B1 => n8914, B2 => 
                           n10964, ZN => n2935);
   U11675 : OAI22_X1 port map( A1 => n13031, A2 => n13293, B1 => n8899, B2 => 
                           n10964, ZN => n2936);
   U11676 : OAI22_X1 port map( A1 => n13031, A2 => n13296, B1 => n8884, B2 => 
                           n10964, ZN => n2937);
   U11677 : OAI22_X1 port map( A1 => n13031, A2 => n13299, B1 => n8869, B2 => 
                           n10964, ZN => n2938);
   U11678 : OAI22_X1 port map( A1 => n13031, A2 => n13302, B1 => n8854, B2 => 
                           n10964, ZN => n2939);
   U11679 : OAI22_X1 port map( A1 => n13032, A2 => n13305, B1 => n8839, B2 => 
                           n10964, ZN => n2940);
   U11680 : OAI22_X1 port map( A1 => n13032, A2 => n13317, B1 => n8824, B2 => 
                           n10964, ZN => n2941);
   U11681 : OAI22_X1 port map( A1 => n12985, A2 => n13288, B1 => n8932, B2 => 
                           n10970, ZN => n2774);
   U11682 : OAI22_X1 port map( A1 => n12986, A2 => n13291, B1 => n8917, B2 => 
                           n10970, ZN => n2775);
   U11683 : OAI22_X1 port map( A1 => n12986, A2 => n13294, B1 => n8902, B2 => 
                           n10970, ZN => n2776);
   U11684 : OAI22_X1 port map( A1 => n12986, A2 => n13297, B1 => n8887, B2 => 
                           n10970, ZN => n2777);
   U11685 : OAI22_X1 port map( A1 => n12986, A2 => n13300, B1 => n8872, B2 => 
                           n10970, ZN => n2778);
   U11686 : OAI22_X1 port map( A1 => n12986, A2 => n13303, B1 => n8857, B2 => 
                           n10970, ZN => n2779);
   U11687 : OAI22_X1 port map( A1 => n12987, A2 => n13306, B1 => n8842, B2 => 
                           n10970, ZN => n2780);
   U11688 : OAI22_X1 port map( A1 => n12987, A2 => n13318, B1 => n8827, B2 => 
                           n10970, ZN => n2781);
   U11689 : OAI22_X1 port map( A1 => n12976, A2 => n13288, B1 => n8931, B2 => 
                           n10971, ZN => n2742);
   U11690 : OAI22_X1 port map( A1 => n12977, A2 => n13291, B1 => n8916, B2 => 
                           n10971, ZN => n2743);
   U11691 : OAI22_X1 port map( A1 => n12977, A2 => n13294, B1 => n8901, B2 => 
                           n10971, ZN => n2744);
   U11692 : OAI22_X1 port map( A1 => n12977, A2 => n13297, B1 => n8886, B2 => 
                           n10971, ZN => n2745);
   U11693 : OAI22_X1 port map( A1 => n12977, A2 => n13300, B1 => n8871, B2 => 
                           n10971, ZN => n2746);
   U11694 : OAI22_X1 port map( A1 => n12977, A2 => n13303, B1 => n8856, B2 => 
                           n10971, ZN => n2747);
   U11695 : OAI22_X1 port map( A1 => n12978, A2 => n13306, B1 => n8841, B2 => 
                           n10971, ZN => n2748);
   U11696 : OAI22_X1 port map( A1 => n12978, A2 => n13318, B1 => n8826, B2 => 
                           n10971, ZN => n2749);
   U11697 : OAI22_X1 port map( A1 => n12949, A2 => n13288, B1 => n8934, B2 => 
                           n10974, ZN => n2646);
   U11698 : OAI22_X1 port map( A1 => n12950, A2 => n13291, B1 => n8919, B2 => 
                           n10974, ZN => n2647);
   U11699 : OAI22_X1 port map( A1 => n12950, A2 => n13294, B1 => n8904, B2 => 
                           n10974, ZN => n2648);
   U11700 : OAI22_X1 port map( A1 => n12950, A2 => n13297, B1 => n8889, B2 => 
                           n10974, ZN => n2649);
   U11701 : OAI22_X1 port map( A1 => n12950, A2 => n13300, B1 => n8874, B2 => 
                           n10974, ZN => n2650);
   U11702 : OAI22_X1 port map( A1 => n12950, A2 => n13303, B1 => n8859, B2 => 
                           n10974, ZN => n2651);
   U11703 : OAI22_X1 port map( A1 => n12951, A2 => n13306, B1 => n8844, B2 => 
                           n10974, ZN => n2652);
   U11704 : OAI22_X1 port map( A1 => n12951, A2 => n13318, B1 => n8829, B2 => 
                           n10974, ZN => n2653);
   U11705 : OAI22_X1 port map( A1 => n13044, A2 => n13215, B1 => n13043, B2 => 
                           n10669, ZN => n2974);
   U11706 : OAI22_X1 port map( A1 => n13044, A2 => n13218, B1 => n13043, B2 => 
                           n10668, ZN => n2975);
   U11707 : OAI22_X1 port map( A1 => n13044, A2 => n13221, B1 => n13043, B2 => 
                           n10667, ZN => n2976);
   U11708 : OAI22_X1 port map( A1 => n13044, A2 => n13224, B1 => n13043, B2 => 
                           n10666, ZN => n2977);
   U11709 : OAI22_X1 port map( A1 => n13044, A2 => n13227, B1 => n13043, B2 => 
                           n10665, ZN => n2978);
   U11710 : OAI22_X1 port map( A1 => n13045, A2 => n13230, B1 => n13043, B2 => 
                           n10664, ZN => n2979);
   U11711 : OAI22_X1 port map( A1 => n13045, A2 => n13233, B1 => n13043, B2 => 
                           n10663, ZN => n2980);
   U11712 : OAI22_X1 port map( A1 => n13045, A2 => n13236, B1 => n13043, B2 => 
                           n10662, ZN => n2981);
   U11713 : OAI22_X1 port map( A1 => n13045, A2 => n13239, B1 => n13043, B2 => 
                           n10661, ZN => n2982);
   U11714 : OAI22_X1 port map( A1 => n13045, A2 => n13242, B1 => n13043, B2 => 
                           n10660, ZN => n2983);
   U11715 : OAI22_X1 port map( A1 => n13046, A2 => n13245, B1 => n13043, B2 => 
                           n10659, ZN => n2984);
   U11716 : OAI22_X1 port map( A1 => n13046, A2 => n13248, B1 => n13043, B2 => 
                           n10658, ZN => n2985);
   U11717 : OAI22_X1 port map( A1 => n13046, A2 => n13251, B1 => n10962, B2 => 
                           n10657, ZN => n2986);
   U11718 : OAI22_X1 port map( A1 => n13046, A2 => n13254, B1 => n10962, B2 => 
                           n10656, ZN => n2987);
   U11719 : OAI22_X1 port map( A1 => n13046, A2 => n13257, B1 => n10962, B2 => 
                           n10655, ZN => n2988);
   U11720 : OAI22_X1 port map( A1 => n13047, A2 => n13260, B1 => n13043, B2 => 
                           n10654, ZN => n2989);
   U11721 : OAI22_X1 port map( A1 => n13047, A2 => n13263, B1 => n13043, B2 => 
                           n10653, ZN => n2990);
   U11722 : OAI22_X1 port map( A1 => n13047, A2 => n13266, B1 => n13043, B2 => 
                           n10652, ZN => n2991);
   U11723 : OAI22_X1 port map( A1 => n13047, A2 => n13269, B1 => n13043, B2 => 
                           n10651, ZN => n2992);
   U11724 : OAI22_X1 port map( A1 => n13047, A2 => n13272, B1 => n13043, B2 => 
                           n10650, ZN => n2993);
   U11725 : OAI22_X1 port map( A1 => n13048, A2 => n13275, B1 => n13043, B2 => 
                           n10649, ZN => n2994);
   U11726 : OAI22_X1 port map( A1 => n13048, A2 => n13278, B1 => n13043, B2 => 
                           n10648, ZN => n2995);
   U11727 : OAI22_X1 port map( A1 => n13048, A2 => n13281, B1 => n13043, B2 => 
                           n10647, ZN => n2996);
   U11728 : OAI22_X1 port map( A1 => n13048, A2 => n13284, B1 => n13043, B2 => 
                           n10646, ZN => n2997);
   U11729 : OAI22_X1 port map( A1 => n9293, A2 => n10975, B1 => n12935, B2 => 
                           n13216, ZN => n2590);
   U11730 : OAI22_X1 port map( A1 => n9278, A2 => n12934, B1 => n12935, B2 => 
                           n13219, ZN => n2591);
   U11731 : OAI22_X1 port map( A1 => n9263, A2 => n12934, B1 => n12935, B2 => 
                           n13222, ZN => n2592);
   U11732 : OAI22_X1 port map( A1 => n9248, A2 => n12934, B1 => n12935, B2 => 
                           n13225, ZN => n2593);
   U11733 : OAI22_X1 port map( A1 => n9233, A2 => n12934, B1 => n12936, B2 => 
                           n13228, ZN => n2594);
   U11734 : OAI22_X1 port map( A1 => n9218, A2 => n12934, B1 => n12936, B2 => 
                           n13231, ZN => n2595);
   U11735 : OAI22_X1 port map( A1 => n9203, A2 => n12934, B1 => n12936, B2 => 
                           n13234, ZN => n2596);
   U11736 : OAI22_X1 port map( A1 => n9188, A2 => n12934, B1 => n12936, B2 => 
                           n13237, ZN => n2597);
   U11737 : OAI22_X1 port map( A1 => n9173, A2 => n12934, B1 => n12937, B2 => 
                           n13240, ZN => n2598);
   U11738 : OAI22_X1 port map( A1 => n9158, A2 => n12934, B1 => n12937, B2 => 
                           n13243, ZN => n2599);
   U11739 : OAI22_X1 port map( A1 => n9143, A2 => n12934, B1 => n12937, B2 => 
                           n13246, ZN => n2600);
   U11740 : OAI22_X1 port map( A1 => n9128, A2 => n12934, B1 => n12937, B2 => 
                           n13249, ZN => n2601);
   U11741 : OAI22_X1 port map( A1 => n9113, A2 => n10975, B1 => n12938, B2 => 
                           n13252, ZN => n2602);
   U11742 : OAI22_X1 port map( A1 => n9098, A2 => n12934, B1 => n12938, B2 => 
                           n13255, ZN => n2603);
   U11743 : OAI22_X1 port map( A1 => n9083, A2 => n10975, B1 => n12938, B2 => 
                           n13258, ZN => n2604);
   U11744 : OAI22_X1 port map( A1 => n9068, A2 => n12934, B1 => n12938, B2 => 
                           n13261, ZN => n2605);
   U11745 : OAI22_X1 port map( A1 => n9053, A2 => n10975, B1 => n12939, B2 => 
                           n13264, ZN => n2606);
   U11746 : OAI22_X1 port map( A1 => n9038, A2 => n12934, B1 => n12939, B2 => 
                           n13267, ZN => n2607);
   U11747 : OAI22_X1 port map( A1 => n9023, A2 => n10975, B1 => n12939, B2 => 
                           n13270, ZN => n2608);
   U11748 : OAI22_X1 port map( A1 => n9008, A2 => n12934, B1 => n12939, B2 => 
                           n13273, ZN => n2609);
   U11749 : OAI22_X1 port map( A1 => n8993, A2 => n10975, B1 => n12940, B2 => 
                           n13276, ZN => n2610);
   U11750 : OAI22_X1 port map( A1 => n8978, A2 => n12934, B1 => n12940, B2 => 
                           n13279, ZN => n2611);
   U11751 : OAI22_X1 port map( A1 => n8963, A2 => n10975, B1 => n12940, B2 => 
                           n13282, ZN => n2612);
   U11752 : OAI22_X1 port map( A1 => n8948, A2 => n12934, B1 => n12940, B2 => 
                           n13285, ZN => n2613);
   U11753 : OAI22_X1 port map( A1 => n8933, A2 => n10975, B1 => n12941, B2 => 
                           n13288, ZN => n2614);
   U11754 : OAI22_X1 port map( A1 => n8918, A2 => n12934, B1 => n12941, B2 => 
                           n13291, ZN => n2615);
   U11755 : OAI22_X1 port map( A1 => n8903, A2 => n10975, B1 => n12941, B2 => 
                           n13294, ZN => n2616);
   U11756 : OAI22_X1 port map( A1 => n8888, A2 => n12934, B1 => n12941, B2 => 
                           n13297, ZN => n2617);
   U11757 : OAI22_X1 port map( A1 => n8873, A2 => n10975, B1 => n12942, B2 => 
                           n13300, ZN => n2618);
   U11758 : OAI22_X1 port map( A1 => n8858, A2 => n12934, B1 => n12942, B2 => 
                           n13303, ZN => n2619);
   U11759 : OAI22_X1 port map( A1 => n8843, A2 => n10975, B1 => n12942, B2 => 
                           n13306, ZN => n2620);
   U11760 : OAI22_X1 port map( A1 => n8828, A2 => n12934, B1 => n12942, B2 => 
                           n13318, ZN => n2621);
   U11761 : OAI22_X1 port map( A1 => n13179, A2 => n13214, B1 => n6599, B2 => 
                           n13178, ZN => n3454);
   U11762 : OAI22_X1 port map( A1 => n13179, A2 => n13217, B1 => n6598, B2 => 
                           n13178, ZN => n3455);
   U11763 : OAI22_X1 port map( A1 => n13179, A2 => n13220, B1 => n6597, B2 => 
                           n13178, ZN => n3456);
   U11764 : OAI22_X1 port map( A1 => n13179, A2 => n13223, B1 => n6596, B2 => 
                           n13178, ZN => n3457);
   U11765 : OAI22_X1 port map( A1 => n13179, A2 => n13226, B1 => n6595, B2 => 
                           n13178, ZN => n3458);
   U11766 : OAI22_X1 port map( A1 => n13180, A2 => n13229, B1 => n6594, B2 => 
                           n13178, ZN => n3459);
   U11767 : OAI22_X1 port map( A1 => n13180, A2 => n13232, B1 => n6593, B2 => 
                           n13178, ZN => n3460);
   U11768 : OAI22_X1 port map( A1 => n13180, A2 => n13235, B1 => n6592, B2 => 
                           n13178, ZN => n3461);
   U11769 : OAI22_X1 port map( A1 => n13180, A2 => n13238, B1 => n6591, B2 => 
                           n13178, ZN => n3462);
   U11770 : OAI22_X1 port map( A1 => n13180, A2 => n13241, B1 => n6590, B2 => 
                           n13178, ZN => n3463);
   U11771 : OAI22_X1 port map( A1 => n13181, A2 => n13244, B1 => n6589, B2 => 
                           n13178, ZN => n3464);
   U11772 : OAI22_X1 port map( A1 => n13181, A2 => n13247, B1 => n6588, B2 => 
                           n13178, ZN => n3465);
   U11773 : OAI22_X1 port map( A1 => n13181, A2 => n13250, B1 => n6587, B2 => 
                           n10940, ZN => n3466);
   U11774 : OAI22_X1 port map( A1 => n13181, A2 => n13253, B1 => n6586, B2 => 
                           n10940, ZN => n3467);
   U11775 : OAI22_X1 port map( A1 => n13181, A2 => n13256, B1 => n6585, B2 => 
                           n10940, ZN => n3468);
   U11776 : OAI22_X1 port map( A1 => n13182, A2 => n13259, B1 => n6584, B2 => 
                           n13178, ZN => n3469);
   U11777 : OAI22_X1 port map( A1 => n13182, A2 => n13262, B1 => n6583, B2 => 
                           n13178, ZN => n3470);
   U11778 : OAI22_X1 port map( A1 => n13182, A2 => n13265, B1 => n6582, B2 => 
                           n13178, ZN => n3471);
   U11779 : OAI22_X1 port map( A1 => n13182, A2 => n13268, B1 => n6581, B2 => 
                           n13178, ZN => n3472);
   U11780 : OAI22_X1 port map( A1 => n13182, A2 => n13271, B1 => n6580, B2 => 
                           n13178, ZN => n3473);
   U11781 : OAI22_X1 port map( A1 => n13183, A2 => n13274, B1 => n6579, B2 => 
                           n13178, ZN => n3474);
   U11782 : OAI22_X1 port map( A1 => n13183, A2 => n13277, B1 => n6578, B2 => 
                           n13178, ZN => n3475);
   U11783 : OAI22_X1 port map( A1 => n13183, A2 => n13280, B1 => n6577, B2 => 
                           n13178, ZN => n3476);
   U11784 : OAI22_X1 port map( A1 => n13183, A2 => n13283, B1 => n6576, B2 => 
                           n13178, ZN => n3477);
   U11785 : OAI22_X1 port map( A1 => n13170, A2 => n13214, B1 => n6631, B2 => 
                           n13169, ZN => n3422);
   U11786 : OAI22_X1 port map( A1 => n13170, A2 => n13217, B1 => n6630, B2 => 
                           n13169, ZN => n3423);
   U11787 : OAI22_X1 port map( A1 => n13170, A2 => n13220, B1 => n6629, B2 => 
                           n13169, ZN => n3424);
   U11788 : OAI22_X1 port map( A1 => n13170, A2 => n13223, B1 => n6628, B2 => 
                           n13169, ZN => n3425);
   U11789 : OAI22_X1 port map( A1 => n13170, A2 => n13226, B1 => n6627, B2 => 
                           n13169, ZN => n3426);
   U11790 : OAI22_X1 port map( A1 => n13171, A2 => n13229, B1 => n6626, B2 => 
                           n13169, ZN => n3427);
   U11791 : OAI22_X1 port map( A1 => n13171, A2 => n13232, B1 => n6625, B2 => 
                           n13169, ZN => n3428);
   U11792 : OAI22_X1 port map( A1 => n13171, A2 => n13235, B1 => n6624, B2 => 
                           n13169, ZN => n3429);
   U11793 : OAI22_X1 port map( A1 => n13171, A2 => n13238, B1 => n6623, B2 => 
                           n13169, ZN => n3430);
   U11794 : OAI22_X1 port map( A1 => n13171, A2 => n13241, B1 => n6622, B2 => 
                           n13169, ZN => n3431);
   U11795 : OAI22_X1 port map( A1 => n13172, A2 => n13244, B1 => n6621, B2 => 
                           n13169, ZN => n3432);
   U11796 : OAI22_X1 port map( A1 => n13172, A2 => n13247, B1 => n6620, B2 => 
                           n13169, ZN => n3433);
   U11797 : OAI22_X1 port map( A1 => n13172, A2 => n13250, B1 => n6619, B2 => 
                           n10942, ZN => n3434);
   U11798 : OAI22_X1 port map( A1 => n13172, A2 => n13253, B1 => n6618, B2 => 
                           n10942, ZN => n3435);
   U11799 : OAI22_X1 port map( A1 => n13172, A2 => n13256, B1 => n6617, B2 => 
                           n10942, ZN => n3436);
   U11800 : OAI22_X1 port map( A1 => n13173, A2 => n13259, B1 => n6616, B2 => 
                           n13169, ZN => n3437);
   U11801 : OAI22_X1 port map( A1 => n13173, A2 => n13262, B1 => n6615, B2 => 
                           n13169, ZN => n3438);
   U11802 : OAI22_X1 port map( A1 => n13173, A2 => n13265, B1 => n6614, B2 => 
                           n13169, ZN => n3439);
   U11803 : OAI22_X1 port map( A1 => n13173, A2 => n13268, B1 => n6613, B2 => 
                           n13169, ZN => n3440);
   U11804 : OAI22_X1 port map( A1 => n13173, A2 => n13271, B1 => n6612, B2 => 
                           n13169, ZN => n3441);
   U11805 : OAI22_X1 port map( A1 => n13174, A2 => n13274, B1 => n6611, B2 => 
                           n13169, ZN => n3442);
   U11806 : OAI22_X1 port map( A1 => n13174, A2 => n13277, B1 => n6610, B2 => 
                           n13169, ZN => n3443);
   U11807 : OAI22_X1 port map( A1 => n13174, A2 => n13280, B1 => n6609, B2 => 
                           n13169, ZN => n3444);
   U11808 : OAI22_X1 port map( A1 => n13174, A2 => n13283, B1 => n6608, B2 => 
                           n13169, ZN => n3445);
   U11809 : OAI22_X1 port map( A1 => n13143, A2 => n13214, B1 => n6663, B2 => 
                           n13142, ZN => n3326);
   U11810 : OAI22_X1 port map( A1 => n13143, A2 => n13217, B1 => n6662, B2 => 
                           n13142, ZN => n3327);
   U11811 : OAI22_X1 port map( A1 => n13143, A2 => n13220, B1 => n6661, B2 => 
                           n13142, ZN => n3328);
   U11812 : OAI22_X1 port map( A1 => n13143, A2 => n13223, B1 => n6660, B2 => 
                           n13142, ZN => n3329);
   U11813 : OAI22_X1 port map( A1 => n13143, A2 => n13226, B1 => n6659, B2 => 
                           n13142, ZN => n3330);
   U11814 : OAI22_X1 port map( A1 => n13144, A2 => n13229, B1 => n6658, B2 => 
                           n13142, ZN => n3331);
   U11815 : OAI22_X1 port map( A1 => n13144, A2 => n13232, B1 => n6657, B2 => 
                           n13142, ZN => n3332);
   U11816 : OAI22_X1 port map( A1 => n13144, A2 => n13235, B1 => n6656, B2 => 
                           n13142, ZN => n3333);
   U11817 : OAI22_X1 port map( A1 => n13144, A2 => n13238, B1 => n6655, B2 => 
                           n13142, ZN => n3334);
   U11818 : OAI22_X1 port map( A1 => n13144, A2 => n13241, B1 => n6654, B2 => 
                           n13142, ZN => n3335);
   U11819 : OAI22_X1 port map( A1 => n13145, A2 => n13244, B1 => n6653, B2 => 
                           n13142, ZN => n3336);
   U11820 : OAI22_X1 port map( A1 => n13145, A2 => n13247, B1 => n6652, B2 => 
                           n13142, ZN => n3337);
   U11821 : OAI22_X1 port map( A1 => n13145, A2 => n13250, B1 => n6651, B2 => 
                           n10949, ZN => n3338);
   U11822 : OAI22_X1 port map( A1 => n13145, A2 => n13253, B1 => n6650, B2 => 
                           n10949, ZN => n3339);
   U11823 : OAI22_X1 port map( A1 => n13145, A2 => n13256, B1 => n6649, B2 => 
                           n10949, ZN => n3340);
   U11824 : OAI22_X1 port map( A1 => n13146, A2 => n13259, B1 => n6648, B2 => 
                           n13142, ZN => n3341);
   U11825 : OAI22_X1 port map( A1 => n13146, A2 => n13262, B1 => n6647, B2 => 
                           n13142, ZN => n3342);
   U11826 : OAI22_X1 port map( A1 => n13146, A2 => n13265, B1 => n6646, B2 => 
                           n13142, ZN => n3343);
   U11827 : OAI22_X1 port map( A1 => n13146, A2 => n13268, B1 => n6645, B2 => 
                           n13142, ZN => n3344);
   U11828 : OAI22_X1 port map( A1 => n13146, A2 => n13271, B1 => n6644, B2 => 
                           n13142, ZN => n3345);
   U11829 : OAI22_X1 port map( A1 => n13147, A2 => n13274, B1 => n6643, B2 => 
                           n13142, ZN => n3346);
   U11830 : OAI22_X1 port map( A1 => n13147, A2 => n13277, B1 => n6642, B2 => 
                           n13142, ZN => n3347);
   U11831 : OAI22_X1 port map( A1 => n13147, A2 => n13280, B1 => n6641, B2 => 
                           n13142, ZN => n3348);
   U11832 : OAI22_X1 port map( A1 => n13147, A2 => n13283, B1 => n6640, B2 => 
                           n13142, ZN => n3349);
   U11833 : OAI22_X1 port map( A1 => n13125, A2 => n13214, B1 => n6727, B2 => 
                           n13124, ZN => n3262);
   U11834 : OAI22_X1 port map( A1 => n13125, A2 => n13217, B1 => n6726, B2 => 
                           n13124, ZN => n3263);
   U11835 : OAI22_X1 port map( A1 => n13125, A2 => n13220, B1 => n6725, B2 => 
                           n13124, ZN => n3264);
   U11836 : OAI22_X1 port map( A1 => n13125, A2 => n13223, B1 => n6724, B2 => 
                           n13124, ZN => n3265);
   U11837 : OAI22_X1 port map( A1 => n13125, A2 => n13226, B1 => n6723, B2 => 
                           n13124, ZN => n3266);
   U11838 : OAI22_X1 port map( A1 => n13126, A2 => n13229, B1 => n6722, B2 => 
                           n13124, ZN => n3267);
   U11839 : OAI22_X1 port map( A1 => n13126, A2 => n13232, B1 => n6721, B2 => 
                           n13124, ZN => n3268);
   U11840 : OAI22_X1 port map( A1 => n13126, A2 => n13235, B1 => n6720, B2 => 
                           n13124, ZN => n3269);
   U11841 : OAI22_X1 port map( A1 => n13126, A2 => n13238, B1 => n6719, B2 => 
                           n13124, ZN => n3270);
   U11842 : OAI22_X1 port map( A1 => n13126, A2 => n13241, B1 => n6718, B2 => 
                           n13124, ZN => n3271);
   U11843 : OAI22_X1 port map( A1 => n13127, A2 => n13244, B1 => n6717, B2 => 
                           n13124, ZN => n3272);
   U11844 : OAI22_X1 port map( A1 => n13127, A2 => n13247, B1 => n6716, B2 => 
                           n13124, ZN => n3273);
   U11845 : OAI22_X1 port map( A1 => n13127, A2 => n13250, B1 => n6715, B2 => 
                           n10952, ZN => n3274);
   U11846 : OAI22_X1 port map( A1 => n13127, A2 => n13253, B1 => n6714, B2 => 
                           n10952, ZN => n3275);
   U11847 : OAI22_X1 port map( A1 => n13127, A2 => n13256, B1 => n6713, B2 => 
                           n10952, ZN => n3276);
   U11848 : OAI22_X1 port map( A1 => n13128, A2 => n13259, B1 => n6712, B2 => 
                           n13124, ZN => n3277);
   U11849 : OAI22_X1 port map( A1 => n13128, A2 => n13262, B1 => n6711, B2 => 
                           n13124, ZN => n3278);
   U11850 : OAI22_X1 port map( A1 => n13128, A2 => n13265, B1 => n6710, B2 => 
                           n13124, ZN => n3279);
   U11851 : OAI22_X1 port map( A1 => n13128, A2 => n13268, B1 => n6709, B2 => 
                           n13124, ZN => n3280);
   U11852 : OAI22_X1 port map( A1 => n13128, A2 => n13271, B1 => n6708, B2 => 
                           n13124, ZN => n3281);
   U11853 : OAI22_X1 port map( A1 => n13129, A2 => n13274, B1 => n6707, B2 => 
                           n13124, ZN => n3282);
   U11854 : OAI22_X1 port map( A1 => n13129, A2 => n13277, B1 => n6706, B2 => 
                           n13124, ZN => n3283);
   U11855 : OAI22_X1 port map( A1 => n13129, A2 => n13280, B1 => n6705, B2 => 
                           n13124, ZN => n3284);
   U11856 : OAI22_X1 port map( A1 => n13129, A2 => n13283, B1 => n6704, B2 => 
                           n13124, ZN => n3285);
   U11857 : OAI22_X1 port map( A1 => n13134, A2 => n13214, B1 => n6695, B2 => 
                           n13133, ZN => n3294);
   U11858 : OAI22_X1 port map( A1 => n13134, A2 => n13217, B1 => n6694, B2 => 
                           n13133, ZN => n3295);
   U11859 : OAI22_X1 port map( A1 => n13134, A2 => n13220, B1 => n6693, B2 => 
                           n13133, ZN => n3296);
   U11860 : OAI22_X1 port map( A1 => n13134, A2 => n13223, B1 => n6692, B2 => 
                           n13133, ZN => n3297);
   U11861 : OAI22_X1 port map( A1 => n13134, A2 => n13226, B1 => n6691, B2 => 
                           n13133, ZN => n3298);
   U11862 : OAI22_X1 port map( A1 => n13135, A2 => n13229, B1 => n6690, B2 => 
                           n13133, ZN => n3299);
   U11863 : OAI22_X1 port map( A1 => n13135, A2 => n13232, B1 => n6689, B2 => 
                           n13133, ZN => n3300);
   U11864 : OAI22_X1 port map( A1 => n13135, A2 => n13235, B1 => n6688, B2 => 
                           n13133, ZN => n3301);
   U11865 : OAI22_X1 port map( A1 => n13135, A2 => n13238, B1 => n6687, B2 => 
                           n13133, ZN => n3302);
   U11866 : OAI22_X1 port map( A1 => n13135, A2 => n13241, B1 => n6686, B2 => 
                           n13133, ZN => n3303);
   U11867 : OAI22_X1 port map( A1 => n13136, A2 => n13244, B1 => n6685, B2 => 
                           n13133, ZN => n3304);
   U11868 : OAI22_X1 port map( A1 => n13136, A2 => n13247, B1 => n6684, B2 => 
                           n13133, ZN => n3305);
   U11869 : OAI22_X1 port map( A1 => n13136, A2 => n13250, B1 => n6683, B2 => 
                           n10951, ZN => n3306);
   U11870 : OAI22_X1 port map( A1 => n13136, A2 => n13253, B1 => n6682, B2 => 
                           n10951, ZN => n3307);
   U11871 : OAI22_X1 port map( A1 => n13136, A2 => n13256, B1 => n6681, B2 => 
                           n10951, ZN => n3308);
   U11872 : OAI22_X1 port map( A1 => n13137, A2 => n13259, B1 => n6680, B2 => 
                           n13133, ZN => n3309);
   U11873 : OAI22_X1 port map( A1 => n13137, A2 => n13262, B1 => n6679, B2 => 
                           n13133, ZN => n3310);
   U11874 : OAI22_X1 port map( A1 => n13137, A2 => n13265, B1 => n6678, B2 => 
                           n13133, ZN => n3311);
   U11875 : OAI22_X1 port map( A1 => n13137, A2 => n13268, B1 => n6677, B2 => 
                           n13133, ZN => n3312);
   U11876 : OAI22_X1 port map( A1 => n13137, A2 => n13271, B1 => n6676, B2 => 
                           n13133, ZN => n3313);
   U11877 : OAI22_X1 port map( A1 => n13138, A2 => n13274, B1 => n6675, B2 => 
                           n13133, ZN => n3314);
   U11878 : OAI22_X1 port map( A1 => n13138, A2 => n13277, B1 => n6674, B2 => 
                           n13133, ZN => n3315);
   U11879 : OAI22_X1 port map( A1 => n13138, A2 => n13280, B1 => n6673, B2 => 
                           n13133, ZN => n3316);
   U11880 : OAI22_X1 port map( A1 => n13138, A2 => n13283, B1 => n6672, B2 => 
                           n13133, ZN => n3317);
   U11881 : OAI22_X1 port map( A1 => n13116, A2 => n13214, B1 => n6759, B2 => 
                           n13115, ZN => n3230);
   U11882 : OAI22_X1 port map( A1 => n13116, A2 => n13217, B1 => n6758, B2 => 
                           n13115, ZN => n3231);
   U11883 : OAI22_X1 port map( A1 => n13116, A2 => n13220, B1 => n6757, B2 => 
                           n13115, ZN => n3232);
   U11884 : OAI22_X1 port map( A1 => n13116, A2 => n13223, B1 => n6756, B2 => 
                           n13115, ZN => n3233);
   U11885 : OAI22_X1 port map( A1 => n13116, A2 => n13226, B1 => n6755, B2 => 
                           n13115, ZN => n3234);
   U11886 : OAI22_X1 port map( A1 => n13117, A2 => n13229, B1 => n6754, B2 => 
                           n13115, ZN => n3235);
   U11887 : OAI22_X1 port map( A1 => n13117, A2 => n13232, B1 => n6753, B2 => 
                           n13115, ZN => n3236);
   U11888 : OAI22_X1 port map( A1 => n13117, A2 => n13235, B1 => n6752, B2 => 
                           n13115, ZN => n3237);
   U11889 : OAI22_X1 port map( A1 => n13117, A2 => n13238, B1 => n6751, B2 => 
                           n13115, ZN => n3238);
   U11890 : OAI22_X1 port map( A1 => n13117, A2 => n13241, B1 => n6750, B2 => 
                           n13115, ZN => n3239);
   U11891 : OAI22_X1 port map( A1 => n13118, A2 => n13244, B1 => n6749, B2 => 
                           n13115, ZN => n3240);
   U11892 : OAI22_X1 port map( A1 => n13118, A2 => n13247, B1 => n6748, B2 => 
                           n13115, ZN => n3241);
   U11893 : OAI22_X1 port map( A1 => n13118, A2 => n13250, B1 => n6747, B2 => 
                           n10953, ZN => n3242);
   U11894 : OAI22_X1 port map( A1 => n13118, A2 => n13253, B1 => n6746, B2 => 
                           n10953, ZN => n3243);
   U11895 : OAI22_X1 port map( A1 => n13118, A2 => n13256, B1 => n6745, B2 => 
                           n10953, ZN => n3244);
   U11896 : OAI22_X1 port map( A1 => n13119, A2 => n13259, B1 => n6744, B2 => 
                           n13115, ZN => n3245);
   U11897 : OAI22_X1 port map( A1 => n13119, A2 => n13262, B1 => n6743, B2 => 
                           n13115, ZN => n3246);
   U11898 : OAI22_X1 port map( A1 => n13119, A2 => n13265, B1 => n6742, B2 => 
                           n13115, ZN => n3247);
   U11899 : OAI22_X1 port map( A1 => n13119, A2 => n13268, B1 => n6741, B2 => 
                           n13115, ZN => n3248);
   U11900 : OAI22_X1 port map( A1 => n13119, A2 => n13271, B1 => n6740, B2 => 
                           n13115, ZN => n3249);
   U11901 : OAI22_X1 port map( A1 => n13120, A2 => n13274, B1 => n6739, B2 => 
                           n13115, ZN => n3250);
   U11902 : OAI22_X1 port map( A1 => n13120, A2 => n13277, B1 => n6738, B2 => 
                           n13115, ZN => n3251);
   U11903 : OAI22_X1 port map( A1 => n13120, A2 => n13280, B1 => n6737, B2 => 
                           n13115, ZN => n3252);
   U11904 : OAI22_X1 port map( A1 => n13120, A2 => n13283, B1 => n6736, B2 => 
                           n13115, ZN => n3253);
   U11905 : OAI22_X1 port map( A1 => n13197, A2 => n13214, B1 => n9281, B2 => 
                           n13196, ZN => n3518);
   U11906 : OAI22_X1 port map( A1 => n13197, A2 => n13217, B1 => n9266, B2 => 
                           n13196, ZN => n3519);
   U11907 : OAI22_X1 port map( A1 => n13197, A2 => n13220, B1 => n9251, B2 => 
                           n13196, ZN => n3520);
   U11908 : OAI22_X1 port map( A1 => n13197, A2 => n13223, B1 => n9236, B2 => 
                           n13196, ZN => n3521);
   U11909 : OAI22_X1 port map( A1 => n13197, A2 => n13226, B1 => n9221, B2 => 
                           n13196, ZN => n3522);
   U11910 : OAI22_X1 port map( A1 => n13198, A2 => n13229, B1 => n9206, B2 => 
                           n13196, ZN => n3523);
   U11911 : OAI22_X1 port map( A1 => n13198, A2 => n13232, B1 => n9191, B2 => 
                           n13196, ZN => n3524);
   U11912 : OAI22_X1 port map( A1 => n13198, A2 => n13235, B1 => n9176, B2 => 
                           n13196, ZN => n3525);
   U11913 : OAI22_X1 port map( A1 => n13198, A2 => n13238, B1 => n9161, B2 => 
                           n13196, ZN => n3526);
   U11914 : OAI22_X1 port map( A1 => n13198, A2 => n13241, B1 => n9146, B2 => 
                           n13196, ZN => n3527);
   U11915 : OAI22_X1 port map( A1 => n13199, A2 => n13244, B1 => n9131, B2 => 
                           n13196, ZN => n3528);
   U11916 : OAI22_X1 port map( A1 => n13199, A2 => n13247, B1 => n9116, B2 => 
                           n13196, ZN => n3529);
   U11917 : OAI22_X1 port map( A1 => n13199, A2 => n13250, B1 => n9101, B2 => 
                           n10936, ZN => n3530);
   U11918 : OAI22_X1 port map( A1 => n13199, A2 => n13253, B1 => n9086, B2 => 
                           n10936, ZN => n3531);
   U11919 : OAI22_X1 port map( A1 => n13199, A2 => n13256, B1 => n9071, B2 => 
                           n10936, ZN => n3532);
   U11920 : OAI22_X1 port map( A1 => n13200, A2 => n13259, B1 => n9056, B2 => 
                           n13196, ZN => n3533);
   U11921 : OAI22_X1 port map( A1 => n13200, A2 => n13262, B1 => n9041, B2 => 
                           n13196, ZN => n3534);
   U11922 : OAI22_X1 port map( A1 => n13200, A2 => n13265, B1 => n9026, B2 => 
                           n13196, ZN => n3535);
   U11923 : OAI22_X1 port map( A1 => n13200, A2 => n13268, B1 => n9011, B2 => 
                           n13196, ZN => n3536);
   U11924 : OAI22_X1 port map( A1 => n13200, A2 => n13271, B1 => n8996, B2 => 
                           n13196, ZN => n3537);
   U11925 : OAI22_X1 port map( A1 => n13201, A2 => n13274, B1 => n8981, B2 => 
                           n13196, ZN => n3538);
   U11926 : OAI22_X1 port map( A1 => n13201, A2 => n13277, B1 => n8966, B2 => 
                           n13196, ZN => n3539);
   U11927 : OAI22_X1 port map( A1 => n13201, A2 => n13280, B1 => n8951, B2 => 
                           n13196, ZN => n3540);
   U11928 : OAI22_X1 port map( A1 => n13201, A2 => n13283, B1 => n8936, B2 => 
                           n13196, ZN => n3541);
   U11929 : OAI22_X1 port map( A1 => n13188, A2 => n13214, B1 => n9282, B2 => 
                           n13187, ZN => n3486);
   U11930 : OAI22_X1 port map( A1 => n13188, A2 => n13217, B1 => n9267, B2 => 
                           n13187, ZN => n3487);
   U11931 : OAI22_X1 port map( A1 => n13188, A2 => n13220, B1 => n9252, B2 => 
                           n13187, ZN => n3488);
   U11932 : OAI22_X1 port map( A1 => n13188, A2 => n13223, B1 => n9237, B2 => 
                           n13187, ZN => n3489);
   U11933 : OAI22_X1 port map( A1 => n13188, A2 => n13226, B1 => n9222, B2 => 
                           n13187, ZN => n3490);
   U11934 : OAI22_X1 port map( A1 => n13189, A2 => n13229, B1 => n9207, B2 => 
                           n13187, ZN => n3491);
   U11935 : OAI22_X1 port map( A1 => n13189, A2 => n13232, B1 => n9192, B2 => 
                           n13187, ZN => n3492);
   U11936 : OAI22_X1 port map( A1 => n13189, A2 => n13235, B1 => n9177, B2 => 
                           n13187, ZN => n3493);
   U11937 : OAI22_X1 port map( A1 => n13189, A2 => n13238, B1 => n9162, B2 => 
                           n13187, ZN => n3494);
   U11938 : OAI22_X1 port map( A1 => n13189, A2 => n13241, B1 => n9147, B2 => 
                           n13187, ZN => n3495);
   U11939 : OAI22_X1 port map( A1 => n13190, A2 => n13244, B1 => n9132, B2 => 
                           n13187, ZN => n3496);
   U11940 : OAI22_X1 port map( A1 => n13190, A2 => n13247, B1 => n9117, B2 => 
                           n13187, ZN => n3497);
   U11941 : OAI22_X1 port map( A1 => n13190, A2 => n13250, B1 => n9102, B2 => 
                           n10938, ZN => n3498);
   U11942 : OAI22_X1 port map( A1 => n13190, A2 => n13253, B1 => n9087, B2 => 
                           n10938, ZN => n3499);
   U11943 : OAI22_X1 port map( A1 => n13190, A2 => n13256, B1 => n9072, B2 => 
                           n10938, ZN => n3500);
   U11944 : OAI22_X1 port map( A1 => n13191, A2 => n13259, B1 => n9057, B2 => 
                           n13187, ZN => n3501);
   U11945 : OAI22_X1 port map( A1 => n13191, A2 => n13262, B1 => n9042, B2 => 
                           n13187, ZN => n3502);
   U11946 : OAI22_X1 port map( A1 => n13191, A2 => n13265, B1 => n9027, B2 => 
                           n13187, ZN => n3503);
   U11947 : OAI22_X1 port map( A1 => n13191, A2 => n13268, B1 => n9012, B2 => 
                           n13187, ZN => n3504);
   U11948 : OAI22_X1 port map( A1 => n13191, A2 => n13271, B1 => n8997, B2 => 
                           n13187, ZN => n3505);
   U11949 : OAI22_X1 port map( A1 => n13192, A2 => n13274, B1 => n8982, B2 => 
                           n13187, ZN => n3506);
   U11950 : OAI22_X1 port map( A1 => n13192, A2 => n13277, B1 => n8967, B2 => 
                           n13187, ZN => n3507);
   U11951 : OAI22_X1 port map( A1 => n13192, A2 => n13280, B1 => n8952, B2 => 
                           n13187, ZN => n3508);
   U11952 : OAI22_X1 port map( A1 => n13192, A2 => n13283, B1 => n8937, B2 => 
                           n13187, ZN => n3509);
   U11953 : OAI22_X1 port map( A1 => n13107, A2 => n13215, B1 => n9286, B2 => 
                           n13106, ZN => n3198);
   U11954 : OAI22_X1 port map( A1 => n13107, A2 => n13218, B1 => n9271, B2 => 
                           n13106, ZN => n3199);
   U11955 : OAI22_X1 port map( A1 => n13107, A2 => n13221, B1 => n9256, B2 => 
                           n13106, ZN => n3200);
   U11956 : OAI22_X1 port map( A1 => n13107, A2 => n13224, B1 => n9241, B2 => 
                           n13106, ZN => n3201);
   U11957 : OAI22_X1 port map( A1 => n13107, A2 => n13227, B1 => n9226, B2 => 
                           n13106, ZN => n3202);
   U11958 : OAI22_X1 port map( A1 => n13108, A2 => n13230, B1 => n9211, B2 => 
                           n13106, ZN => n3203);
   U11959 : OAI22_X1 port map( A1 => n13108, A2 => n13233, B1 => n9196, B2 => 
                           n13106, ZN => n3204);
   U11960 : OAI22_X1 port map( A1 => n13108, A2 => n13236, B1 => n9181, B2 => 
                           n13106, ZN => n3205);
   U11961 : OAI22_X1 port map( A1 => n13108, A2 => n13239, B1 => n9166, B2 => 
                           n13106, ZN => n3206);
   U11962 : OAI22_X1 port map( A1 => n13108, A2 => n13242, B1 => n9151, B2 => 
                           n13106, ZN => n3207);
   U11963 : OAI22_X1 port map( A1 => n13109, A2 => n13245, B1 => n9136, B2 => 
                           n13106, ZN => n3208);
   U11964 : OAI22_X1 port map( A1 => n13109, A2 => n13248, B1 => n9121, B2 => 
                           n13106, ZN => n3209);
   U11965 : OAI22_X1 port map( A1 => n13109, A2 => n13251, B1 => n9106, B2 => 
                           n10954, ZN => n3210);
   U11966 : OAI22_X1 port map( A1 => n13109, A2 => n13254, B1 => n9091, B2 => 
                           n10954, ZN => n3211);
   U11967 : OAI22_X1 port map( A1 => n13109, A2 => n13257, B1 => n9076, B2 => 
                           n10954, ZN => n3212);
   U11968 : OAI22_X1 port map( A1 => n13110, A2 => n13260, B1 => n9061, B2 => 
                           n13106, ZN => n3213);
   U11969 : OAI22_X1 port map( A1 => n13110, A2 => n13263, B1 => n9046, B2 => 
                           n13106, ZN => n3214);
   U11970 : OAI22_X1 port map( A1 => n13110, A2 => n13266, B1 => n9031, B2 => 
                           n13106, ZN => n3215);
   U11971 : OAI22_X1 port map( A1 => n13110, A2 => n13269, B1 => n9016, B2 => 
                           n13106, ZN => n3216);
   U11972 : OAI22_X1 port map( A1 => n13110, A2 => n13272, B1 => n9001, B2 => 
                           n13106, ZN => n3217);
   U11973 : OAI22_X1 port map( A1 => n13111, A2 => n13275, B1 => n8986, B2 => 
                           n13106, ZN => n3218);
   U11974 : OAI22_X1 port map( A1 => n13111, A2 => n13278, B1 => n8971, B2 => 
                           n13106, ZN => n3219);
   U11975 : OAI22_X1 port map( A1 => n13111, A2 => n13281, B1 => n8956, B2 => 
                           n13106, ZN => n3220);
   U11976 : OAI22_X1 port map( A1 => n13111, A2 => n13284, B1 => n8941, B2 => 
                           n13106, ZN => n3221);
   U11977 : OAI22_X1 port map( A1 => n13098, A2 => n13215, B1 => n9285, B2 => 
                           n13097, ZN => n3166);
   U11978 : OAI22_X1 port map( A1 => n13098, A2 => n13218, B1 => n9270, B2 => 
                           n13097, ZN => n3167);
   U11979 : OAI22_X1 port map( A1 => n13098, A2 => n13221, B1 => n9255, B2 => 
                           n13097, ZN => n3168);
   U11980 : OAI22_X1 port map( A1 => n13098, A2 => n13224, B1 => n9240, B2 => 
                           n13097, ZN => n3169);
   U11981 : OAI22_X1 port map( A1 => n13098, A2 => n13227, B1 => n9225, B2 => 
                           n13097, ZN => n3170);
   U11982 : OAI22_X1 port map( A1 => n13099, A2 => n13230, B1 => n9210, B2 => 
                           n13097, ZN => n3171);
   U11983 : OAI22_X1 port map( A1 => n13099, A2 => n13233, B1 => n9195, B2 => 
                           n13097, ZN => n3172);
   U11984 : OAI22_X1 port map( A1 => n13099, A2 => n13236, B1 => n9180, B2 => 
                           n13097, ZN => n3173);
   U11985 : OAI22_X1 port map( A1 => n13099, A2 => n13239, B1 => n9165, B2 => 
                           n13097, ZN => n3174);
   U11986 : OAI22_X1 port map( A1 => n13099, A2 => n13242, B1 => n9150, B2 => 
                           n13097, ZN => n3175);
   U11987 : OAI22_X1 port map( A1 => n13100, A2 => n13245, B1 => n9135, B2 => 
                           n13097, ZN => n3176);
   U11988 : OAI22_X1 port map( A1 => n13100, A2 => n13248, B1 => n9120, B2 => 
                           n13097, ZN => n3177);
   U11989 : OAI22_X1 port map( A1 => n13100, A2 => n13251, B1 => n9105, B2 => 
                           n10955, ZN => n3178);
   U11990 : OAI22_X1 port map( A1 => n13100, A2 => n13254, B1 => n9090, B2 => 
                           n10955, ZN => n3179);
   U11991 : OAI22_X1 port map( A1 => n13100, A2 => n13257, B1 => n9075, B2 => 
                           n10955, ZN => n3180);
   U11992 : OAI22_X1 port map( A1 => n13101, A2 => n13260, B1 => n9060, B2 => 
                           n13097, ZN => n3181);
   U11993 : OAI22_X1 port map( A1 => n13101, A2 => n13263, B1 => n9045, B2 => 
                           n13097, ZN => n3182);
   U11994 : OAI22_X1 port map( A1 => n13101, A2 => n13266, B1 => n9030, B2 => 
                           n13097, ZN => n3183);
   U11995 : OAI22_X1 port map( A1 => n13101, A2 => n13269, B1 => n9015, B2 => 
                           n13097, ZN => n3184);
   U11996 : OAI22_X1 port map( A1 => n13101, A2 => n13272, B1 => n9000, B2 => 
                           n13097, ZN => n3185);
   U11997 : OAI22_X1 port map( A1 => n13102, A2 => n13275, B1 => n8985, B2 => 
                           n13097, ZN => n3186);
   U11998 : OAI22_X1 port map( A1 => n13102, A2 => n13278, B1 => n8970, B2 => 
                           n13097, ZN => n3187);
   U11999 : OAI22_X1 port map( A1 => n13102, A2 => n13281, B1 => n8955, B2 => 
                           n13097, ZN => n3188);
   U12000 : OAI22_X1 port map( A1 => n13102, A2 => n13284, B1 => n8940, B2 => 
                           n13097, ZN => n3189);
   U12001 : OAI22_X1 port map( A1 => n13071, A2 => n13215, B1 => n9288, B2 => 
                           n13070, ZN => n3070);
   U12002 : OAI22_X1 port map( A1 => n13071, A2 => n13218, B1 => n9273, B2 => 
                           n13070, ZN => n3071);
   U12003 : OAI22_X1 port map( A1 => n13071, A2 => n13221, B1 => n9258, B2 => 
                           n13070, ZN => n3072);
   U12004 : OAI22_X1 port map( A1 => n13071, A2 => n13224, B1 => n9243, B2 => 
                           n13070, ZN => n3073);
   U12005 : OAI22_X1 port map( A1 => n13071, A2 => n13227, B1 => n9228, B2 => 
                           n13070, ZN => n3074);
   U12006 : OAI22_X1 port map( A1 => n13072, A2 => n13230, B1 => n9213, B2 => 
                           n13070, ZN => n3075);
   U12007 : OAI22_X1 port map( A1 => n13072, A2 => n13233, B1 => n9198, B2 => 
                           n13070, ZN => n3076);
   U12008 : OAI22_X1 port map( A1 => n13072, A2 => n13236, B1 => n9183, B2 => 
                           n13070, ZN => n3077);
   U12009 : OAI22_X1 port map( A1 => n13072, A2 => n13239, B1 => n9168, B2 => 
                           n13070, ZN => n3078);
   U12010 : OAI22_X1 port map( A1 => n13072, A2 => n13242, B1 => n9153, B2 => 
                           n13070, ZN => n3079);
   U12011 : OAI22_X1 port map( A1 => n13073, A2 => n13245, B1 => n9138, B2 => 
                           n13070, ZN => n3080);
   U12012 : OAI22_X1 port map( A1 => n13073, A2 => n13248, B1 => n9123, B2 => 
                           n13070, ZN => n3081);
   U12013 : OAI22_X1 port map( A1 => n13073, A2 => n13251, B1 => n9108, B2 => 
                           n10958, ZN => n3082);
   U12014 : OAI22_X1 port map( A1 => n13073, A2 => n13254, B1 => n9093, B2 => 
                           n10958, ZN => n3083);
   U12015 : OAI22_X1 port map( A1 => n13073, A2 => n13257, B1 => n9078, B2 => 
                           n10958, ZN => n3084);
   U12016 : OAI22_X1 port map( A1 => n13074, A2 => n13260, B1 => n9063, B2 => 
                           n13070, ZN => n3085);
   U12017 : OAI22_X1 port map( A1 => n13074, A2 => n13263, B1 => n9048, B2 => 
                           n13070, ZN => n3086);
   U12018 : OAI22_X1 port map( A1 => n13074, A2 => n13266, B1 => n9033, B2 => 
                           n13070, ZN => n3087);
   U12019 : OAI22_X1 port map( A1 => n13074, A2 => n13269, B1 => n9018, B2 => 
                           n13070, ZN => n3088);
   U12020 : OAI22_X1 port map( A1 => n13074, A2 => n13272, B1 => n9003, B2 => 
                           n13070, ZN => n3089);
   U12021 : OAI22_X1 port map( A1 => n13075, A2 => n13275, B1 => n8988, B2 => 
                           n13070, ZN => n3090);
   U12022 : OAI22_X1 port map( A1 => n13075, A2 => n13278, B1 => n8973, B2 => 
                           n13070, ZN => n3091);
   U12023 : OAI22_X1 port map( A1 => n13075, A2 => n13281, B1 => n8958, B2 => 
                           n13070, ZN => n3092);
   U12024 : OAI22_X1 port map( A1 => n13075, A2 => n13284, B1 => n8943, B2 => 
                           n13070, ZN => n3093);
   U12025 : OAI22_X1 port map( A1 => n13062, A2 => n13215, B1 => n9287, B2 => 
                           n13061, ZN => n3038);
   U12026 : OAI22_X1 port map( A1 => n13062, A2 => n13218, B1 => n9272, B2 => 
                           n13061, ZN => n3039);
   U12027 : OAI22_X1 port map( A1 => n13062, A2 => n13221, B1 => n9257, B2 => 
                           n13061, ZN => n3040);
   U12028 : OAI22_X1 port map( A1 => n13062, A2 => n13224, B1 => n9242, B2 => 
                           n13061, ZN => n3041);
   U12029 : OAI22_X1 port map( A1 => n13062, A2 => n13227, B1 => n9227, B2 => 
                           n13061, ZN => n3042);
   U12030 : OAI22_X1 port map( A1 => n13063, A2 => n13230, B1 => n9212, B2 => 
                           n13061, ZN => n3043);
   U12031 : OAI22_X1 port map( A1 => n13063, A2 => n13233, B1 => n9197, B2 => 
                           n13061, ZN => n3044);
   U12032 : OAI22_X1 port map( A1 => n13063, A2 => n13236, B1 => n9182, B2 => 
                           n13061, ZN => n3045);
   U12033 : OAI22_X1 port map( A1 => n13063, A2 => n13239, B1 => n9167, B2 => 
                           n13061, ZN => n3046);
   U12034 : OAI22_X1 port map( A1 => n13063, A2 => n13242, B1 => n9152, B2 => 
                           n13061, ZN => n3047);
   U12035 : OAI22_X1 port map( A1 => n13064, A2 => n13245, B1 => n9137, B2 => 
                           n13061, ZN => n3048);
   U12036 : OAI22_X1 port map( A1 => n13064, A2 => n13248, B1 => n9122, B2 => 
                           n13061, ZN => n3049);
   U12037 : OAI22_X1 port map( A1 => n13064, A2 => n13251, B1 => n9107, B2 => 
                           n10960, ZN => n3050);
   U12038 : OAI22_X1 port map( A1 => n13064, A2 => n13254, B1 => n9092, B2 => 
                           n10960, ZN => n3051);
   U12039 : OAI22_X1 port map( A1 => n13064, A2 => n13257, B1 => n9077, B2 => 
                           n10960, ZN => n3052);
   U12040 : OAI22_X1 port map( A1 => n13065, A2 => n13260, B1 => n9062, B2 => 
                           n13061, ZN => n3053);
   U12041 : OAI22_X1 port map( A1 => n13065, A2 => n13263, B1 => n9047, B2 => 
                           n13061, ZN => n3054);
   U12042 : OAI22_X1 port map( A1 => n13065, A2 => n13266, B1 => n9032, B2 => 
                           n13061, ZN => n3055);
   U12043 : OAI22_X1 port map( A1 => n13065, A2 => n13269, B1 => n9017, B2 => 
                           n13061, ZN => n3056);
   U12044 : OAI22_X1 port map( A1 => n13065, A2 => n13272, B1 => n9002, B2 => 
                           n13061, ZN => n3057);
   U12045 : OAI22_X1 port map( A1 => n13066, A2 => n13275, B1 => n8987, B2 => 
                           n13061, ZN => n3058);
   U12046 : OAI22_X1 port map( A1 => n13066, A2 => n13278, B1 => n8972, B2 => 
                           n13061, ZN => n3059);
   U12047 : OAI22_X1 port map( A1 => n13066, A2 => n13281, B1 => n8957, B2 => 
                           n13061, ZN => n3060);
   U12048 : OAI22_X1 port map( A1 => n13066, A2 => n13284, B1 => n8942, B2 => 
                           n13061, ZN => n3061);
   U12049 : OAI22_X1 port map( A1 => n13035, A2 => n13215, B1 => n9290, B2 => 
                           n13034, ZN => n2942);
   U12050 : OAI22_X1 port map( A1 => n13035, A2 => n13218, B1 => n9275, B2 => 
                           n13034, ZN => n2943);
   U12051 : OAI22_X1 port map( A1 => n13035, A2 => n13221, B1 => n9260, B2 => 
                           n13034, ZN => n2944);
   U12052 : OAI22_X1 port map( A1 => n13035, A2 => n13224, B1 => n9245, B2 => 
                           n13034, ZN => n2945);
   U12053 : OAI22_X1 port map( A1 => n13035, A2 => n13227, B1 => n9230, B2 => 
                           n13034, ZN => n2946);
   U12054 : OAI22_X1 port map( A1 => n13036, A2 => n13230, B1 => n9215, B2 => 
                           n13034, ZN => n2947);
   U12055 : OAI22_X1 port map( A1 => n13036, A2 => n13233, B1 => n9200, B2 => 
                           n13034, ZN => n2948);
   U12056 : OAI22_X1 port map( A1 => n13036, A2 => n13236, B1 => n9185, B2 => 
                           n13034, ZN => n2949);
   U12057 : OAI22_X1 port map( A1 => n13036, A2 => n13239, B1 => n9170, B2 => 
                           n13034, ZN => n2950);
   U12058 : OAI22_X1 port map( A1 => n13036, A2 => n13242, B1 => n9155, B2 => 
                           n13034, ZN => n2951);
   U12059 : OAI22_X1 port map( A1 => n13037, A2 => n13245, B1 => n9140, B2 => 
                           n13034, ZN => n2952);
   U12060 : OAI22_X1 port map( A1 => n13037, A2 => n13248, B1 => n9125, B2 => 
                           n13034, ZN => n2953);
   U12061 : OAI22_X1 port map( A1 => n13037, A2 => n13251, B1 => n9110, B2 => 
                           n10963, ZN => n2954);
   U12062 : OAI22_X1 port map( A1 => n13037, A2 => n13254, B1 => n9095, B2 => 
                           n10963, ZN => n2955);
   U12063 : OAI22_X1 port map( A1 => n13037, A2 => n13257, B1 => n9080, B2 => 
                           n10963, ZN => n2956);
   U12064 : OAI22_X1 port map( A1 => n13038, A2 => n13260, B1 => n9065, B2 => 
                           n13034, ZN => n2957);
   U12065 : OAI22_X1 port map( A1 => n13038, A2 => n13263, B1 => n9050, B2 => 
                           n13034, ZN => n2958);
   U12066 : OAI22_X1 port map( A1 => n13038, A2 => n13266, B1 => n9035, B2 => 
                           n13034, ZN => n2959);
   U12067 : OAI22_X1 port map( A1 => n13038, A2 => n13269, B1 => n9020, B2 => 
                           n13034, ZN => n2960);
   U12068 : OAI22_X1 port map( A1 => n13038, A2 => n13272, B1 => n9005, B2 => 
                           n13034, ZN => n2961);
   U12069 : OAI22_X1 port map( A1 => n13039, A2 => n13275, B1 => n8990, B2 => 
                           n13034, ZN => n2962);
   U12070 : OAI22_X1 port map( A1 => n13039, A2 => n13278, B1 => n8975, B2 => 
                           n13034, ZN => n2963);
   U12071 : OAI22_X1 port map( A1 => n13039, A2 => n13281, B1 => n8960, B2 => 
                           n13034, ZN => n2964);
   U12072 : OAI22_X1 port map( A1 => n13039, A2 => n13284, B1 => n8945, B2 => 
                           n13034, ZN => n2965);
   U12073 : OAI22_X1 port map( A1 => n13026, A2 => n13215, B1 => n9289, B2 => 
                           n13025, ZN => n2910);
   U12074 : OAI22_X1 port map( A1 => n13026, A2 => n13218, B1 => n9274, B2 => 
                           n13025, ZN => n2911);
   U12075 : OAI22_X1 port map( A1 => n13026, A2 => n13221, B1 => n9259, B2 => 
                           n13025, ZN => n2912);
   U12076 : OAI22_X1 port map( A1 => n13026, A2 => n13224, B1 => n9244, B2 => 
                           n13025, ZN => n2913);
   U12077 : OAI22_X1 port map( A1 => n13026, A2 => n13227, B1 => n9229, B2 => 
                           n13025, ZN => n2914);
   U12078 : OAI22_X1 port map( A1 => n13027, A2 => n13230, B1 => n9214, B2 => 
                           n13025, ZN => n2915);
   U12079 : OAI22_X1 port map( A1 => n13027, A2 => n13233, B1 => n9199, B2 => 
                           n13025, ZN => n2916);
   U12080 : OAI22_X1 port map( A1 => n13027, A2 => n13236, B1 => n9184, B2 => 
                           n13025, ZN => n2917);
   U12081 : OAI22_X1 port map( A1 => n13027, A2 => n13239, B1 => n9169, B2 => 
                           n13025, ZN => n2918);
   U12082 : OAI22_X1 port map( A1 => n13027, A2 => n13242, B1 => n9154, B2 => 
                           n13025, ZN => n2919);
   U12083 : OAI22_X1 port map( A1 => n13028, A2 => n13245, B1 => n9139, B2 => 
                           n13025, ZN => n2920);
   U12084 : OAI22_X1 port map( A1 => n13028, A2 => n13248, B1 => n9124, B2 => 
                           n13025, ZN => n2921);
   U12085 : OAI22_X1 port map( A1 => n13028, A2 => n13251, B1 => n9109, B2 => 
                           n10964, ZN => n2922);
   U12086 : OAI22_X1 port map( A1 => n13028, A2 => n13254, B1 => n9094, B2 => 
                           n10964, ZN => n2923);
   U12087 : OAI22_X1 port map( A1 => n13028, A2 => n13257, B1 => n9079, B2 => 
                           n10964, ZN => n2924);
   U12088 : OAI22_X1 port map( A1 => n13029, A2 => n13260, B1 => n9064, B2 => 
                           n13025, ZN => n2925);
   U12089 : OAI22_X1 port map( A1 => n13029, A2 => n13263, B1 => n9049, B2 => 
                           n13025, ZN => n2926);
   U12090 : OAI22_X1 port map( A1 => n13029, A2 => n13266, B1 => n9034, B2 => 
                           n13025, ZN => n2927);
   U12091 : OAI22_X1 port map( A1 => n13029, A2 => n13269, B1 => n9019, B2 => 
                           n13025, ZN => n2928);
   U12092 : OAI22_X1 port map( A1 => n13029, A2 => n13272, B1 => n9004, B2 => 
                           n13025, ZN => n2929);
   U12093 : OAI22_X1 port map( A1 => n13030, A2 => n13275, B1 => n8989, B2 => 
                           n13025, ZN => n2930);
   U12094 : OAI22_X1 port map( A1 => n13030, A2 => n13278, B1 => n8974, B2 => 
                           n13025, ZN => n2931);
   U12095 : OAI22_X1 port map( A1 => n13030, A2 => n13281, B1 => n8959, B2 => 
                           n13025, ZN => n2932);
   U12096 : OAI22_X1 port map( A1 => n13030, A2 => n13284, B1 => n8944, B2 => 
                           n13025, ZN => n2933);
   U12097 : OAI22_X1 port map( A1 => n12981, A2 => n13216, B1 => n9292, B2 => 
                           n12980, ZN => n2750);
   U12098 : OAI22_X1 port map( A1 => n12981, A2 => n13219, B1 => n9277, B2 => 
                           n12980, ZN => n2751);
   U12099 : OAI22_X1 port map( A1 => n12981, A2 => n13222, B1 => n9262, B2 => 
                           n12980, ZN => n2752);
   U12100 : OAI22_X1 port map( A1 => n12981, A2 => n13225, B1 => n9247, B2 => 
                           n12980, ZN => n2753);
   U12101 : OAI22_X1 port map( A1 => n12981, A2 => n13228, B1 => n9232, B2 => 
                           n12980, ZN => n2754);
   U12102 : OAI22_X1 port map( A1 => n12982, A2 => n13231, B1 => n9217, B2 => 
                           n12980, ZN => n2755);
   U12103 : OAI22_X1 port map( A1 => n12982, A2 => n13234, B1 => n9202, B2 => 
                           n12980, ZN => n2756);
   U12104 : OAI22_X1 port map( A1 => n12982, A2 => n13237, B1 => n9187, B2 => 
                           n12980, ZN => n2757);
   U12105 : OAI22_X1 port map( A1 => n12982, A2 => n13240, B1 => n9172, B2 => 
                           n12980, ZN => n2758);
   U12106 : OAI22_X1 port map( A1 => n12982, A2 => n13243, B1 => n9157, B2 => 
                           n12980, ZN => n2759);
   U12107 : OAI22_X1 port map( A1 => n12983, A2 => n13246, B1 => n9142, B2 => 
                           n12980, ZN => n2760);
   U12108 : OAI22_X1 port map( A1 => n12983, A2 => n13249, B1 => n9127, B2 => 
                           n12980, ZN => n2761);
   U12109 : OAI22_X1 port map( A1 => n12983, A2 => n13252, B1 => n9112, B2 => 
                           n10970, ZN => n2762);
   U12110 : OAI22_X1 port map( A1 => n12983, A2 => n13255, B1 => n9097, B2 => 
                           n10970, ZN => n2763);
   U12111 : OAI22_X1 port map( A1 => n12983, A2 => n13258, B1 => n9082, B2 => 
                           n10970, ZN => n2764);
   U12112 : OAI22_X1 port map( A1 => n12984, A2 => n13261, B1 => n9067, B2 => 
                           n12980, ZN => n2765);
   U12113 : OAI22_X1 port map( A1 => n12984, A2 => n13264, B1 => n9052, B2 => 
                           n12980, ZN => n2766);
   U12114 : OAI22_X1 port map( A1 => n12984, A2 => n13267, B1 => n9037, B2 => 
                           n12980, ZN => n2767);
   U12115 : OAI22_X1 port map( A1 => n12984, A2 => n13270, B1 => n9022, B2 => 
                           n12980, ZN => n2768);
   U12116 : OAI22_X1 port map( A1 => n12984, A2 => n13273, B1 => n9007, B2 => 
                           n12980, ZN => n2769);
   U12117 : OAI22_X1 port map( A1 => n12985, A2 => n13276, B1 => n8992, B2 => 
                           n12980, ZN => n2770);
   U12118 : OAI22_X1 port map( A1 => n12985, A2 => n13279, B1 => n8977, B2 => 
                           n12980, ZN => n2771);
   U12119 : OAI22_X1 port map( A1 => n12985, A2 => n13282, B1 => n8962, B2 => 
                           n12980, ZN => n2772);
   U12120 : OAI22_X1 port map( A1 => n12985, A2 => n13285, B1 => n8947, B2 => 
                           n12980, ZN => n2773);
   U12121 : OAI22_X1 port map( A1 => n12972, A2 => n13216, B1 => n9291, B2 => 
                           n12971, ZN => n2718);
   U12122 : OAI22_X1 port map( A1 => n12972, A2 => n13219, B1 => n9276, B2 => 
                           n12971, ZN => n2719);
   U12123 : OAI22_X1 port map( A1 => n12972, A2 => n13222, B1 => n9261, B2 => 
                           n12971, ZN => n2720);
   U12124 : OAI22_X1 port map( A1 => n12972, A2 => n13225, B1 => n9246, B2 => 
                           n12971, ZN => n2721);
   U12125 : OAI22_X1 port map( A1 => n12972, A2 => n13228, B1 => n9231, B2 => 
                           n12971, ZN => n2722);
   U12126 : OAI22_X1 port map( A1 => n12973, A2 => n13231, B1 => n9216, B2 => 
                           n12971, ZN => n2723);
   U12127 : OAI22_X1 port map( A1 => n12973, A2 => n13234, B1 => n9201, B2 => 
                           n12971, ZN => n2724);
   U12128 : OAI22_X1 port map( A1 => n12973, A2 => n13237, B1 => n9186, B2 => 
                           n12971, ZN => n2725);
   U12129 : OAI22_X1 port map( A1 => n12973, A2 => n13240, B1 => n9171, B2 => 
                           n12971, ZN => n2726);
   U12130 : OAI22_X1 port map( A1 => n12973, A2 => n13243, B1 => n9156, B2 => 
                           n12971, ZN => n2727);
   U12131 : OAI22_X1 port map( A1 => n12974, A2 => n13246, B1 => n9141, B2 => 
                           n12971, ZN => n2728);
   U12132 : OAI22_X1 port map( A1 => n12974, A2 => n13249, B1 => n9126, B2 => 
                           n12971, ZN => n2729);
   U12133 : OAI22_X1 port map( A1 => n12974, A2 => n13252, B1 => n9111, B2 => 
                           n10971, ZN => n2730);
   U12134 : OAI22_X1 port map( A1 => n12974, A2 => n13255, B1 => n9096, B2 => 
                           n10971, ZN => n2731);
   U12135 : OAI22_X1 port map( A1 => n12974, A2 => n13258, B1 => n9081, B2 => 
                           n10971, ZN => n2732);
   U12136 : OAI22_X1 port map( A1 => n12975, A2 => n13261, B1 => n9066, B2 => 
                           n12971, ZN => n2733);
   U12137 : OAI22_X1 port map( A1 => n12975, A2 => n13264, B1 => n9051, B2 => 
                           n12971, ZN => n2734);
   U12138 : OAI22_X1 port map( A1 => n12975, A2 => n13267, B1 => n9036, B2 => 
                           n12971, ZN => n2735);
   U12139 : OAI22_X1 port map( A1 => n12975, A2 => n13270, B1 => n9021, B2 => 
                           n12971, ZN => n2736);
   U12140 : OAI22_X1 port map( A1 => n12975, A2 => n13273, B1 => n9006, B2 => 
                           n12971, ZN => n2737);
   U12141 : OAI22_X1 port map( A1 => n12976, A2 => n13276, B1 => n8991, B2 => 
                           n12971, ZN => n2738);
   U12142 : OAI22_X1 port map( A1 => n12976, A2 => n13279, B1 => n8976, B2 => 
                           n12971, ZN => n2739);
   U12143 : OAI22_X1 port map( A1 => n12976, A2 => n13282, B1 => n8961, B2 => 
                           n12971, ZN => n2740);
   U12144 : OAI22_X1 port map( A1 => n12976, A2 => n13285, B1 => n8946, B2 => 
                           n12971, ZN => n2741);
   U12145 : OAI22_X1 port map( A1 => n12945, A2 => n13216, B1 => n9294, B2 => 
                           n12944, ZN => n2622);
   U12146 : OAI22_X1 port map( A1 => n12945, A2 => n13219, B1 => n9279, B2 => 
                           n12944, ZN => n2623);
   U12147 : OAI22_X1 port map( A1 => n12945, A2 => n13222, B1 => n9264, B2 => 
                           n12944, ZN => n2624);
   U12148 : OAI22_X1 port map( A1 => n12945, A2 => n13225, B1 => n9249, B2 => 
                           n12944, ZN => n2625);
   U12149 : OAI22_X1 port map( A1 => n12945, A2 => n13228, B1 => n9234, B2 => 
                           n12944, ZN => n2626);
   U12150 : OAI22_X1 port map( A1 => n12946, A2 => n13231, B1 => n9219, B2 => 
                           n12944, ZN => n2627);
   U12151 : OAI22_X1 port map( A1 => n12946, A2 => n13234, B1 => n9204, B2 => 
                           n12944, ZN => n2628);
   U12152 : OAI22_X1 port map( A1 => n12946, A2 => n13237, B1 => n9189, B2 => 
                           n12944, ZN => n2629);
   U12153 : OAI22_X1 port map( A1 => n12946, A2 => n13240, B1 => n9174, B2 => 
                           n12944, ZN => n2630);
   U12154 : OAI22_X1 port map( A1 => n12946, A2 => n13243, B1 => n9159, B2 => 
                           n12944, ZN => n2631);
   U12155 : OAI22_X1 port map( A1 => n12947, A2 => n13246, B1 => n9144, B2 => 
                           n12944, ZN => n2632);
   U12156 : OAI22_X1 port map( A1 => n12947, A2 => n13249, B1 => n9129, B2 => 
                           n12944, ZN => n2633);
   U12157 : OAI22_X1 port map( A1 => n12947, A2 => n13252, B1 => n9114, B2 => 
                           n10974, ZN => n2634);
   U12158 : OAI22_X1 port map( A1 => n12947, A2 => n13255, B1 => n9099, B2 => 
                           n10974, ZN => n2635);
   U12159 : OAI22_X1 port map( A1 => n12947, A2 => n13258, B1 => n9084, B2 => 
                           n10974, ZN => n2636);
   U12160 : OAI22_X1 port map( A1 => n12948, A2 => n13261, B1 => n9069, B2 => 
                           n12944, ZN => n2637);
   U12161 : OAI22_X1 port map( A1 => n12948, A2 => n13264, B1 => n9054, B2 => 
                           n12944, ZN => n2638);
   U12162 : OAI22_X1 port map( A1 => n12948, A2 => n13267, B1 => n9039, B2 => 
                           n12944, ZN => n2639);
   U12163 : OAI22_X1 port map( A1 => n12948, A2 => n13270, B1 => n9024, B2 => 
                           n12944, ZN => n2640);
   U12164 : OAI22_X1 port map( A1 => n12948, A2 => n13273, B1 => n9009, B2 => 
                           n12944, ZN => n2641);
   U12165 : OAI22_X1 port map( A1 => n12949, A2 => n13276, B1 => n8994, B2 => 
                           n12944, ZN => n2642);
   U12166 : OAI22_X1 port map( A1 => n12949, A2 => n13279, B1 => n8979, B2 => 
                           n12944, ZN => n2643);
   U12167 : OAI22_X1 port map( A1 => n12949, A2 => n13282, B1 => n8964, B2 => 
                           n12944, ZN => n2644);
   U12168 : OAI22_X1 port map( A1 => n12949, A2 => n13285, B1 => n8949, B2 => 
                           n12944, ZN => n2645);
   U12169 : OAI21_X1 port map( B1 => n9280, B2 => n12828, A => n12251, ZN => 
                           n2526);
   U12170 : OAI21_X1 port map( B1 => n12252, B2 => n12253, A => n12831, ZN => 
                           n12251);
   U12171 : NAND4_X1 port map( A1 => n12270, A2 => n12271, A3 => n12272, A4 => 
                           n12273, ZN => n12252);
   U12172 : NAND4_X1 port map( A1 => n12254, A2 => n12255, A3 => n12256, A4 => 
                           n12257, ZN => n12253);
   U12173 : OAI21_X1 port map( B1 => n9265, B2 => n12828, A => n12232, ZN => 
                           n2527);
   U12174 : OAI21_X1 port map( B1 => n12233, B2 => n12234, A => n12831, ZN => 
                           n12232);
   U12175 : NAND4_X1 port map( A1 => n12243, A2 => n12244, A3 => n12245, A4 => 
                           n12246, ZN => n12233);
   U12176 : NAND4_X1 port map( A1 => n12235, A2 => n12236, A3 => n12237, A4 => 
                           n12238, ZN => n12234);
   U12177 : OAI21_X1 port map( B1 => n9250, B2 => n12828, A => n12213, ZN => 
                           n2528);
   U12178 : OAI21_X1 port map( B1 => n12214, B2 => n12215, A => n12830, ZN => 
                           n12213);
   U12179 : NAND4_X1 port map( A1 => n12224, A2 => n12225, A3 => n12226, A4 => 
                           n12227, ZN => n12214);
   U12180 : NAND4_X1 port map( A1 => n12216, A2 => n12217, A3 => n12218, A4 => 
                           n12219, ZN => n12215);
   U12181 : OAI21_X1 port map( B1 => n9235, B2 => n12828, A => n12194, ZN => 
                           n2529);
   U12182 : OAI21_X1 port map( B1 => n12195, B2 => n12196, A => n12830, ZN => 
                           n12194);
   U12183 : NAND4_X1 port map( A1 => n12205, A2 => n12206, A3 => n12207, A4 => 
                           n12208, ZN => n12195);
   U12184 : NAND4_X1 port map( A1 => n12197, A2 => n12198, A3 => n12199, A4 => 
                           n12200, ZN => n12196);
   U12185 : OAI21_X1 port map( B1 => n9220, B2 => n12828, A => n12175, ZN => 
                           n2530);
   U12186 : OAI21_X1 port map( B1 => n12176, B2 => n12177, A => n12830, ZN => 
                           n12175);
   U12187 : NAND4_X1 port map( A1 => n12186, A2 => n12187, A3 => n12188, A4 => 
                           n12189, ZN => n12176);
   U12188 : NAND4_X1 port map( A1 => n12178, A2 => n12179, A3 => n12180, A4 => 
                           n12181, ZN => n12177);
   U12189 : OAI21_X1 port map( B1 => n9205, B2 => n12828, A => n12156, ZN => 
                           n2531);
   U12190 : OAI21_X1 port map( B1 => n12157, B2 => n12158, A => n12829, ZN => 
                           n12156);
   U12191 : NAND4_X1 port map( A1 => n12167, A2 => n12168, A3 => n12169, A4 => 
                           n12170, ZN => n12157);
   U12192 : NAND4_X1 port map( A1 => n12159, A2 => n12160, A3 => n12161, A4 => 
                           n12162, ZN => n12158);
   U12193 : OAI21_X1 port map( B1 => n9190, B2 => n12828, A => n12137, ZN => 
                           n2532);
   U12194 : OAI21_X1 port map( B1 => n12138, B2 => n12139, A => n12830, ZN => 
                           n12137);
   U12195 : NAND4_X1 port map( A1 => n12148, A2 => n12149, A3 => n12150, A4 => 
                           n12151, ZN => n12138);
   U12196 : NAND4_X1 port map( A1 => n12140, A2 => n12141, A3 => n12142, A4 => 
                           n12143, ZN => n12139);
   U12197 : OAI21_X1 port map( B1 => n9160, B2 => n12828, A => n12099, ZN => 
                           n2534);
   U12198 : OAI21_X1 port map( B1 => n12100, B2 => n12101, A => n12829, ZN => 
                           n12099);
   U12199 : NAND4_X1 port map( A1 => n12110, A2 => n12111, A3 => n12112, A4 => 
                           n12113, ZN => n12100);
   U12200 : NAND4_X1 port map( A1 => n12102, A2 => n12103, A3 => n12104, A4 => 
                           n12105, ZN => n12101);
   U12201 : OAI21_X1 port map( B1 => n8814, B2 => n12930, A => n11598, ZN => 
                           n2558);
   U12202 : OAI21_X1 port map( B1 => n11599, B2 => n11600, A => n12933, ZN => 
                           n11598);
   U12203 : NAND4_X1 port map( A1 => n11617, A2 => n11618, A3 => n11619, A4 => 
                           n11620, ZN => n11599);
   U12204 : NAND4_X1 port map( A1 => n11601, A2 => n11602, A3 => n11603, A4 => 
                           n11604, ZN => n11600);
   U12205 : OAI21_X1 port map( B1 => n8813, B2 => n12930, A => n11579, ZN => 
                           n2559);
   U12206 : OAI21_X1 port map( B1 => n11580, B2 => n11581, A => n12933, ZN => 
                           n11579);
   U12207 : NAND4_X1 port map( A1 => n11590, A2 => n11591, A3 => n11592, A4 => 
                           n11593, ZN => n11580);
   U12208 : NAND4_X1 port map( A1 => n11582, A2 => n11583, A3 => n11584, A4 => 
                           n11585, ZN => n11581);
   U12209 : OAI21_X1 port map( B1 => n8812, B2 => n12930, A => n11560, ZN => 
                           n2560);
   U12210 : OAI21_X1 port map( B1 => n11561, B2 => n11562, A => n12932, ZN => 
                           n11560);
   U12211 : NAND4_X1 port map( A1 => n11571, A2 => n11572, A3 => n11573, A4 => 
                           n11574, ZN => n11561);
   U12212 : NAND4_X1 port map( A1 => n11563, A2 => n11564, A3 => n11565, A4 => 
                           n11566, ZN => n11562);
   U12213 : OAI21_X1 port map( B1 => n8811, B2 => n12930, A => n11541, ZN => 
                           n2561);
   U12214 : OAI21_X1 port map( B1 => n11542, B2 => n11543, A => n12932, ZN => 
                           n11541);
   U12215 : NAND4_X1 port map( A1 => n11552, A2 => n11553, A3 => n11554, A4 => 
                           n11555, ZN => n11542);
   U12216 : NAND4_X1 port map( A1 => n11544, A2 => n11545, A3 => n11546, A4 => 
                           n11547, ZN => n11543);
   U12217 : OAI21_X1 port map( B1 => n8810, B2 => n12930, A => n11522, ZN => 
                           n2562);
   U12218 : OAI21_X1 port map( B1 => n11523, B2 => n11524, A => n12932, ZN => 
                           n11522);
   U12219 : NAND4_X1 port map( A1 => n11533, A2 => n11534, A3 => n11535, A4 => 
                           n11536, ZN => n11523);
   U12220 : NAND4_X1 port map( A1 => n11525, A2 => n11526, A3 => n11527, A4 => 
                           n11528, ZN => n11524);
   U12221 : OAI21_X1 port map( B1 => n8809, B2 => n12930, A => n11503, ZN => 
                           n2563);
   U12222 : OAI21_X1 port map( B1 => n11504, B2 => n11505, A => n12931, ZN => 
                           n11503);
   U12223 : NAND4_X1 port map( A1 => n11514, A2 => n11515, A3 => n11516, A4 => 
                           n11517, ZN => n11504);
   U12224 : NAND4_X1 port map( A1 => n11506, A2 => n11507, A3 => n11508, A4 => 
                           n11509, ZN => n11505);
   U12225 : OAI21_X1 port map( B1 => n8808, B2 => n12930, A => n11484, ZN => 
                           n2564);
   U12226 : OAI21_X1 port map( B1 => n11485, B2 => n11486, A => n12932, ZN => 
                           n11484);
   U12227 : NAND4_X1 port map( A1 => n11495, A2 => n11496, A3 => n11497, A4 => 
                           n11498, ZN => n11485);
   U12228 : NAND4_X1 port map( A1 => n11487, A2 => n11488, A3 => n11489, A4 => 
                           n11490, ZN => n11486);
   U12229 : OAI21_X1 port map( B1 => n8806, B2 => n12930, A => n11446, ZN => 
                           n2566);
   U12230 : OAI21_X1 port map( B1 => n11447, B2 => n11448, A => n12931, ZN => 
                           n11446);
   U12231 : NAND4_X1 port map( A1 => n11457, A2 => n11458, A3 => n11459, A4 => 
                           n11460, ZN => n11447);
   U12232 : NAND4_X1 port map( A1 => n11449, A2 => n11450, A3 => n11451, A4 => 
                           n11452, ZN => n11448);
   U12233 : OAI21_X1 port map( B1 => n9175, B2 => n12827, A => n12118, ZN => 
                           n2533);
   U12234 : OAI21_X1 port map( B1 => n12119, B2 => n12120, A => n12829, ZN => 
                           n12118);
   U12235 : NAND4_X1 port map( A1 => n12129, A2 => n12130, A3 => n12131, A4 => 
                           n12132, ZN => n12119);
   U12236 : NAND4_X1 port map( A1 => n12121, A2 => n12122, A3 => n12123, A4 => 
                           n12124, ZN => n12120);
   U12237 : OAI21_X1 port map( B1 => n9145, B2 => n12827, A => n12080, ZN => 
                           n2535);
   U12238 : OAI21_X1 port map( B1 => n12081, B2 => n12082, A => n12829, ZN => 
                           n12080);
   U12239 : NAND4_X1 port map( A1 => n12091, A2 => n12092, A3 => n12093, A4 => 
                           n12094, ZN => n12081);
   U12240 : NAND4_X1 port map( A1 => n12083, A2 => n12084, A3 => n12085, A4 => 
                           n12086, ZN => n12082);
   U12241 : OAI21_X1 port map( B1 => n9130, B2 => n12827, A => n12061, ZN => 
                           n2536);
   U12242 : OAI21_X1 port map( B1 => n12062, B2 => n12063, A => n12828, ZN => 
                           n12061);
   U12243 : NAND4_X1 port map( A1 => n12072, A2 => n12073, A3 => n12074, A4 => 
                           n12075, ZN => n12062);
   U12244 : NAND4_X1 port map( A1 => n12064, A2 => n12065, A3 => n12066, A4 => 
                           n12067, ZN => n12063);
   U12245 : OAI21_X1 port map( B1 => n9115, B2 => n12827, A => n12042, ZN => 
                           n2537);
   U12246 : OAI21_X1 port map( B1 => n12043, B2 => n12044, A => n12828, ZN => 
                           n12042);
   U12247 : NAND4_X1 port map( A1 => n12053, A2 => n12054, A3 => n12055, A4 => 
                           n12056, ZN => n12043);
   U12248 : NAND4_X1 port map( A1 => n12045, A2 => n12046, A3 => n12047, A4 => 
                           n12048, ZN => n12044);
   U12249 : OAI21_X1 port map( B1 => n9100, B2 => n12827, A => n12023, ZN => 
                           n2538);
   U12250 : OAI21_X1 port map( B1 => n12024, B2 => n12025, A => n12829, ZN => 
                           n12023);
   U12251 : NAND4_X1 port map( A1 => n12034, A2 => n12035, A3 => n12036, A4 => 
                           n12037, ZN => n12024);
   U12252 : NAND4_X1 port map( A1 => n12026, A2 => n12027, A3 => n12028, A4 => 
                           n12029, ZN => n12025);
   U12253 : OAI21_X1 port map( B1 => n9085, B2 => n12827, A => n12004, ZN => 
                           n2539);
   U12254 : OAI21_X1 port map( B1 => n12005, B2 => n12006, A => n12828, ZN => 
                           n12004);
   U12255 : NAND4_X1 port map( A1 => n12015, A2 => n12016, A3 => n12017, A4 => 
                           n12018, ZN => n12005);
   U12256 : NAND4_X1 port map( A1 => n12007, A2 => n12008, A3 => n12009, A4 => 
                           n12010, ZN => n12006);
   U12257 : OAI21_X1 port map( B1 => n9070, B2 => n12827, A => n11985, ZN => 
                           n2540);
   U12258 : OAI21_X1 port map( B1 => n11986, B2 => n11987, A => n12828, ZN => 
                           n11985);
   U12259 : NAND4_X1 port map( A1 => n11996, A2 => n11997, A3 => n11998, A4 => 
                           n11999, ZN => n11986);
   U12260 : NAND4_X1 port map( A1 => n11988, A2 => n11989, A3 => n11990, A4 => 
                           n11991, ZN => n11987);
   U12261 : OAI21_X1 port map( B1 => n9055, B2 => n12827, A => n11966, ZN => 
                           n2541);
   U12262 : OAI21_X1 port map( B1 => n11967, B2 => n11968, A => n12829, ZN => 
                           n11966);
   U12263 : NAND4_X1 port map( A1 => n11977, A2 => n11978, A3 => n11979, A4 => 
                           n11980, ZN => n11967);
   U12264 : NAND4_X1 port map( A1 => n11969, A2 => n11970, A3 => n11971, A4 => 
                           n11972, ZN => n11968);
   U12265 : OAI21_X1 port map( B1 => n9040, B2 => n12827, A => n11947, ZN => 
                           n2542);
   U12266 : OAI21_X1 port map( B1 => n11948, B2 => n11949, A => n12829, ZN => 
                           n11947);
   U12267 : NAND4_X1 port map( A1 => n11958, A2 => n11959, A3 => n11960, A4 => 
                           n11961, ZN => n11948);
   U12268 : NAND4_X1 port map( A1 => n11950, A2 => n11951, A3 => n11952, A4 => 
                           n11953, ZN => n11949);
   U12269 : OAI21_X1 port map( B1 => n9025, B2 => n12827, A => n11928, ZN => 
                           n2543);
   U12270 : OAI21_X1 port map( B1 => n11929, B2 => n11930, A => n12829, ZN => 
                           n11928);
   U12271 : NAND4_X1 port map( A1 => n11939, A2 => n11940, A3 => n11941, A4 => 
                           n11942, ZN => n11929);
   U12272 : NAND4_X1 port map( A1 => n11931, A2 => n11932, A3 => n11933, A4 => 
                           n11934, ZN => n11930);
   U12273 : OAI21_X1 port map( B1 => n9010, B2 => n12827, A => n11909, ZN => 
                           n2544);
   U12274 : OAI21_X1 port map( B1 => n11910, B2 => n11911, A => n12829, ZN => 
                           n11909);
   U12275 : NAND4_X1 port map( A1 => n11920, A2 => n11921, A3 => n11922, A4 => 
                           n11923, ZN => n11910);
   U12276 : NAND4_X1 port map( A1 => n11912, A2 => n11913, A3 => n11914, A4 => 
                           n11915, ZN => n11911);
   U12277 : OAI21_X1 port map( B1 => n8995, B2 => n12826, A => n11890, ZN => 
                           n2545);
   U12278 : OAI21_X1 port map( B1 => n11891, B2 => n11892, A => n12829, ZN => 
                           n11890);
   U12279 : NAND4_X1 port map( A1 => n11901, A2 => n11902, A3 => n11903, A4 => 
                           n11904, ZN => n11891);
   U12280 : NAND4_X1 port map( A1 => n11893, A2 => n11894, A3 => n11895, A4 => 
                           n11896, ZN => n11892);
   U12281 : OAI21_X1 port map( B1 => n8980, B2 => n12826, A => n11871, ZN => 
                           n2546);
   U12282 : OAI21_X1 port map( B1 => n11872, B2 => n11873, A => n12829, ZN => 
                           n11871);
   U12283 : NAND4_X1 port map( A1 => n11882, A2 => n11883, A3 => n11884, A4 => 
                           n11885, ZN => n11872);
   U12284 : NAND4_X1 port map( A1 => n11874, A2 => n11875, A3 => n11876, A4 => 
                           n11877, ZN => n11873);
   U12285 : OAI21_X1 port map( B1 => n8965, B2 => n12826, A => n11852, ZN => 
                           n2547);
   U12286 : OAI21_X1 port map( B1 => n11853, B2 => n11854, A => n12830, ZN => 
                           n11852);
   U12287 : NAND4_X1 port map( A1 => n11863, A2 => n11864, A3 => n11865, A4 => 
                           n11866, ZN => n11853);
   U12288 : NAND4_X1 port map( A1 => n11855, A2 => n11856, A3 => n11857, A4 => 
                           n11858, ZN => n11854);
   U12289 : OAI21_X1 port map( B1 => n8950, B2 => n12826, A => n11833, ZN => 
                           n2548);
   U12290 : OAI21_X1 port map( B1 => n11834, B2 => n11835, A => n12829, ZN => 
                           n11833);
   U12291 : NAND4_X1 port map( A1 => n11844, A2 => n11845, A3 => n11846, A4 => 
                           n11847, ZN => n11834);
   U12292 : NAND4_X1 port map( A1 => n11836, A2 => n11837, A3 => n11838, A4 => 
                           n11839, ZN => n11835);
   U12293 : OAI21_X1 port map( B1 => n8935, B2 => n12826, A => n11814, ZN => 
                           n2549);
   U12294 : OAI21_X1 port map( B1 => n11815, B2 => n11816, A => n12830, ZN => 
                           n11814);
   U12295 : NAND4_X1 port map( A1 => n11825, A2 => n11826, A3 => n11827, A4 => 
                           n11828, ZN => n11815);
   U12296 : NAND4_X1 port map( A1 => n11817, A2 => n11818, A3 => n11819, A4 => 
                           n11820, ZN => n11816);
   U12297 : OAI21_X1 port map( B1 => n8920, B2 => n12826, A => n11795, ZN => 
                           n2550);
   U12298 : OAI21_X1 port map( B1 => n11796, B2 => n11797, A => n12830, ZN => 
                           n11795);
   U12299 : NAND4_X1 port map( A1 => n11806, A2 => n11807, A3 => n11808, A4 => 
                           n11809, ZN => n11796);
   U12300 : NAND4_X1 port map( A1 => n11798, A2 => n11799, A3 => n11800, A4 => 
                           n11801, ZN => n11797);
   U12301 : OAI21_X1 port map( B1 => n8905, B2 => n12826, A => n11776, ZN => 
                           n2551);
   U12302 : OAI21_X1 port map( B1 => n11777, B2 => n11778, A => n12830, ZN => 
                           n11776);
   U12303 : NAND4_X1 port map( A1 => n11787, A2 => n11788, A3 => n11789, A4 => 
                           n11790, ZN => n11777);
   U12304 : NAND4_X1 port map( A1 => n11779, A2 => n11780, A3 => n11781, A4 => 
                           n11782, ZN => n11778);
   U12305 : OAI21_X1 port map( B1 => n8890, B2 => n12826, A => n11757, ZN => 
                           n2552);
   U12306 : OAI21_X1 port map( B1 => n11758, B2 => n11759, A => n12830, ZN => 
                           n11757);
   U12307 : NAND4_X1 port map( A1 => n11768, A2 => n11769, A3 => n11770, A4 => 
                           n11771, ZN => n11758);
   U12308 : NAND4_X1 port map( A1 => n11760, A2 => n11761, A3 => n11762, A4 => 
                           n11763, ZN => n11759);
   U12309 : OAI21_X1 port map( B1 => n8875, B2 => n12826, A => n11738, ZN => 
                           n2553);
   U12310 : OAI21_X1 port map( B1 => n11739, B2 => n11740, A => n12830, ZN => 
                           n11738);
   U12311 : NAND4_X1 port map( A1 => n11749, A2 => n11750, A3 => n11751, A4 => 
                           n11752, ZN => n11739);
   U12312 : NAND4_X1 port map( A1 => n11741, A2 => n11742, A3 => n11743, A4 => 
                           n11744, ZN => n11740);
   U12313 : OAI21_X1 port map( B1 => n8860, B2 => n12826, A => n11719, ZN => 
                           n2554);
   U12314 : OAI21_X1 port map( B1 => n11720, B2 => n11721, A => n12830, ZN => 
                           n11719);
   U12315 : NAND4_X1 port map( A1 => n11730, A2 => n11731, A3 => n11732, A4 => 
                           n11733, ZN => n11720);
   U12316 : NAND4_X1 port map( A1 => n11722, A2 => n11723, A3 => n11724, A4 => 
                           n11725, ZN => n11721);
   U12317 : OAI21_X1 port map( B1 => n8845, B2 => n12826, A => n11700, ZN => 
                           n2555);
   U12318 : OAI21_X1 port map( B1 => n11701, B2 => n11702, A => n12830, ZN => 
                           n11700);
   U12319 : NAND4_X1 port map( A1 => n11711, A2 => n11712, A3 => n11713, A4 => 
                           n11714, ZN => n11701);
   U12320 : NAND4_X1 port map( A1 => n11703, A2 => n11704, A3 => n11705, A4 => 
                           n11706, ZN => n11702);
   U12321 : OAI21_X1 port map( B1 => n8830, B2 => n12826, A => n11681, ZN => 
                           n2556);
   U12322 : OAI21_X1 port map( B1 => n11682, B2 => n11683, A => n12831, ZN => 
                           n11681);
   U12323 : NAND4_X1 port map( A1 => n11692, A2 => n11693, A3 => n11694, A4 => 
                           n11695, ZN => n11682);
   U12324 : NAND4_X1 port map( A1 => n11684, A2 => n11685, A3 => n11686, A4 => 
                           n11687, ZN => n11683);
   U12325 : OAI21_X1 port map( B1 => n8815, B2 => n12827, A => n11630, ZN => 
                           n2557);
   U12326 : OAI21_X1 port map( B1 => n11631, B2 => n11632, A => n12831, ZN => 
                           n11630);
   U12327 : NAND4_X1 port map( A1 => n11657, A2 => n11658, A3 => n11659, A4 => 
                           n11660, ZN => n11631);
   U12328 : NAND4_X1 port map( A1 => n11633, A2 => n11634, A3 => n11635, A4 => 
                           n11636, ZN => n11632);
   U12329 : OAI21_X1 port map( B1 => n8807, B2 => n12929, A => n11465, ZN => 
                           n2565);
   U12330 : OAI21_X1 port map( B1 => n11466, B2 => n11467, A => n12931, ZN => 
                           n11465);
   U12331 : NAND4_X1 port map( A1 => n11476, A2 => n11477, A3 => n11478, A4 => 
                           n11479, ZN => n11466);
   U12332 : NAND4_X1 port map( A1 => n11468, A2 => n11469, A3 => n11470, A4 => 
                           n11471, ZN => n11467);
   U12333 : OAI21_X1 port map( B1 => n8805, B2 => n12929, A => n11427, ZN => 
                           n2567);
   U12334 : OAI21_X1 port map( B1 => n11428, B2 => n11429, A => n12931, ZN => 
                           n11427);
   U12335 : NAND4_X1 port map( A1 => n11438, A2 => n11439, A3 => n11440, A4 => 
                           n11441, ZN => n11428);
   U12336 : NAND4_X1 port map( A1 => n11430, A2 => n11431, A3 => n11432, A4 => 
                           n11433, ZN => n11429);
   U12337 : OAI21_X1 port map( B1 => n8804, B2 => n12929, A => n11408, ZN => 
                           n2568);
   U12338 : OAI21_X1 port map( B1 => n11409, B2 => n11410, A => n12930, ZN => 
                           n11408);
   U12339 : NAND4_X1 port map( A1 => n11419, A2 => n11420, A3 => n11421, A4 => 
                           n11422, ZN => n11409);
   U12340 : NAND4_X1 port map( A1 => n11411, A2 => n11412, A3 => n11413, A4 => 
                           n11414, ZN => n11410);
   U12341 : OAI21_X1 port map( B1 => n8803, B2 => n12929, A => n11389, ZN => 
                           n2569);
   U12342 : OAI21_X1 port map( B1 => n11390, B2 => n11391, A => n12930, ZN => 
                           n11389);
   U12343 : NAND4_X1 port map( A1 => n11400, A2 => n11401, A3 => n11402, A4 => 
                           n11403, ZN => n11390);
   U12344 : NAND4_X1 port map( A1 => n11392, A2 => n11393, A3 => n11394, A4 => 
                           n11395, ZN => n11391);
   U12345 : OAI21_X1 port map( B1 => n8802, B2 => n12929, A => n11370, ZN => 
                           n2570);
   U12346 : OAI21_X1 port map( B1 => n11371, B2 => n11372, A => n12931, ZN => 
                           n11370);
   U12347 : NAND4_X1 port map( A1 => n11381, A2 => n11382, A3 => n11383, A4 => 
                           n11384, ZN => n11371);
   U12348 : NAND4_X1 port map( A1 => n11373, A2 => n11374, A3 => n11375, A4 => 
                           n11376, ZN => n11372);
   U12349 : OAI21_X1 port map( B1 => n8801, B2 => n12929, A => n11351, ZN => 
                           n2571);
   U12350 : OAI21_X1 port map( B1 => n11352, B2 => n11353, A => n12930, ZN => 
                           n11351);
   U12351 : NAND4_X1 port map( A1 => n11362, A2 => n11363, A3 => n11364, A4 => 
                           n11365, ZN => n11352);
   U12352 : NAND4_X1 port map( A1 => n11354, A2 => n11355, A3 => n11356, A4 => 
                           n11357, ZN => n11353);
   U12353 : OAI21_X1 port map( B1 => n8800, B2 => n12929, A => n11332, ZN => 
                           n2572);
   U12354 : OAI21_X1 port map( B1 => n11333, B2 => n11334, A => n12930, ZN => 
                           n11332);
   U12355 : NAND4_X1 port map( A1 => n11343, A2 => n11344, A3 => n11345, A4 => 
                           n11346, ZN => n11333);
   U12356 : NAND4_X1 port map( A1 => n11335, A2 => n11336, A3 => n11337, A4 => 
                           n11338, ZN => n11334);
   U12357 : OAI21_X1 port map( B1 => n8799, B2 => n12929, A => n11313, ZN => 
                           n2573);
   U12358 : OAI21_X1 port map( B1 => n11314, B2 => n11315, A => n12931, ZN => 
                           n11313);
   U12359 : NAND4_X1 port map( A1 => n11324, A2 => n11325, A3 => n11326, A4 => 
                           n11327, ZN => n11314);
   U12360 : NAND4_X1 port map( A1 => n11316, A2 => n11317, A3 => n11318, A4 => 
                           n11319, ZN => n11315);
   U12361 : OAI21_X1 port map( B1 => n8798, B2 => n12929, A => n11294, ZN => 
                           n2574);
   U12362 : OAI21_X1 port map( B1 => n11295, B2 => n11296, A => n12931, ZN => 
                           n11294);
   U12363 : NAND4_X1 port map( A1 => n11305, A2 => n11306, A3 => n11307, A4 => 
                           n11308, ZN => n11295);
   U12364 : NAND4_X1 port map( A1 => n11297, A2 => n11298, A3 => n11299, A4 => 
                           n11300, ZN => n11296);
   U12365 : OAI21_X1 port map( B1 => n8797, B2 => n12929, A => n11275, ZN => 
                           n2575);
   U12366 : OAI21_X1 port map( B1 => n11276, B2 => n11277, A => n12931, ZN => 
                           n11275);
   U12367 : NAND4_X1 port map( A1 => n11286, A2 => n11287, A3 => n11288, A4 => 
                           n11289, ZN => n11276);
   U12368 : NAND4_X1 port map( A1 => n11278, A2 => n11279, A3 => n11280, A4 => 
                           n11281, ZN => n11277);
   U12369 : OAI21_X1 port map( B1 => n8796, B2 => n12929, A => n11256, ZN => 
                           n2576);
   U12370 : OAI21_X1 port map( B1 => n11257, B2 => n11258, A => n12931, ZN => 
                           n11256);
   U12371 : NAND4_X1 port map( A1 => n11267, A2 => n11268, A3 => n11269, A4 => 
                           n11270, ZN => n11257);
   U12372 : NAND4_X1 port map( A1 => n11259, A2 => n11260, A3 => n11261, A4 => 
                           n11262, ZN => n11258);
   U12373 : OAI21_X1 port map( B1 => n8795, B2 => n12928, A => n11237, ZN => 
                           n2577);
   U12374 : OAI21_X1 port map( B1 => n11238, B2 => n11239, A => n12931, ZN => 
                           n11237);
   U12375 : NAND4_X1 port map( A1 => n11248, A2 => n11249, A3 => n11250, A4 => 
                           n11251, ZN => n11238);
   U12376 : NAND4_X1 port map( A1 => n11240, A2 => n11241, A3 => n11242, A4 => 
                           n11243, ZN => n11239);
   U12377 : OAI21_X1 port map( B1 => n8794, B2 => n12928, A => n11218, ZN => 
                           n2578);
   U12378 : OAI21_X1 port map( B1 => n11219, B2 => n11220, A => n12931, ZN => 
                           n11218);
   U12379 : NAND4_X1 port map( A1 => n11229, A2 => n11230, A3 => n11231, A4 => 
                           n11232, ZN => n11219);
   U12380 : NAND4_X1 port map( A1 => n11221, A2 => n11222, A3 => n11223, A4 => 
                           n11224, ZN => n11220);
   U12381 : OAI21_X1 port map( B1 => n8793, B2 => n12928, A => n11199, ZN => 
                           n2579);
   U12382 : OAI21_X1 port map( B1 => n11200, B2 => n11201, A => n12932, ZN => 
                           n11199);
   U12383 : NAND4_X1 port map( A1 => n11210, A2 => n11211, A3 => n11212, A4 => 
                           n11213, ZN => n11200);
   U12384 : NAND4_X1 port map( A1 => n11202, A2 => n11203, A3 => n11204, A4 => 
                           n11205, ZN => n11201);
   U12385 : OAI21_X1 port map( B1 => n8792, B2 => n12928, A => n11180, ZN => 
                           n2580);
   U12386 : OAI21_X1 port map( B1 => n11181, B2 => n11182, A => n12931, ZN => 
                           n11180);
   U12387 : NAND4_X1 port map( A1 => n11191, A2 => n11192, A3 => n11193, A4 => 
                           n11194, ZN => n11181);
   U12388 : NAND4_X1 port map( A1 => n11183, A2 => n11184, A3 => n11185, A4 => 
                           n11186, ZN => n11182);
   U12389 : OAI21_X1 port map( B1 => n8791, B2 => n12928, A => n11161, ZN => 
                           n2581);
   U12390 : OAI21_X1 port map( B1 => n11162, B2 => n11163, A => n12932, ZN => 
                           n11161);
   U12391 : NAND4_X1 port map( A1 => n11172, A2 => n11173, A3 => n11174, A4 => 
                           n11175, ZN => n11162);
   U12392 : NAND4_X1 port map( A1 => n11164, A2 => n11165, A3 => n11166, A4 => 
                           n11167, ZN => n11163);
   U12393 : OAI21_X1 port map( B1 => n8790, B2 => n12928, A => n11142, ZN => 
                           n2582);
   U12394 : OAI21_X1 port map( B1 => n11143, B2 => n11144, A => n12932, ZN => 
                           n11142);
   U12395 : NAND4_X1 port map( A1 => n11153, A2 => n11154, A3 => n11155, A4 => 
                           n11156, ZN => n11143);
   U12396 : NAND4_X1 port map( A1 => n11145, A2 => n11146, A3 => n11147, A4 => 
                           n11148, ZN => n11144);
   U12397 : OAI21_X1 port map( B1 => n8789, B2 => n12928, A => n11123, ZN => 
                           n2583);
   U12398 : OAI21_X1 port map( B1 => n11124, B2 => n11125, A => n12932, ZN => 
                           n11123);
   U12399 : NAND4_X1 port map( A1 => n11134, A2 => n11135, A3 => n11136, A4 => 
                           n11137, ZN => n11124);
   U12400 : NAND4_X1 port map( A1 => n11126, A2 => n11127, A3 => n11128, A4 => 
                           n11129, ZN => n11125);
   U12401 : OAI21_X1 port map( B1 => n8788, B2 => n12928, A => n11104, ZN => 
                           n2584);
   U12402 : OAI21_X1 port map( B1 => n11105, B2 => n11106, A => n12932, ZN => 
                           n11104);
   U12403 : NAND4_X1 port map( A1 => n11115, A2 => n11116, A3 => n11117, A4 => 
                           n11118, ZN => n11105);
   U12404 : NAND4_X1 port map( A1 => n11107, A2 => n11108, A3 => n11109, A4 => 
                           n11110, ZN => n11106);
   U12405 : OAI21_X1 port map( B1 => n8787, B2 => n12928, A => n11085, ZN => 
                           n2585);
   U12406 : OAI21_X1 port map( B1 => n11086, B2 => n11087, A => n12932, ZN => 
                           n11085);
   U12407 : NAND4_X1 port map( A1 => n11096, A2 => n11097, A3 => n11098, A4 => 
                           n11099, ZN => n11086);
   U12408 : NAND4_X1 port map( A1 => n11088, A2 => n11089, A3 => n11090, A4 => 
                           n11091, ZN => n11087);
   U12409 : OAI21_X1 port map( B1 => n8786, B2 => n12928, A => n11066, ZN => 
                           n2586);
   U12410 : OAI21_X1 port map( B1 => n11067, B2 => n11068, A => n12932, ZN => 
                           n11066);
   U12411 : NAND4_X1 port map( A1 => n11077, A2 => n11078, A3 => n11079, A4 => 
                           n11080, ZN => n11067);
   U12412 : NAND4_X1 port map( A1 => n11069, A2 => n11070, A3 => n11071, A4 => 
                           n11072, ZN => n11068);
   U12413 : OAI21_X1 port map( B1 => n8785, B2 => n12928, A => n11047, ZN => 
                           n2587);
   U12414 : OAI21_X1 port map( B1 => n11048, B2 => n11049, A => n12932, ZN => 
                           n11047);
   U12415 : NAND4_X1 port map( A1 => n11058, A2 => n11059, A3 => n11060, A4 => 
                           n11061, ZN => n11048);
   U12416 : NAND4_X1 port map( A1 => n11050, A2 => n11051, A3 => n11052, A4 => 
                           n11053, ZN => n11049);
   U12417 : OAI21_X1 port map( B1 => n8784, B2 => n12928, A => n11028, ZN => 
                           n2588);
   U12418 : OAI21_X1 port map( B1 => n11029, B2 => n11030, A => n12933, ZN => 
                           n11028);
   U12419 : NAND4_X1 port map( A1 => n11039, A2 => n11040, A3 => n11041, A4 => 
                           n11042, ZN => n11029);
   U12420 : NAND4_X1 port map( A1 => n11031, A2 => n11032, A3 => n11033, A4 => 
                           n11034, ZN => n11030);
   U12421 : OAI21_X1 port map( B1 => n8783, B2 => n12929, A => n10977, ZN => 
                           n2589);
   U12422 : OAI21_X1 port map( B1 => n10978, B2 => n10979, A => n12933, ZN => 
                           n10977);
   U12423 : NAND4_X1 port map( A1 => n11004, A2 => n11005, A3 => n11006, A4 => 
                           n11007, ZN => n10978);
   U12424 : NAND4_X1 port map( A1 => n10980, A2 => n10981, A3 => n10982, A4 => 
                           n10983, ZN => n10979);
   U12425 : OAI22_X1 port map( A1 => n13053, A2 => n13215, B1 => n13052, B2 => 
                           n10542, ZN => n3006);
   U12426 : OAI22_X1 port map( A1 => n13053, A2 => n13218, B1 => n13052, B2 => 
                           n10541, ZN => n3007);
   U12427 : OAI22_X1 port map( A1 => n13053, A2 => n13221, B1 => n13052, B2 => 
                           n10540, ZN => n3008);
   U12428 : OAI22_X1 port map( A1 => n13053, A2 => n13224, B1 => n13052, B2 => 
                           n10539, ZN => n3009);
   U12429 : OAI22_X1 port map( A1 => n13053, A2 => n13227, B1 => n13052, B2 => 
                           n10538, ZN => n3010);
   U12430 : OAI22_X1 port map( A1 => n13054, A2 => n13230, B1 => n13052, B2 => 
                           n10537, ZN => n3011);
   U12431 : OAI22_X1 port map( A1 => n13054, A2 => n13233, B1 => n13052, B2 => 
                           n10536, ZN => n3012);
   U12432 : OAI22_X1 port map( A1 => n13054, A2 => n13236, B1 => n13052, B2 => 
                           n10535, ZN => n3013);
   U12433 : OAI22_X1 port map( A1 => n13054, A2 => n13239, B1 => n13052, B2 => 
                           n10534, ZN => n3014);
   U12434 : OAI22_X1 port map( A1 => n13054, A2 => n13242, B1 => n13052, B2 => 
                           n10533, ZN => n3015);
   U12435 : OAI22_X1 port map( A1 => n13055, A2 => n13245, B1 => n13052, B2 => 
                           n10532, ZN => n3016);
   U12436 : OAI22_X1 port map( A1 => n13055, A2 => n13248, B1 => n13052, B2 => 
                           n10531, ZN => n3017);
   U12437 : OAI22_X1 port map( A1 => n13055, A2 => n13251, B1 => n10961, B2 => 
                           n10530, ZN => n3018);
   U12438 : OAI22_X1 port map( A1 => n13055, A2 => n13254, B1 => n10961, B2 => 
                           n10529, ZN => n3019);
   U12439 : OAI22_X1 port map( A1 => n13055, A2 => n13257, B1 => n10961, B2 => 
                           n10528, ZN => n3020);
   U12440 : OAI22_X1 port map( A1 => n13056, A2 => n13260, B1 => n13052, B2 => 
                           n10527, ZN => n3021);
   U12441 : OAI22_X1 port map( A1 => n13056, A2 => n13263, B1 => n13052, B2 => 
                           n10526, ZN => n3022);
   U12442 : OAI22_X1 port map( A1 => n13056, A2 => n13266, B1 => n13052, B2 => 
                           n10525, ZN => n3023);
   U12443 : OAI22_X1 port map( A1 => n13056, A2 => n13269, B1 => n13052, B2 => 
                           n10524, ZN => n3024);
   U12444 : OAI22_X1 port map( A1 => n13056, A2 => n13272, B1 => n13052, B2 => 
                           n10523, ZN => n3025);
   U12445 : OAI22_X1 port map( A1 => n13057, A2 => n13275, B1 => n13052, B2 => 
                           n10522, ZN => n3026);
   U12446 : OAI22_X1 port map( A1 => n13057, A2 => n13278, B1 => n13052, B2 => 
                           n10521, ZN => n3027);
   U12447 : OAI22_X1 port map( A1 => n13057, A2 => n13281, B1 => n13052, B2 => 
                           n10520, ZN => n3028);
   U12448 : OAI22_X1 port map( A1 => n13057, A2 => n13284, B1 => n13052, B2 => 
                           n10519, ZN => n3029);
   U12449 : OAI22_X1 port map( A1 => n13057, A2 => n13287, B1 => n10961, B2 => 
                           n10386, ZN => n3030);
   U12450 : OAI22_X1 port map( A1 => n13058, A2 => n13290, B1 => n10961, B2 => 
                           n10385, ZN => n3031);
   U12451 : OAI22_X1 port map( A1 => n13058, A2 => n13293, B1 => n10961, B2 => 
                           n10384, ZN => n3032);
   U12452 : OAI22_X1 port map( A1 => n13058, A2 => n13296, B1 => n10961, B2 => 
                           n10383, ZN => n3033);
   U12453 : OAI22_X1 port map( A1 => n13058, A2 => n13299, B1 => n10961, B2 => 
                           n10382, ZN => n3034);
   U12454 : OAI22_X1 port map( A1 => n13058, A2 => n13302, B1 => n10961, B2 => 
                           n10381, ZN => n3035);
   U12455 : OAI22_X1 port map( A1 => n13059, A2 => n13305, B1 => n10961, B2 => 
                           n10380, ZN => n3036);
   U12456 : OAI22_X1 port map( A1 => n13059, A2 => n13317, B1 => n10961, B2 => 
                           n10379, ZN => n3037);
   U12457 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(3), A3 => n9929, 
                           ZN => n12275);
   U12458 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(3), A3 => n9934, 
                           ZN => n11622);
   U12459 : NOR3_X1 port map( A1 => n9929, A2 => ADD_RD1(3), A3 => n9933, ZN =>
                           n12276);
   U12460 : NOR3_X1 port map( A1 => n9934, A2 => ADD_RD2(3), A3 => n9938, ZN =>
                           n11623);
   U12461 : NOR2_X1 port map( A1 => n9937, A2 => ADD_RD2(2), ZN => n11609);
   U12462 : NOR2_X1 port map( A1 => n9931, A2 => ADD_RD1(1), ZN => n12265);
   U12463 : NOR2_X1 port map( A1 => n9936, A2 => ADD_RD2(1), ZN => n11612);
   U12464 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => 
                           ADD_RD1(0), ZN => n12261);
   U12465 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => 
                           ADD_RD2(0), ZN => n11608);
   U12466 : NOR3_X1 port map( A1 => n9933, A2 => ADD_RD1(4), A3 => n9930, ZN =>
                           n12268);
   U12467 : NOR3_X1 port map( A1 => n9929, A2 => ADD_RD1(0), A3 => n9930, ZN =>
                           n12279);
   U12468 : NOR3_X1 port map( A1 => n9938, A2 => ADD_RD2(4), A3 => n9935, ZN =>
                           n11615);
   U12469 : NOR3_X1 port map( A1 => n9934, A2 => ADD_RD2(0), A3 => n9935, ZN =>
                           n11626);
   U12470 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => n9933, 
                           ZN => n12259);
   U12471 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(4), A3 => n9930, 
                           ZN => n12267);
   U12472 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => n9938, 
                           ZN => n11606);
   U12473 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(4), A3 => n9935, 
                           ZN => n11614);
   U12474 : NOR2_X1 port map( A1 => n9932, A2 => ADD_RD1(2), ZN => n12262);
   U12475 : INV_X1 port map( A => RESET, ZN => n9923);
   U12476 : AND3_X1 port map( A1 => ENABLE, A2 => n13324, A3 => RD1, ZN => 
                           n11629);
   U12477 : AND3_X1 port map( A1 => ENABLE, A2 => n13324, A3 => RD2, ZN => 
                           n10976);
   U12478 : INV_X1 port map( A => ADD_RD1(3), ZN => n9930);
   U12479 : INV_X1 port map( A => ADD_RD2(3), ZN => n9935);
   U12480 : INV_X1 port map( A => ADD_RD1(0), ZN => n9933);
   U12481 : INV_X1 port map( A => ADD_RD2(0), ZN => n9938);
   U12482 : INV_X1 port map( A => ADD_RD1(4), ZN => n9929);
   U12483 : INV_X1 port map( A => ADD_RD2(4), ZN => n9934);
   U12484 : NAND2_X1 port map( A1 => DATAIN(31), A2 => n13319, ZN => n10899);
   U12485 : NAND2_X1 port map( A1 => DATAIN(20), A2 => n13319, ZN => n10911);
   U12486 : NAND2_X1 port map( A1 => DATAIN(21), A2 => n13319, ZN => n10910);
   U12487 : NAND2_X1 port map( A1 => DATAIN(22), A2 => n13319, ZN => n10909);
   U12488 : NAND2_X1 port map( A1 => DATAIN(28), A2 => n13319, ZN => n10903);
   U12489 : NAND2_X1 port map( A1 => DATAIN(29), A2 => n13319, ZN => n10902);
   U12490 : NAND2_X1 port map( A1 => DATAIN(30), A2 => n13319, ZN => n10901);
   U12491 : NAND2_X1 port map( A1 => DATAIN(8), A2 => n13320, ZN => n10923);
   U12492 : NAND2_X1 port map( A1 => DATAIN(9), A2 => n13320, ZN => n10922);
   U12493 : NAND2_X1 port map( A1 => DATAIN(10), A2 => n13320, ZN => n10921);
   U12494 : NAND2_X1 port map( A1 => DATAIN(11), A2 => n13320, ZN => n10920);
   U12495 : NAND2_X1 port map( A1 => DATAIN(12), A2 => n13320, ZN => n10919);
   U12496 : NAND2_X1 port map( A1 => DATAIN(13), A2 => n13320, ZN => n10918);
   U12497 : NAND2_X1 port map( A1 => DATAIN(14), A2 => n13320, ZN => n10917);
   U12498 : NAND2_X1 port map( A1 => DATAIN(15), A2 => n13320, ZN => n10916);
   U12499 : NAND2_X1 port map( A1 => DATAIN(16), A2 => n13320, ZN => n10915);
   U12500 : NAND2_X1 port map( A1 => DATAIN(17), A2 => n13320, ZN => n10914);
   U12501 : NAND2_X1 port map( A1 => DATAIN(18), A2 => n13320, ZN => n10913);
   U12502 : NAND2_X1 port map( A1 => DATAIN(19), A2 => n13320, ZN => n10912);
   U12503 : NAND2_X1 port map( A1 => DATAIN(23), A2 => n13319, ZN => n10908);
   U12504 : NAND2_X1 port map( A1 => DATAIN(24), A2 => n13319, ZN => n10907);
   U12505 : NAND2_X1 port map( A1 => DATAIN(25), A2 => n13319, ZN => n10906);
   U12506 : NAND2_X1 port map( A1 => DATAIN(26), A2 => n13319, ZN => n10905);
   U12507 : NAND2_X1 port map( A1 => DATAIN(27), A2 => n13319, ZN => n10904);
   U12508 : NAND2_X1 port map( A1 => DATAIN(0), A2 => n13321, ZN => n10931);
   U12509 : NAND2_X1 port map( A1 => DATAIN(1), A2 => n13321, ZN => n10930);
   U12510 : NAND2_X1 port map( A1 => DATAIN(2), A2 => n13321, ZN => n10929);
   U12511 : NAND2_X1 port map( A1 => DATAIN(3), A2 => n13321, ZN => n10928);
   U12512 : NAND2_X1 port map( A1 => DATAIN(4), A2 => n13321, ZN => n10927);
   U12513 : NAND2_X1 port map( A1 => DATAIN(5), A2 => n13321, ZN => n10926);
   U12514 : NAND2_X1 port map( A1 => DATAIN(6), A2 => n13321, ZN => n10925);
   U12515 : NAND2_X1 port map( A1 => DATAIN(7), A2 => n13321, ZN => n10924);
   U12516 : AND2_X1 port map( A1 => WR, A2 => ENABLE, ZN => n10948);
   U12517 : INV_X1 port map( A => ADD_WR(2), ZN => n9926);
   U12518 : INV_X1 port map( A => ADD_WR(0), ZN => n9928);
   U12519 : INV_X1 port map( A => ADD_WR(1), ZN => n9927);
   U12520 : INV_X1 port map( A => ADD_RD1(1), ZN => n9932);
   U12521 : INV_X1 port map( A => ADD_RD2(1), ZN => n9937);
   U12522 : INV_X1 port map( A => ADD_RD1(2), ZN => n9931);
   U12523 : INV_X1 port map( A => ADD_RD2(2), ZN => n9936);
   U12524 : INV_X1 port map( A => ADD_WR(4), ZN => n9924);
   U12525 : INV_X1 port map( A => ADD_WR(3), ZN => n9925);
   U12526 : CLKBUF_X1 port map( A => n11629, Z => n12831);
   U12527 : CLKBUF_X1 port map( A => n10976, Z => n12933);
   U12528 : CLKBUF_X1 port map( A => n9923, Z => n13324);

end SYN_Behavioural;
