
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_RF_ADDR_W5_DATA_W32 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_RF_ADDR_W5_DATA_W32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_RF_ADDR_W5_DATA_W32.all;

entity RF_ADDR_W5_DATA_W32 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end RF_ADDR_W5_DATA_W32;

architecture SYN_Behavioural of RF_ADDR_W5_DATA_W32 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7, n8, n9, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
      n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n2526, n2527, n2528, 
      n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, 
      n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, 
      n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, 
      n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, 
      n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, 
      n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, 
      n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, 
      n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, 
      n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, 
      n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, 
      n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, 
      n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, 
      n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, 
      n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, 
      n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, 
      n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, 
      n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, 
      n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, 
      n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, 
      n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, 
      n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, 
      n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, 
      n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, 
      n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, 
      n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, 
      n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, 
      n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, 
      n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, 
      n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, 
      n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, 
      n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, 
      n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, 
      n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, 
      n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, 
      n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, 
      n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, 
      n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, 
      n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, 
      n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, 
      n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, 
      n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, 
      n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, 
      n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, 
      n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, 
      n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, 
      n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, 
      n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, 
      n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, 
      n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, 
      n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, 
      n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, 
      n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, 
      n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, 
      n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, 
      n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, 
      n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, 
      n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, 
      n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, 
      n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, 
      n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, 
      n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, 
      n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, 
      n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, 
      n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, 
      n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, 
      n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, 
      n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, 
      n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, 
      n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, 
      n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, 
      n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, 
      n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, 
      n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, 
      n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, 
      n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, 
      n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, 
      n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, 
      n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, 
      n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, 
      n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, 
      n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, 
      n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, 
      n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, 
      n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, 
      n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, 
      n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, 
      n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, 
      n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, 
      n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, 
      n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, 
      n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, 
      n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, 
      n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, 
      n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, 
      n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, 
      n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, 
      n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, 
      n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, 
      n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, 
      n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, 
      n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, 
      n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, 
      n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, 
      n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, 
      n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, 
      n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, 
      n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, 
      n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, 
      n3609, n3610, n3611, n3612, n3613, n3934, n3935, n3936, n3937, n3938, 
      n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, 
      n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, 
      n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, 
      n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, 
      n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, 
      n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n4318, 
      n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, 
      n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, 
      n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, 
      n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, 
      n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, 
      n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, 
      n4379, n4380, n4381, n4414, n4415, n4416, n4417, n4418, n4419, n4420, 
      n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, 
      n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, 
      n4441, n4442, n4443, n4444, n4445, n4478, n4479, n4480, n4481, n4482, 
      n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, 
      n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, 
      n4503, n4504, n4505, n4506, n4507, n4508, n4509, n6451, n6452, n6453, 
      n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, 
      n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, 
      n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, 
      n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, 
      n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, 
      n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, 
      n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, 
      n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, 
      n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, 
      n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, 
      n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, 
      n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, 
      n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, 
      n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, 
      n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, 
      n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, 
      n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, 
      n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, 
      n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, 
      n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, 
      n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, 
      n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, 
      n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, 
      n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, 
      n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, 
      n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, 
      n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, 
      n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, 
      n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, 
      n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, 
      n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, 
      n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, 
      n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, 
      n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, 
      n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, 
      n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, 
      n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, 
      n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, 
      n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, 
      n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, 
      n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, 
      n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, 
      n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, 
      n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, 
      n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, 
      n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, 
      n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, 
      n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, 
      n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, 
      n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, 
      n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, 
      n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, 
      n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, 
      n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, 
      n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, 
      n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, 
      n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, 
      n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, 
      n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, 
      n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, 
      n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, 
      n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, 
      n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, 
      n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, 
      n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, 
      n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, 
      n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, 
      n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, 
      n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, 
      n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, 
      n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, 
      n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, 
      n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, 
      n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, 
      n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, 
      n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, 
      n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, 
      n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, 
      n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, 
      n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, 
      n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, 
      n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, 
      n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, 
      n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, 
      n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, 
      n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, 
      n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, 
      n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, 
      n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, 
      n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, 
      n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, 
      n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, 
      n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, 
      n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, 
      n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, 
      n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, 
      n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, 
      n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, 
      n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, 
      n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, 
      n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, 
      n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, 
      n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, 
      n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, 
      n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, 
      n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, 
      n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, 
      n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, 
      n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, 
      n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, 
      n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, 
      n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, 
      n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, 
      n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, 
      n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, 
      n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, 
      n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, 
      n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, 
      n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, 
      n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, 
      n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, 
      n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, 
      n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, 
      n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, 
      n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, 
      n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, 
      n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, 
      n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, 
      n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, 
      n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, 
      n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, 
      n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, 
      n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, 
      n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, 
      n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, 
      n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, 
      n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, 
      n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, 
      n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, 
      n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, 
      n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, 
      n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, 
      n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, 
      n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, 
      n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, 
      n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, 
      n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, 
      n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, 
      n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, 
      n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, 
      n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, 
      n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, 
      n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, 
      n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, 
      n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, 
      n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, 
      n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, 
      n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, 
      n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, 
      n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, 
      n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, 
      n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, 
      n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, 
      n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, 
      n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, 
      n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, 
      n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, 
      n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, 
      n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, 
      n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, 
      n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, 
      n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, 
      n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, 
      n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, 
      n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, 
      n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, 
      n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, 
      n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, 
      n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, 
      n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, 
      n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, 
      n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, 
      n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, 
      n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, 
      n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, 
      n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, 
      n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, 
      n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, 
      n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, 
      n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, 
      n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, 
      n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, 
      n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, 
      n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, 
      n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, 
      n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, 
      n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, 
      n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, 
      n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, 
      n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, 
      n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, 
      n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, 
      n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, 
      n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, 
      n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, 
      n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, 
      n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, 
      n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, 
      n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, 
      n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, 
      n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, 
      n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, 
      n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, 
      n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, 
      n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, 
      n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, 
      n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, 
      n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, 
      n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, 
      n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, 
      n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, 
      n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, 
      n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, 
      n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, 
      n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, 
      n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, 
      n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, 
      n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, 
      n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, 
      n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, 
      n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, 
      n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, 
      n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, 
      n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, 
      n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, 
      n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, 
      n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, 
      n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, 
      n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, 
      n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, 
      n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, 
      n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, 
      n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, 
      n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, 
      n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, 
      n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, 
      n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, 
      n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, 
      n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, 
      n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, 
      n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, 
      n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, 
      n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, 
      n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, 
      n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, 
      n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, 
      n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, 
      n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, 
      n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, 
      n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, 
      n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, 
      n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, 
      n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, 
      n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, 
      n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, 
      n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, 
      n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, 
      n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, 
      n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, 
      n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, 
      n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, 
      n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, 
      n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, 
      n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, 
      n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, 
      n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, 
      n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, 
      n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, 
      n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, 
      n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, 
      n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, 
      n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, 
      n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, 
      n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, 
      n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, 
      n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, 
      n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, 
      n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, 
      n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, 
      n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, 
      n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, 
      n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, 
      n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, 
      n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, 
      n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, 
      n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, 
      n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, 
      n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, 
      n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, 
      n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, 
      n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, 
      n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, 
      n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, 
      n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, 
      n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, 
      n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, 
      n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, 
      n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, 
      n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, 
      n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, 
      n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, 
      n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, 
      n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, 
      n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, 
      n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, 
      n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, 
      n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, 
      n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, 
      n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, 
      n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, 
      n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, 
      n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, 
      n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, 
      n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, 
      n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, 
      n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, 
      n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, 
      n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, 
      n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, 
      n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, 
      n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, 
      n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, 
      n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, 
      n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, 
      n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, 
      n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, 
      n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, 
      n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, 
      n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, 
      n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, 
      n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, 
      n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, 
      n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, 
      n9884, n9885, n9886, n9887, n9888, n9889, n9890, n_1000, n_1001, n_1002, 
      n_1003, n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, n_1011, 
      n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, 
      n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, 
      n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, 
      n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, 
      n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, 
      n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, 
      n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, 
      n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, 
      n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, 
      n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, 
      n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, 
      n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, 
      n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, 
      n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, 
      n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, 
      n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, 
      n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, 
      n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, 
      n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, 
      n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, 
      n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, 
      n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, 
      n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, 
      n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, 
      n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, 
      n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, 
      n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, 
      n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, 
      n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, 
      n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, 
      n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, 
      n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, 
      n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, 
      n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, 
      n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, 
      n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, 
      n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, 
      n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, 
      n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, 
      n_1363, n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, 
      n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, 
      n_1381, n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, 
      n_1390, n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, 
      n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, 
      n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, 
      n_1417, n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, 
      n_1426, n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, 
      n_1435, n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, 
      n_1444, n_1445, n_1446, n_1447 : std_logic;

begin
   
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n3609, CK => CLK, Q => 
                           n_1000, QN => n5);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n3608, CK => CLK, Q => 
                           n_1001, QN => n6);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n3607, CK => CLK, Q => 
                           n_1002, QN => n7);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n3606, CK => CLK, Q => 
                           n_1003, QN => n8);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n3605, CK => CLK, Q => 
                           n_1004, QN => n9);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n3569, CK => CLK, Q => 
                           n_1005, QN => n45);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n3568, CK => CLK, Q => 
                           n_1006, QN => n46);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n3567, CK => CLK, Q => 
                           n_1007, QN => n47);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n3566, CK => CLK, Q => 
                           n_1008, QN => n48);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n3565, CK => CLK, Q => 
                           n_1009, QN => n49);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n3564, CK => CLK, Q => 
                           n_1010, QN => n50);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n3563, CK => CLK, Q => 
                           n_1011, QN => n51);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n3562, CK => CLK, Q => 
                           n_1012, QN => n52);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n3561, CK => CLK, Q => 
                           n_1013, QN => n53);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n3560, CK => CLK, Q => 
                           n_1014, QN => n54);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n3559, CK => CLK, Q => n_1015
                           , QN => n55);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n3558, CK => CLK, Q => n_1016
                           , QN => n56);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n3557, CK => CLK, Q => n_1017
                           , QN => n57);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n3556, CK => CLK, Q => n_1018
                           , QN => n58);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n3555, CK => CLK, Q => n_1019
                           , QN => n59);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n3554, CK => CLK, Q => n_1020
                           , QN => n60);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n3553, CK => CLK, Q => n_1021
                           , QN => n61);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n3552, CK => CLK, Q => n_1022
                           , QN => n62);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n3551, CK => CLK, Q => n_1023
                           , QN => n63);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n3550, CK => CLK, Q => n_1024
                           , QN => n64);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n3420, CK => CLK, Q => 
                           n_1025, QN => n8833);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n3419, CK => CLK, Q => 
                           n_1026, QN => n8848);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n3418, CK => CLK, Q => 
                           n_1027, QN => n8863);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n3417, CK => CLK, Q => 
                           n_1028, QN => n8878);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n3416, CK => CLK, Q => 
                           n_1029, QN => n8893);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n3415, CK => CLK, Q => 
                           n_1030, QN => n8908);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n3414, CK => CLK, Q => 
                           n_1031, QN => n8923);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n3413, CK => CLK, Q => 
                           n_1032, QN => n8938);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n3412, CK => CLK, Q => 
                           n_1033, QN => n8953);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n3411, CK => CLK, Q => 
                           n_1034, QN => n8968);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n3410, CK => CLK, Q => 
                           n_1035, QN => n8983);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n3409, CK => CLK, Q => 
                           n_1036, QN => n8998);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n3408, CK => CLK, Q => 
                           n_1037, QN => n9013);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n3407, CK => CLK, Q => 
                           n_1038, QN => n9028);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n3406, CK => CLK, Q => 
                           n_1039, QN => n9043);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n3405, CK => CLK, Q => 
                           n_1040, QN => n9058);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n3404, CK => CLK, Q => 
                           n_1041, QN => n9073);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n3403, CK => CLK, Q => 
                           n_1042, QN => n9088);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n3402, CK => CLK, Q => 
                           n_1043, QN => n9103);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n3401, CK => CLK, Q => 
                           n_1044, QN => n9118);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n3400, CK => CLK, Q => 
                           n_1045, QN => n9133);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n3399, CK => CLK, Q => n_1046
                           , QN => n9148);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n3398, CK => CLK, Q => n_1047
                           , QN => n9163);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n3397, CK => CLK, Q => n_1048
                           , QN => n9178);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n3396, CK => CLK, Q => n_1049
                           , QN => n9193);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n3395, CK => CLK, Q => n_1050
                           , QN => n9208);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n3394, CK => CLK, Q => n_1051
                           , QN => n9223);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n3393, CK => CLK, Q => n_1052
                           , QN => n9238);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n3392, CK => CLK, Q => n_1053
                           , QN => n9253);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n3391, CK => CLK, Q => n_1054
                           , QN => n9268);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n3390, CK => CLK, Q => n_1055
                           , QN => n9283);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n3389, CK => CLK, Q => 
                           n_1056, QN => n8819);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n3388, CK => CLK, Q => 
                           n_1057, QN => n8834);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n3387, CK => CLK, Q => 
                           n_1058, QN => n8849);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n3386, CK => CLK, Q => 
                           n_1059, QN => n8864);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n3385, CK => CLK, Q => 
                           n_1060, QN => n8879);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n3384, CK => CLK, Q => 
                           n_1061, QN => n8894);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n3383, CK => CLK, Q => 
                           n_1062, QN => n8909);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n3382, CK => CLK, Q => 
                           n_1063, QN => n8924);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n3381, CK => CLK, Q => 
                           n_1064, QN => n8939);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n3380, CK => CLK, Q => 
                           n_1065, QN => n8954);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n3379, CK => CLK, Q => 
                           n_1066, QN => n8969);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n3378, CK => CLK, Q => 
                           n_1067, QN => n8984);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n3377, CK => CLK, Q => 
                           n_1068, QN => n8999);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n3376, CK => CLK, Q => 
                           n_1069, QN => n9014);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n3375, CK => CLK, Q => 
                           n_1070, QN => n9029);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n3374, CK => CLK, Q => 
                           n_1071, QN => n9044);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n3373, CK => CLK, Q => 
                           n_1072, QN => n9059);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n3372, CK => CLK, Q => 
                           n_1073, QN => n9074);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n3371, CK => CLK, Q => 
                           n_1074, QN => n9089);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n3370, CK => CLK, Q => 
                           n_1075, QN => n9104);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n3369, CK => CLK, Q => 
                           n_1076, QN => n9119);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n3368, CK => CLK, Q => 
                           n_1077, QN => n9134);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n3367, CK => CLK, Q => n_1078
                           , QN => n9149);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n3366, CK => CLK, Q => n_1079
                           , QN => n9164);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n3365, CK => CLK, Q => n_1080
                           , QN => n9179);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n3364, CK => CLK, Q => n_1081
                           , QN => n9194);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n3363, CK => CLK, Q => n_1082
                           , QN => n9209);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n3362, CK => CLK, Q => n_1083
                           , QN => n9224);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n3361, CK => CLK, Q => n_1084
                           , QN => n9239);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n3360, CK => CLK, Q => n_1085
                           , QN => n9254);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n3359, CK => CLK, Q => n_1086
                           , QN => n9269);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n3358, CK => CLK, Q => n_1087
                           , QN => n9284);
   OUT2_reg_31_inst : DFF_X1 port map( D => n2589, CK => CLK, Q => OUT2(31), QN
                           => n8783);
   OUT2_reg_30_inst : DFF_X1 port map( D => n2588, CK => CLK, Q => OUT2(30), QN
                           => n8784);
   OUT2_reg_29_inst : DFF_X1 port map( D => n2587, CK => CLK, Q => OUT2(29), QN
                           => n8785);
   OUT2_reg_28_inst : DFF_X1 port map( D => n2586, CK => CLK, Q => OUT2(28), QN
                           => n8786);
   OUT2_reg_27_inst : DFF_X1 port map( D => n2585, CK => CLK, Q => OUT2(27), QN
                           => n8787);
   OUT2_reg_26_inst : DFF_X1 port map( D => n2584, CK => CLK, Q => OUT2(26), QN
                           => n8788);
   OUT2_reg_25_inst : DFF_X1 port map( D => n2583, CK => CLK, Q => OUT2(25), QN
                           => n8789);
   OUT2_reg_24_inst : DFF_X1 port map( D => n2582, CK => CLK, Q => OUT2(24), QN
                           => n8790);
   OUT2_reg_23_inst : DFF_X1 port map( D => n2581, CK => CLK, Q => OUT2(23), QN
                           => n8791);
   OUT2_reg_22_inst : DFF_X1 port map( D => n2580, CK => CLK, Q => OUT2(22), QN
                           => n8792);
   OUT2_reg_21_inst : DFF_X1 port map( D => n2579, CK => CLK, Q => OUT2(21), QN
                           => n8793);
   OUT2_reg_20_inst : DFF_X1 port map( D => n2578, CK => CLK, Q => OUT2(20), QN
                           => n8794);
   OUT2_reg_19_inst : DFF_X1 port map( D => n2577, CK => CLK, Q => OUT2(19), QN
                           => n8795);
   OUT2_reg_18_inst : DFF_X1 port map( D => n2576, CK => CLK, Q => OUT2(18), QN
                           => n8796);
   OUT2_reg_17_inst : DFF_X1 port map( D => n2575, CK => CLK, Q => OUT2(17), QN
                           => n8797);
   OUT2_reg_16_inst : DFF_X1 port map( D => n2574, CK => CLK, Q => OUT2(16), QN
                           => n8798);
   OUT2_reg_15_inst : DFF_X1 port map( D => n2573, CK => CLK, Q => OUT2(15), QN
                           => n8799);
   OUT2_reg_14_inst : DFF_X1 port map( D => n2572, CK => CLK, Q => OUT2(14), QN
                           => n8800);
   OUT2_reg_13_inst : DFF_X1 port map( D => n2571, CK => CLK, Q => OUT2(13), QN
                           => n8801);
   OUT2_reg_12_inst : DFF_X1 port map( D => n2570, CK => CLK, Q => OUT2(12), QN
                           => n8802);
   OUT2_reg_11_inst : DFF_X1 port map( D => n2569, CK => CLK, Q => OUT2(11), QN
                           => n8803);
   OUT2_reg_10_inst : DFF_X1 port map( D => n2568, CK => CLK, Q => OUT2(10), QN
                           => n8804);
   OUT2_reg_9_inst : DFF_X1 port map( D => n2567, CK => CLK, Q => OUT2(9), QN 
                           => n8805);
   OUT2_reg_8_inst : DFF_X1 port map( D => n2566, CK => CLK, Q => OUT2(8), QN 
                           => n8806);
   OUT2_reg_7_inst : DFF_X1 port map( D => n2565, CK => CLK, Q => OUT2(7), QN 
                           => n8807);
   OUT2_reg_6_inst : DFF_X1 port map( D => n2564, CK => CLK, Q => OUT2(6), QN 
                           => n8808);
   OUT2_reg_5_inst : DFF_X1 port map( D => n2563, CK => CLK, Q => OUT2(5), QN 
                           => n8809);
   OUT2_reg_4_inst : DFF_X1 port map( D => n2562, CK => CLK, Q => OUT2(4), QN 
                           => n8810);
   OUT2_reg_3_inst : DFF_X1 port map( D => n2561, CK => CLK, Q => OUT2(3), QN 
                           => n8811);
   OUT2_reg_2_inst : DFF_X1 port map( D => n2560, CK => CLK, Q => OUT2(2), QN 
                           => n8812);
   OUT2_reg_1_inst : DFF_X1 port map( D => n2559, CK => CLK, Q => OUT2(1), QN 
                           => n8813);
   OUT2_reg_0_inst : DFF_X1 port map( D => n2558, CK => CLK, Q => OUT2(0), QN 
                           => n8814);
   OUT1_reg_31_inst : DFF_X1 port map( D => n2557, CK => CLK, Q => OUT1(31), QN
                           => n8815);
   OUT1_reg_30_inst : DFF_X1 port map( D => n2556, CK => CLK, Q => OUT1(30), QN
                           => n8830);
   OUT1_reg_29_inst : DFF_X1 port map( D => n2555, CK => CLK, Q => OUT1(29), QN
                           => n8845);
   OUT1_reg_28_inst : DFF_X1 port map( D => n2554, CK => CLK, Q => OUT1(28), QN
                           => n8860);
   OUT1_reg_27_inst : DFF_X1 port map( D => n2553, CK => CLK, Q => OUT1(27), QN
                           => n8875);
   OUT1_reg_26_inst : DFF_X1 port map( D => n2552, CK => CLK, Q => OUT1(26), QN
                           => n8890);
   OUT1_reg_25_inst : DFF_X1 port map( D => n2551, CK => CLK, Q => OUT1(25), QN
                           => n8905);
   OUT1_reg_24_inst : DFF_X1 port map( D => n2550, CK => CLK, Q => OUT1(24), QN
                           => n8920);
   OUT1_reg_23_inst : DFF_X1 port map( D => n2549, CK => CLK, Q => OUT1(23), QN
                           => n8935);
   OUT1_reg_22_inst : DFF_X1 port map( D => n2548, CK => CLK, Q => OUT1(22), QN
                           => n8950);
   OUT1_reg_21_inst : DFF_X1 port map( D => n2547, CK => CLK, Q => OUT1(21), QN
                           => n8965);
   OUT1_reg_20_inst : DFF_X1 port map( D => n2546, CK => CLK, Q => OUT1(20), QN
                           => n8980);
   OUT1_reg_19_inst : DFF_X1 port map( D => n2545, CK => CLK, Q => OUT1(19), QN
                           => n8995);
   OUT1_reg_18_inst : DFF_X1 port map( D => n2544, CK => CLK, Q => OUT1(18), QN
                           => n9010);
   OUT1_reg_17_inst : DFF_X1 port map( D => n2543, CK => CLK, Q => OUT1(17), QN
                           => n9025);
   OUT1_reg_16_inst : DFF_X1 port map( D => n2542, CK => CLK, Q => OUT1(16), QN
                           => n9040);
   OUT1_reg_15_inst : DFF_X1 port map( D => n2541, CK => CLK, Q => OUT1(15), QN
                           => n9055);
   OUT1_reg_14_inst : DFF_X1 port map( D => n2540, CK => CLK, Q => OUT1(14), QN
                           => n9070);
   OUT1_reg_13_inst : DFF_X1 port map( D => n2539, CK => CLK, Q => OUT1(13), QN
                           => n9085);
   OUT1_reg_12_inst : DFF_X1 port map( D => n2538, CK => CLK, Q => OUT1(12), QN
                           => n9100);
   OUT1_reg_11_inst : DFF_X1 port map( D => n2537, CK => CLK, Q => OUT1(11), QN
                           => n9115);
   OUT1_reg_10_inst : DFF_X1 port map( D => n2536, CK => CLK, Q => OUT1(10), QN
                           => n9130);
   OUT1_reg_9_inst : DFF_X1 port map( D => n2535, CK => CLK, Q => OUT1(9), QN 
                           => n9145);
   OUT1_reg_8_inst : DFF_X1 port map( D => n2534, CK => CLK, Q => OUT1(8), QN 
                           => n9160);
   OUT1_reg_7_inst : DFF_X1 port map( D => n2533, CK => CLK, Q => OUT1(7), QN 
                           => n9175);
   OUT1_reg_6_inst : DFF_X1 port map( D => n2532, CK => CLK, Q => OUT1(6), QN 
                           => n9190);
   OUT1_reg_5_inst : DFF_X1 port map( D => n2531, CK => CLK, Q => OUT1(5), QN 
                           => n9205);
   OUT1_reg_4_inst : DFF_X1 port map( D => n2530, CK => CLK, Q => OUT1(4), QN 
                           => n9220);
   OUT1_reg_3_inst : DFF_X1 port map( D => n2529, CK => CLK, Q => OUT1(3), QN 
                           => n9235);
   OUT1_reg_2_inst : DFF_X1 port map( D => n2528, CK => CLK, Q => OUT1(2), QN 
                           => n9250);
   OUT1_reg_1_inst : DFF_X1 port map( D => n2527, CK => CLK, Q => OUT1(1), QN 
                           => n9265);
   OUT1_reg_0_inst : DFF_X1 port map( D => n2526, CK => CLK, Q => OUT1(0), QN 
                           => n9280);
   U5968 : NAND3_X1 port map( A1 => n6453, A2 => n6452, A3 => n7449, ZN => 
                           n7433);
   U5969 : NAND3_X1 port map( A1 => n7449, A2 => n6452, A3 => ADD_WR(3), ZN => 
                           n7451);
   U5970 : NAND3_X1 port map( A1 => n7449, A2 => n6453, A3 => ADD_WR(4), ZN => 
                           n7460);
   U5971 : NAND3_X1 port map( A1 => n6455, A2 => n6454, A3 => n6456, ZN => 
                           n7434);
   U5972 : NAND3_X1 port map( A1 => n6455, A2 => n6454, A3 => ADD_WR(0), ZN => 
                           n7436);
   U5973 : NAND3_X1 port map( A1 => n6456, A2 => n6454, A3 => ADD_WR(1), ZN => 
                           n7438);
   U5974 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n6454, A3 => ADD_WR(1), ZN
                           => n7440);
   U5975 : NAND3_X1 port map( A1 => n6456, A2 => n6455, A3 => ADD_WR(2), ZN => 
                           n7442);
   U5976 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n6455, A3 => ADD_WR(2), ZN
                           => n7444);
   U5977 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => n6456, A3 => ADD_WR(2), ZN
                           => n7446);
   U5978 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => n7449, A3 => ADD_WR(4), ZN
                           => n7469);
   U5979 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), A3 => ADD_WR(2)
                           , ZN => n7448);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n2621, CK => CLK, Q => 
                           n7368, QN => n8828);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n2620, CK => CLK, Q => 
                           n7369, QN => n8843);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n2619, CK => CLK, Q => 
                           n7370, QN => n8858);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n2618, CK => CLK, Q => 
                           n7371, QN => n8873);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n2617, CK => CLK, Q => 
                           n7372, QN => n8888);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n2616, CK => CLK, Q => 
                           n7373, QN => n8903);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n2615, CK => CLK, Q => 
                           n7374, QN => n8918);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n2614, CK => CLK, Q => 
                           n7375, QN => n8933);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n2613, CK => CLK, Q => 
                           n7376, QN => n8948);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n2612, CK => CLK, Q => 
                           n7377, QN => n8963);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n2611, CK => CLK, Q => 
                           n7378, QN => n8978);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n2610, CK => CLK, Q => 
                           n7379, QN => n8993);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n2609, CK => CLK, Q => 
                           n7380, QN => n9008);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n2608, CK => CLK, Q => 
                           n7381, QN => n9023);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n2607, CK => CLK, Q => 
                           n7382, QN => n9038);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n2606, CK => CLK, Q => 
                           n7383, QN => n9053);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n2605, CK => CLK, Q => 
                           n7384, QN => n9068);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n2604, CK => CLK, Q => 
                           n7385, QN => n9083);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n2603, CK => CLK, Q => 
                           n7386, QN => n9098);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n2602, CK => CLK, Q => 
                           n7387, QN => n9113);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n2601, CK => CLK, Q => 
                           n7388, QN => n9128);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n2600, CK => CLK, Q => 
                           n7389, QN => n9143);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n2599, CK => CLK, Q => n7390
                           , QN => n9158);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n2598, CK => CLK, Q => n7391
                           , QN => n9173);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n2597, CK => CLK, Q => n7392
                           , QN => n9188);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n2596, CK => CLK, Q => n7393
                           , QN => n9203);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n2595, CK => CLK, Q => n7394
                           , QN => n9218);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n2594, CK => CLK, Q => n7395
                           , QN => n9233);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n2593, CK => CLK, Q => n7396
                           , QN => n9248);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n2592, CK => CLK, Q => n7397
                           , QN => n9263);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n2591, CK => CLK, Q => n7398
                           , QN => n9278);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n2590, CK => CLK, Q => n7399
                           , QN => n9293);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n2653, CK => CLK, Q => 
                           n7336, QN => n8829);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n2652, CK => CLK, Q => 
                           n7337, QN => n8844);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n2651, CK => CLK, Q => 
                           n7338, QN => n8859);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n2650, CK => CLK, Q => 
                           n7339, QN => n8874);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n2649, CK => CLK, Q => 
                           n7340, QN => n8889);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n2648, CK => CLK, Q => 
                           n7341, QN => n8904);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n2647, CK => CLK, Q => 
                           n7342, QN => n8919);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n2646, CK => CLK, Q => 
                           n7343, QN => n8934);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n2749, CK => CLK, Q => 
                           n7240, QN => n8826);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n2748, CK => CLK, Q => 
                           n7241, QN => n8841);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n2747, CK => CLK, Q => 
                           n7242, QN => n8856);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n2746, CK => CLK, Q => 
                           n7243, QN => n8871);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n2745, CK => CLK, Q => 
                           n7244, QN => n8886);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n2744, CK => CLK, Q => 
                           n7245, QN => n8901);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n2743, CK => CLK, Q => 
                           n7246, QN => n8916);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n2742, CK => CLK, Q => 
                           n7247, QN => n8931);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n2781, CK => CLK, Q => 
                           n7208, QN => n8827);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n2780, CK => CLK, Q => 
                           n7209, QN => n8842);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n2779, CK => CLK, Q => 
                           n7210, QN => n8857);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n2778, CK => CLK, Q => 
                           n7211, QN => n8872);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n2777, CK => CLK, Q => 
                           n7212, QN => n8887);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n2776, CK => CLK, Q => 
                           n7213, QN => n8902);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n2775, CK => CLK, Q => 
                           n7214, QN => n8917);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n2774, CK => CLK, Q => 
                           n7215, QN => n8932);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n2941, CK => CLK, Q => 
                           n7048, QN => n8824);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n2940, CK => CLK, Q => 
                           n7049, QN => n8839);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n2939, CK => CLK, Q => 
                           n7050, QN => n8854);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n2938, CK => CLK, Q => 
                           n7051, QN => n8869);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n2937, CK => CLK, Q => 
                           n7052, QN => n8884);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n2936, CK => CLK, Q => 
                           n7053, QN => n8899);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n2935, CK => CLK, Q => 
                           n7054, QN => n8914);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n2934, CK => CLK, Q => 
                           n7055, QN => n8929);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n2973, CK => CLK, Q => 
                           n7016, QN => n8825);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n2972, CK => CLK, Q => 
                           n7017, QN => n8840);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n2971, CK => CLK, Q => 
                           n7018, QN => n8855);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n2970, CK => CLK, Q => 
                           n7019, QN => n8870);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n2969, CK => CLK, Q => 
                           n7020, QN => n8885);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n2968, CK => CLK, Q => 
                           n7021, QN => n8900);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n2967, CK => CLK, Q => 
                           n7022, QN => n8915);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n2966, CK => CLK, Q => 
                           n7023, QN => n8930);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n3069, CK => CLK, Q => 
                           n6920, QN => n8822);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n3068, CK => CLK, Q => 
                           n6921, QN => n8837);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n3067, CK => CLK, Q => 
                           n6922, QN => n8852);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n3066, CK => CLK, Q => 
                           n6923, QN => n8867);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n3065, CK => CLK, Q => 
                           n6924, QN => n8882);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n3064, CK => CLK, Q => 
                           n6925, QN => n8897);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n3063, CK => CLK, Q => 
                           n6926, QN => n8912);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n3062, CK => CLK, Q => 
                           n6927, QN => n8927);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n3101, CK => CLK, Q => 
                           n6888, QN => n8823);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n3100, CK => CLK, Q => 
                           n6889, QN => n8838);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n3099, CK => CLK, Q => 
                           n6890, QN => n8853);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n3098, CK => CLK, Q => 
                           n6891, QN => n8868);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n3097, CK => CLK, Q => 
                           n6892, QN => n8883);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n3096, CK => CLK, Q => 
                           n6893, QN => n8898);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n3095, CK => CLK, Q => 
                           n6894, QN => n8913);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n3094, CK => CLK, Q => 
                           n6895, QN => n8928);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n3197, CK => CLK, Q => 
                           n6792, QN => n8820);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n3196, CK => CLK, Q => 
                           n6793, QN => n8835);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n3195, CK => CLK, Q => 
                           n6794, QN => n8850);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n3194, CK => CLK, Q => 
                           n6795, QN => n8865);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n3193, CK => CLK, Q => 
                           n6796, QN => n8880);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n3192, CK => CLK, Q => 
                           n6797, QN => n8895);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n3191, CK => CLK, Q => 
                           n6798, QN => n8910);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n3190, CK => CLK, Q => 
                           n6799, QN => n8925);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n3229, CK => CLK, Q => 
                           n6760, QN => n8821);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n3228, CK => CLK, Q => 
                           n6761, QN => n8836);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n3227, CK => CLK, Q => 
                           n6762, QN => n8851);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n3226, CK => CLK, Q => 
                           n6763, QN => n8866);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n3225, CK => CLK, Q => 
                           n6764, QN => n8881);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n3224, CK => CLK, Q => 
                           n6765, QN => n8896);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n3223, CK => CLK, Q => 
                           n6766, QN => n8911);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n3222, CK => CLK, Q => 
                           n6767, QN => n8926);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n3517, CK => CLK, Q => n6536
                           , QN => n8817);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n3516, CK => CLK, Q => n6537
                           , QN => n8832);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n3515, CK => CLK, Q => n6538
                           , QN => n8847);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n3514, CK => CLK, Q => n6539
                           , QN => n8862);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n3513, CK => CLK, Q => n6540
                           , QN => n8877);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n3512, CK => CLK, Q => n6541
                           , QN => n8892);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n3511, CK => CLK, Q => n6542
                           , QN => n8907);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n3510, CK => CLK, Q => n6543
                           , QN => n8922);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n3549, CK => CLK, Q => n6504
                           , QN => n8816);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n3548, CK => CLK, Q => n6505
                           , QN => n8831);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n3547, CK => CLK, Q => n6506
                           , QN => n8846);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n3546, CK => CLK, Q => n6507
                           , QN => n8861);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n3545, CK => CLK, Q => n6508
                           , QN => n8876);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n3544, CK => CLK, Q => n6509
                           , QN => n8891);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n3543, CK => CLK, Q => n6510
                           , QN => n8906);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n3542, CK => CLK, Q => n6511
                           , QN => n8921);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n2645, CK => CLK, Q => 
                           n7344, QN => n8949);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n2644, CK => CLK, Q => 
                           n7345, QN => n8964);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n2643, CK => CLK, Q => 
                           n7346, QN => n8979);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n2642, CK => CLK, Q => 
                           n7347, QN => n8994);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n2641, CK => CLK, Q => 
                           n7348, QN => n9009);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n2640, CK => CLK, Q => 
                           n7349, QN => n9024);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n2639, CK => CLK, Q => 
                           n7350, QN => n9039);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n2638, CK => CLK, Q => 
                           n7351, QN => n9054);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n2637, CK => CLK, Q => 
                           n7352, QN => n9069);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n2636, CK => CLK, Q => 
                           n7353, QN => n9084);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n2635, CK => CLK, Q => 
                           n7354, QN => n9099);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n2634, CK => CLK, Q => 
                           n7355, QN => n9114);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n2633, CK => CLK, Q => 
                           n7356, QN => n9129);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n2632, CK => CLK, Q => 
                           n7357, QN => n9144);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n2631, CK => CLK, Q => n7358
                           , QN => n9159);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n2630, CK => CLK, Q => n7359
                           , QN => n9174);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n2629, CK => CLK, Q => n7360
                           , QN => n9189);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n2628, CK => CLK, Q => n7361
                           , QN => n9204);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n2627, CK => CLK, Q => n7362
                           , QN => n9219);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n2626, CK => CLK, Q => n7363
                           , QN => n9234);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n2625, CK => CLK, Q => n7364
                           , QN => n9249);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n2624, CK => CLK, Q => n7365
                           , QN => n9264);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n2623, CK => CLK, Q => n7366
                           , QN => n9279);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n2622, CK => CLK, Q => n7367
                           , QN => n9294);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n2741, CK => CLK, Q => 
                           n7248, QN => n8946);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n2740, CK => CLK, Q => 
                           n7249, QN => n8961);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n2739, CK => CLK, Q => 
                           n7250, QN => n8976);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n2738, CK => CLK, Q => 
                           n7251, QN => n8991);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n2737, CK => CLK, Q => 
                           n7252, QN => n9006);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n2736, CK => CLK, Q => 
                           n7253, QN => n9021);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n2735, CK => CLK, Q => 
                           n7254, QN => n9036);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n2734, CK => CLK, Q => 
                           n7255, QN => n9051);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n2733, CK => CLK, Q => 
                           n7256, QN => n9066);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n2732, CK => CLK, Q => 
                           n7257, QN => n9081);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n2731, CK => CLK, Q => 
                           n7258, QN => n9096);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n2730, CK => CLK, Q => 
                           n7259, QN => n9111);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n2729, CK => CLK, Q => 
                           n7260, QN => n9126);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n2728, CK => CLK, Q => 
                           n7261, QN => n9141);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n2727, CK => CLK, Q => n7262
                           , QN => n9156);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n2726, CK => CLK, Q => n7263
                           , QN => n9171);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n2725, CK => CLK, Q => n7264
                           , QN => n9186);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n2724, CK => CLK, Q => n7265
                           , QN => n9201);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n2723, CK => CLK, Q => n7266
                           , QN => n9216);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n2722, CK => CLK, Q => n7267
                           , QN => n9231);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n2721, CK => CLK, Q => n7268
                           , QN => n9246);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n2720, CK => CLK, Q => n7269
                           , QN => n9261);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n2719, CK => CLK, Q => n7270
                           , QN => n9276);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n2718, CK => CLK, Q => n7271
                           , QN => n9291);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n2773, CK => CLK, Q => 
                           n7216, QN => n8947);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n2772, CK => CLK, Q => 
                           n7217, QN => n8962);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n2771, CK => CLK, Q => 
                           n7218, QN => n8977);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n2770, CK => CLK, Q => 
                           n7219, QN => n8992);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n2769, CK => CLK, Q => 
                           n7220, QN => n9007);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n2768, CK => CLK, Q => 
                           n7221, QN => n9022);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n2767, CK => CLK, Q => 
                           n7222, QN => n9037);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n2766, CK => CLK, Q => 
                           n7223, QN => n9052);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n2765, CK => CLK, Q => 
                           n7224, QN => n9067);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n2764, CK => CLK, Q => 
                           n7225, QN => n9082);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n2763, CK => CLK, Q => 
                           n7226, QN => n9097);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n2762, CK => CLK, Q => 
                           n7227, QN => n9112);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n2761, CK => CLK, Q => 
                           n7228, QN => n9127);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n2760, CK => CLK, Q => 
                           n7229, QN => n9142);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n2759, CK => CLK, Q => n7230
                           , QN => n9157);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n2758, CK => CLK, Q => n7231
                           , QN => n9172);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n2757, CK => CLK, Q => n7232
                           , QN => n9187);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n2756, CK => CLK, Q => n7233
                           , QN => n9202);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n2755, CK => CLK, Q => n7234
                           , QN => n9217);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n2754, CK => CLK, Q => n7235
                           , QN => n9232);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n2753, CK => CLK, Q => n7236
                           , QN => n9247);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n2752, CK => CLK, Q => n7237
                           , QN => n9262);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n2751, CK => CLK, Q => n7238
                           , QN => n9277);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n2750, CK => CLK, Q => n7239
                           , QN => n9292);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n2933, CK => CLK, Q => 
                           n7056, QN => n8944);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n2932, CK => CLK, Q => 
                           n7057, QN => n8959);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n2931, CK => CLK, Q => 
                           n7058, QN => n8974);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n2930, CK => CLK, Q => 
                           n7059, QN => n8989);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n2929, CK => CLK, Q => 
                           n7060, QN => n9004);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n2928, CK => CLK, Q => 
                           n7061, QN => n9019);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n2927, CK => CLK, Q => 
                           n7062, QN => n9034);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n2926, CK => CLK, Q => 
                           n7063, QN => n9049);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n2925, CK => CLK, Q => 
                           n7064, QN => n9064);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n2924, CK => CLK, Q => 
                           n7065, QN => n9079);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n2923, CK => CLK, Q => 
                           n7066, QN => n9094);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n2922, CK => CLK, Q => 
                           n7067, QN => n9109);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n2921, CK => CLK, Q => 
                           n7068, QN => n9124);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n2920, CK => CLK, Q => 
                           n7069, QN => n9139);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n2919, CK => CLK, Q => n7070
                           , QN => n9154);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n2918, CK => CLK, Q => n7071
                           , QN => n9169);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n2917, CK => CLK, Q => n7072
                           , QN => n9184);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n2916, CK => CLK, Q => n7073
                           , QN => n9199);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n2915, CK => CLK, Q => n7074
                           , QN => n9214);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n2914, CK => CLK, Q => n7075
                           , QN => n9229);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n2913, CK => CLK, Q => n7076
                           , QN => n9244);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n2912, CK => CLK, Q => n7077
                           , QN => n9259);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n2911, CK => CLK, Q => n7078
                           , QN => n9274);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n2910, CK => CLK, Q => n7079
                           , QN => n9289);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n2965, CK => CLK, Q => 
                           n7024, QN => n8945);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n2964, CK => CLK, Q => 
                           n7025, QN => n8960);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n2963, CK => CLK, Q => 
                           n7026, QN => n8975);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n2962, CK => CLK, Q => 
                           n7027, QN => n8990);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n2961, CK => CLK, Q => 
                           n7028, QN => n9005);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n2960, CK => CLK, Q => 
                           n7029, QN => n9020);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n2959, CK => CLK, Q => 
                           n7030, QN => n9035);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n2958, CK => CLK, Q => 
                           n7031, QN => n9050);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n2957, CK => CLK, Q => 
                           n7032, QN => n9065);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n2956, CK => CLK, Q => 
                           n7033, QN => n9080);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n2955, CK => CLK, Q => 
                           n7034, QN => n9095);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n2954, CK => CLK, Q => 
                           n7035, QN => n9110);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n2953, CK => CLK, Q => 
                           n7036, QN => n9125);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n2952, CK => CLK, Q => 
                           n7037, QN => n9140);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n2951, CK => CLK, Q => n7038
                           , QN => n9155);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n2950, CK => CLK, Q => n7039
                           , QN => n9170);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n2949, CK => CLK, Q => n7040
                           , QN => n9185);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n2948, CK => CLK, Q => n7041
                           , QN => n9200);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n2947, CK => CLK, Q => n7042
                           , QN => n9215);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n2946, CK => CLK, Q => n7043
                           , QN => n9230);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n2945, CK => CLK, Q => n7044
                           , QN => n9245);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n2944, CK => CLK, Q => n7045
                           , QN => n9260);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n2943, CK => CLK, Q => n7046
                           , QN => n9275);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n2942, CK => CLK, Q => n7047
                           , QN => n9290);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n3061, CK => CLK, Q => 
                           n6928, QN => n8942);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n3060, CK => CLK, Q => 
                           n6929, QN => n8957);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n3059, CK => CLK, Q => 
                           n6930, QN => n8972);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n3058, CK => CLK, Q => 
                           n6931, QN => n8987);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n3057, CK => CLK, Q => 
                           n6932, QN => n9002);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n3056, CK => CLK, Q => 
                           n6933, QN => n9017);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n3055, CK => CLK, Q => 
                           n6934, QN => n9032);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n3054, CK => CLK, Q => 
                           n6935, QN => n9047);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n3053, CK => CLK, Q => 
                           n6936, QN => n9062);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n3052, CK => CLK, Q => 
                           n6937, QN => n9077);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n3051, CK => CLK, Q => 
                           n6938, QN => n9092);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n3050, CK => CLK, Q => 
                           n6939, QN => n9107);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n3049, CK => CLK, Q => 
                           n6940, QN => n9122);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n3048, CK => CLK, Q => 
                           n6941, QN => n9137);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n3047, CK => CLK, Q => n6942
                           , QN => n9152);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n3046, CK => CLK, Q => n6943
                           , QN => n9167);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n3045, CK => CLK, Q => n6944
                           , QN => n9182);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n3044, CK => CLK, Q => n6945
                           , QN => n9197);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n3043, CK => CLK, Q => n6946
                           , QN => n9212);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n3042, CK => CLK, Q => n6947
                           , QN => n9227);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n3041, CK => CLK, Q => n6948
                           , QN => n9242);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n3040, CK => CLK, Q => n6949
                           , QN => n9257);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n3039, CK => CLK, Q => n6950
                           , QN => n9272);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n3038, CK => CLK, Q => n6951
                           , QN => n9287);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n3093, CK => CLK, Q => 
                           n6896, QN => n8943);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n3092, CK => CLK, Q => 
                           n6897, QN => n8958);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n3091, CK => CLK, Q => 
                           n6898, QN => n8973);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n3090, CK => CLK, Q => 
                           n6899, QN => n8988);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n3089, CK => CLK, Q => 
                           n6900, QN => n9003);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n3088, CK => CLK, Q => 
                           n6901, QN => n9018);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n3087, CK => CLK, Q => 
                           n6902, QN => n9033);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n3086, CK => CLK, Q => 
                           n6903, QN => n9048);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n3085, CK => CLK, Q => 
                           n6904, QN => n9063);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n3084, CK => CLK, Q => 
                           n6905, QN => n9078);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n3083, CK => CLK, Q => 
                           n6906, QN => n9093);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n3082, CK => CLK, Q => 
                           n6907, QN => n9108);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n3081, CK => CLK, Q => 
                           n6908, QN => n9123);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n3080, CK => CLK, Q => 
                           n6909, QN => n9138);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n3079, CK => CLK, Q => n6910
                           , QN => n9153);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n3078, CK => CLK, Q => n6911
                           , QN => n9168);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n3077, CK => CLK, Q => n6912
                           , QN => n9183);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n3076, CK => CLK, Q => n6913
                           , QN => n9198);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n3075, CK => CLK, Q => n6914
                           , QN => n9213);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n3074, CK => CLK, Q => n6915
                           , QN => n9228);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n3073, CK => CLK, Q => n6916
                           , QN => n9243);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n3072, CK => CLK, Q => n6917
                           , QN => n9258);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n3071, CK => CLK, Q => n6918
                           , QN => n9273);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n3070, CK => CLK, Q => n6919
                           , QN => n9288);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n3189, CK => CLK, Q => 
                           n6800, QN => n8940);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n3188, CK => CLK, Q => 
                           n6801, QN => n8955);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n3187, CK => CLK, Q => 
                           n6802, QN => n8970);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n3186, CK => CLK, Q => 
                           n6803, QN => n8985);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n3185, CK => CLK, Q => 
                           n6804, QN => n9000);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n3184, CK => CLK, Q => 
                           n6805, QN => n9015);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n3183, CK => CLK, Q => 
                           n6806, QN => n9030);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n3182, CK => CLK, Q => 
                           n6807, QN => n9045);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n3181, CK => CLK, Q => 
                           n6808, QN => n9060);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n3180, CK => CLK, Q => 
                           n6809, QN => n9075);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n3179, CK => CLK, Q => 
                           n6810, QN => n9090);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n3178, CK => CLK, Q => 
                           n6811, QN => n9105);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n3177, CK => CLK, Q => 
                           n6812, QN => n9120);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n3176, CK => CLK, Q => 
                           n6813, QN => n9135);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n3175, CK => CLK, Q => n6814
                           , QN => n9150);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n3174, CK => CLK, Q => n6815
                           , QN => n9165);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n3173, CK => CLK, Q => n6816
                           , QN => n9180);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n3172, CK => CLK, Q => n6817
                           , QN => n9195);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n3171, CK => CLK, Q => n6818
                           , QN => n9210);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n3170, CK => CLK, Q => n6819
                           , QN => n9225);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n3169, CK => CLK, Q => n6820
                           , QN => n9240);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n3168, CK => CLK, Q => n6821
                           , QN => n9255);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n3167, CK => CLK, Q => n6822
                           , QN => n9270);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n3166, CK => CLK, Q => n6823
                           , QN => n9285);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n3221, CK => CLK, Q => 
                           n6768, QN => n8941);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n3220, CK => CLK, Q => 
                           n6769, QN => n8956);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n3219, CK => CLK, Q => 
                           n6770, QN => n8971);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n3218, CK => CLK, Q => 
                           n6771, QN => n8986);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n3217, CK => CLK, Q => 
                           n6772, QN => n9001);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n3216, CK => CLK, Q => 
                           n6773, QN => n9016);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n3215, CK => CLK, Q => 
                           n6774, QN => n9031);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n3214, CK => CLK, Q => 
                           n6775, QN => n9046);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n3213, CK => CLK, Q => 
                           n6776, QN => n9061);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n3212, CK => CLK, Q => 
                           n6777, QN => n9076);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n3211, CK => CLK, Q => 
                           n6778, QN => n9091);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n3210, CK => CLK, Q => 
                           n6779, QN => n9106);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n3209, CK => CLK, Q => 
                           n6780, QN => n9121);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n3208, CK => CLK, Q => 
                           n6781, QN => n9136);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n3207, CK => CLK, Q => n6782
                           , QN => n9151);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n3206, CK => CLK, Q => n6783
                           , QN => n9166);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n3205, CK => CLK, Q => n6784
                           , QN => n9181);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n3204, CK => CLK, Q => n6785
                           , QN => n9196);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n3203, CK => CLK, Q => n6786
                           , QN => n9211);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n3202, CK => CLK, Q => n6787
                           , QN => n9226);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n3201, CK => CLK, Q => n6788
                           , QN => n9241);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n3200, CK => CLK, Q => n6789
                           , QN => n9256);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n3199, CK => CLK, Q => n6790
                           , QN => n9271);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n3198, CK => CLK, Q => n6791
                           , QN => n9286);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n3509, CK => CLK, Q => n6544
                           , QN => n8937);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n3508, CK => CLK, Q => n6545
                           , QN => n8952);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n3507, CK => CLK, Q => n6546
                           , QN => n8967);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n3506, CK => CLK, Q => n6547
                           , QN => n8982);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n3505, CK => CLK, Q => n6548
                           , QN => n8997);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n3504, CK => CLK, Q => n6549
                           , QN => n9012);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n3503, CK => CLK, Q => n6550
                           , QN => n9027);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n3502, CK => CLK, Q => n6551
                           , QN => n9042);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n3501, CK => CLK, Q => n6552
                           , QN => n9057);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n3500, CK => CLK, Q => n6553
                           , QN => n9072);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n3499, CK => CLK, Q => n6554
                           , QN => n9087);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n3498, CK => CLK, Q => n6555
                           , QN => n9102);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n3497, CK => CLK, Q => n6556
                           , QN => n9117);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n3496, CK => CLK, Q => n6557
                           , QN => n9132);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n3495, CK => CLK, Q => n6558,
                           QN => n9147);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n3494, CK => CLK, Q => n6559,
                           QN => n9162);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n3493, CK => CLK, Q => n6560,
                           QN => n9177);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n3492, CK => CLK, Q => n6561,
                           QN => n9192);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n3491, CK => CLK, Q => n6562,
                           QN => n9207);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n3490, CK => CLK, Q => n6563,
                           QN => n9222);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n3489, CK => CLK, Q => n6564,
                           QN => n9237);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n3488, CK => CLK, Q => n6565,
                           QN => n9252);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n3487, CK => CLK, Q => n6566,
                           QN => n9267);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n3486, CK => CLK, Q => n6567,
                           QN => n9282);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n3541, CK => CLK, Q => n6512
                           , QN => n8936);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n3540, CK => CLK, Q => n6513
                           , QN => n8951);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n3539, CK => CLK, Q => n6514
                           , QN => n8966);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n3538, CK => CLK, Q => n6515
                           , QN => n8981);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n3537, CK => CLK, Q => n6516
                           , QN => n8996);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n3536, CK => CLK, Q => n6517
                           , QN => n9011);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n3535, CK => CLK, Q => n6518
                           , QN => n9026);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n3534, CK => CLK, Q => n6519
                           , QN => n9041);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n3533, CK => CLK, Q => n6520
                           , QN => n9056);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n3532, CK => CLK, Q => n6521
                           , QN => n9071);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n3531, CK => CLK, Q => n6522
                           , QN => n9086);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n3530, CK => CLK, Q => n6523
                           , QN => n9101);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n3529, CK => CLK, Q => n6524
                           , QN => n9116);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n3528, CK => CLK, Q => n6525
                           , QN => n9131);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n3527, CK => CLK, Q => n6526,
                           QN => n9146);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n3526, CK => CLK, Q => n6527,
                           QN => n9161);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n3525, CK => CLK, Q => n6528,
                           QN => n9176);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n3524, CK => CLK, Q => n6529,
                           QN => n9191);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n3523, CK => CLK, Q => n6530,
                           QN => n9206);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n3522, CK => CLK, Q => n6531,
                           QN => n9221);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n3521, CK => CLK, Q => n6532,
                           QN => n9236);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n3520, CK => CLK, Q => n6533,
                           QN => n9251);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n3519, CK => CLK, Q => n6534,
                           QN => n9266);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n3518, CK => CLK, Q => n6535,
                           QN => n9281);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n3421, CK => CLK, Q => 
                           n_1088, QN => n8818);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n3589, CK => CLK, Q => n_1089
                           , QN => n6484);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n3588, CK => CLK, Q => n_1090
                           , QN => n6485);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n3587, CK => CLK, Q => n_1091
                           , QN => n6486);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n3586, CK => CLK, Q => n_1092
                           , QN => n6487);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n3585, CK => CLK, Q => n_1093
                           , QN => n6488);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n3584, CK => CLK, Q => n_1094
                           , QN => n6489);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n3583, CK => CLK, Q => n_1095
                           , QN => n6490);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n2717, CK => CLK, Q => 
                           n_1096, QN => n7272);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n2716, CK => CLK, Q => 
                           n_1097, QN => n7273);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n2715, CK => CLK, Q => 
                           n_1098, QN => n7274);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n2714, CK => CLK, Q => 
                           n_1099, QN => n7275);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n2713, CK => CLK, Q => 
                           n_1100, QN => n7276);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n2712, CK => CLK, Q => 
                           n_1101, QN => n7277);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n2711, CK => CLK, Q => 
                           n_1102, QN => n7278);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n2710, CK => CLK, Q => 
                           n_1103, QN => n7279);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n2845, CK => CLK, Q => 
                           n_1104, QN => n7144);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n2844, CK => CLK, Q => 
                           n_1105, QN => n7145);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n2843, CK => CLK, Q => 
                           n_1106, QN => n7146);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n2842, CK => CLK, Q => 
                           n_1107, QN => n7147);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n2841, CK => CLK, Q => 
                           n_1108, QN => n7148);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n2840, CK => CLK, Q => 
                           n_1109, QN => n7149);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n2839, CK => CLK, Q => 
                           n_1110, QN => n7150);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n2838, CK => CLK, Q => 
                           n_1111, QN => n7151);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n2909, CK => CLK, Q => 
                           n_1112, QN => n7080);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n2908, CK => CLK, Q => 
                           n_1113, QN => n7081);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n2907, CK => CLK, Q => 
                           n_1114, QN => n7082);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n2906, CK => CLK, Q => 
                           n_1115, QN => n7083);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n2905, CK => CLK, Q => 
                           n_1116, QN => n7084);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n2904, CK => CLK, Q => 
                           n_1117, QN => n7085);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n2903, CK => CLK, Q => 
                           n_1118, QN => n7086);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n2902, CK => CLK, Q => 
                           n_1119, QN => n7087);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n3037, CK => CLK, Q => 
                           n_1120, QN => n6952);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n3036, CK => CLK, Q => 
                           n_1121, QN => n6953);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n3035, CK => CLK, Q => 
                           n_1122, QN => n6954);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n3034, CK => CLK, Q => 
                           n_1123, QN => n6955);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n3033, CK => CLK, Q => 
                           n_1124, QN => n6956);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n3032, CK => CLK, Q => 
                           n_1125, QN => n6957);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n3031, CK => CLK, Q => 
                           n_1126, QN => n6958);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n3030, CK => CLK, Q => 
                           n_1127, QN => n6959);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n3165, CK => CLK, Q => 
                           n_1128, QN => n6824);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n3164, CK => CLK, Q => 
                           n_1129, QN => n6825);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n3163, CK => CLK, Q => 
                           n_1130, QN => n6826);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n3162, CK => CLK, Q => 
                           n_1131, QN => n6827);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n3161, CK => CLK, Q => 
                           n_1132, QN => n6828);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n3160, CK => CLK, Q => 
                           n_1133, QN => n6829);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n3159, CK => CLK, Q => 
                           n_1134, QN => n6830);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n3158, CK => CLK, Q => 
                           n_1135, QN => n6831);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n3581, CK => CLK, Q => 
                           n_1136, QN => n6492);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n3580, CK => CLK, Q => 
                           n_1137, QN => n6493);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n3579, CK => CLK, Q => 
                           n_1138, QN => n6494);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n3578, CK => CLK, Q => 
                           n_1139, QN => n6495);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n3577, CK => CLK, Q => 
                           n_1140, QN => n6496);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n3576, CK => CLK, Q => 
                           n_1141, QN => n6497);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n3575, CK => CLK, Q => 
                           n_1142, QN => n6498);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n3574, CK => CLK, Q => 
                           n_1143, QN => n6499);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n2685, CK => CLK, Q => 
                           n_1144, QN => n7304);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n2684, CK => CLK, Q => 
                           n_1145, QN => n7305);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n2683, CK => CLK, Q => 
                           n_1146, QN => n7306);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n2682, CK => CLK, Q => 
                           n_1147, QN => n7307);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n2681, CK => CLK, Q => 
                           n_1148, QN => n7308);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n2680, CK => CLK, Q => 
                           n_1149, QN => n7309);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n2679, CK => CLK, Q => 
                           n_1150, QN => n7310);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n2678, CK => CLK, Q => 
                           n_1151, QN => n7311);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n2813, CK => CLK, Q => 
                           n_1152, QN => n7176);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n2812, CK => CLK, Q => 
                           n_1153, QN => n7177);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n2811, CK => CLK, Q => 
                           n_1154, QN => n7178);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n2810, CK => CLK, Q => 
                           n_1155, QN => n7179);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n2809, CK => CLK, Q => 
                           n_1156, QN => n7180);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n2808, CK => CLK, Q => 
                           n_1157, QN => n7181);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n2807, CK => CLK, Q => 
                           n_1158, QN => n7182);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n2806, CK => CLK, Q => 
                           n_1159, QN => n7183);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n2877, CK => CLK, Q => 
                           n_1160, QN => n7112);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n2876, CK => CLK, Q => 
                           n_1161, QN => n7113);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n2875, CK => CLK, Q => 
                           n_1162, QN => n7114);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n2874, CK => CLK, Q => 
                           n_1163, QN => n7115);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n2873, CK => CLK, Q => 
                           n_1164, QN => n7116);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n2872, CK => CLK, Q => 
                           n_1165, QN => n7117);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n2871, CK => CLK, Q => 
                           n_1166, QN => n7118);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n2870, CK => CLK, Q => 
                           n_1167, QN => n7119);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n3005, CK => CLK, Q => 
                           n_1168, QN => n6984);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n3004, CK => CLK, Q => 
                           n_1169, QN => n6985);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n3003, CK => CLK, Q => 
                           n_1170, QN => n6986);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n3002, CK => CLK, Q => 
                           n_1171, QN => n6987);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n3001, CK => CLK, Q => 
                           n_1172, QN => n6988);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n3000, CK => CLK, Q => 
                           n_1173, QN => n6989);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n2999, CK => CLK, Q => 
                           n_1174, QN => n6990);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n2998, CK => CLK, Q => 
                           n_1175, QN => n6991);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n3133, CK => CLK, Q => 
                           n_1176, QN => n6856);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n3132, CK => CLK, Q => 
                           n_1177, QN => n6857);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n3131, CK => CLK, Q => 
                           n_1178, QN => n6858);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n3130, CK => CLK, Q => 
                           n_1179, QN => n6859);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n3129, CK => CLK, Q => 
                           n_1180, QN => n6860);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n3128, CK => CLK, Q => 
                           n_1181, QN => n6861);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n3127, CK => CLK, Q => 
                           n_1182, QN => n6862);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n3126, CK => CLK, Q => 
                           n_1183, QN => n6863);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n3573, CK => CLK, Q => 
                           n_1184, QN => n6500);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n3572, CK => CLK, Q => 
                           n_1185, QN => n6501);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n3571, CK => CLK, Q => 
                           n_1186, QN => n6502);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n3570, CK => CLK, Q => 
                           n_1187, QN => n6503);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n2709, CK => CLK, Q => 
                           n_1188, QN => n7280);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n2708, CK => CLK, Q => 
                           n_1189, QN => n7281);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n2707, CK => CLK, Q => 
                           n_1190, QN => n7282);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n2706, CK => CLK, Q => 
                           n_1191, QN => n7283);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n2705, CK => CLK, Q => 
                           n_1192, QN => n7284);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n2704, CK => CLK, Q => 
                           n_1193, QN => n7285);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n2703, CK => CLK, Q => 
                           n_1194, QN => n7286);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n2702, CK => CLK, Q => 
                           n_1195, QN => n7287);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n2701, CK => CLK, Q => 
                           n_1196, QN => n7288);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n2700, CK => CLK, Q => 
                           n_1197, QN => n7289);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n2699, CK => CLK, Q => 
                           n_1198, QN => n7290);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n2698, CK => CLK, Q => 
                           n_1199, QN => n7291);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n2697, CK => CLK, Q => 
                           n_1200, QN => n7292);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n2696, CK => CLK, Q => 
                           n_1201, QN => n7293);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n2695, CK => CLK, Q => 
                           n_1202, QN => n7294);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n2694, CK => CLK, Q => 
                           n_1203, QN => n7295);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n2693, CK => CLK, Q => 
                           n_1204, QN => n7296);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n2692, CK => CLK, Q => 
                           n_1205, QN => n7297);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n2691, CK => CLK, Q => 
                           n_1206, QN => n7298);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n2690, CK => CLK, Q => 
                           n_1207, QN => n7299);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n2689, CK => CLK, Q => 
                           n_1208, QN => n7300);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n2688, CK => CLK, Q => 
                           n_1209, QN => n7301);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n2687, CK => CLK, Q => 
                           n_1210, QN => n7302);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n2686, CK => CLK, Q => 
                           n_1211, QN => n7303);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n2837, CK => CLK, Q => 
                           n_1212, QN => n7152);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n2836, CK => CLK, Q => 
                           n_1213, QN => n7153);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n2835, CK => CLK, Q => 
                           n_1214, QN => n7154);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n2834, CK => CLK, Q => 
                           n_1215, QN => n7155);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n2833, CK => CLK, Q => 
                           n_1216, QN => n7156);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n2832, CK => CLK, Q => 
                           n_1217, QN => n7157);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n2831, CK => CLK, Q => 
                           n_1218, QN => n7158);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n2830, CK => CLK, Q => 
                           n_1219, QN => n7159);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n2829, CK => CLK, Q => 
                           n_1220, QN => n7160);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n2828, CK => CLK, Q => 
                           n_1221, QN => n7161);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n2827, CK => CLK, Q => 
                           n_1222, QN => n7162);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n2826, CK => CLK, Q => 
                           n_1223, QN => n7163);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n2825, CK => CLK, Q => 
                           n_1224, QN => n7164);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n2824, CK => CLK, Q => 
                           n_1225, QN => n7165);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n2823, CK => CLK, Q => 
                           n_1226, QN => n7166);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n2822, CK => CLK, Q => 
                           n_1227, QN => n7167);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n2821, CK => CLK, Q => 
                           n_1228, QN => n7168);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n2820, CK => CLK, Q => 
                           n_1229, QN => n7169);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n2819, CK => CLK, Q => 
                           n_1230, QN => n7170);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n2818, CK => CLK, Q => 
                           n_1231, QN => n7171);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n2817, CK => CLK, Q => 
                           n_1232, QN => n7172);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n2816, CK => CLK, Q => 
                           n_1233, QN => n7173);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n2815, CK => CLK, Q => 
                           n_1234, QN => n7174);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n2814, CK => CLK, Q => 
                           n_1235, QN => n7175);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n2901, CK => CLK, Q => 
                           n_1236, QN => n7088);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n2900, CK => CLK, Q => 
                           n_1237, QN => n7089);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n2899, CK => CLK, Q => 
                           n_1238, QN => n7090);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n2898, CK => CLK, Q => 
                           n_1239, QN => n7091);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n2897, CK => CLK, Q => 
                           n_1240, QN => n7092);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n2896, CK => CLK, Q => 
                           n_1241, QN => n7093);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n2895, CK => CLK, Q => 
                           n_1242, QN => n7094);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n2894, CK => CLK, Q => 
                           n_1243, QN => n7095);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n2893, CK => CLK, Q => 
                           n_1244, QN => n7096);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n2892, CK => CLK, Q => 
                           n_1245, QN => n7097);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n2891, CK => CLK, Q => 
                           n_1246, QN => n7098);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n2890, CK => CLK, Q => 
                           n_1247, QN => n7099);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n2889, CK => CLK, Q => 
                           n_1248, QN => n7100);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n2888, CK => CLK, Q => 
                           n_1249, QN => n7101);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n2887, CK => CLK, Q => 
                           n_1250, QN => n7102);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n2886, CK => CLK, Q => 
                           n_1251, QN => n7103);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n2885, CK => CLK, Q => 
                           n_1252, QN => n7104);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n2884, CK => CLK, Q => 
                           n_1253, QN => n7105);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n2883, CK => CLK, Q => 
                           n_1254, QN => n7106);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n2882, CK => CLK, Q => 
                           n_1255, QN => n7107);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n2881, CK => CLK, Q => 
                           n_1256, QN => n7108);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n2880, CK => CLK, Q => 
                           n_1257, QN => n7109);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n2879, CK => CLK, Q => 
                           n_1258, QN => n7110);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n2878, CK => CLK, Q => 
                           n_1259, QN => n7111);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n3029, CK => CLK, Q => 
                           n_1260, QN => n6960);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n3028, CK => CLK, Q => 
                           n_1261, QN => n6961);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n3027, CK => CLK, Q => 
                           n_1262, QN => n6962);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n3026, CK => CLK, Q => 
                           n_1263, QN => n6963);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n3025, CK => CLK, Q => 
                           n_1264, QN => n6964);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n3024, CK => CLK, Q => 
                           n_1265, QN => n6965);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n3023, CK => CLK, Q => 
                           n_1266, QN => n6966);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n3022, CK => CLK, Q => 
                           n_1267, QN => n6967);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n3021, CK => CLK, Q => 
                           n_1268, QN => n6968);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n3020, CK => CLK, Q => 
                           n_1269, QN => n6969);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n3019, CK => CLK, Q => 
                           n_1270, QN => n6970);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n3018, CK => CLK, Q => 
                           n_1271, QN => n6971);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n3017, CK => CLK, Q => 
                           n_1272, QN => n6972);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n3016, CK => CLK, Q => 
                           n_1273, QN => n6973);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n3015, CK => CLK, Q => 
                           n_1274, QN => n6974);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n3014, CK => CLK, Q => 
                           n_1275, QN => n6975);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n3013, CK => CLK, Q => 
                           n_1276, QN => n6976);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n3012, CK => CLK, Q => 
                           n_1277, QN => n6977);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n3011, CK => CLK, Q => 
                           n_1278, QN => n6978);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n3010, CK => CLK, Q => 
                           n_1279, QN => n6979);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n3009, CK => CLK, Q => 
                           n_1280, QN => n6980);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n3008, CK => CLK, Q => 
                           n_1281, QN => n6981);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n3007, CK => CLK, Q => 
                           n_1282, QN => n6982);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n3006, CK => CLK, Q => 
                           n_1283, QN => n6983);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n3157, CK => CLK, Q => 
                           n_1284, QN => n6832);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n3156, CK => CLK, Q => 
                           n_1285, QN => n6833);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n3155, CK => CLK, Q => 
                           n_1286, QN => n6834);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n3154, CK => CLK, Q => 
                           n_1287, QN => n6835);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n3153, CK => CLK, Q => 
                           n_1288, QN => n6836);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n3152, CK => CLK, Q => 
                           n_1289, QN => n6837);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n3151, CK => CLK, Q => 
                           n_1290, QN => n6838);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n3150, CK => CLK, Q => 
                           n_1291, QN => n6839);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n3149, CK => CLK, Q => 
                           n_1292, QN => n6840);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n3148, CK => CLK, Q => 
                           n_1293, QN => n6841);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n3147, CK => CLK, Q => 
                           n_1294, QN => n6842);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n3146, CK => CLK, Q => 
                           n_1295, QN => n6843);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n3145, CK => CLK, Q => 
                           n_1296, QN => n6844);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n3144, CK => CLK, Q => 
                           n_1297, QN => n6845);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n3143, CK => CLK, Q => 
                           n_1298, QN => n6846);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n3142, CK => CLK, Q => 
                           n_1299, QN => n6847);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n3141, CK => CLK, Q => 
                           n_1300, QN => n6848);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n3140, CK => CLK, Q => 
                           n_1301, QN => n6849);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n3139, CK => CLK, Q => 
                           n_1302, QN => n6850);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n3138, CK => CLK, Q => 
                           n_1303, QN => n6851);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n3137, CK => CLK, Q => 
                           n_1304, QN => n6852);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n3136, CK => CLK, Q => 
                           n_1305, QN => n6853);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n3135, CK => CLK, Q => 
                           n_1306, QN => n6854);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n3134, CK => CLK, Q => 
                           n_1307, QN => n6855);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n3613, CK => CLK, Q => 
                           n_1308, QN => n6465);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n3612, CK => CLK, Q => 
                           n_1309, QN => n6466);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n3611, CK => CLK, Q => 
                           n_1310, QN => n6467);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n3610, CK => CLK, Q => 
                           n_1311, QN => n6468);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n3604, CK => CLK, Q => 
                           n_1312, QN => n6469);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n3603, CK => CLK, Q => 
                           n_1313, QN => n6470);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n3602, CK => CLK, Q => 
                           n_1314, QN => n6471);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n2677, CK => CLK, Q => 
                           n_1315, QN => n7312);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n2676, CK => CLK, Q => 
                           n_1316, QN => n7313);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n2675, CK => CLK, Q => 
                           n_1317, QN => n7314);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n2674, CK => CLK, Q => 
                           n_1318, QN => n7315);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n2673, CK => CLK, Q => 
                           n_1319, QN => n7316);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n2672, CK => CLK, Q => 
                           n_1320, QN => n7317);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n2671, CK => CLK, Q => 
                           n_1321, QN => n7318);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n2670, CK => CLK, Q => 
                           n_1322, QN => n7319);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n2669, CK => CLK, Q => 
                           n_1323, QN => n7320);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n2668, CK => CLK, Q => 
                           n_1324, QN => n7321);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n2667, CK => CLK, Q => 
                           n_1325, QN => n7322);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n2666, CK => CLK, Q => 
                           n_1326, QN => n7323);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n2665, CK => CLK, Q => 
                           n_1327, QN => n7324);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n2664, CK => CLK, Q => 
                           n_1328, QN => n7325);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n2663, CK => CLK, Q => 
                           n_1329, QN => n7326);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n2662, CK => CLK, Q => 
                           n_1330, QN => n7327);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n2661, CK => CLK, Q => 
                           n_1331, QN => n7328);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n2660, CK => CLK, Q => 
                           n_1332, QN => n7329);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n2659, CK => CLK, Q => 
                           n_1333, QN => n7330);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n2658, CK => CLK, Q => 
                           n_1334, QN => n7331);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n2657, CK => CLK, Q => 
                           n_1335, QN => n7332);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n2656, CK => CLK, Q => 
                           n_1336, QN => n7333);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n2655, CK => CLK, Q => 
                           n_1337, QN => n7334);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n2654, CK => CLK, Q => 
                           n_1338, QN => n7335);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n2805, CK => CLK, Q => 
                           n_1339, QN => n7184);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n2804, CK => CLK, Q => 
                           n_1340, QN => n7185);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n2803, CK => CLK, Q => 
                           n_1341, QN => n7186);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n2802, CK => CLK, Q => 
                           n_1342, QN => n7187);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n2801, CK => CLK, Q => 
                           n_1343, QN => n7188);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n2800, CK => CLK, Q => 
                           n_1344, QN => n7189);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n2799, CK => CLK, Q => 
                           n_1345, QN => n7190);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n2798, CK => CLK, Q => 
                           n_1346, QN => n7191);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n2797, CK => CLK, Q => 
                           n_1347, QN => n7192);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n2796, CK => CLK, Q => 
                           n_1348, QN => n7193);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n2795, CK => CLK, Q => 
                           n_1349, QN => n7194);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n2794, CK => CLK, Q => 
                           n_1350, QN => n7195);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n2793, CK => CLK, Q => 
                           n_1351, QN => n7196);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n2792, CK => CLK, Q => 
                           n_1352, QN => n7197);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n2791, CK => CLK, Q => 
                           n_1353, QN => n7198);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n2790, CK => CLK, Q => 
                           n_1354, QN => n7199);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n2789, CK => CLK, Q => 
                           n_1355, QN => n7200);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n2788, CK => CLK, Q => 
                           n_1356, QN => n7201);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n2787, CK => CLK, Q => 
                           n_1357, QN => n7202);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n2786, CK => CLK, Q => 
                           n_1358, QN => n7203);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n2785, CK => CLK, Q => 
                           n_1359, QN => n7204);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n2784, CK => CLK, Q => 
                           n_1360, QN => n7205);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n2783, CK => CLK, Q => 
                           n_1361, QN => n7206);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n2782, CK => CLK, Q => 
                           n_1362, QN => n7207);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n2869, CK => CLK, Q => 
                           n_1363, QN => n7120);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n2868, CK => CLK, Q => 
                           n_1364, QN => n7121);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n2867, CK => CLK, Q => 
                           n_1365, QN => n7122);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n2866, CK => CLK, Q => 
                           n_1366, QN => n7123);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n2865, CK => CLK, Q => 
                           n_1367, QN => n7124);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n2864, CK => CLK, Q => 
                           n_1368, QN => n7125);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n2863, CK => CLK, Q => 
                           n_1369, QN => n7126);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n2862, CK => CLK, Q => 
                           n_1370, QN => n7127);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n2861, CK => CLK, Q => 
                           n_1371, QN => n7128);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n2860, CK => CLK, Q => 
                           n_1372, QN => n7129);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n2859, CK => CLK, Q => 
                           n_1373, QN => n7130);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n2858, CK => CLK, Q => 
                           n_1374, QN => n7131);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n2857, CK => CLK, Q => 
                           n_1375, QN => n7132);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n2856, CK => CLK, Q => 
                           n_1376, QN => n7133);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n2855, CK => CLK, Q => 
                           n_1377, QN => n7134);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n2854, CK => CLK, Q => 
                           n_1378, QN => n7135);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n2853, CK => CLK, Q => 
                           n_1379, QN => n7136);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n2852, CK => CLK, Q => 
                           n_1380, QN => n7137);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n2851, CK => CLK, Q => 
                           n_1381, QN => n7138);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n2850, CK => CLK, Q => 
                           n_1382, QN => n7139);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n2849, CK => CLK, Q => 
                           n_1383, QN => n7140);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n2848, CK => CLK, Q => 
                           n_1384, QN => n7141);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n2847, CK => CLK, Q => 
                           n_1385, QN => n7142);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n2846, CK => CLK, Q => 
                           n_1386, QN => n7143);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n2997, CK => CLK, Q => 
                           n_1387, QN => n6992);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n2996, CK => CLK, Q => 
                           n_1388, QN => n6993);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n2995, CK => CLK, Q => 
                           n_1389, QN => n6994);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n2994, CK => CLK, Q => 
                           n_1390, QN => n6995);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n2993, CK => CLK, Q => 
                           n_1391, QN => n6996);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n2992, CK => CLK, Q => 
                           n_1392, QN => n6997);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n2991, CK => CLK, Q => 
                           n_1393, QN => n6998);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n2990, CK => CLK, Q => 
                           n_1394, QN => n6999);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n2989, CK => CLK, Q => 
                           n_1395, QN => n7000);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n2988, CK => CLK, Q => 
                           n_1396, QN => n7001);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n2987, CK => CLK, Q => 
                           n_1397, QN => n7002);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n2986, CK => CLK, Q => 
                           n_1398, QN => n7003);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n2985, CK => CLK, Q => 
                           n_1399, QN => n7004);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n2984, CK => CLK, Q => 
                           n_1400, QN => n7005);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n2983, CK => CLK, Q => 
                           n_1401, QN => n7006);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n2982, CK => CLK, Q => 
                           n_1402, QN => n7007);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n2981, CK => CLK, Q => 
                           n_1403, QN => n7008);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n2980, CK => CLK, Q => 
                           n_1404, QN => n7009);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n2979, CK => CLK, Q => 
                           n_1405, QN => n7010);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n2978, CK => CLK, Q => 
                           n_1406, QN => n7011);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n2977, CK => CLK, Q => 
                           n_1407, QN => n7012);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n2976, CK => CLK, Q => 
                           n_1408, QN => n7013);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n2975, CK => CLK, Q => 
                           n_1409, QN => n7014);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n2974, CK => CLK, Q => 
                           n_1410, QN => n7015);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n3125, CK => CLK, Q => 
                           n_1411, QN => n6864);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n3124, CK => CLK, Q => 
                           n_1412, QN => n6865);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n3123, CK => CLK, Q => 
                           n_1413, QN => n6866);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n3122, CK => CLK, Q => 
                           n_1414, QN => n6867);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n3121, CK => CLK, Q => 
                           n_1415, QN => n6868);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n3120, CK => CLK, Q => 
                           n_1416, QN => n6869);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n3119, CK => CLK, Q => 
                           n_1417, QN => n6870);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n3118, CK => CLK, Q => 
                           n_1418, QN => n6871);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n3117, CK => CLK, Q => 
                           n_1419, QN => n6872);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n3116, CK => CLK, Q => 
                           n_1420, QN => n6873);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n3115, CK => CLK, Q => 
                           n_1421, QN => n6874);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n3114, CK => CLK, Q => 
                           n_1422, QN => n6875);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n3113, CK => CLK, Q => 
                           n_1423, QN => n6876);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n3112, CK => CLK, Q => 
                           n_1424, QN => n6877);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n3111, CK => CLK, Q => 
                           n_1425, QN => n6878);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n3110, CK => CLK, Q => 
                           n_1426, QN => n6879);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n3109, CK => CLK, Q => 
                           n_1427, QN => n6880);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n3108, CK => CLK, Q => 
                           n_1428, QN => n6881);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n3107, CK => CLK, Q => 
                           n_1429, QN => n6882);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n3106, CK => CLK, Q => 
                           n_1430, QN => n6883);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n3105, CK => CLK, Q => 
                           n_1431, QN => n6884);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n3104, CK => CLK, Q => 
                           n_1432, QN => n6885);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n3103, CK => CLK, Q => 
                           n_1433, QN => n6886);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n3102, CK => CLK, Q => 
                           n_1434, QN => n6887);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n3601, CK => CLK, Q => 
                           n_1435, QN => n6472);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n3600, CK => CLK, Q => 
                           n_1436, QN => n6473);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n3599, CK => CLK, Q => 
                           n_1437, QN => n6474);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n3598, CK => CLK, Q => 
                           n_1438, QN => n6475);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n3597, CK => CLK, Q => 
                           n_1439, QN => n6476);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n3596, CK => CLK, Q => 
                           n_1440, QN => n6477);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n3595, CK => CLK, Q => 
                           n_1441, QN => n6478);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n3594, CK => CLK, Q => 
                           n_1442, QN => n6479);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n3593, CK => CLK, Q => 
                           n_1443, QN => n6480);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n3592, CK => CLK, Q => 
                           n_1444, QN => n6481);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n3591, CK => CLK, Q => n_1445
                           , QN => n6482);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n3590, CK => CLK, Q => n_1446
                           , QN => n6483);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n3582, CK => CLK, Q => n_1447
                           , QN => n6491);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n3261, CK => CLK, Q => 
                           n4350, QN => n6728);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n3260, CK => CLK, Q => 
                           n4351, QN => n6729);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n3259, CK => CLK, Q => 
                           n4352, QN => n6730);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n3258, CK => CLK, Q => 
                           n4353, QN => n6731);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n3257, CK => CLK, Q => 
                           n4354, QN => n6732);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n3256, CK => CLK, Q => 
                           n4355, QN => n6733);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n3255, CK => CLK, Q => 
                           n4356, QN => n6734);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n3254, CK => CLK, Q => 
                           n4357, QN => n6735);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n3325, CK => CLK, Q => n4318
                           , QN => n6664);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n3324, CK => CLK, Q => n4319
                           , QN => n6665);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n3323, CK => CLK, Q => n4320
                           , QN => n6666);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n3322, CK => CLK, Q => n4321
                           , QN => n6667);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n3321, CK => CLK, Q => n4322
                           , QN => n6668);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n3320, CK => CLK, Q => n4323
                           , QN => n6669);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n3319, CK => CLK, Q => n4324
                           , QN => n6670);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n3318, CK => CLK, Q => n4325
                           , QN => n6671);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n3253, CK => CLK, Q => 
                           n4358, QN => n6736);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n3252, CK => CLK, Q => 
                           n4359, QN => n6737);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n3251, CK => CLK, Q => 
                           n4360, QN => n6738);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n3250, CK => CLK, Q => 
                           n4361, QN => n6739);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n3249, CK => CLK, Q => 
                           n4362, QN => n6740);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n3248, CK => CLK, Q => 
                           n4363, QN => n6741);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n3247, CK => CLK, Q => 
                           n4364, QN => n6742);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n3246, CK => CLK, Q => 
                           n4365, QN => n6743);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n3245, CK => CLK, Q => 
                           n4366, QN => n6744);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n3244, CK => CLK, Q => 
                           n4367, QN => n6745);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n3243, CK => CLK, Q => 
                           n4368, QN => n6746);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n3242, CK => CLK, Q => 
                           n4369, QN => n6747);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n3241, CK => CLK, Q => 
                           n4370, QN => n6748);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n3240, CK => CLK, Q => 
                           n4371, QN => n6749);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n3239, CK => CLK, Q => n4372
                           , QN => n6750);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n3238, CK => CLK, Q => n4373
                           , QN => n6751);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n3237, CK => CLK, Q => n4374
                           , QN => n6752);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n3236, CK => CLK, Q => n4375
                           , QN => n6753);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n3235, CK => CLK, Q => n4376
                           , QN => n6754);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n3234, CK => CLK, Q => n4377
                           , QN => n6755);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n3233, CK => CLK, Q => n4378
                           , QN => n6756);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n3232, CK => CLK, Q => n4379
                           , QN => n6757);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n3231, CK => CLK, Q => n4380
                           , QN => n6758);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n3230, CK => CLK, Q => n4381
                           , QN => n6759);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n3317, CK => CLK, Q => n4326
                           , QN => n6672);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n3316, CK => CLK, Q => n4327
                           , QN => n6673);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n3315, CK => CLK, Q => n4328
                           , QN => n6674);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n3314, CK => CLK, Q => n4329
                           , QN => n6675);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n3313, CK => CLK, Q => n4330
                           , QN => n6676);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n3312, CK => CLK, Q => n4331
                           , QN => n6677);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n3311, CK => CLK, Q => n4332
                           , QN => n6678);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n3310, CK => CLK, Q => n4333
                           , QN => n6679);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n3309, CK => CLK, Q => n4334
                           , QN => n6680);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n3308, CK => CLK, Q => n4335
                           , QN => n6681);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n3307, CK => CLK, Q => n4336
                           , QN => n6682);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n3306, CK => CLK, Q => n4337
                           , QN => n6683);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n3305, CK => CLK, Q => n4338
                           , QN => n6684);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n3304, CK => CLK, Q => n4339
                           , QN => n6685);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n3303, CK => CLK, Q => n4340,
                           QN => n6686);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n3302, CK => CLK, Q => n4341,
                           QN => n6687);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n3301, CK => CLK, Q => n4342,
                           QN => n6688);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n3300, CK => CLK, Q => n4343,
                           QN => n6689);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n3299, CK => CLK, Q => n4344,
                           QN => n6690);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n3298, CK => CLK, Q => n4345,
                           QN => n6691);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n3297, CK => CLK, Q => n4346,
                           QN => n6692);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n3296, CK => CLK, Q => n4347,
                           QN => n6693);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n3295, CK => CLK, Q => n4348,
                           QN => n6694);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n3294, CK => CLK, Q => n4349,
                           QN => n6695);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n3293, CK => CLK, Q => 
                           n3966, QN => n6696);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n3292, CK => CLK, Q => 
                           n3967, QN => n6697);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n3291, CK => CLK, Q => 
                           n3968, QN => n6698);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n3290, CK => CLK, Q => 
                           n3969, QN => n6699);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n3289, CK => CLK, Q => 
                           n3970, QN => n6700);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n3288, CK => CLK, Q => 
                           n3971, QN => n6701);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n3287, CK => CLK, Q => 
                           n3972, QN => n6702);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n3286, CK => CLK, Q => 
                           n3973, QN => n6703);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n3357, CK => CLK, Q => n3934
                           , QN => n6632);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n3356, CK => CLK, Q => n3935
                           , QN => n6633);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n3355, CK => CLK, Q => n3936
                           , QN => n6634);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n3354, CK => CLK, Q => n3937
                           , QN => n6635);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n3353, CK => CLK, Q => n3938
                           , QN => n6636);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n3352, CK => CLK, Q => n3939
                           , QN => n6637);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n3351, CK => CLK, Q => n3940
                           , QN => n6638);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n3350, CK => CLK, Q => n3941
                           , QN => n6639);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n3285, CK => CLK, Q => 
                           n3974, QN => n6704);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n3284, CK => CLK, Q => 
                           n3975, QN => n6705);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n3283, CK => CLK, Q => 
                           n3976, QN => n6706);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n3282, CK => CLK, Q => 
                           n3977, QN => n6707);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n3281, CK => CLK, Q => 
                           n3978, QN => n6708);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n3280, CK => CLK, Q => 
                           n3979, QN => n6709);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n3279, CK => CLK, Q => 
                           n3980, QN => n6710);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n3278, CK => CLK, Q => 
                           n3981, QN => n6711);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n3277, CK => CLK, Q => 
                           n3982, QN => n6712);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n3276, CK => CLK, Q => 
                           n3983, QN => n6713);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n3275, CK => CLK, Q => 
                           n3984, QN => n6714);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n3274, CK => CLK, Q => 
                           n3985, QN => n6715);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n3273, CK => CLK, Q => 
                           n3986, QN => n6716);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n3272, CK => CLK, Q => 
                           n3987, QN => n6717);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n3271, CK => CLK, Q => n3988
                           , QN => n6718);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n3270, CK => CLK, Q => n3989
                           , QN => n6719);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n3269, CK => CLK, Q => n3990
                           , QN => n6720);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n3268, CK => CLK, Q => n3991
                           , QN => n6721);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n3267, CK => CLK, Q => n3992
                           , QN => n6722);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n3266, CK => CLK, Q => n3993
                           , QN => n6723);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n3265, CK => CLK, Q => n3994
                           , QN => n6724);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n3264, CK => CLK, Q => n3995
                           , QN => n6725);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n3263, CK => CLK, Q => n3996
                           , QN => n6726);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n3262, CK => CLK, Q => n3997
                           , QN => n6727);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n3349, CK => CLK, Q => n3942
                           , QN => n6640);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n3348, CK => CLK, Q => n3943
                           , QN => n6641);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n3347, CK => CLK, Q => n3944
                           , QN => n6642);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n3346, CK => CLK, Q => n3945
                           , QN => n6643);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n3345, CK => CLK, Q => n3946
                           , QN => n6644);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n3344, CK => CLK, Q => n3947
                           , QN => n6645);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n3343, CK => CLK, Q => n3948
                           , QN => n6646);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n3342, CK => CLK, Q => n3949
                           , QN => n6647);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n3341, CK => CLK, Q => n3950
                           , QN => n6648);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n3340, CK => CLK, Q => n3951
                           , QN => n6649);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n3339, CK => CLK, Q => n3952
                           , QN => n6650);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n3338, CK => CLK, Q => n3953
                           , QN => n6651);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n3337, CK => CLK, Q => n3954
                           , QN => n6652);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n3336, CK => CLK, Q => n3955
                           , QN => n6653);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n3335, CK => CLK, Q => n3956,
                           QN => n6654);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n3334, CK => CLK, Q => n3957,
                           QN => n6655);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n3333, CK => CLK, Q => n3958,
                           QN => n6656);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n3332, CK => CLK, Q => n3959,
                           QN => n6657);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n3331, CK => CLK, Q => n3960,
                           QN => n6658);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n3330, CK => CLK, Q => n3961,
                           QN => n6659);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n3329, CK => CLK, Q => n3962,
                           QN => n6660);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n3328, CK => CLK, Q => n3963,
                           QN => n6661);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n3327, CK => CLK, Q => n3964,
                           QN => n6662);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n3326, CK => CLK, Q => n3965,
                           QN => n6663);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n3453, CK => CLK, Q => n4478
                           , QN => n6600);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n3452, CK => CLK, Q => n4479
                           , QN => n6601);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n3451, CK => CLK, Q => n4480
                           , QN => n6602);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n3450, CK => CLK, Q => n4481
                           , QN => n6603);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n3449, CK => CLK, Q => n4482
                           , QN => n6604);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n3448, CK => CLK, Q => n4483
                           , QN => n6605);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n3447, CK => CLK, Q => n4484
                           , QN => n6606);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n3446, CK => CLK, Q => n4485
                           , QN => n6607);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n3445, CK => CLK, Q => n4486
                           , QN => n6608);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n3444, CK => CLK, Q => n4487
                           , QN => n6609);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n3443, CK => CLK, Q => n4488
                           , QN => n6610);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n3442, CK => CLK, Q => n4489
                           , QN => n6611);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n3441, CK => CLK, Q => n4490
                           , QN => n6612);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n3440, CK => CLK, Q => n4491
                           , QN => n6613);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n3439, CK => CLK, Q => n4492
                           , QN => n6614);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n3438, CK => CLK, Q => n4493
                           , QN => n6615);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n3437, CK => CLK, Q => n4494
                           , QN => n6616);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n3436, CK => CLK, Q => n4495
                           , QN => n6617);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n3435, CK => CLK, Q => n4496
                           , QN => n6618);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n3434, CK => CLK, Q => n4497
                           , QN => n6619);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n3433, CK => CLK, Q => n4498
                           , QN => n6620);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n3432, CK => CLK, Q => n4499
                           , QN => n6621);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n3431, CK => CLK, Q => n4500,
                           QN => n6622);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n3430, CK => CLK, Q => n4501,
                           QN => n6623);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n3429, CK => CLK, Q => n4502,
                           QN => n6624);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n3428, CK => CLK, Q => n4503,
                           QN => n6625);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n3427, CK => CLK, Q => n4504,
                           QN => n6626);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n3426, CK => CLK, Q => n4505,
                           QN => n6627);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n3425, CK => CLK, Q => n4506,
                           QN => n6628);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n3424, CK => CLK, Q => n4507,
                           QN => n6629);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n3423, CK => CLK, Q => n4508,
                           QN => n6630);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n3422, CK => CLK, Q => n4509,
                           QN => n6631);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n3485, CK => CLK, Q => n4414
                           , QN => n6568);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n3484, CK => CLK, Q => n4415
                           , QN => n6569);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n3483, CK => CLK, Q => n4416
                           , QN => n6570);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n3482, CK => CLK, Q => n4417
                           , QN => n6571);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n3481, CK => CLK, Q => n4418
                           , QN => n6572);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n3480, CK => CLK, Q => n4419
                           , QN => n6573);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n3479, CK => CLK, Q => n4420
                           , QN => n6574);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n3478, CK => CLK, Q => n4421
                           , QN => n6575);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n3477, CK => CLK, Q => n4422
                           , QN => n6576);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n3476, CK => CLK, Q => n4423
                           , QN => n6577);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n3475, CK => CLK, Q => n4424
                           , QN => n6578);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n3474, CK => CLK, Q => n4425
                           , QN => n6579);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n3473, CK => CLK, Q => n4426
                           , QN => n6580);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n3472, CK => CLK, Q => n4427
                           , QN => n6581);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n3471, CK => CLK, Q => n4428
                           , QN => n6582);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n3470, CK => CLK, Q => n4429
                           , QN => n6583);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n3469, CK => CLK, Q => n4430
                           , QN => n6584);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n3468, CK => CLK, Q => n4431
                           , QN => n6585);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n3467, CK => CLK, Q => n4432
                           , QN => n6586);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n3466, CK => CLK, Q => n4433
                           , QN => n6587);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n3465, CK => CLK, Q => n4434
                           , QN => n6588);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n3464, CK => CLK, Q => n4435
                           , QN => n6589);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n3463, CK => CLK, Q => n4436,
                           QN => n6590);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n3462, CK => CLK, Q => n4437,
                           QN => n6591);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n3461, CK => CLK, Q => n4438,
                           QN => n6592);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n3460, CK => CLK, Q => n4439,
                           QN => n6593);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n3459, CK => CLK, Q => n4440,
                           QN => n6594);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n3458, CK => CLK, Q => n4441,
                           QN => n6595);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n3457, CK => CLK, Q => n4442,
                           QN => n6596);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n3456, CK => CLK, Q => n4443,
                           QN => n6597);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n3455, CK => CLK, Q => n4444,
                           QN => n6598);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n3454, CK => CLK, Q => n4445,
                           QN => n6599);
   U5980 : NOR2_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), ZN => n8763);
   U5981 : INV_X1 port map( A => n9880, ZN => n9873);
   U5982 : INV_X1 port map( A => n9517, ZN => n9510);
   U5983 : INV_X1 port map( A => n9544, ZN => n9537);
   U5984 : INV_X1 port map( A => n9553, ZN => n9546);
   U5985 : INV_X1 port map( A => n9598, ZN => n9591);
   U5986 : INV_X1 port map( A => n9607, ZN => n9600);
   U5987 : INV_X1 port map( A => n9634, ZN => n9627);
   U5988 : INV_X1 port map( A => n9643, ZN => n9636);
   U5989 : INV_X1 port map( A => n9670, ZN => n9663);
   U5990 : INV_X1 port map( A => n9679, ZN => n9672);
   U5991 : INV_X1 port map( A => n9724, ZN => n9717);
   U5992 : INV_X1 port map( A => n9733, ZN => n9726);
   U5993 : INV_X1 port map( A => n9760, ZN => n9753);
   U5994 : INV_X1 port map( A => n9769, ZN => n9762);
   U5995 : INV_X1 port map( A => n9778, ZN => n9771);
   U5996 : INV_X1 port map( A => n9526, ZN => n9519);
   U5997 : INV_X1 port map( A => n9535, ZN => n9528);
   U5998 : INV_X1 port map( A => n9562, ZN => n9555);
   U5999 : INV_X1 port map( A => n9571, ZN => n9564);
   U6000 : INV_X1 port map( A => n9580, ZN => n9573);
   U6001 : INV_X1 port map( A => n9589, ZN => n9582);
   U6002 : INV_X1 port map( A => n9616, ZN => n9609);
   U6003 : INV_X1 port map( A => n9625, ZN => n9618);
   U6004 : INV_X1 port map( A => n9652, ZN => n9645);
   U6005 : INV_X1 port map( A => n9661, ZN => n9654);
   U6006 : INV_X1 port map( A => n9688, ZN => n9681);
   U6007 : INV_X1 port map( A => n9697, ZN => n9690);
   U6008 : INV_X1 port map( A => n9706, ZN => n9699);
   U6009 : INV_X1 port map( A => n9715, ZN => n9708);
   U6010 : INV_X1 port map( A => n9742, ZN => n9735);
   U6011 : INV_X1 port map( A => n9751, ZN => n9744);
   U6012 : BUF_X1 port map( A => n9881, Z => n9874);
   U6013 : BUF_X1 port map( A => n9881, Z => n9875);
   U6014 : BUF_X1 port map( A => n9881, Z => n9876);
   U6015 : BUF_X1 port map( A => n9881, Z => n9877);
   U6016 : BUF_X1 port map( A => n9881, Z => n9878);
   U6017 : BUF_X1 port map( A => n9881, Z => n9879);
   U6018 : BUF_X1 port map( A => n9881, Z => n9880);
   U6019 : BUF_X1 port map( A => n9509, Z => n9508);
   U6020 : BUF_X1 port map( A => n9509, Z => n9506);
   U6021 : BUF_X1 port map( A => n9509, Z => n9505);
   U6022 : BUF_X1 port map( A => n9508, Z => n9504);
   U6023 : BUF_X1 port map( A => n9502, Z => n9503);
   U6024 : BUF_X1 port map( A => n9509, Z => n9502);
   U6025 : BUF_X1 port map( A => n9508, Z => n9501);
   U6026 : BUF_X1 port map( A => n9509, Z => n9500);
   U6027 : BUF_X1 port map( A => n9509, Z => n9507);
   U6028 : BUF_X1 port map( A => n8141, Z => n9382);
   U6029 : BUF_X1 port map( A => n8146, Z => n9370);
   U6030 : BUF_X1 port map( A => n8151, Z => n9358);
   U6031 : BUF_X1 port map( A => n8156, Z => n9346);
   U6032 : BUF_X1 port map( A => n8175, Z => n9310);
   U6033 : BUF_X1 port map( A => n8165, Z => n9334);
   U6034 : BUF_X1 port map( A => n8180, Z => n9298);
   U6035 : BUF_X1 port map( A => n8170, Z => n9322);
   U6036 : BUF_X1 port map( A => n8141, Z => n9383);
   U6037 : BUF_X1 port map( A => n8146, Z => n9371);
   U6038 : BUF_X1 port map( A => n8151, Z => n9359);
   U6039 : BUF_X1 port map( A => n8156, Z => n9347);
   U6040 : BUF_X1 port map( A => n8165, Z => n9335);
   U6041 : BUF_X1 port map( A => n8175, Z => n9311);
   U6042 : BUF_X1 port map( A => n8180, Z => n9299);
   U6043 : BUF_X1 port map( A => n8170, Z => n9323);
   U6044 : BUF_X1 port map( A => n7488, Z => n9484);
   U6045 : BUF_X1 port map( A => n7493, Z => n9472);
   U6046 : BUF_X1 port map( A => n7498, Z => n9460);
   U6047 : BUF_X1 port map( A => n7503, Z => n9448);
   U6048 : BUF_X1 port map( A => n7522, Z => n9412);
   U6049 : BUF_X1 port map( A => n7512, Z => n9436);
   U6050 : BUF_X1 port map( A => n7527, Z => n9400);
   U6051 : BUF_X1 port map( A => n7517, Z => n9424);
   U6052 : BUF_X1 port map( A => n7488, Z => n9485);
   U6053 : BUF_X1 port map( A => n7493, Z => n9473);
   U6054 : BUF_X1 port map( A => n7498, Z => n9461);
   U6055 : BUF_X1 port map( A => n7503, Z => n9449);
   U6056 : BUF_X1 port map( A => n7512, Z => n9437);
   U6057 : BUF_X1 port map( A => n7522, Z => n9413);
   U6058 : BUF_X1 port map( A => n7527, Z => n9401);
   U6059 : BUF_X1 port map( A => n7517, Z => n9425);
   U6060 : BUF_X1 port map( A => n8142, Z => n9379);
   U6061 : BUF_X1 port map( A => n8147, Z => n9367);
   U6062 : BUF_X1 port map( A => n8152, Z => n9355);
   U6063 : BUF_X1 port map( A => n8157, Z => n9343);
   U6064 : BUF_X1 port map( A => n8176, Z => n9307);
   U6065 : BUF_X1 port map( A => n8166, Z => n9331);
   U6066 : BUF_X1 port map( A => n8181, Z => n9295);
   U6067 : BUF_X1 port map( A => n8171, Z => n9319);
   U6068 : BUF_X1 port map( A => n8142, Z => n9380);
   U6069 : BUF_X1 port map( A => n8147, Z => n9368);
   U6070 : BUF_X1 port map( A => n8152, Z => n9356);
   U6071 : BUF_X1 port map( A => n8157, Z => n9344);
   U6072 : BUF_X1 port map( A => n8166, Z => n9332);
   U6073 : BUF_X1 port map( A => n8176, Z => n9308);
   U6074 : BUF_X1 port map( A => n8181, Z => n9296);
   U6075 : BUF_X1 port map( A => n8171, Z => n9320);
   U6076 : BUF_X1 port map( A => n7489, Z => n9481);
   U6077 : BUF_X1 port map( A => n7494, Z => n9469);
   U6078 : BUF_X1 port map( A => n7499, Z => n9457);
   U6079 : BUF_X1 port map( A => n7504, Z => n9445);
   U6080 : BUF_X1 port map( A => n7523, Z => n9409);
   U6081 : BUF_X1 port map( A => n7513, Z => n9433);
   U6082 : BUF_X1 port map( A => n7528, Z => n9397);
   U6083 : BUF_X1 port map( A => n7518, Z => n9421);
   U6084 : BUF_X1 port map( A => n7489, Z => n9482);
   U6085 : BUF_X1 port map( A => n7494, Z => n9470);
   U6086 : BUF_X1 port map( A => n7499, Z => n9458);
   U6087 : BUF_X1 port map( A => n7504, Z => n9446);
   U6088 : BUF_X1 port map( A => n7513, Z => n9434);
   U6089 : BUF_X1 port map( A => n7523, Z => n9410);
   U6090 : BUF_X1 port map( A => n7528, Z => n9398);
   U6091 : BUF_X1 port map( A => n7518, Z => n9422);
   U6092 : BUF_X1 port map( A => n8138, Z => n9388);
   U6093 : BUF_X1 port map( A => n8143, Z => n9376);
   U6094 : BUF_X1 port map( A => n8148, Z => n9364);
   U6095 : BUF_X1 port map( A => n8153, Z => n9352);
   U6096 : BUF_X1 port map( A => n8172, Z => n9316);
   U6097 : BUF_X1 port map( A => n8162, Z => n9340);
   U6098 : BUF_X1 port map( A => n8177, Z => n9304);
   U6099 : BUF_X1 port map( A => n8167, Z => n9328);
   U6100 : BUF_X1 port map( A => n8138, Z => n9389);
   U6101 : BUF_X1 port map( A => n8143, Z => n9377);
   U6102 : BUF_X1 port map( A => n8148, Z => n9365);
   U6103 : BUF_X1 port map( A => n8153, Z => n9353);
   U6104 : BUF_X1 port map( A => n8162, Z => n9341);
   U6105 : BUF_X1 port map( A => n8172, Z => n9317);
   U6106 : BUF_X1 port map( A => n8177, Z => n9305);
   U6107 : BUF_X1 port map( A => n8167, Z => n9329);
   U6108 : BUF_X1 port map( A => n7485, Z => n9490);
   U6109 : BUF_X1 port map( A => n7490, Z => n9478);
   U6110 : BUF_X1 port map( A => n7495, Z => n9466);
   U6111 : BUF_X1 port map( A => n7500, Z => n9454);
   U6112 : BUF_X1 port map( A => n7519, Z => n9418);
   U6113 : BUF_X1 port map( A => n7509, Z => n9442);
   U6114 : BUF_X1 port map( A => n7524, Z => n9406);
   U6115 : BUF_X1 port map( A => n7514, Z => n9430);
   U6116 : BUF_X1 port map( A => n7485, Z => n9491);
   U6117 : BUF_X1 port map( A => n7490, Z => n9479);
   U6118 : BUF_X1 port map( A => n7495, Z => n9467);
   U6119 : BUF_X1 port map( A => n7500, Z => n9455);
   U6120 : BUF_X1 port map( A => n7509, Z => n9443);
   U6121 : BUF_X1 port map( A => n7519, Z => n9419);
   U6122 : BUF_X1 port map( A => n7524, Z => n9407);
   U6123 : BUF_X1 port map( A => n7514, Z => n9431);
   U6124 : BUF_X1 port map( A => n8139, Z => n9385);
   U6125 : BUF_X1 port map( A => n8144, Z => n9373);
   U6126 : BUF_X1 port map( A => n8149, Z => n9361);
   U6127 : BUF_X1 port map( A => n8154, Z => n9349);
   U6128 : BUF_X1 port map( A => n8173, Z => n9313);
   U6129 : BUF_X1 port map( A => n8163, Z => n9337);
   U6130 : BUF_X1 port map( A => n8178, Z => n9301);
   U6131 : BUF_X1 port map( A => n8168, Z => n9325);
   U6132 : BUF_X1 port map( A => n8139, Z => n9386);
   U6133 : BUF_X1 port map( A => n8144, Z => n9374);
   U6134 : BUF_X1 port map( A => n8149, Z => n9362);
   U6135 : BUF_X1 port map( A => n8154, Z => n9350);
   U6136 : BUF_X1 port map( A => n8163, Z => n9338);
   U6137 : BUF_X1 port map( A => n8173, Z => n9314);
   U6138 : BUF_X1 port map( A => n8178, Z => n9302);
   U6139 : BUF_X1 port map( A => n8168, Z => n9326);
   U6140 : BUF_X1 port map( A => n7486, Z => n9487);
   U6141 : BUF_X1 port map( A => n7491, Z => n9475);
   U6142 : BUF_X1 port map( A => n7496, Z => n9463);
   U6143 : BUF_X1 port map( A => n7501, Z => n9451);
   U6144 : BUF_X1 port map( A => n7520, Z => n9415);
   U6145 : BUF_X1 port map( A => n7510, Z => n9439);
   U6146 : BUF_X1 port map( A => n7525, Z => n9403);
   U6147 : BUF_X1 port map( A => n7515, Z => n9427);
   U6148 : BUF_X1 port map( A => n7486, Z => n9488);
   U6149 : BUF_X1 port map( A => n7491, Z => n9476);
   U6150 : BUF_X1 port map( A => n7496, Z => n9464);
   U6151 : BUF_X1 port map( A => n7501, Z => n9452);
   U6152 : BUF_X1 port map( A => n7510, Z => n9440);
   U6153 : BUF_X1 port map( A => n7520, Z => n9416);
   U6154 : BUF_X1 port map( A => n7525, Z => n9404);
   U6155 : BUF_X1 port map( A => n7515, Z => n9428);
   U6156 : BUF_X1 port map( A => n8141, Z => n9384);
   U6157 : BUF_X1 port map( A => n8146, Z => n9372);
   U6158 : BUF_X1 port map( A => n8151, Z => n9360);
   U6159 : BUF_X1 port map( A => n8156, Z => n9348);
   U6160 : BUF_X1 port map( A => n8165, Z => n9336);
   U6161 : BUF_X1 port map( A => n8175, Z => n9312);
   U6162 : BUF_X1 port map( A => n8180, Z => n9300);
   U6163 : BUF_X1 port map( A => n8170, Z => n9324);
   U6164 : BUF_X1 port map( A => n7488, Z => n9486);
   U6165 : BUF_X1 port map( A => n7493, Z => n9474);
   U6166 : BUF_X1 port map( A => n7498, Z => n9462);
   U6167 : BUF_X1 port map( A => n7503, Z => n9450);
   U6168 : BUF_X1 port map( A => n7512, Z => n9438);
   U6169 : BUF_X1 port map( A => n7522, Z => n9414);
   U6170 : BUF_X1 port map( A => n7527, Z => n9402);
   U6171 : BUF_X1 port map( A => n7517, Z => n9426);
   U6172 : BUF_X1 port map( A => n8142, Z => n9381);
   U6173 : BUF_X1 port map( A => n8147, Z => n9369);
   U6174 : BUF_X1 port map( A => n8152, Z => n9357);
   U6175 : BUF_X1 port map( A => n8157, Z => n9345);
   U6176 : BUF_X1 port map( A => n8166, Z => n9333);
   U6177 : BUF_X1 port map( A => n8176, Z => n9309);
   U6178 : BUF_X1 port map( A => n8181, Z => n9297);
   U6179 : BUF_X1 port map( A => n8171, Z => n9321);
   U6180 : BUF_X1 port map( A => n7489, Z => n9483);
   U6181 : BUF_X1 port map( A => n7494, Z => n9471);
   U6182 : BUF_X1 port map( A => n7499, Z => n9459);
   U6183 : BUF_X1 port map( A => n7504, Z => n9447);
   U6184 : BUF_X1 port map( A => n7513, Z => n9435);
   U6185 : BUF_X1 port map( A => n7523, Z => n9411);
   U6186 : BUF_X1 port map( A => n7528, Z => n9399);
   U6187 : BUF_X1 port map( A => n7518, Z => n9423);
   U6188 : BUF_X1 port map( A => n8138, Z => n9390);
   U6189 : BUF_X1 port map( A => n8143, Z => n9378);
   U6190 : BUF_X1 port map( A => n8148, Z => n9366);
   U6191 : BUF_X1 port map( A => n8153, Z => n9354);
   U6192 : BUF_X1 port map( A => n8162, Z => n9342);
   U6193 : BUF_X1 port map( A => n8172, Z => n9318);
   U6194 : BUF_X1 port map( A => n8177, Z => n9306);
   U6195 : BUF_X1 port map( A => n8167, Z => n9330);
   U6196 : BUF_X1 port map( A => n7485, Z => n9492);
   U6197 : BUF_X1 port map( A => n7490, Z => n9480);
   U6198 : BUF_X1 port map( A => n7495, Z => n9468);
   U6199 : BUF_X1 port map( A => n7500, Z => n9456);
   U6200 : BUF_X1 port map( A => n7509, Z => n9444);
   U6201 : BUF_X1 port map( A => n7519, Z => n9420);
   U6202 : BUF_X1 port map( A => n7524, Z => n9408);
   U6203 : BUF_X1 port map( A => n7514, Z => n9432);
   U6204 : BUF_X1 port map( A => n8139, Z => n9387);
   U6205 : BUF_X1 port map( A => n8144, Z => n9375);
   U6206 : BUF_X1 port map( A => n8149, Z => n9363);
   U6207 : BUF_X1 port map( A => n8154, Z => n9351);
   U6208 : BUF_X1 port map( A => n8163, Z => n9339);
   U6209 : BUF_X1 port map( A => n8173, Z => n9315);
   U6210 : BUF_X1 port map( A => n8178, Z => n9303);
   U6211 : BUF_X1 port map( A => n8168, Z => n9327);
   U6212 : BUF_X1 port map( A => n7486, Z => n9489);
   U6213 : BUF_X1 port map( A => n7491, Z => n9477);
   U6214 : BUF_X1 port map( A => n7496, Z => n9465);
   U6215 : BUF_X1 port map( A => n7501, Z => n9453);
   U6216 : BUF_X1 port map( A => n7510, Z => n9441);
   U6217 : BUF_X1 port map( A => n7520, Z => n9417);
   U6218 : BUF_X1 port map( A => n7525, Z => n9405);
   U6219 : BUF_X1 port map( A => n7515, Z => n9429);
   U6220 : BUF_X1 port map( A => n9518, Z => n9511);
   U6221 : BUF_X1 port map( A => n9518, Z => n9512);
   U6222 : BUF_X1 port map( A => n9518, Z => n9513);
   U6223 : BUF_X1 port map( A => n9518, Z => n9514);
   U6224 : BUF_X1 port map( A => n9518, Z => n9515);
   U6225 : BUF_X1 port map( A => n9518, Z => n9516);
   U6226 : BUF_X1 port map( A => n9527, Z => n9520);
   U6227 : BUF_X1 port map( A => n9527, Z => n9521);
   U6228 : BUF_X1 port map( A => n9527, Z => n9522);
   U6229 : BUF_X1 port map( A => n9527, Z => n9523);
   U6230 : BUF_X1 port map( A => n9527, Z => n9524);
   U6231 : BUF_X1 port map( A => n9527, Z => n9525);
   U6232 : BUF_X1 port map( A => n9536, Z => n9529);
   U6233 : BUF_X1 port map( A => n9536, Z => n9530);
   U6234 : BUF_X1 port map( A => n9536, Z => n9531);
   U6235 : BUF_X1 port map( A => n9536, Z => n9532);
   U6236 : BUF_X1 port map( A => n9536, Z => n9533);
   U6237 : BUF_X1 port map( A => n9536, Z => n9534);
   U6238 : BUF_X1 port map( A => n9545, Z => n9538);
   U6239 : BUF_X1 port map( A => n9545, Z => n9539);
   U6240 : BUF_X1 port map( A => n9545, Z => n9540);
   U6241 : BUF_X1 port map( A => n9545, Z => n9541);
   U6242 : BUF_X1 port map( A => n9545, Z => n9542);
   U6243 : BUF_X1 port map( A => n9545, Z => n9543);
   U6244 : BUF_X1 port map( A => n9554, Z => n9547);
   U6245 : BUF_X1 port map( A => n9554, Z => n9548);
   U6246 : BUF_X1 port map( A => n9554, Z => n9549);
   U6247 : BUF_X1 port map( A => n9554, Z => n9550);
   U6248 : BUF_X1 port map( A => n9554, Z => n9551);
   U6249 : BUF_X1 port map( A => n9554, Z => n9552);
   U6250 : BUF_X1 port map( A => n9563, Z => n9556);
   U6251 : BUF_X1 port map( A => n9563, Z => n9557);
   U6252 : BUF_X1 port map( A => n9563, Z => n9558);
   U6253 : BUF_X1 port map( A => n9563, Z => n9559);
   U6254 : BUF_X1 port map( A => n9563, Z => n9560);
   U6255 : BUF_X1 port map( A => n9563, Z => n9561);
   U6256 : BUF_X1 port map( A => n9572, Z => n9565);
   U6257 : BUF_X1 port map( A => n9572, Z => n9566);
   U6258 : BUF_X1 port map( A => n9572, Z => n9567);
   U6259 : BUF_X1 port map( A => n9572, Z => n9568);
   U6260 : BUF_X1 port map( A => n9572, Z => n9569);
   U6261 : BUF_X1 port map( A => n9572, Z => n9570);
   U6262 : BUF_X1 port map( A => n9581, Z => n9574);
   U6263 : BUF_X1 port map( A => n9581, Z => n9575);
   U6264 : BUF_X1 port map( A => n9581, Z => n9576);
   U6265 : BUF_X1 port map( A => n9581, Z => n9577);
   U6266 : BUF_X1 port map( A => n9581, Z => n9578);
   U6267 : BUF_X1 port map( A => n9581, Z => n9579);
   U6268 : BUF_X1 port map( A => n9590, Z => n9583);
   U6269 : BUF_X1 port map( A => n9590, Z => n9584);
   U6270 : BUF_X1 port map( A => n9590, Z => n9585);
   U6271 : BUF_X1 port map( A => n9590, Z => n9586);
   U6272 : BUF_X1 port map( A => n9590, Z => n9587);
   U6273 : BUF_X1 port map( A => n9590, Z => n9588);
   U6274 : BUF_X1 port map( A => n9599, Z => n9592);
   U6275 : BUF_X1 port map( A => n9599, Z => n9593);
   U6276 : BUF_X1 port map( A => n9599, Z => n9594);
   U6277 : BUF_X1 port map( A => n9599, Z => n9595);
   U6278 : BUF_X1 port map( A => n9599, Z => n9596);
   U6279 : BUF_X1 port map( A => n9599, Z => n9597);
   U6280 : BUF_X1 port map( A => n9608, Z => n9601);
   U6281 : BUF_X1 port map( A => n9608, Z => n9602);
   U6282 : BUF_X1 port map( A => n9608, Z => n9603);
   U6283 : BUF_X1 port map( A => n9608, Z => n9604);
   U6284 : BUF_X1 port map( A => n9608, Z => n9605);
   U6285 : BUF_X1 port map( A => n9608, Z => n9606);
   U6286 : BUF_X1 port map( A => n9617, Z => n9610);
   U6287 : BUF_X1 port map( A => n9617, Z => n9611);
   U6288 : BUF_X1 port map( A => n9617, Z => n9612);
   U6289 : BUF_X1 port map( A => n9617, Z => n9613);
   U6290 : BUF_X1 port map( A => n9617, Z => n9614);
   U6291 : BUF_X1 port map( A => n9617, Z => n9615);
   U6292 : BUF_X1 port map( A => n9626, Z => n9619);
   U6293 : BUF_X1 port map( A => n9626, Z => n9620);
   U6294 : BUF_X1 port map( A => n9626, Z => n9621);
   U6295 : BUF_X1 port map( A => n9626, Z => n9622);
   U6296 : BUF_X1 port map( A => n9626, Z => n9623);
   U6297 : BUF_X1 port map( A => n9626, Z => n9624);
   U6298 : BUF_X1 port map( A => n9635, Z => n9628);
   U6299 : BUF_X1 port map( A => n9635, Z => n9629);
   U6300 : BUF_X1 port map( A => n9635, Z => n9630);
   U6301 : BUF_X1 port map( A => n9635, Z => n9631);
   U6302 : BUF_X1 port map( A => n9635, Z => n9632);
   U6303 : BUF_X1 port map( A => n9635, Z => n9633);
   U6304 : BUF_X1 port map( A => n9644, Z => n9637);
   U6305 : BUF_X1 port map( A => n9644, Z => n9638);
   U6306 : BUF_X1 port map( A => n9644, Z => n9639);
   U6307 : BUF_X1 port map( A => n9644, Z => n9640);
   U6308 : BUF_X1 port map( A => n9644, Z => n9641);
   U6309 : BUF_X1 port map( A => n9644, Z => n9642);
   U6310 : BUF_X1 port map( A => n9653, Z => n9646);
   U6311 : BUF_X1 port map( A => n9653, Z => n9647);
   U6312 : BUF_X1 port map( A => n9653, Z => n9648);
   U6313 : BUF_X1 port map( A => n9653, Z => n9649);
   U6314 : BUF_X1 port map( A => n9653, Z => n9650);
   U6315 : BUF_X1 port map( A => n9653, Z => n9651);
   U6316 : BUF_X1 port map( A => n9662, Z => n9655);
   U6317 : BUF_X1 port map( A => n9662, Z => n9656);
   U6318 : BUF_X1 port map( A => n9662, Z => n9657);
   U6319 : BUF_X1 port map( A => n9662, Z => n9658);
   U6320 : BUF_X1 port map( A => n9662, Z => n9659);
   U6321 : BUF_X1 port map( A => n9662, Z => n9660);
   U6322 : BUF_X1 port map( A => n9671, Z => n9664);
   U6323 : BUF_X1 port map( A => n9671, Z => n9665);
   U6324 : BUF_X1 port map( A => n9671, Z => n9666);
   U6325 : BUF_X1 port map( A => n9671, Z => n9667);
   U6326 : BUF_X1 port map( A => n9671, Z => n9668);
   U6327 : BUF_X1 port map( A => n9671, Z => n9669);
   U6328 : BUF_X1 port map( A => n9680, Z => n9673);
   U6329 : BUF_X1 port map( A => n9680, Z => n9674);
   U6330 : BUF_X1 port map( A => n9680, Z => n9675);
   U6331 : BUF_X1 port map( A => n9680, Z => n9676);
   U6332 : BUF_X1 port map( A => n9680, Z => n9677);
   U6333 : BUF_X1 port map( A => n9680, Z => n9678);
   U6334 : BUF_X1 port map( A => n9689, Z => n9682);
   U6335 : BUF_X1 port map( A => n9689, Z => n9683);
   U6336 : BUF_X1 port map( A => n9689, Z => n9684);
   U6337 : BUF_X1 port map( A => n9689, Z => n9685);
   U6338 : BUF_X1 port map( A => n9689, Z => n9686);
   U6339 : BUF_X1 port map( A => n9689, Z => n9687);
   U6340 : BUF_X1 port map( A => n9698, Z => n9691);
   U6341 : BUF_X1 port map( A => n9698, Z => n9692);
   U6342 : BUF_X1 port map( A => n9698, Z => n9693);
   U6343 : BUF_X1 port map( A => n9698, Z => n9694);
   U6344 : BUF_X1 port map( A => n9698, Z => n9695);
   U6345 : BUF_X1 port map( A => n9698, Z => n9696);
   U6346 : BUF_X1 port map( A => n9707, Z => n9700);
   U6347 : BUF_X1 port map( A => n9707, Z => n9701);
   U6348 : BUF_X1 port map( A => n9707, Z => n9702);
   U6349 : BUF_X1 port map( A => n9707, Z => n9703);
   U6350 : BUF_X1 port map( A => n9707, Z => n9704);
   U6351 : BUF_X1 port map( A => n9707, Z => n9705);
   U6352 : BUF_X1 port map( A => n9716, Z => n9709);
   U6353 : BUF_X1 port map( A => n9716, Z => n9710);
   U6354 : BUF_X1 port map( A => n9716, Z => n9711);
   U6355 : BUF_X1 port map( A => n9716, Z => n9712);
   U6356 : BUF_X1 port map( A => n9716, Z => n9713);
   U6357 : BUF_X1 port map( A => n9716, Z => n9714);
   U6358 : BUF_X1 port map( A => n9725, Z => n9718);
   U6359 : BUF_X1 port map( A => n9725, Z => n9719);
   U6360 : BUF_X1 port map( A => n9725, Z => n9720);
   U6361 : BUF_X1 port map( A => n9725, Z => n9721);
   U6362 : BUF_X1 port map( A => n9725, Z => n9722);
   U6363 : BUF_X1 port map( A => n9725, Z => n9723);
   U6364 : BUF_X1 port map( A => n9734, Z => n9727);
   U6365 : BUF_X1 port map( A => n9734, Z => n9728);
   U6366 : BUF_X1 port map( A => n9734, Z => n9729);
   U6367 : BUF_X1 port map( A => n9734, Z => n9730);
   U6368 : BUF_X1 port map( A => n9734, Z => n9731);
   U6369 : BUF_X1 port map( A => n9734, Z => n9732);
   U6370 : BUF_X1 port map( A => n9743, Z => n9736);
   U6371 : BUF_X1 port map( A => n9743, Z => n9737);
   U6372 : BUF_X1 port map( A => n9743, Z => n9738);
   U6373 : BUF_X1 port map( A => n9743, Z => n9739);
   U6374 : BUF_X1 port map( A => n9743, Z => n9740);
   U6375 : BUF_X1 port map( A => n9743, Z => n9741);
   U6376 : BUF_X1 port map( A => n9752, Z => n9745);
   U6377 : BUF_X1 port map( A => n9752, Z => n9746);
   U6378 : BUF_X1 port map( A => n9752, Z => n9747);
   U6379 : BUF_X1 port map( A => n9752, Z => n9748);
   U6380 : BUF_X1 port map( A => n9752, Z => n9749);
   U6381 : BUF_X1 port map( A => n9752, Z => n9750);
   U6382 : BUF_X1 port map( A => n9761, Z => n9754);
   U6383 : BUF_X1 port map( A => n9761, Z => n9755);
   U6384 : BUF_X1 port map( A => n9761, Z => n9756);
   U6385 : BUF_X1 port map( A => n9761, Z => n9757);
   U6386 : BUF_X1 port map( A => n9761, Z => n9758);
   U6387 : BUF_X1 port map( A => n9761, Z => n9759);
   U6388 : BUF_X1 port map( A => n9770, Z => n9763);
   U6389 : BUF_X1 port map( A => n9770, Z => n9764);
   U6390 : BUF_X1 port map( A => n9770, Z => n9765);
   U6391 : BUF_X1 port map( A => n9770, Z => n9766);
   U6392 : BUF_X1 port map( A => n9770, Z => n9767);
   U6393 : BUF_X1 port map( A => n9770, Z => n9768);
   U6394 : BUF_X1 port map( A => n9779, Z => n9772);
   U6395 : BUF_X1 port map( A => n9779, Z => n9773);
   U6396 : BUF_X1 port map( A => n9779, Z => n9774);
   U6397 : BUF_X1 port map( A => n9779, Z => n9775);
   U6398 : BUF_X1 port map( A => n9779, Z => n9776);
   U6399 : BUF_X1 port map( A => n9779, Z => n9777);
   U6400 : BUF_X1 port map( A => n9518, Z => n9517);
   U6401 : BUF_X1 port map( A => n9527, Z => n9526);
   U6402 : BUF_X1 port map( A => n9536, Z => n9535);
   U6403 : BUF_X1 port map( A => n9545, Z => n9544);
   U6404 : BUF_X1 port map( A => n9554, Z => n9553);
   U6405 : BUF_X1 port map( A => n9563, Z => n9562);
   U6406 : BUF_X1 port map( A => n9572, Z => n9571);
   U6407 : BUF_X1 port map( A => n9581, Z => n9580);
   U6408 : BUF_X1 port map( A => n9590, Z => n9589);
   U6409 : BUF_X1 port map( A => n9599, Z => n9598);
   U6410 : BUF_X1 port map( A => n9608, Z => n9607);
   U6411 : BUF_X1 port map( A => n9617, Z => n9616);
   U6412 : BUF_X1 port map( A => n9626, Z => n9625);
   U6413 : BUF_X1 port map( A => n9635, Z => n9634);
   U6414 : BUF_X1 port map( A => n9644, Z => n9643);
   U6415 : BUF_X1 port map( A => n9653, Z => n9652);
   U6416 : BUF_X1 port map( A => n9662, Z => n9661);
   U6417 : BUF_X1 port map( A => n9671, Z => n9670);
   U6418 : BUF_X1 port map( A => n9680, Z => n9679);
   U6419 : BUF_X1 port map( A => n9689, Z => n9688);
   U6420 : BUF_X1 port map( A => n9698, Z => n9697);
   U6421 : BUF_X1 port map( A => n9707, Z => n9706);
   U6422 : BUF_X1 port map( A => n9716, Z => n9715);
   U6423 : BUF_X1 port map( A => n9725, Z => n9724);
   U6424 : BUF_X1 port map( A => n9734, Z => n9733);
   U6425 : BUF_X1 port map( A => n9743, Z => n9742);
   U6426 : BUF_X1 port map( A => n9752, Z => n9751);
   U6427 : BUF_X1 port map( A => n9761, Z => n9760);
   U6428 : BUF_X1 port map( A => n9770, Z => n9769);
   U6429 : BUF_X1 port map( A => n9779, Z => n9778);
   U6430 : INV_X1 port map( A => n7401, ZN => n9881);
   U6431 : OAI21_X1 port map( B1 => n7433, B2 => n7434, A => n9887, ZN => n7401
                           );
   U6432 : INV_X1 port map( A => n9499, ZN => n9509);
   U6433 : AOI221_X1 port map( B1 => n9388, B2 => n6951, C1 => n9385, C2 => 
                           n6919, A => n8759, ZN => n8758);
   U6434 : OAI22_X1 port map( A1 => n7015, A2 => n9382, B1 => n6983, B2 => 
                           n9379, ZN => n8759);
   U6435 : AOI221_X1 port map( B1 => n9388, B2 => n6950, C1 => n9385, C2 => 
                           n6918, A => n8740, ZN => n8739);
   U6436 : OAI22_X1 port map( A1 => n7014, A2 => n9382, B1 => n6982, B2 => 
                           n9379, ZN => n8740);
   U6437 : AOI221_X1 port map( B1 => n9388, B2 => n6949, C1 => n9385, C2 => 
                           n6917, A => n8721, ZN => n8720);
   U6438 : OAI22_X1 port map( A1 => n7013, A2 => n9382, B1 => n6981, B2 => 
                           n9379, ZN => n8721);
   U6439 : AOI221_X1 port map( B1 => n9388, B2 => n6948, C1 => n9385, C2 => 
                           n6916, A => n8702, ZN => n8701);
   U6440 : OAI22_X1 port map( A1 => n7012, A2 => n9382, B1 => n6980, B2 => 
                           n9379, ZN => n8702);
   U6441 : AOI221_X1 port map( B1 => n9388, B2 => n6947, C1 => n9385, C2 => 
                           n6915, A => n8683, ZN => n8682);
   U6442 : OAI22_X1 port map( A1 => n7011, A2 => n9382, B1 => n6979, B2 => 
                           n9379, ZN => n8683);
   U6443 : AOI221_X1 port map( B1 => n9388, B2 => n6946, C1 => n9385, C2 => 
                           n6914, A => n8664, ZN => n8663);
   U6444 : OAI22_X1 port map( A1 => n7010, A2 => n9382, B1 => n6978, B2 => 
                           n9379, ZN => n8664);
   U6445 : AOI221_X1 port map( B1 => n9388, B2 => n6945, C1 => n9385, C2 => 
                           n6913, A => n8645, ZN => n8644);
   U6446 : OAI22_X1 port map( A1 => n7009, A2 => n9382, B1 => n6977, B2 => 
                           n9379, ZN => n8645);
   U6447 : AOI221_X1 port map( B1 => n9388, B2 => n6944, C1 => n9385, C2 => 
                           n6912, A => n8626, ZN => n8625);
   U6448 : OAI22_X1 port map( A1 => n7008, A2 => n9382, B1 => n6976, B2 => 
                           n9379, ZN => n8626);
   U6449 : AOI221_X1 port map( B1 => n9388, B2 => n6943, C1 => n9385, C2 => 
                           n6911, A => n8607, ZN => n8606);
   U6450 : OAI22_X1 port map( A1 => n7007, A2 => n9382, B1 => n6975, B2 => 
                           n9379, ZN => n8607);
   U6451 : AOI221_X1 port map( B1 => n9388, B2 => n6942, C1 => n9385, C2 => 
                           n6910, A => n8588, ZN => n8587);
   U6452 : OAI22_X1 port map( A1 => n7006, A2 => n9382, B1 => n6974, B2 => 
                           n9379, ZN => n8588);
   U6453 : AOI221_X1 port map( B1 => n9388, B2 => n6941, C1 => n9385, C2 => 
                           n6909, A => n8569, ZN => n8568);
   U6454 : OAI22_X1 port map( A1 => n7005, A2 => n9382, B1 => n6973, B2 => 
                           n9379, ZN => n8569);
   U6455 : AOI221_X1 port map( B1 => n9388, B2 => n6940, C1 => n9385, C2 => 
                           n6908, A => n8550, ZN => n8549);
   U6456 : OAI22_X1 port map( A1 => n7004, A2 => n9382, B1 => n6972, B2 => 
                           n9379, ZN => n8550);
   U6457 : AOI221_X1 port map( B1 => n9389, B2 => n6939, C1 => n9386, C2 => 
                           n6907, A => n8531, ZN => n8530);
   U6458 : OAI22_X1 port map( A1 => n7003, A2 => n9383, B1 => n6971, B2 => 
                           n9380, ZN => n8531);
   U6459 : AOI221_X1 port map( B1 => n9389, B2 => n6938, C1 => n9386, C2 => 
                           n6906, A => n8512, ZN => n8511);
   U6460 : OAI22_X1 port map( A1 => n7002, A2 => n9383, B1 => n6970, B2 => 
                           n9380, ZN => n8512);
   U6461 : AOI221_X1 port map( B1 => n9389, B2 => n6937, C1 => n9386, C2 => 
                           n6905, A => n8493, ZN => n8492);
   U6462 : OAI22_X1 port map( A1 => n7001, A2 => n9383, B1 => n6969, B2 => 
                           n9380, ZN => n8493);
   U6463 : AOI221_X1 port map( B1 => n9389, B2 => n6936, C1 => n9386, C2 => 
                           n6904, A => n8474, ZN => n8473);
   U6464 : OAI22_X1 port map( A1 => n7000, A2 => n9383, B1 => n6968, B2 => 
                           n9380, ZN => n8474);
   U6465 : AOI221_X1 port map( B1 => n9389, B2 => n6935, C1 => n9386, C2 => 
                           n6903, A => n8455, ZN => n8454);
   U6466 : OAI22_X1 port map( A1 => n6999, A2 => n9383, B1 => n6967, B2 => 
                           n9380, ZN => n8455);
   U6467 : AOI221_X1 port map( B1 => n9389, B2 => n6934, C1 => n9386, C2 => 
                           n6902, A => n8436, ZN => n8435);
   U6468 : OAI22_X1 port map( A1 => n6998, A2 => n9383, B1 => n6966, B2 => 
                           n9380, ZN => n8436);
   U6469 : AOI221_X1 port map( B1 => n9389, B2 => n6933, C1 => n9386, C2 => 
                           n6901, A => n8417, ZN => n8416);
   U6470 : OAI22_X1 port map( A1 => n6997, A2 => n9383, B1 => n6965, B2 => 
                           n9380, ZN => n8417);
   U6471 : AOI221_X1 port map( B1 => n9389, B2 => n6932, C1 => n9386, C2 => 
                           n6900, A => n8398, ZN => n8397);
   U6472 : OAI22_X1 port map( A1 => n6996, A2 => n9383, B1 => n6964, B2 => 
                           n9380, ZN => n8398);
   U6473 : AOI221_X1 port map( B1 => n9389, B2 => n6931, C1 => n9386, C2 => 
                           n6899, A => n8379, ZN => n8378);
   U6474 : OAI22_X1 port map( A1 => n6995, A2 => n9383, B1 => n6963, B2 => 
                           n9380, ZN => n8379);
   U6475 : AOI221_X1 port map( B1 => n9341, B2 => n6515, C1 => n9338, C2 => 
                           n6547, A => n8387, ZN => n8386);
   U6476 : OAI22_X1 port map( A1 => n6471, A2 => n9335, B1 => n6503, B2 => 
                           n9332, ZN => n8387);
   U6477 : AOI221_X1 port map( B1 => n9389, B2 => n6930, C1 => n9386, C2 => 
                           n6898, A => n8360, ZN => n8359);
   U6478 : OAI22_X1 port map( A1 => n6994, A2 => n9383, B1 => n6962, B2 => 
                           n9380, ZN => n8360);
   U6479 : AOI221_X1 port map( B1 => n9341, B2 => n6514, C1 => n9338, C2 => 
                           n6546, A => n8368, ZN => n8367);
   U6480 : OAI22_X1 port map( A1 => n6470, A2 => n9335, B1 => n6502, B2 => 
                           n9332, ZN => n8368);
   U6481 : AOI221_X1 port map( B1 => n9389, B2 => n6929, C1 => n9386, C2 => 
                           n6897, A => n8341, ZN => n8340);
   U6482 : OAI22_X1 port map( A1 => n6993, A2 => n9383, B1 => n6961, B2 => 
                           n9380, ZN => n8341);
   U6483 : AOI221_X1 port map( B1 => n9341, B2 => n6513, C1 => n9338, C2 => 
                           n6545, A => n8349, ZN => n8348);
   U6484 : OAI22_X1 port map( A1 => n6469, A2 => n9335, B1 => n6501, B2 => 
                           n9332, ZN => n8349);
   U6485 : AOI221_X1 port map( B1 => n9389, B2 => n6928, C1 => n9386, C2 => 
                           n6896, A => n8322, ZN => n8321);
   U6486 : OAI22_X1 port map( A1 => n6992, A2 => n9383, B1 => n6960, B2 => 
                           n9380, ZN => n8322);
   U6487 : AOI221_X1 port map( B1 => n9390, B2 => n6927, C1 => n9387, C2 => 
                           n6895, A => n8303, ZN => n8302);
   U6488 : OAI22_X1 port map( A1 => n6991, A2 => n9384, B1 => n6959, B2 => 
                           n9381, ZN => n8303);
   U6489 : AOI221_X1 port map( B1 => n9390, B2 => n6926, C1 => n9387, C2 => 
                           n6894, A => n8284, ZN => n8283);
   U6490 : OAI22_X1 port map( A1 => n6990, A2 => n9384, B1 => n6958, B2 => 
                           n9381, ZN => n8284);
   U6491 : AOI221_X1 port map( B1 => n9390, B2 => n6925, C1 => n9387, C2 => 
                           n6893, A => n8265, ZN => n8264);
   U6492 : OAI22_X1 port map( A1 => n6989, A2 => n9384, B1 => n6957, B2 => 
                           n9381, ZN => n8265);
   U6493 : AOI221_X1 port map( B1 => n9390, B2 => n6924, C1 => n9387, C2 => 
                           n6892, A => n8246, ZN => n8245);
   U6494 : OAI22_X1 port map( A1 => n6988, A2 => n9384, B1 => n6956, B2 => 
                           n9381, ZN => n8246);
   U6495 : AOI221_X1 port map( B1 => n9390, B2 => n6923, C1 => n9387, C2 => 
                           n6891, A => n8227, ZN => n8226);
   U6496 : OAI22_X1 port map( A1 => n6987, A2 => n9384, B1 => n6955, B2 => 
                           n9381, ZN => n8227);
   U6497 : AOI221_X1 port map( B1 => n9342, B2 => n6507, C1 => n9339, C2 => 
                           n6539, A => n8235, ZN => n8234);
   U6498 : OAI22_X1 port map( A1 => n6468, A2 => n9336, B1 => n6495, B2 => 
                           n9333, ZN => n8235);
   U6499 : AOI221_X1 port map( B1 => n9390, B2 => n6922, C1 => n9387, C2 => 
                           n6890, A => n8208, ZN => n8207);
   U6500 : OAI22_X1 port map( A1 => n6986, A2 => n9384, B1 => n6954, B2 => 
                           n9381, ZN => n8208);
   U6501 : AOI221_X1 port map( B1 => n9342, B2 => n6506, C1 => n9339, C2 => 
                           n6538, A => n8216, ZN => n8215);
   U6502 : OAI22_X1 port map( A1 => n6467, A2 => n9336, B1 => n6494, B2 => 
                           n9333, ZN => n8216);
   U6503 : AOI221_X1 port map( B1 => n9390, B2 => n6921, C1 => n9387, C2 => 
                           n6889, A => n8189, ZN => n8188);
   U6504 : OAI22_X1 port map( A1 => n6985, A2 => n9384, B1 => n6953, B2 => 
                           n9381, ZN => n8189);
   U6505 : AOI221_X1 port map( B1 => n9342, B2 => n6505, C1 => n9339, C2 => 
                           n6537, A => n8197, ZN => n8196);
   U6506 : OAI22_X1 port map( A1 => n6466, A2 => n9336, B1 => n6493, B2 => 
                           n9333, ZN => n8197);
   U6507 : AOI221_X1 port map( B1 => n9390, B2 => n6920, C1 => n9387, C2 => 
                           n6888, A => n8140, ZN => n8137);
   U6508 : OAI22_X1 port map( A1 => n6984, A2 => n9384, B1 => n6952, B2 => 
                           n9381, ZN => n8140);
   U6509 : AOI221_X1 port map( B1 => n9342, B2 => n6504, C1 => n9339, C2 => 
                           n6536, A => n8164, ZN => n8161);
   U6510 : OAI22_X1 port map( A1 => n6465, A2 => n9336, B1 => n6492, B2 => 
                           n9333, ZN => n8164);
   U6511 : AOI221_X1 port map( B1 => n9490, B2 => n6951, C1 => n9487, C2 => 
                           n6919, A => n8106, ZN => n8105);
   U6512 : OAI22_X1 port map( A1 => n7015, A2 => n9484, B1 => n6983, B2 => 
                           n9481, ZN => n8106);
   U6513 : AOI221_X1 port map( B1 => n9490, B2 => n6950, C1 => n9487, C2 => 
                           n6918, A => n8087, ZN => n8086);
   U6514 : OAI22_X1 port map( A1 => n7014, A2 => n9484, B1 => n6982, B2 => 
                           n9481, ZN => n8087);
   U6515 : AOI221_X1 port map( B1 => n9490, B2 => n6949, C1 => n9487, C2 => 
                           n6917, A => n8068, ZN => n8067);
   U6516 : OAI22_X1 port map( A1 => n7013, A2 => n9484, B1 => n6981, B2 => 
                           n9481, ZN => n8068);
   U6517 : AOI221_X1 port map( B1 => n9490, B2 => n6948, C1 => n9487, C2 => 
                           n6916, A => n8049, ZN => n8048);
   U6518 : OAI22_X1 port map( A1 => n7012, A2 => n9484, B1 => n6980, B2 => 
                           n9481, ZN => n8049);
   U6519 : AOI221_X1 port map( B1 => n9490, B2 => n6947, C1 => n9487, C2 => 
                           n6915, A => n8030, ZN => n8029);
   U6520 : OAI22_X1 port map( A1 => n7011, A2 => n9484, B1 => n6979, B2 => 
                           n9481, ZN => n8030);
   U6521 : AOI221_X1 port map( B1 => n9490, B2 => n6946, C1 => n9487, C2 => 
                           n6914, A => n8011, ZN => n8010);
   U6522 : OAI22_X1 port map( A1 => n7010, A2 => n9484, B1 => n6978, B2 => 
                           n9481, ZN => n8011);
   U6523 : AOI221_X1 port map( B1 => n9490, B2 => n6945, C1 => n9487, C2 => 
                           n6913, A => n7992, ZN => n7991);
   U6524 : OAI22_X1 port map( A1 => n7009, A2 => n9484, B1 => n6977, B2 => 
                           n9481, ZN => n7992);
   U6525 : AOI221_X1 port map( B1 => n9490, B2 => n6944, C1 => n9487, C2 => 
                           n6912, A => n7973, ZN => n7972);
   U6526 : OAI22_X1 port map( A1 => n7008, A2 => n9484, B1 => n6976, B2 => 
                           n9481, ZN => n7973);
   U6527 : AOI221_X1 port map( B1 => n9490, B2 => n6943, C1 => n9487, C2 => 
                           n6911, A => n7954, ZN => n7953);
   U6528 : OAI22_X1 port map( A1 => n7007, A2 => n9484, B1 => n6975, B2 => 
                           n9481, ZN => n7954);
   U6529 : AOI221_X1 port map( B1 => n9490, B2 => n6942, C1 => n9487, C2 => 
                           n6910, A => n7935, ZN => n7934);
   U6530 : OAI22_X1 port map( A1 => n7006, A2 => n9484, B1 => n6974, B2 => 
                           n9481, ZN => n7935);
   U6531 : AOI221_X1 port map( B1 => n9490, B2 => n6941, C1 => n9487, C2 => 
                           n6909, A => n7916, ZN => n7915);
   U6532 : OAI22_X1 port map( A1 => n7005, A2 => n9484, B1 => n6973, B2 => 
                           n9481, ZN => n7916);
   U6533 : AOI221_X1 port map( B1 => n9490, B2 => n6940, C1 => n9487, C2 => 
                           n6908, A => n7897, ZN => n7896);
   U6534 : OAI22_X1 port map( A1 => n7004, A2 => n9484, B1 => n6972, B2 => 
                           n9481, ZN => n7897);
   U6535 : AOI221_X1 port map( B1 => n9491, B2 => n6939, C1 => n9488, C2 => 
                           n6907, A => n7878, ZN => n7877);
   U6536 : OAI22_X1 port map( A1 => n7003, A2 => n9485, B1 => n6971, B2 => 
                           n9482, ZN => n7878);
   U6537 : AOI221_X1 port map( B1 => n9491, B2 => n6938, C1 => n9488, C2 => 
                           n6906, A => n7859, ZN => n7858);
   U6538 : OAI22_X1 port map( A1 => n7002, A2 => n9485, B1 => n6970, B2 => 
                           n9482, ZN => n7859);
   U6539 : AOI221_X1 port map( B1 => n9491, B2 => n6937, C1 => n9488, C2 => 
                           n6905, A => n7840, ZN => n7839);
   U6540 : OAI22_X1 port map( A1 => n7001, A2 => n9485, B1 => n6969, B2 => 
                           n9482, ZN => n7840);
   U6541 : AOI221_X1 port map( B1 => n9491, B2 => n6936, C1 => n9488, C2 => 
                           n6904, A => n7821, ZN => n7820);
   U6542 : OAI22_X1 port map( A1 => n7000, A2 => n9485, B1 => n6968, B2 => 
                           n9482, ZN => n7821);
   U6543 : AOI221_X1 port map( B1 => n9491, B2 => n6935, C1 => n9488, C2 => 
                           n6903, A => n7802, ZN => n7801);
   U6544 : OAI22_X1 port map( A1 => n6999, A2 => n9485, B1 => n6967, B2 => 
                           n9482, ZN => n7802);
   U6545 : AOI221_X1 port map( B1 => n9491, B2 => n6934, C1 => n9488, C2 => 
                           n6902, A => n7783, ZN => n7782);
   U6546 : OAI22_X1 port map( A1 => n6998, A2 => n9485, B1 => n6966, B2 => 
                           n9482, ZN => n7783);
   U6547 : AOI221_X1 port map( B1 => n9491, B2 => n6933, C1 => n9488, C2 => 
                           n6901, A => n7764, ZN => n7763);
   U6548 : OAI22_X1 port map( A1 => n6997, A2 => n9485, B1 => n6965, B2 => 
                           n9482, ZN => n7764);
   U6549 : AOI221_X1 port map( B1 => n9491, B2 => n6932, C1 => n9488, C2 => 
                           n6900, A => n7745, ZN => n7744);
   U6550 : OAI22_X1 port map( A1 => n6996, A2 => n9485, B1 => n6964, B2 => 
                           n9482, ZN => n7745);
   U6551 : AOI221_X1 port map( B1 => n9491, B2 => n6931, C1 => n9488, C2 => 
                           n6899, A => n7726, ZN => n7725);
   U6552 : OAI22_X1 port map( A1 => n6995, A2 => n9485, B1 => n6963, B2 => 
                           n9482, ZN => n7726);
   U6553 : AOI221_X1 port map( B1 => n9443, B2 => n6515, C1 => n9440, C2 => 
                           n6547, A => n7734, ZN => n7733);
   U6554 : OAI22_X1 port map( A1 => n6471, A2 => n9437, B1 => n6503, B2 => 
                           n9434, ZN => n7734);
   U6555 : AOI221_X1 port map( B1 => n9491, B2 => n6930, C1 => n9488, C2 => 
                           n6898, A => n7707, ZN => n7706);
   U6556 : OAI22_X1 port map( A1 => n6994, A2 => n9485, B1 => n6962, B2 => 
                           n9482, ZN => n7707);
   U6557 : AOI221_X1 port map( B1 => n9443, B2 => n6514, C1 => n9440, C2 => 
                           n6546, A => n7715, ZN => n7714);
   U6558 : OAI22_X1 port map( A1 => n6470, A2 => n9437, B1 => n6502, B2 => 
                           n9434, ZN => n7715);
   U6559 : AOI221_X1 port map( B1 => n9491, B2 => n6929, C1 => n9488, C2 => 
                           n6897, A => n7688, ZN => n7687);
   U6560 : OAI22_X1 port map( A1 => n6993, A2 => n9485, B1 => n6961, B2 => 
                           n9482, ZN => n7688);
   U6561 : AOI221_X1 port map( B1 => n9443, B2 => n6513, C1 => n9440, C2 => 
                           n6545, A => n7696, ZN => n7695);
   U6562 : OAI22_X1 port map( A1 => n6469, A2 => n9437, B1 => n6501, B2 => 
                           n9434, ZN => n7696);
   U6563 : AOI221_X1 port map( B1 => n9491, B2 => n6928, C1 => n9488, C2 => 
                           n6896, A => n7669, ZN => n7668);
   U6564 : OAI22_X1 port map( A1 => n6992, A2 => n9485, B1 => n6960, B2 => 
                           n9482, ZN => n7669);
   U6565 : AOI221_X1 port map( B1 => n9492, B2 => n6927, C1 => n9489, C2 => 
                           n6895, A => n7650, ZN => n7649);
   U6566 : OAI22_X1 port map( A1 => n6991, A2 => n9486, B1 => n6959, B2 => 
                           n9483, ZN => n7650);
   U6567 : AOI221_X1 port map( B1 => n9492, B2 => n6926, C1 => n9489, C2 => 
                           n6894, A => n7631, ZN => n7630);
   U6568 : OAI22_X1 port map( A1 => n6990, A2 => n9486, B1 => n6958, B2 => 
                           n9483, ZN => n7631);
   U6569 : AOI221_X1 port map( B1 => n9492, B2 => n6925, C1 => n9489, C2 => 
                           n6893, A => n7612, ZN => n7611);
   U6570 : OAI22_X1 port map( A1 => n6989, A2 => n9486, B1 => n6957, B2 => 
                           n9483, ZN => n7612);
   U6571 : AOI221_X1 port map( B1 => n9492, B2 => n6924, C1 => n9489, C2 => 
                           n6892, A => n7593, ZN => n7592);
   U6572 : OAI22_X1 port map( A1 => n6988, A2 => n9486, B1 => n6956, B2 => 
                           n9483, ZN => n7593);
   U6573 : AOI221_X1 port map( B1 => n9492, B2 => n6923, C1 => n9489, C2 => 
                           n6891, A => n7574, ZN => n7573);
   U6574 : OAI22_X1 port map( A1 => n6987, A2 => n9486, B1 => n6955, B2 => 
                           n9483, ZN => n7574);
   U6575 : AOI221_X1 port map( B1 => n9444, B2 => n6507, C1 => n9441, C2 => 
                           n6539, A => n7582, ZN => n7581);
   U6576 : OAI22_X1 port map( A1 => n6468, A2 => n9438, B1 => n6495, B2 => 
                           n9435, ZN => n7582);
   U6577 : AOI221_X1 port map( B1 => n9492, B2 => n6922, C1 => n9489, C2 => 
                           n6890, A => n7555, ZN => n7554);
   U6578 : OAI22_X1 port map( A1 => n6986, A2 => n9486, B1 => n6954, B2 => 
                           n9483, ZN => n7555);
   U6579 : AOI221_X1 port map( B1 => n9444, B2 => n6506, C1 => n9441, C2 => 
                           n6538, A => n7563, ZN => n7562);
   U6580 : OAI22_X1 port map( A1 => n6467, A2 => n9438, B1 => n6494, B2 => 
                           n9435, ZN => n7563);
   U6581 : AOI221_X1 port map( B1 => n9492, B2 => n6921, C1 => n9489, C2 => 
                           n6889, A => n7536, ZN => n7535);
   U6582 : OAI22_X1 port map( A1 => n6985, A2 => n9486, B1 => n6953, B2 => 
                           n9483, ZN => n7536);
   U6583 : AOI221_X1 port map( B1 => n9444, B2 => n6505, C1 => n9441, C2 => 
                           n6537, A => n7544, ZN => n7543);
   U6584 : OAI22_X1 port map( A1 => n6466, A2 => n9438, B1 => n6493, B2 => 
                           n9435, ZN => n7544);
   U6585 : AOI221_X1 port map( B1 => n9492, B2 => n6920, C1 => n9489, C2 => 
                           n6888, A => n7487, ZN => n7484);
   U6586 : OAI22_X1 port map( A1 => n6984, A2 => n9486, B1 => n6952, B2 => 
                           n9483, ZN => n7487);
   U6587 : AOI221_X1 port map( B1 => n9444, B2 => n6504, C1 => n9441, C2 => 
                           n6536, A => n7511, ZN => n7508);
   U6588 : OAI22_X1 port map( A1 => n6465, A2 => n9438, B1 => n6492, B2 => 
                           n9435, ZN => n7511);
   U6589 : AOI221_X1 port map( B1 => n9376, B2 => n7079, C1 => n9373, C2 => 
                           n7047, A => n8764, ZN => n8757);
   U6590 : OAI22_X1 port map( A1 => n7143, A2 => n9370, B1 => n7111, B2 => 
                           n9367, ZN => n8764);
   U6591 : AOI221_X1 port map( B1 => n9376, B2 => n7078, C1 => n9373, C2 => 
                           n7046, A => n8741, ZN => n8738);
   U6592 : OAI22_X1 port map( A1 => n7142, A2 => n9370, B1 => n7110, B2 => 
                           n9367, ZN => n8741);
   U6593 : AOI221_X1 port map( B1 => n9376, B2 => n7077, C1 => n9373, C2 => 
                           n7045, A => n8722, ZN => n8719);
   U6594 : OAI22_X1 port map( A1 => n7141, A2 => n9370, B1 => n7109, B2 => 
                           n9367, ZN => n8722);
   U6595 : AOI221_X1 port map( B1 => n9376, B2 => n7076, C1 => n9373, C2 => 
                           n7044, A => n8703, ZN => n8700);
   U6596 : OAI22_X1 port map( A1 => n7140, A2 => n9370, B1 => n7108, B2 => 
                           n9367, ZN => n8703);
   U6597 : AOI221_X1 port map( B1 => n9376, B2 => n7075, C1 => n9373, C2 => 
                           n7043, A => n8684, ZN => n8681);
   U6598 : OAI22_X1 port map( A1 => n7139, A2 => n9370, B1 => n7107, B2 => 
                           n9367, ZN => n8684);
   U6599 : AOI221_X1 port map( B1 => n9376, B2 => n7074, C1 => n9373, C2 => 
                           n7042, A => n8665, ZN => n8662);
   U6600 : OAI22_X1 port map( A1 => n7138, A2 => n9370, B1 => n7106, B2 => 
                           n9367, ZN => n8665);
   U6601 : AOI221_X1 port map( B1 => n9376, B2 => n7073, C1 => n9373, C2 => 
                           n7041, A => n8646, ZN => n8643);
   U6602 : OAI22_X1 port map( A1 => n7137, A2 => n9370, B1 => n7105, B2 => 
                           n9367, ZN => n8646);
   U6603 : AOI221_X1 port map( B1 => n9376, B2 => n7072, C1 => n9373, C2 => 
                           n7040, A => n8627, ZN => n8624);
   U6604 : OAI22_X1 port map( A1 => n7136, A2 => n9370, B1 => n7104, B2 => 
                           n9367, ZN => n8627);
   U6605 : AOI221_X1 port map( B1 => n9376, B2 => n7071, C1 => n9373, C2 => 
                           n7039, A => n8608, ZN => n8605);
   U6606 : OAI22_X1 port map( A1 => n7135, A2 => n9370, B1 => n7103, B2 => 
                           n9367, ZN => n8608);
   U6607 : AOI221_X1 port map( B1 => n9376, B2 => n7070, C1 => n9373, C2 => 
                           n7038, A => n8589, ZN => n8586);
   U6608 : OAI22_X1 port map( A1 => n7134, A2 => n9370, B1 => n7102, B2 => 
                           n9367, ZN => n8589);
   U6609 : AOI221_X1 port map( B1 => n9376, B2 => n7069, C1 => n9373, C2 => 
                           n7037, A => n8570, ZN => n8567);
   U6610 : OAI22_X1 port map( A1 => n7133, A2 => n9370, B1 => n7101, B2 => 
                           n9367, ZN => n8570);
   U6611 : AOI221_X1 port map( B1 => n9376, B2 => n7068, C1 => n9373, C2 => 
                           n7036, A => n8551, ZN => n8548);
   U6612 : OAI22_X1 port map( A1 => n7132, A2 => n9370, B1 => n7100, B2 => 
                           n9367, ZN => n8551);
   U6613 : AOI221_X1 port map( B1 => n9377, B2 => n7067, C1 => n9374, C2 => 
                           n7035, A => n8532, ZN => n8529);
   U6614 : OAI22_X1 port map( A1 => n7131, A2 => n9371, B1 => n7099, B2 => 
                           n9368, ZN => n8532);
   U6615 : AOI221_X1 port map( B1 => n9377, B2 => n7066, C1 => n9374, C2 => 
                           n7034, A => n8513, ZN => n8510);
   U6616 : OAI22_X1 port map( A1 => n7130, A2 => n9371, B1 => n7098, B2 => 
                           n9368, ZN => n8513);
   U6617 : AOI221_X1 port map( B1 => n9377, B2 => n7065, C1 => n9374, C2 => 
                           n7033, A => n8494, ZN => n8491);
   U6618 : OAI22_X1 port map( A1 => n7129, A2 => n9371, B1 => n7097, B2 => 
                           n9368, ZN => n8494);
   U6619 : AOI221_X1 port map( B1 => n9377, B2 => n7064, C1 => n9374, C2 => 
                           n7032, A => n8475, ZN => n8472);
   U6620 : OAI22_X1 port map( A1 => n7128, A2 => n9371, B1 => n7096, B2 => 
                           n9368, ZN => n8475);
   U6621 : AOI221_X1 port map( B1 => n9377, B2 => n7063, C1 => n9374, C2 => 
                           n7031, A => n8456, ZN => n8453);
   U6622 : OAI22_X1 port map( A1 => n7127, A2 => n9371, B1 => n7095, B2 => 
                           n9368, ZN => n8456);
   U6623 : AOI221_X1 port map( B1 => n9377, B2 => n7062, C1 => n9374, C2 => 
                           n7030, A => n8437, ZN => n8434);
   U6624 : OAI22_X1 port map( A1 => n7126, A2 => n9371, B1 => n7094, B2 => 
                           n9368, ZN => n8437);
   U6625 : AOI221_X1 port map( B1 => n9377, B2 => n7061, C1 => n9374, C2 => 
                           n7029, A => n8418, ZN => n8415);
   U6626 : OAI22_X1 port map( A1 => n7125, A2 => n9371, B1 => n7093, B2 => 
                           n9368, ZN => n8418);
   U6627 : AOI221_X1 port map( B1 => n9377, B2 => n7060, C1 => n9374, C2 => 
                           n7028, A => n8399, ZN => n8396);
   U6628 : OAI22_X1 port map( A1 => n7124, A2 => n9371, B1 => n7092, B2 => 
                           n9368, ZN => n8399);
   U6629 : AOI221_X1 port map( B1 => n9377, B2 => n7059, C1 => n9374, C2 => 
                           n7027, A => n8380, ZN => n8377);
   U6630 : OAI22_X1 port map( A1 => n7123, A2 => n9371, B1 => n7091, B2 => 
                           n9368, ZN => n8380);
   U6631 : AOI221_X1 port map( B1 => n9377, B2 => n7058, C1 => n9374, C2 => 
                           n7026, A => n8361, ZN => n8358);
   U6632 : OAI22_X1 port map( A1 => n7122, A2 => n9371, B1 => n7090, B2 => 
                           n9368, ZN => n8361);
   U6633 : AOI221_X1 port map( B1 => n9377, B2 => n7057, C1 => n9374, C2 => 
                           n7025, A => n8342, ZN => n8339);
   U6634 : OAI22_X1 port map( A1 => n7121, A2 => n9371, B1 => n7089, B2 => 
                           n9368, ZN => n8342);
   U6635 : AOI221_X1 port map( B1 => n9377, B2 => n7056, C1 => n9374, C2 => 
                           n7024, A => n8323, ZN => n8320);
   U6636 : OAI22_X1 port map( A1 => n7120, A2 => n9371, B1 => n7088, B2 => 
                           n9368, ZN => n8323);
   U6637 : AOI221_X1 port map( B1 => n9478, B2 => n7079, C1 => n9475, C2 => 
                           n7047, A => n8111, ZN => n8104);
   U6638 : OAI22_X1 port map( A1 => n7143, A2 => n9472, B1 => n7111, B2 => 
                           n9469, ZN => n8111);
   U6639 : AOI221_X1 port map( B1 => n9478, B2 => n7078, C1 => n9475, C2 => 
                           n7046, A => n8088, ZN => n8085);
   U6640 : OAI22_X1 port map( A1 => n7142, A2 => n9472, B1 => n7110, B2 => 
                           n9469, ZN => n8088);
   U6641 : AOI221_X1 port map( B1 => n9478, B2 => n7077, C1 => n9475, C2 => 
                           n7045, A => n8069, ZN => n8066);
   U6642 : OAI22_X1 port map( A1 => n7141, A2 => n9472, B1 => n7109, B2 => 
                           n9469, ZN => n8069);
   U6643 : AOI221_X1 port map( B1 => n9478, B2 => n7076, C1 => n9475, C2 => 
                           n7044, A => n8050, ZN => n8047);
   U6644 : OAI22_X1 port map( A1 => n7140, A2 => n9472, B1 => n7108, B2 => 
                           n9469, ZN => n8050);
   U6645 : AOI221_X1 port map( B1 => n9478, B2 => n7075, C1 => n9475, C2 => 
                           n7043, A => n8031, ZN => n8028);
   U6646 : OAI22_X1 port map( A1 => n7139, A2 => n9472, B1 => n7107, B2 => 
                           n9469, ZN => n8031);
   U6647 : AOI221_X1 port map( B1 => n9478, B2 => n7074, C1 => n9475, C2 => 
                           n7042, A => n8012, ZN => n8009);
   U6648 : OAI22_X1 port map( A1 => n7138, A2 => n9472, B1 => n7106, B2 => 
                           n9469, ZN => n8012);
   U6649 : AOI221_X1 port map( B1 => n9478, B2 => n7073, C1 => n9475, C2 => 
                           n7041, A => n7993, ZN => n7990);
   U6650 : OAI22_X1 port map( A1 => n7137, A2 => n9472, B1 => n7105, B2 => 
                           n9469, ZN => n7993);
   U6651 : AOI221_X1 port map( B1 => n9478, B2 => n7072, C1 => n9475, C2 => 
                           n7040, A => n7974, ZN => n7971);
   U6652 : OAI22_X1 port map( A1 => n7136, A2 => n9472, B1 => n7104, B2 => 
                           n9469, ZN => n7974);
   U6653 : AOI221_X1 port map( B1 => n9478, B2 => n7071, C1 => n9475, C2 => 
                           n7039, A => n7955, ZN => n7952);
   U6654 : OAI22_X1 port map( A1 => n7135, A2 => n9472, B1 => n7103, B2 => 
                           n9469, ZN => n7955);
   U6655 : AOI221_X1 port map( B1 => n9478, B2 => n7070, C1 => n9475, C2 => 
                           n7038, A => n7936, ZN => n7933);
   U6656 : OAI22_X1 port map( A1 => n7134, A2 => n9472, B1 => n7102, B2 => 
                           n9469, ZN => n7936);
   U6657 : AOI221_X1 port map( B1 => n9478, B2 => n7069, C1 => n9475, C2 => 
                           n7037, A => n7917, ZN => n7914);
   U6658 : OAI22_X1 port map( A1 => n7133, A2 => n9472, B1 => n7101, B2 => 
                           n9469, ZN => n7917);
   U6659 : AOI221_X1 port map( B1 => n9478, B2 => n7068, C1 => n9475, C2 => 
                           n7036, A => n7898, ZN => n7895);
   U6660 : OAI22_X1 port map( A1 => n7132, A2 => n9472, B1 => n7100, B2 => 
                           n9469, ZN => n7898);
   U6661 : AOI221_X1 port map( B1 => n9479, B2 => n7067, C1 => n9476, C2 => 
                           n7035, A => n7879, ZN => n7876);
   U6662 : OAI22_X1 port map( A1 => n7131, A2 => n9473, B1 => n7099, B2 => 
                           n9470, ZN => n7879);
   U6663 : AOI221_X1 port map( B1 => n9479, B2 => n7066, C1 => n9476, C2 => 
                           n7034, A => n7860, ZN => n7857);
   U6664 : OAI22_X1 port map( A1 => n7130, A2 => n9473, B1 => n7098, B2 => 
                           n9470, ZN => n7860);
   U6665 : AOI221_X1 port map( B1 => n9479, B2 => n7065, C1 => n9476, C2 => 
                           n7033, A => n7841, ZN => n7838);
   U6666 : OAI22_X1 port map( A1 => n7129, A2 => n9473, B1 => n7097, B2 => 
                           n9470, ZN => n7841);
   U6667 : AOI221_X1 port map( B1 => n9479, B2 => n7064, C1 => n9476, C2 => 
                           n7032, A => n7822, ZN => n7819);
   U6668 : OAI22_X1 port map( A1 => n7128, A2 => n9473, B1 => n7096, B2 => 
                           n9470, ZN => n7822);
   U6669 : AOI221_X1 port map( B1 => n9479, B2 => n7063, C1 => n9476, C2 => 
                           n7031, A => n7803, ZN => n7800);
   U6670 : OAI22_X1 port map( A1 => n7127, A2 => n9473, B1 => n7095, B2 => 
                           n9470, ZN => n7803);
   U6671 : AOI221_X1 port map( B1 => n9479, B2 => n7062, C1 => n9476, C2 => 
                           n7030, A => n7784, ZN => n7781);
   U6672 : OAI22_X1 port map( A1 => n7126, A2 => n9473, B1 => n7094, B2 => 
                           n9470, ZN => n7784);
   U6673 : AOI221_X1 port map( B1 => n9479, B2 => n7061, C1 => n9476, C2 => 
                           n7029, A => n7765, ZN => n7762);
   U6674 : OAI22_X1 port map( A1 => n7125, A2 => n9473, B1 => n7093, B2 => 
                           n9470, ZN => n7765);
   U6675 : AOI221_X1 port map( B1 => n9479, B2 => n7060, C1 => n9476, C2 => 
                           n7028, A => n7746, ZN => n7743);
   U6676 : OAI22_X1 port map( A1 => n7124, A2 => n9473, B1 => n7092, B2 => 
                           n9470, ZN => n7746);
   U6677 : AOI221_X1 port map( B1 => n9479, B2 => n7059, C1 => n9476, C2 => 
                           n7027, A => n7727, ZN => n7724);
   U6678 : OAI22_X1 port map( A1 => n7123, A2 => n9473, B1 => n7091, B2 => 
                           n9470, ZN => n7727);
   U6679 : AOI221_X1 port map( B1 => n9479, B2 => n7058, C1 => n9476, C2 => 
                           n7026, A => n7708, ZN => n7705);
   U6680 : OAI22_X1 port map( A1 => n7122, A2 => n9473, B1 => n7090, B2 => 
                           n9470, ZN => n7708);
   U6681 : AOI221_X1 port map( B1 => n9479, B2 => n7057, C1 => n9476, C2 => 
                           n7025, A => n7689, ZN => n7686);
   U6682 : OAI22_X1 port map( A1 => n7121, A2 => n9473, B1 => n7089, B2 => 
                           n9470, ZN => n7689);
   U6683 : AOI221_X1 port map( B1 => n9479, B2 => n7056, C1 => n9476, C2 => 
                           n7024, A => n7670, ZN => n7667);
   U6684 : OAI22_X1 port map( A1 => n7120, A2 => n9473, B1 => n7088, B2 => 
                           n9470, ZN => n7670);
   U6685 : AOI221_X1 port map( B1 => n9364, B2 => n7271, C1 => n9361, C2 => 
                           n7239, A => n8767, ZN => n8756);
   U6686 : OAI22_X1 port map( A1 => n7207, A2 => n9358, B1 => n7175, B2 => 
                           n9355, ZN => n8767);
   U6687 : AOI221_X1 port map( B1 => n9364, B2 => n7270, C1 => n9361, C2 => 
                           n7238, A => n8742, ZN => n8737);
   U6688 : OAI22_X1 port map( A1 => n7206, A2 => n9358, B1 => n7174, B2 => 
                           n9355, ZN => n8742);
   U6689 : AOI221_X1 port map( B1 => n9364, B2 => n7269, C1 => n9361, C2 => 
                           n7237, A => n8723, ZN => n8718);
   U6690 : OAI22_X1 port map( A1 => n7205, A2 => n9358, B1 => n7173, B2 => 
                           n9355, ZN => n8723);
   U6691 : AOI221_X1 port map( B1 => n9364, B2 => n7268, C1 => n9361, C2 => 
                           n7236, A => n8704, ZN => n8699);
   U6692 : OAI22_X1 port map( A1 => n7204, A2 => n9358, B1 => n7172, B2 => 
                           n9355, ZN => n8704);
   U6693 : AOI221_X1 port map( B1 => n9364, B2 => n7267, C1 => n9361, C2 => 
                           n7235, A => n8685, ZN => n8680);
   U6694 : OAI22_X1 port map( A1 => n7203, A2 => n9358, B1 => n7171, B2 => 
                           n9355, ZN => n8685);
   U6695 : AOI221_X1 port map( B1 => n9364, B2 => n7266, C1 => n9361, C2 => 
                           n7234, A => n8666, ZN => n8661);
   U6696 : OAI22_X1 port map( A1 => n7202, A2 => n9358, B1 => n7170, B2 => 
                           n9355, ZN => n8666);
   U6697 : AOI221_X1 port map( B1 => n9364, B2 => n7265, C1 => n9361, C2 => 
                           n7233, A => n8647, ZN => n8642);
   U6698 : OAI22_X1 port map( A1 => n7201, A2 => n9358, B1 => n7169, B2 => 
                           n9355, ZN => n8647);
   U6699 : AOI221_X1 port map( B1 => n9364, B2 => n7264, C1 => n9361, C2 => 
                           n7232, A => n8628, ZN => n8623);
   U6700 : OAI22_X1 port map( A1 => n7200, A2 => n9358, B1 => n7168, B2 => 
                           n9355, ZN => n8628);
   U6701 : AOI221_X1 port map( B1 => n9364, B2 => n7263, C1 => n9361, C2 => 
                           n7231, A => n8609, ZN => n8604);
   U6702 : OAI22_X1 port map( A1 => n7199, A2 => n9358, B1 => n7167, B2 => 
                           n9355, ZN => n8609);
   U6703 : AOI221_X1 port map( B1 => n9364, B2 => n7262, C1 => n9361, C2 => 
                           n7230, A => n8590, ZN => n8585);
   U6704 : OAI22_X1 port map( A1 => n7198, A2 => n9358, B1 => n7166, B2 => 
                           n9355, ZN => n8590);
   U6705 : AOI221_X1 port map( B1 => n9364, B2 => n7261, C1 => n9361, C2 => 
                           n7229, A => n8571, ZN => n8566);
   U6706 : OAI22_X1 port map( A1 => n7197, A2 => n9358, B1 => n7165, B2 => 
                           n9355, ZN => n8571);
   U6707 : AOI221_X1 port map( B1 => n9364, B2 => n7260, C1 => n9361, C2 => 
                           n7228, A => n8552, ZN => n8547);
   U6708 : OAI22_X1 port map( A1 => n7196, A2 => n9358, B1 => n7164, B2 => 
                           n9355, ZN => n8552);
   U6709 : AOI221_X1 port map( B1 => n9365, B2 => n7259, C1 => n9362, C2 => 
                           n7227, A => n8533, ZN => n8528);
   U6710 : OAI22_X1 port map( A1 => n7195, A2 => n9359, B1 => n7163, B2 => 
                           n9356, ZN => n8533);
   U6711 : AOI221_X1 port map( B1 => n9365, B2 => n7258, C1 => n9362, C2 => 
                           n7226, A => n8514, ZN => n8509);
   U6712 : OAI22_X1 port map( A1 => n7194, A2 => n9359, B1 => n7162, B2 => 
                           n9356, ZN => n8514);
   U6713 : AOI221_X1 port map( B1 => n9365, B2 => n7257, C1 => n9362, C2 => 
                           n7225, A => n8495, ZN => n8490);
   U6714 : OAI22_X1 port map( A1 => n7193, A2 => n9359, B1 => n7161, B2 => 
                           n9356, ZN => n8495);
   U6715 : AOI221_X1 port map( B1 => n9365, B2 => n7256, C1 => n9362, C2 => 
                           n7224, A => n8476, ZN => n8471);
   U6716 : OAI22_X1 port map( A1 => n7192, A2 => n9359, B1 => n7160, B2 => 
                           n9356, ZN => n8476);
   U6717 : AOI221_X1 port map( B1 => n9365, B2 => n7255, C1 => n9362, C2 => 
                           n7223, A => n8457, ZN => n8452);
   U6718 : OAI22_X1 port map( A1 => n7191, A2 => n9359, B1 => n7159, B2 => 
                           n9356, ZN => n8457);
   U6719 : AOI221_X1 port map( B1 => n9365, B2 => n7254, C1 => n9362, C2 => 
                           n7222, A => n8438, ZN => n8433);
   U6720 : OAI22_X1 port map( A1 => n7190, A2 => n9359, B1 => n7158, B2 => 
                           n9356, ZN => n8438);
   U6721 : AOI221_X1 port map( B1 => n9365, B2 => n7253, C1 => n9362, C2 => 
                           n7221, A => n8419, ZN => n8414);
   U6722 : OAI22_X1 port map( A1 => n7189, A2 => n9359, B1 => n7157, B2 => 
                           n9356, ZN => n8419);
   U6723 : AOI221_X1 port map( B1 => n9365, B2 => n7252, C1 => n9362, C2 => 
                           n7220, A => n8400, ZN => n8395);
   U6724 : OAI22_X1 port map( A1 => n7188, A2 => n9359, B1 => n7156, B2 => 
                           n9356, ZN => n8400);
   U6725 : AOI221_X1 port map( B1 => n9365, B2 => n7251, C1 => n9362, C2 => 
                           n7219, A => n8381, ZN => n8376);
   U6726 : OAI22_X1 port map( A1 => n7187, A2 => n9359, B1 => n7155, B2 => 
                           n9356, ZN => n8381);
   U6727 : AOI221_X1 port map( B1 => n9365, B2 => n7250, C1 => n9362, C2 => 
                           n7218, A => n8362, ZN => n8357);
   U6728 : OAI22_X1 port map( A1 => n7186, A2 => n9359, B1 => n7154, B2 => 
                           n9356, ZN => n8362);
   U6729 : AOI221_X1 port map( B1 => n9365, B2 => n7249, C1 => n9362, C2 => 
                           n7217, A => n8343, ZN => n8338);
   U6730 : OAI22_X1 port map( A1 => n7185, A2 => n9359, B1 => n7153, B2 => 
                           n9356, ZN => n8343);
   U6731 : AOI221_X1 port map( B1 => n9365, B2 => n7248, C1 => n9362, C2 => 
                           n7216, A => n8324, ZN => n8319);
   U6732 : OAI22_X1 port map( A1 => n7184, A2 => n9359, B1 => n7152, B2 => 
                           n9356, ZN => n8324);
   U6733 : AOI221_X1 port map( B1 => n9366, B2 => n7247, C1 => n9363, C2 => 
                           n7215, A => n8305, ZN => n8300);
   U6734 : OAI22_X1 port map( A1 => n7183, A2 => n9360, B1 => n7151, B2 => 
                           n9357, ZN => n8305);
   U6735 : AOI221_X1 port map( B1 => n9366, B2 => n7246, C1 => n9363, C2 => 
                           n7214, A => n8286, ZN => n8281);
   U6736 : OAI22_X1 port map( A1 => n7182, A2 => n9360, B1 => n7150, B2 => 
                           n9357, ZN => n8286);
   U6737 : AOI221_X1 port map( B1 => n9366, B2 => n7245, C1 => n9363, C2 => 
                           n7213, A => n8267, ZN => n8262);
   U6738 : OAI22_X1 port map( A1 => n7181, A2 => n9360, B1 => n7149, B2 => 
                           n9357, ZN => n8267);
   U6739 : AOI221_X1 port map( B1 => n9366, B2 => n7244, C1 => n9363, C2 => 
                           n7212, A => n8248, ZN => n8243);
   U6740 : OAI22_X1 port map( A1 => n7180, A2 => n9360, B1 => n7148, B2 => 
                           n9357, ZN => n8248);
   U6741 : AOI221_X1 port map( B1 => n9366, B2 => n7243, C1 => n9363, C2 => 
                           n7211, A => n8229, ZN => n8224);
   U6742 : OAI22_X1 port map( A1 => n7179, A2 => n9360, B1 => n7147, B2 => 
                           n9357, ZN => n8229);
   U6743 : AOI221_X1 port map( B1 => n9366, B2 => n7242, C1 => n9363, C2 => 
                           n7210, A => n8210, ZN => n8205);
   U6744 : OAI22_X1 port map( A1 => n7178, A2 => n9360, B1 => n7146, B2 => 
                           n9357, ZN => n8210);
   U6745 : AOI221_X1 port map( B1 => n9366, B2 => n7241, C1 => n9363, C2 => 
                           n7209, A => n8191, ZN => n8186);
   U6746 : OAI22_X1 port map( A1 => n7177, A2 => n9360, B1 => n7145, B2 => 
                           n9357, ZN => n8191);
   U6747 : AOI221_X1 port map( B1 => n9366, B2 => n7240, C1 => n9363, C2 => 
                           n7208, A => n8150, ZN => n8135);
   U6748 : OAI22_X1 port map( A1 => n7176, A2 => n9360, B1 => n7144, B2 => 
                           n9357, ZN => n8150);
   U6749 : AOI221_X1 port map( B1 => n9466, B2 => n7271, C1 => n9463, C2 => 
                           n7239, A => n8114, ZN => n8103);
   U6750 : OAI22_X1 port map( A1 => n7207, A2 => n9460, B1 => n7175, B2 => 
                           n9457, ZN => n8114);
   U6751 : AOI221_X1 port map( B1 => n9466, B2 => n7270, C1 => n9463, C2 => 
                           n7238, A => n8089, ZN => n8084);
   U6752 : OAI22_X1 port map( A1 => n7206, A2 => n9460, B1 => n7174, B2 => 
                           n9457, ZN => n8089);
   U6753 : AOI221_X1 port map( B1 => n9466, B2 => n7269, C1 => n9463, C2 => 
                           n7237, A => n8070, ZN => n8065);
   U6754 : OAI22_X1 port map( A1 => n7205, A2 => n9460, B1 => n7173, B2 => 
                           n9457, ZN => n8070);
   U6755 : AOI221_X1 port map( B1 => n9466, B2 => n7268, C1 => n9463, C2 => 
                           n7236, A => n8051, ZN => n8046);
   U6756 : OAI22_X1 port map( A1 => n7204, A2 => n9460, B1 => n7172, B2 => 
                           n9457, ZN => n8051);
   U6757 : AOI221_X1 port map( B1 => n9466, B2 => n7267, C1 => n9463, C2 => 
                           n7235, A => n8032, ZN => n8027);
   U6758 : OAI22_X1 port map( A1 => n7203, A2 => n9460, B1 => n7171, B2 => 
                           n9457, ZN => n8032);
   U6759 : AOI221_X1 port map( B1 => n9466, B2 => n7266, C1 => n9463, C2 => 
                           n7234, A => n8013, ZN => n8008);
   U6760 : OAI22_X1 port map( A1 => n7202, A2 => n9460, B1 => n7170, B2 => 
                           n9457, ZN => n8013);
   U6761 : AOI221_X1 port map( B1 => n9466, B2 => n7265, C1 => n9463, C2 => 
                           n7233, A => n7994, ZN => n7989);
   U6762 : OAI22_X1 port map( A1 => n7201, A2 => n9460, B1 => n7169, B2 => 
                           n9457, ZN => n7994);
   U6763 : AOI221_X1 port map( B1 => n9466, B2 => n7264, C1 => n9463, C2 => 
                           n7232, A => n7975, ZN => n7970);
   U6764 : OAI22_X1 port map( A1 => n7200, A2 => n9460, B1 => n7168, B2 => 
                           n9457, ZN => n7975);
   U6765 : AOI221_X1 port map( B1 => n9466, B2 => n7263, C1 => n9463, C2 => 
                           n7231, A => n7956, ZN => n7951);
   U6766 : OAI22_X1 port map( A1 => n7199, A2 => n9460, B1 => n7167, B2 => 
                           n9457, ZN => n7956);
   U6767 : AOI221_X1 port map( B1 => n9466, B2 => n7262, C1 => n9463, C2 => 
                           n7230, A => n7937, ZN => n7932);
   U6768 : OAI22_X1 port map( A1 => n7198, A2 => n9460, B1 => n7166, B2 => 
                           n9457, ZN => n7937);
   U6769 : AOI221_X1 port map( B1 => n9466, B2 => n7261, C1 => n9463, C2 => 
                           n7229, A => n7918, ZN => n7913);
   U6770 : OAI22_X1 port map( A1 => n7197, A2 => n9460, B1 => n7165, B2 => 
                           n9457, ZN => n7918);
   U6771 : AOI221_X1 port map( B1 => n9466, B2 => n7260, C1 => n9463, C2 => 
                           n7228, A => n7899, ZN => n7894);
   U6772 : OAI22_X1 port map( A1 => n7196, A2 => n9460, B1 => n7164, B2 => 
                           n9457, ZN => n7899);
   U6773 : AOI221_X1 port map( B1 => n9467, B2 => n7259, C1 => n9464, C2 => 
                           n7227, A => n7880, ZN => n7875);
   U6774 : OAI22_X1 port map( A1 => n7195, A2 => n9461, B1 => n7163, B2 => 
                           n9458, ZN => n7880);
   U6775 : AOI221_X1 port map( B1 => n9467, B2 => n7258, C1 => n9464, C2 => 
                           n7226, A => n7861, ZN => n7856);
   U6776 : OAI22_X1 port map( A1 => n7194, A2 => n9461, B1 => n7162, B2 => 
                           n9458, ZN => n7861);
   U6777 : AOI221_X1 port map( B1 => n9467, B2 => n7257, C1 => n9464, C2 => 
                           n7225, A => n7842, ZN => n7837);
   U6778 : OAI22_X1 port map( A1 => n7193, A2 => n9461, B1 => n7161, B2 => 
                           n9458, ZN => n7842);
   U6779 : AOI221_X1 port map( B1 => n9467, B2 => n7256, C1 => n9464, C2 => 
                           n7224, A => n7823, ZN => n7818);
   U6780 : OAI22_X1 port map( A1 => n7192, A2 => n9461, B1 => n7160, B2 => 
                           n9458, ZN => n7823);
   U6781 : AOI221_X1 port map( B1 => n9467, B2 => n7255, C1 => n9464, C2 => 
                           n7223, A => n7804, ZN => n7799);
   U6782 : OAI22_X1 port map( A1 => n7191, A2 => n9461, B1 => n7159, B2 => 
                           n9458, ZN => n7804);
   U6783 : AOI221_X1 port map( B1 => n9467, B2 => n7254, C1 => n9464, C2 => 
                           n7222, A => n7785, ZN => n7780);
   U6784 : OAI22_X1 port map( A1 => n7190, A2 => n9461, B1 => n7158, B2 => 
                           n9458, ZN => n7785);
   U6785 : AOI221_X1 port map( B1 => n9467, B2 => n7253, C1 => n9464, C2 => 
                           n7221, A => n7766, ZN => n7761);
   U6786 : OAI22_X1 port map( A1 => n7189, A2 => n9461, B1 => n7157, B2 => 
                           n9458, ZN => n7766);
   U6787 : AOI221_X1 port map( B1 => n9467, B2 => n7252, C1 => n9464, C2 => 
                           n7220, A => n7747, ZN => n7742);
   U6788 : OAI22_X1 port map( A1 => n7188, A2 => n9461, B1 => n7156, B2 => 
                           n9458, ZN => n7747);
   U6789 : AOI221_X1 port map( B1 => n9467, B2 => n7251, C1 => n9464, C2 => 
                           n7219, A => n7728, ZN => n7723);
   U6790 : OAI22_X1 port map( A1 => n7187, A2 => n9461, B1 => n7155, B2 => 
                           n9458, ZN => n7728);
   U6791 : AOI221_X1 port map( B1 => n9467, B2 => n7250, C1 => n9464, C2 => 
                           n7218, A => n7709, ZN => n7704);
   U6792 : OAI22_X1 port map( A1 => n7186, A2 => n9461, B1 => n7154, B2 => 
                           n9458, ZN => n7709);
   U6793 : AOI221_X1 port map( B1 => n9467, B2 => n7249, C1 => n9464, C2 => 
                           n7217, A => n7690, ZN => n7685);
   U6794 : OAI22_X1 port map( A1 => n7185, A2 => n9461, B1 => n7153, B2 => 
                           n9458, ZN => n7690);
   U6795 : AOI221_X1 port map( B1 => n9467, B2 => n7248, C1 => n9464, C2 => 
                           n7216, A => n7671, ZN => n7666);
   U6796 : OAI22_X1 port map( A1 => n7184, A2 => n9461, B1 => n7152, B2 => 
                           n9458, ZN => n7671);
   U6797 : AOI221_X1 port map( B1 => n9468, B2 => n7247, C1 => n9465, C2 => 
                           n7215, A => n7652, ZN => n7647);
   U6798 : OAI22_X1 port map( A1 => n7183, A2 => n9462, B1 => n7151, B2 => 
                           n9459, ZN => n7652);
   U6799 : AOI221_X1 port map( B1 => n9468, B2 => n7246, C1 => n9465, C2 => 
                           n7214, A => n7633, ZN => n7628);
   U6800 : OAI22_X1 port map( A1 => n7182, A2 => n9462, B1 => n7150, B2 => 
                           n9459, ZN => n7633);
   U6801 : AOI221_X1 port map( B1 => n9468, B2 => n7245, C1 => n9465, C2 => 
                           n7213, A => n7614, ZN => n7609);
   U6802 : OAI22_X1 port map( A1 => n7181, A2 => n9462, B1 => n7149, B2 => 
                           n9459, ZN => n7614);
   U6803 : AOI221_X1 port map( B1 => n9468, B2 => n7244, C1 => n9465, C2 => 
                           n7212, A => n7595, ZN => n7590);
   U6804 : OAI22_X1 port map( A1 => n7180, A2 => n9462, B1 => n7148, B2 => 
                           n9459, ZN => n7595);
   U6805 : AOI221_X1 port map( B1 => n9468, B2 => n7243, C1 => n9465, C2 => 
                           n7211, A => n7576, ZN => n7571);
   U6806 : OAI22_X1 port map( A1 => n7179, A2 => n9462, B1 => n7147, B2 => 
                           n9459, ZN => n7576);
   U6807 : AOI221_X1 port map( B1 => n9468, B2 => n7242, C1 => n9465, C2 => 
                           n7210, A => n7557, ZN => n7552);
   U6808 : OAI22_X1 port map( A1 => n7178, A2 => n9462, B1 => n7146, B2 => 
                           n9459, ZN => n7557);
   U6809 : AOI221_X1 port map( B1 => n9468, B2 => n7241, C1 => n9465, C2 => 
                           n7209, A => n7538, ZN => n7533);
   U6810 : OAI22_X1 port map( A1 => n7177, A2 => n9462, B1 => n7145, B2 => 
                           n9459, ZN => n7538);
   U6811 : AOI221_X1 port map( B1 => n9468, B2 => n7240, C1 => n9465, C2 => 
                           n7208, A => n7497, ZN => n7482);
   U6812 : OAI22_X1 port map( A1 => n7176, A2 => n9462, B1 => n7144, B2 => 
                           n9459, ZN => n7497);
   U6813 : AOI221_X1 port map( B1 => n9352, B2 => n7399, C1 => n9349, C2 => 
                           n7367, A => n8770, ZN => n8755);
   U6814 : OAI22_X1 port map( A1 => n7335, A2 => n9346, B1 => n7303, B2 => 
                           n9343, ZN => n8770);
   U6815 : AOI221_X1 port map( B1 => n9304, B2 => n6823, C1 => n9301, C2 => 
                           n6791, A => n8782, ZN => n8771);
   U6816 : OAI22_X1 port map( A1 => n6887, A2 => n9298, B1 => n6855, B2 => 
                           n9295, ZN => n8782);
   U6817 : AOI221_X1 port map( B1 => n9352, B2 => n7398, C1 => n9349, C2 => 
                           n7366, A => n8743, ZN => n8736);
   U6818 : OAI22_X1 port map( A1 => n7334, A2 => n9346, B1 => n7302, B2 => 
                           n9343, ZN => n8743);
   U6819 : AOI221_X1 port map( B1 => n9304, B2 => n6822, C1 => n9301, C2 => 
                           n6790, A => n8751, ZN => n8744);
   U6820 : OAI22_X1 port map( A1 => n6886, A2 => n9298, B1 => n6854, B2 => 
                           n9295, ZN => n8751);
   U6821 : AOI221_X1 port map( B1 => n9352, B2 => n7397, C1 => n9349, C2 => 
                           n7365, A => n8724, ZN => n8717);
   U6822 : OAI22_X1 port map( A1 => n7333, A2 => n9346, B1 => n7301, B2 => 
                           n9343, ZN => n8724);
   U6823 : AOI221_X1 port map( B1 => n9304, B2 => n6821, C1 => n9301, C2 => 
                           n6789, A => n8732, ZN => n8725);
   U6824 : OAI22_X1 port map( A1 => n6885, A2 => n9298, B1 => n6853, B2 => 
                           n9295, ZN => n8732);
   U6825 : AOI221_X1 port map( B1 => n9352, B2 => n7396, C1 => n9349, C2 => 
                           n7364, A => n8705, ZN => n8698);
   U6826 : OAI22_X1 port map( A1 => n7332, A2 => n9346, B1 => n7300, B2 => 
                           n9343, ZN => n8705);
   U6827 : AOI221_X1 port map( B1 => n9304, B2 => n6820, C1 => n9301, C2 => 
                           n6788, A => n8713, ZN => n8706);
   U6828 : OAI22_X1 port map( A1 => n6884, A2 => n9298, B1 => n6852, B2 => 
                           n9295, ZN => n8713);
   U6829 : AOI221_X1 port map( B1 => n9352, B2 => n7395, C1 => n9349, C2 => 
                           n7363, A => n8686, ZN => n8679);
   U6830 : OAI22_X1 port map( A1 => n7331, A2 => n9346, B1 => n7299, B2 => 
                           n9343, ZN => n8686);
   U6831 : AOI221_X1 port map( B1 => n9304, B2 => n6819, C1 => n9301, C2 => 
                           n6787, A => n8694, ZN => n8687);
   U6832 : OAI22_X1 port map( A1 => n6883, A2 => n9298, B1 => n6851, B2 => 
                           n9295, ZN => n8694);
   U6833 : AOI221_X1 port map( B1 => n9352, B2 => n7394, C1 => n9349, C2 => 
                           n7362, A => n8667, ZN => n8660);
   U6834 : OAI22_X1 port map( A1 => n7330, A2 => n9346, B1 => n7298, B2 => 
                           n9343, ZN => n8667);
   U6835 : AOI221_X1 port map( B1 => n9304, B2 => n6818, C1 => n9301, C2 => 
                           n6786, A => n8675, ZN => n8668);
   U6836 : OAI22_X1 port map( A1 => n6882, A2 => n9298, B1 => n6850, B2 => 
                           n9295, ZN => n8675);
   U6837 : AOI221_X1 port map( B1 => n9352, B2 => n7393, C1 => n9349, C2 => 
                           n7361, A => n8648, ZN => n8641);
   U6838 : OAI22_X1 port map( A1 => n7329, A2 => n9346, B1 => n7297, B2 => 
                           n9343, ZN => n8648);
   U6839 : AOI221_X1 port map( B1 => n9304, B2 => n6817, C1 => n9301, C2 => 
                           n6785, A => n8656, ZN => n8649);
   U6840 : OAI22_X1 port map( A1 => n6881, A2 => n9298, B1 => n6849, B2 => 
                           n9295, ZN => n8656);
   U6841 : AOI221_X1 port map( B1 => n9352, B2 => n7392, C1 => n9349, C2 => 
                           n7360, A => n8629, ZN => n8622);
   U6842 : OAI22_X1 port map( A1 => n7328, A2 => n9346, B1 => n7296, B2 => 
                           n9343, ZN => n8629);
   U6843 : AOI221_X1 port map( B1 => n9304, B2 => n6816, C1 => n9301, C2 => 
                           n6784, A => n8637, ZN => n8630);
   U6844 : OAI22_X1 port map( A1 => n6880, A2 => n9298, B1 => n6848, B2 => 
                           n9295, ZN => n8637);
   U6845 : AOI221_X1 port map( B1 => n9352, B2 => n7391, C1 => n9349, C2 => 
                           n7359, A => n8610, ZN => n8603);
   U6846 : OAI22_X1 port map( A1 => n7327, A2 => n9346, B1 => n7295, B2 => 
                           n9343, ZN => n8610);
   U6847 : AOI221_X1 port map( B1 => n9304, B2 => n6815, C1 => n9301, C2 => 
                           n6783, A => n8618, ZN => n8611);
   U6848 : OAI22_X1 port map( A1 => n6879, A2 => n9298, B1 => n6847, B2 => 
                           n9295, ZN => n8618);
   U6849 : AOI221_X1 port map( B1 => n9352, B2 => n7390, C1 => n9349, C2 => 
                           n7358, A => n8591, ZN => n8584);
   U6850 : OAI22_X1 port map( A1 => n7326, A2 => n9346, B1 => n7294, B2 => 
                           n9343, ZN => n8591);
   U6851 : AOI221_X1 port map( B1 => n9304, B2 => n6814, C1 => n9301, C2 => 
                           n6782, A => n8599, ZN => n8592);
   U6852 : OAI22_X1 port map( A1 => n6878, A2 => n9298, B1 => n6846, B2 => 
                           n9295, ZN => n8599);
   U6853 : AOI221_X1 port map( B1 => n9352, B2 => n7389, C1 => n9349, C2 => 
                           n7357, A => n8572, ZN => n8565);
   U6854 : OAI22_X1 port map( A1 => n7325, A2 => n9346, B1 => n7293, B2 => 
                           n9343, ZN => n8572);
   U6855 : AOI221_X1 port map( B1 => n9304, B2 => n6813, C1 => n9301, C2 => 
                           n6781, A => n8580, ZN => n8573);
   U6856 : OAI22_X1 port map( A1 => n6877, A2 => n9298, B1 => n6845, B2 => 
                           n9295, ZN => n8580);
   U6857 : AOI221_X1 port map( B1 => n9352, B2 => n7388, C1 => n9349, C2 => 
                           n7356, A => n8553, ZN => n8546);
   U6858 : OAI22_X1 port map( A1 => n7324, A2 => n9346, B1 => n7292, B2 => 
                           n9343, ZN => n8553);
   U6859 : AOI221_X1 port map( B1 => n9304, B2 => n6812, C1 => n9301, C2 => 
                           n6780, A => n8561, ZN => n8554);
   U6860 : OAI22_X1 port map( A1 => n6876, A2 => n9298, B1 => n6844, B2 => 
                           n9295, ZN => n8561);
   U6861 : AOI221_X1 port map( B1 => n9353, B2 => n7387, C1 => n9350, C2 => 
                           n7355, A => n8534, ZN => n8527);
   U6862 : OAI22_X1 port map( A1 => n7323, A2 => n9347, B1 => n7291, B2 => 
                           n9344, ZN => n8534);
   U6863 : AOI221_X1 port map( B1 => n9305, B2 => n6811, C1 => n9302, C2 => 
                           n6779, A => n8542, ZN => n8535);
   U6864 : OAI22_X1 port map( A1 => n6875, A2 => n9299, B1 => n6843, B2 => 
                           n9296, ZN => n8542);
   U6865 : AOI221_X1 port map( B1 => n9353, B2 => n7386, C1 => n9350, C2 => 
                           n7354, A => n8515, ZN => n8508);
   U6866 : OAI22_X1 port map( A1 => n7322, A2 => n9347, B1 => n7290, B2 => 
                           n9344, ZN => n8515);
   U6867 : AOI221_X1 port map( B1 => n9305, B2 => n6810, C1 => n9302, C2 => 
                           n6778, A => n8523, ZN => n8516);
   U6868 : OAI22_X1 port map( A1 => n6874, A2 => n9299, B1 => n6842, B2 => 
                           n9296, ZN => n8523);
   U6869 : AOI221_X1 port map( B1 => n9353, B2 => n7385, C1 => n9350, C2 => 
                           n7353, A => n8496, ZN => n8489);
   U6870 : OAI22_X1 port map( A1 => n7321, A2 => n9347, B1 => n7289, B2 => 
                           n9344, ZN => n8496);
   U6871 : AOI221_X1 port map( B1 => n9305, B2 => n6809, C1 => n9302, C2 => 
                           n6777, A => n8504, ZN => n8497);
   U6872 : OAI22_X1 port map( A1 => n6873, A2 => n9299, B1 => n6841, B2 => 
                           n9296, ZN => n8504);
   U6873 : AOI221_X1 port map( B1 => n9353, B2 => n7384, C1 => n9350, C2 => 
                           n7352, A => n8477, ZN => n8470);
   U6874 : OAI22_X1 port map( A1 => n7320, A2 => n9347, B1 => n7288, B2 => 
                           n9344, ZN => n8477);
   U6875 : AOI221_X1 port map( B1 => n9305, B2 => n6808, C1 => n9302, C2 => 
                           n6776, A => n8485, ZN => n8478);
   U6876 : OAI22_X1 port map( A1 => n6872, A2 => n9299, B1 => n6840, B2 => 
                           n9296, ZN => n8485);
   U6877 : AOI221_X1 port map( B1 => n9353, B2 => n7383, C1 => n9350, C2 => 
                           n7351, A => n8458, ZN => n8451);
   U6878 : OAI22_X1 port map( A1 => n7319, A2 => n9347, B1 => n7287, B2 => 
                           n9344, ZN => n8458);
   U6879 : AOI221_X1 port map( B1 => n9305, B2 => n6807, C1 => n9302, C2 => 
                           n6775, A => n8466, ZN => n8459);
   U6880 : OAI22_X1 port map( A1 => n6871, A2 => n9299, B1 => n6839, B2 => 
                           n9296, ZN => n8466);
   U6881 : AOI221_X1 port map( B1 => n9353, B2 => n7382, C1 => n9350, C2 => 
                           n7350, A => n8439, ZN => n8432);
   U6882 : OAI22_X1 port map( A1 => n7318, A2 => n9347, B1 => n7286, B2 => 
                           n9344, ZN => n8439);
   U6883 : AOI221_X1 port map( B1 => n9305, B2 => n6806, C1 => n9302, C2 => 
                           n6774, A => n8447, ZN => n8440);
   U6884 : OAI22_X1 port map( A1 => n6870, A2 => n9299, B1 => n6838, B2 => 
                           n9296, ZN => n8447);
   U6885 : AOI221_X1 port map( B1 => n9353, B2 => n7381, C1 => n9350, C2 => 
                           n7349, A => n8420, ZN => n8413);
   U6886 : OAI22_X1 port map( A1 => n7317, A2 => n9347, B1 => n7285, B2 => 
                           n9344, ZN => n8420);
   U6887 : AOI221_X1 port map( B1 => n9305, B2 => n6805, C1 => n9302, C2 => 
                           n6773, A => n8428, ZN => n8421);
   U6888 : OAI22_X1 port map( A1 => n6869, A2 => n9299, B1 => n6837, B2 => 
                           n9296, ZN => n8428);
   U6889 : AOI221_X1 port map( B1 => n9353, B2 => n7380, C1 => n9350, C2 => 
                           n7348, A => n8401, ZN => n8394);
   U6890 : OAI22_X1 port map( A1 => n7316, A2 => n9347, B1 => n7284, B2 => 
                           n9344, ZN => n8401);
   U6891 : AOI221_X1 port map( B1 => n9305, B2 => n6804, C1 => n9302, C2 => 
                           n6772, A => n8409, ZN => n8402);
   U6892 : OAI22_X1 port map( A1 => n6868, A2 => n9299, B1 => n6836, B2 => 
                           n9296, ZN => n8409);
   U6893 : AOI221_X1 port map( B1 => n9353, B2 => n7379, C1 => n9350, C2 => 
                           n7347, A => n8382, ZN => n8375);
   U6894 : OAI22_X1 port map( A1 => n7315, A2 => n9347, B1 => n7283, B2 => 
                           n9344, ZN => n8382);
   U6895 : AOI221_X1 port map( B1 => n9305, B2 => n6803, C1 => n9302, C2 => 
                           n6771, A => n8390, ZN => n8383);
   U6896 : OAI22_X1 port map( A1 => n6867, A2 => n9299, B1 => n6835, B2 => 
                           n9296, ZN => n8390);
   U6897 : AOI221_X1 port map( B1 => n9353, B2 => n7378, C1 => n9350, C2 => 
                           n7346, A => n8363, ZN => n8356);
   U6898 : OAI22_X1 port map( A1 => n7314, A2 => n9347, B1 => n7282, B2 => 
                           n9344, ZN => n8363);
   U6899 : AOI221_X1 port map( B1 => n9305, B2 => n6802, C1 => n9302, C2 => 
                           n6770, A => n8371, ZN => n8364);
   U6900 : OAI22_X1 port map( A1 => n6866, A2 => n9299, B1 => n6834, B2 => 
                           n9296, ZN => n8371);
   U6901 : AOI221_X1 port map( B1 => n9353, B2 => n7377, C1 => n9350, C2 => 
                           n7345, A => n8344, ZN => n8337);
   U6902 : OAI22_X1 port map( A1 => n7313, A2 => n9347, B1 => n7281, B2 => 
                           n9344, ZN => n8344);
   U6903 : AOI221_X1 port map( B1 => n9305, B2 => n6801, C1 => n9302, C2 => 
                           n6769, A => n8352, ZN => n8345);
   U6904 : OAI22_X1 port map( A1 => n6865, A2 => n9299, B1 => n6833, B2 => 
                           n9296, ZN => n8352);
   U6905 : AOI221_X1 port map( B1 => n9353, B2 => n7376, C1 => n9350, C2 => 
                           n7344, A => n8325, ZN => n8318);
   U6906 : OAI22_X1 port map( A1 => n7312, A2 => n9347, B1 => n7280, B2 => 
                           n9344, ZN => n8325);
   U6907 : AOI221_X1 port map( B1 => n9305, B2 => n6800, C1 => n9302, C2 => 
                           n6768, A => n8333, ZN => n8326);
   U6908 : OAI22_X1 port map( A1 => n6864, A2 => n9299, B1 => n6832, B2 => 
                           n9296, ZN => n8333);
   U6909 : AOI221_X1 port map( B1 => n9354, B2 => n7375, C1 => n9351, C2 => 
                           n7343, A => n8306, ZN => n8299);
   U6910 : OAI22_X1 port map( A1 => n7311, A2 => n9348, B1 => n7279, B2 => 
                           n9345, ZN => n8306);
   U6911 : AOI221_X1 port map( B1 => n9306, B2 => n6799, C1 => n9303, C2 => 
                           n6767, A => n8314, ZN => n8307);
   U6912 : OAI22_X1 port map( A1 => n6863, A2 => n9300, B1 => n6831, B2 => 
                           n9297, ZN => n8314);
   U6913 : AOI221_X1 port map( B1 => n9354, B2 => n7374, C1 => n9351, C2 => 
                           n7342, A => n8287, ZN => n8280);
   U6914 : OAI22_X1 port map( A1 => n7310, A2 => n9348, B1 => n7278, B2 => 
                           n9345, ZN => n8287);
   U6915 : AOI221_X1 port map( B1 => n9306, B2 => n6798, C1 => n9303, C2 => 
                           n6766, A => n8295, ZN => n8288);
   U6916 : OAI22_X1 port map( A1 => n6862, A2 => n9300, B1 => n6830, B2 => 
                           n9297, ZN => n8295);
   U6917 : AOI221_X1 port map( B1 => n9354, B2 => n7373, C1 => n9351, C2 => 
                           n7341, A => n8268, ZN => n8261);
   U6918 : OAI22_X1 port map( A1 => n7309, A2 => n9348, B1 => n7277, B2 => 
                           n9345, ZN => n8268);
   U6919 : AOI221_X1 port map( B1 => n9306, B2 => n6797, C1 => n9303, C2 => 
                           n6765, A => n8276, ZN => n8269);
   U6920 : OAI22_X1 port map( A1 => n6861, A2 => n9300, B1 => n6829, B2 => 
                           n9297, ZN => n8276);
   U6921 : AOI221_X1 port map( B1 => n9354, B2 => n7372, C1 => n9351, C2 => 
                           n7340, A => n8249, ZN => n8242);
   U6922 : OAI22_X1 port map( A1 => n7308, A2 => n9348, B1 => n7276, B2 => 
                           n9345, ZN => n8249);
   U6923 : AOI221_X1 port map( B1 => n9306, B2 => n6796, C1 => n9303, C2 => 
                           n6764, A => n8257, ZN => n8250);
   U6924 : OAI22_X1 port map( A1 => n6860, A2 => n9300, B1 => n6828, B2 => 
                           n9297, ZN => n8257);
   U6925 : AOI221_X1 port map( B1 => n9354, B2 => n7371, C1 => n9351, C2 => 
                           n7339, A => n8230, ZN => n8223);
   U6926 : OAI22_X1 port map( A1 => n7307, A2 => n9348, B1 => n7275, B2 => 
                           n9345, ZN => n8230);
   U6927 : AOI221_X1 port map( B1 => n9306, B2 => n6795, C1 => n9303, C2 => 
                           n6763, A => n8238, ZN => n8231);
   U6928 : OAI22_X1 port map( A1 => n6859, A2 => n9300, B1 => n6827, B2 => 
                           n9297, ZN => n8238);
   U6929 : AOI221_X1 port map( B1 => n9354, B2 => n7370, C1 => n9351, C2 => 
                           n7338, A => n8211, ZN => n8204);
   U6930 : OAI22_X1 port map( A1 => n7306, A2 => n9348, B1 => n7274, B2 => 
                           n9345, ZN => n8211);
   U6931 : AOI221_X1 port map( B1 => n9306, B2 => n6794, C1 => n9303, C2 => 
                           n6762, A => n8219, ZN => n8212);
   U6932 : OAI22_X1 port map( A1 => n6858, A2 => n9300, B1 => n6826, B2 => 
                           n9297, ZN => n8219);
   U6933 : AOI221_X1 port map( B1 => n9354, B2 => n7369, C1 => n9351, C2 => 
                           n7337, A => n8192, ZN => n8185);
   U6934 : OAI22_X1 port map( A1 => n7305, A2 => n9348, B1 => n7273, B2 => 
                           n9345, ZN => n8192);
   U6935 : AOI221_X1 port map( B1 => n9306, B2 => n6793, C1 => n9303, C2 => 
                           n6761, A => n8200, ZN => n8193);
   U6936 : OAI22_X1 port map( A1 => n6857, A2 => n9300, B1 => n6825, B2 => 
                           n9297, ZN => n8200);
   U6937 : AOI221_X1 port map( B1 => n9354, B2 => n7368, C1 => n9351, C2 => 
                           n7336, A => n8155, ZN => n8134);
   U6938 : OAI22_X1 port map( A1 => n7304, A2 => n9348, B1 => n7272, B2 => 
                           n9345, ZN => n8155);
   U6939 : AOI221_X1 port map( B1 => n9306, B2 => n6792, C1 => n9303, C2 => 
                           n6760, A => n8179, ZN => n8158);
   U6940 : OAI22_X1 port map( A1 => n6856, A2 => n9300, B1 => n6824, B2 => 
                           n9297, ZN => n8179);
   U6941 : AOI221_X1 port map( B1 => n9454, B2 => n7399, C1 => n9451, C2 => 
                           n7367, A => n8117, ZN => n8102);
   U6942 : OAI22_X1 port map( A1 => n7335, A2 => n9448, B1 => n7303, B2 => 
                           n9445, ZN => n8117);
   U6943 : AOI221_X1 port map( B1 => n9406, B2 => n6823, C1 => n9403, C2 => 
                           n6791, A => n8129, ZN => n8118);
   U6944 : OAI22_X1 port map( A1 => n6887, A2 => n9400, B1 => n6855, B2 => 
                           n9397, ZN => n8129);
   U6945 : AOI221_X1 port map( B1 => n9454, B2 => n7398, C1 => n9451, C2 => 
                           n7366, A => n8090, ZN => n8083);
   U6946 : OAI22_X1 port map( A1 => n7334, A2 => n9448, B1 => n7302, B2 => 
                           n9445, ZN => n8090);
   U6947 : AOI221_X1 port map( B1 => n9406, B2 => n6822, C1 => n9403, C2 => 
                           n6790, A => n8098, ZN => n8091);
   U6948 : OAI22_X1 port map( A1 => n6886, A2 => n9400, B1 => n6854, B2 => 
                           n9397, ZN => n8098);
   U6949 : AOI221_X1 port map( B1 => n9454, B2 => n7397, C1 => n9451, C2 => 
                           n7365, A => n8071, ZN => n8064);
   U6950 : OAI22_X1 port map( A1 => n7333, A2 => n9448, B1 => n7301, B2 => 
                           n9445, ZN => n8071);
   U6951 : AOI221_X1 port map( B1 => n9406, B2 => n6821, C1 => n9403, C2 => 
                           n6789, A => n8079, ZN => n8072);
   U6952 : OAI22_X1 port map( A1 => n6885, A2 => n9400, B1 => n6853, B2 => 
                           n9397, ZN => n8079);
   U6953 : AOI221_X1 port map( B1 => n9454, B2 => n7396, C1 => n9451, C2 => 
                           n7364, A => n8052, ZN => n8045);
   U6954 : OAI22_X1 port map( A1 => n7332, A2 => n9448, B1 => n7300, B2 => 
                           n9445, ZN => n8052);
   U6955 : AOI221_X1 port map( B1 => n9406, B2 => n6820, C1 => n9403, C2 => 
                           n6788, A => n8060, ZN => n8053);
   U6956 : OAI22_X1 port map( A1 => n6884, A2 => n9400, B1 => n6852, B2 => 
                           n9397, ZN => n8060);
   U6957 : AOI221_X1 port map( B1 => n9454, B2 => n7395, C1 => n9451, C2 => 
                           n7363, A => n8033, ZN => n8026);
   U6958 : OAI22_X1 port map( A1 => n7331, A2 => n9448, B1 => n7299, B2 => 
                           n9445, ZN => n8033);
   U6959 : AOI221_X1 port map( B1 => n9406, B2 => n6819, C1 => n9403, C2 => 
                           n6787, A => n8041, ZN => n8034);
   U6960 : OAI22_X1 port map( A1 => n6883, A2 => n9400, B1 => n6851, B2 => 
                           n9397, ZN => n8041);
   U6961 : AOI221_X1 port map( B1 => n9454, B2 => n7394, C1 => n9451, C2 => 
                           n7362, A => n8014, ZN => n8007);
   U6962 : OAI22_X1 port map( A1 => n7330, A2 => n9448, B1 => n7298, B2 => 
                           n9445, ZN => n8014);
   U6963 : AOI221_X1 port map( B1 => n9406, B2 => n6818, C1 => n9403, C2 => 
                           n6786, A => n8022, ZN => n8015);
   U6964 : OAI22_X1 port map( A1 => n6882, A2 => n9400, B1 => n6850, B2 => 
                           n9397, ZN => n8022);
   U6965 : AOI221_X1 port map( B1 => n9454, B2 => n7393, C1 => n9451, C2 => 
                           n7361, A => n7995, ZN => n7988);
   U6966 : OAI22_X1 port map( A1 => n7329, A2 => n9448, B1 => n7297, B2 => 
                           n9445, ZN => n7995);
   U6967 : AOI221_X1 port map( B1 => n9406, B2 => n6817, C1 => n9403, C2 => 
                           n6785, A => n8003, ZN => n7996);
   U6968 : OAI22_X1 port map( A1 => n6881, A2 => n9400, B1 => n6849, B2 => 
                           n9397, ZN => n8003);
   U6969 : AOI221_X1 port map( B1 => n9454, B2 => n7392, C1 => n9451, C2 => 
                           n7360, A => n7976, ZN => n7969);
   U6970 : OAI22_X1 port map( A1 => n7328, A2 => n9448, B1 => n7296, B2 => 
                           n9445, ZN => n7976);
   U6971 : AOI221_X1 port map( B1 => n9406, B2 => n6816, C1 => n9403, C2 => 
                           n6784, A => n7984, ZN => n7977);
   U6972 : OAI22_X1 port map( A1 => n6880, A2 => n9400, B1 => n6848, B2 => 
                           n9397, ZN => n7984);
   U6973 : AOI221_X1 port map( B1 => n9454, B2 => n7391, C1 => n9451, C2 => 
                           n7359, A => n7957, ZN => n7950);
   U6974 : OAI22_X1 port map( A1 => n7327, A2 => n9448, B1 => n7295, B2 => 
                           n9445, ZN => n7957);
   U6975 : AOI221_X1 port map( B1 => n9406, B2 => n6815, C1 => n9403, C2 => 
                           n6783, A => n7965, ZN => n7958);
   U6976 : OAI22_X1 port map( A1 => n6879, A2 => n9400, B1 => n6847, B2 => 
                           n9397, ZN => n7965);
   U6977 : AOI221_X1 port map( B1 => n9454, B2 => n7390, C1 => n9451, C2 => 
                           n7358, A => n7938, ZN => n7931);
   U6978 : OAI22_X1 port map( A1 => n7326, A2 => n9448, B1 => n7294, B2 => 
                           n9445, ZN => n7938);
   U6979 : AOI221_X1 port map( B1 => n9406, B2 => n6814, C1 => n9403, C2 => 
                           n6782, A => n7946, ZN => n7939);
   U6980 : OAI22_X1 port map( A1 => n6878, A2 => n9400, B1 => n6846, B2 => 
                           n9397, ZN => n7946);
   U6981 : AOI221_X1 port map( B1 => n9454, B2 => n7389, C1 => n9451, C2 => 
                           n7357, A => n7919, ZN => n7912);
   U6982 : OAI22_X1 port map( A1 => n7325, A2 => n9448, B1 => n7293, B2 => 
                           n9445, ZN => n7919);
   U6983 : AOI221_X1 port map( B1 => n9406, B2 => n6813, C1 => n9403, C2 => 
                           n6781, A => n7927, ZN => n7920);
   U6984 : OAI22_X1 port map( A1 => n6877, A2 => n9400, B1 => n6845, B2 => 
                           n9397, ZN => n7927);
   U6985 : AOI221_X1 port map( B1 => n9454, B2 => n7388, C1 => n9451, C2 => 
                           n7356, A => n7900, ZN => n7893);
   U6986 : OAI22_X1 port map( A1 => n7324, A2 => n9448, B1 => n7292, B2 => 
                           n9445, ZN => n7900);
   U6987 : AOI221_X1 port map( B1 => n9406, B2 => n6812, C1 => n9403, C2 => 
                           n6780, A => n7908, ZN => n7901);
   U6988 : OAI22_X1 port map( A1 => n6876, A2 => n9400, B1 => n6844, B2 => 
                           n9397, ZN => n7908);
   U6989 : AOI221_X1 port map( B1 => n9455, B2 => n7387, C1 => n9452, C2 => 
                           n7355, A => n7881, ZN => n7874);
   U6990 : OAI22_X1 port map( A1 => n7323, A2 => n9449, B1 => n7291, B2 => 
                           n9446, ZN => n7881);
   U6991 : AOI221_X1 port map( B1 => n9407, B2 => n6811, C1 => n9404, C2 => 
                           n6779, A => n7889, ZN => n7882);
   U6992 : OAI22_X1 port map( A1 => n6875, A2 => n9401, B1 => n6843, B2 => 
                           n9398, ZN => n7889);
   U6993 : AOI221_X1 port map( B1 => n9455, B2 => n7386, C1 => n9452, C2 => 
                           n7354, A => n7862, ZN => n7855);
   U6994 : OAI22_X1 port map( A1 => n7322, A2 => n9449, B1 => n7290, B2 => 
                           n9446, ZN => n7862);
   U6995 : AOI221_X1 port map( B1 => n9407, B2 => n6810, C1 => n9404, C2 => 
                           n6778, A => n7870, ZN => n7863);
   U6996 : OAI22_X1 port map( A1 => n6874, A2 => n9401, B1 => n6842, B2 => 
                           n9398, ZN => n7870);
   U6997 : AOI221_X1 port map( B1 => n9455, B2 => n7385, C1 => n9452, C2 => 
                           n7353, A => n7843, ZN => n7836);
   U6998 : OAI22_X1 port map( A1 => n7321, A2 => n9449, B1 => n7289, B2 => 
                           n9446, ZN => n7843);
   U6999 : AOI221_X1 port map( B1 => n9407, B2 => n6809, C1 => n9404, C2 => 
                           n6777, A => n7851, ZN => n7844);
   U7000 : OAI22_X1 port map( A1 => n6873, A2 => n9401, B1 => n6841, B2 => 
                           n9398, ZN => n7851);
   U7001 : AOI221_X1 port map( B1 => n9455, B2 => n7384, C1 => n9452, C2 => 
                           n7352, A => n7824, ZN => n7817);
   U7002 : OAI22_X1 port map( A1 => n7320, A2 => n9449, B1 => n7288, B2 => 
                           n9446, ZN => n7824);
   U7003 : AOI221_X1 port map( B1 => n9407, B2 => n6808, C1 => n9404, C2 => 
                           n6776, A => n7832, ZN => n7825);
   U7004 : OAI22_X1 port map( A1 => n6872, A2 => n9401, B1 => n6840, B2 => 
                           n9398, ZN => n7832);
   U7005 : AOI221_X1 port map( B1 => n9455, B2 => n7383, C1 => n9452, C2 => 
                           n7351, A => n7805, ZN => n7798);
   U7006 : OAI22_X1 port map( A1 => n7319, A2 => n9449, B1 => n7287, B2 => 
                           n9446, ZN => n7805);
   U7007 : AOI221_X1 port map( B1 => n9407, B2 => n6807, C1 => n9404, C2 => 
                           n6775, A => n7813, ZN => n7806);
   U7008 : OAI22_X1 port map( A1 => n6871, A2 => n9401, B1 => n6839, B2 => 
                           n9398, ZN => n7813);
   U7009 : AOI221_X1 port map( B1 => n9455, B2 => n7382, C1 => n9452, C2 => 
                           n7350, A => n7786, ZN => n7779);
   U7010 : OAI22_X1 port map( A1 => n7318, A2 => n9449, B1 => n7286, B2 => 
                           n9446, ZN => n7786);
   U7011 : AOI221_X1 port map( B1 => n9407, B2 => n6806, C1 => n9404, C2 => 
                           n6774, A => n7794, ZN => n7787);
   U7012 : OAI22_X1 port map( A1 => n6870, A2 => n9401, B1 => n6838, B2 => 
                           n9398, ZN => n7794);
   U7013 : AOI221_X1 port map( B1 => n9455, B2 => n7381, C1 => n9452, C2 => 
                           n7349, A => n7767, ZN => n7760);
   U7014 : OAI22_X1 port map( A1 => n7317, A2 => n9449, B1 => n7285, B2 => 
                           n9446, ZN => n7767);
   U7015 : AOI221_X1 port map( B1 => n9407, B2 => n6805, C1 => n9404, C2 => 
                           n6773, A => n7775, ZN => n7768);
   U7016 : OAI22_X1 port map( A1 => n6869, A2 => n9401, B1 => n6837, B2 => 
                           n9398, ZN => n7775);
   U7017 : AOI221_X1 port map( B1 => n9455, B2 => n7380, C1 => n9452, C2 => 
                           n7348, A => n7748, ZN => n7741);
   U7018 : OAI22_X1 port map( A1 => n7316, A2 => n9449, B1 => n7284, B2 => 
                           n9446, ZN => n7748);
   U7019 : AOI221_X1 port map( B1 => n9407, B2 => n6804, C1 => n9404, C2 => 
                           n6772, A => n7756, ZN => n7749);
   U7020 : OAI22_X1 port map( A1 => n6868, A2 => n9401, B1 => n6836, B2 => 
                           n9398, ZN => n7756);
   U7021 : AOI221_X1 port map( B1 => n9455, B2 => n7379, C1 => n9452, C2 => 
                           n7347, A => n7729, ZN => n7722);
   U7022 : OAI22_X1 port map( A1 => n7315, A2 => n9449, B1 => n7283, B2 => 
                           n9446, ZN => n7729);
   U7023 : AOI221_X1 port map( B1 => n9407, B2 => n6803, C1 => n9404, C2 => 
                           n6771, A => n7737, ZN => n7730);
   U7024 : OAI22_X1 port map( A1 => n6867, A2 => n9401, B1 => n6835, B2 => 
                           n9398, ZN => n7737);
   U7025 : AOI221_X1 port map( B1 => n9455, B2 => n7378, C1 => n9452, C2 => 
                           n7346, A => n7710, ZN => n7703);
   U7026 : OAI22_X1 port map( A1 => n7314, A2 => n9449, B1 => n7282, B2 => 
                           n9446, ZN => n7710);
   U7027 : AOI221_X1 port map( B1 => n9407, B2 => n6802, C1 => n9404, C2 => 
                           n6770, A => n7718, ZN => n7711);
   U7028 : OAI22_X1 port map( A1 => n6866, A2 => n9401, B1 => n6834, B2 => 
                           n9398, ZN => n7718);
   U7029 : AOI221_X1 port map( B1 => n9455, B2 => n7377, C1 => n9452, C2 => 
                           n7345, A => n7691, ZN => n7684);
   U7030 : OAI22_X1 port map( A1 => n7313, A2 => n9449, B1 => n7281, B2 => 
                           n9446, ZN => n7691);
   U7031 : AOI221_X1 port map( B1 => n9407, B2 => n6801, C1 => n9404, C2 => 
                           n6769, A => n7699, ZN => n7692);
   U7032 : OAI22_X1 port map( A1 => n6865, A2 => n9401, B1 => n6833, B2 => 
                           n9398, ZN => n7699);
   U7033 : AOI221_X1 port map( B1 => n9455, B2 => n7376, C1 => n9452, C2 => 
                           n7344, A => n7672, ZN => n7665);
   U7034 : OAI22_X1 port map( A1 => n7312, A2 => n9449, B1 => n7280, B2 => 
                           n9446, ZN => n7672);
   U7035 : AOI221_X1 port map( B1 => n9407, B2 => n6800, C1 => n9404, C2 => 
                           n6768, A => n7680, ZN => n7673);
   U7036 : OAI22_X1 port map( A1 => n6864, A2 => n9401, B1 => n6832, B2 => 
                           n9398, ZN => n7680);
   U7037 : AOI221_X1 port map( B1 => n9456, B2 => n7375, C1 => n9453, C2 => 
                           n7343, A => n7653, ZN => n7646);
   U7038 : OAI22_X1 port map( A1 => n7311, A2 => n9450, B1 => n7279, B2 => 
                           n9447, ZN => n7653);
   U7039 : AOI221_X1 port map( B1 => n9408, B2 => n6799, C1 => n9405, C2 => 
                           n6767, A => n7661, ZN => n7654);
   U7040 : OAI22_X1 port map( A1 => n6863, A2 => n9402, B1 => n6831, B2 => 
                           n9399, ZN => n7661);
   U7041 : AOI221_X1 port map( B1 => n9456, B2 => n7374, C1 => n9453, C2 => 
                           n7342, A => n7634, ZN => n7627);
   U7042 : OAI22_X1 port map( A1 => n7310, A2 => n9450, B1 => n7278, B2 => 
                           n9447, ZN => n7634);
   U7043 : AOI221_X1 port map( B1 => n9408, B2 => n6798, C1 => n9405, C2 => 
                           n6766, A => n7642, ZN => n7635);
   U7044 : OAI22_X1 port map( A1 => n6862, A2 => n9402, B1 => n6830, B2 => 
                           n9399, ZN => n7642);
   U7045 : AOI221_X1 port map( B1 => n9456, B2 => n7373, C1 => n9453, C2 => 
                           n7341, A => n7615, ZN => n7608);
   U7046 : OAI22_X1 port map( A1 => n7309, A2 => n9450, B1 => n7277, B2 => 
                           n9447, ZN => n7615);
   U7047 : AOI221_X1 port map( B1 => n9408, B2 => n6797, C1 => n9405, C2 => 
                           n6765, A => n7623, ZN => n7616);
   U7048 : OAI22_X1 port map( A1 => n6861, A2 => n9402, B1 => n6829, B2 => 
                           n9399, ZN => n7623);
   U7049 : AOI221_X1 port map( B1 => n9456, B2 => n7372, C1 => n9453, C2 => 
                           n7340, A => n7596, ZN => n7589);
   U7050 : OAI22_X1 port map( A1 => n7308, A2 => n9450, B1 => n7276, B2 => 
                           n9447, ZN => n7596);
   U7051 : AOI221_X1 port map( B1 => n9408, B2 => n6796, C1 => n9405, C2 => 
                           n6764, A => n7604, ZN => n7597);
   U7052 : OAI22_X1 port map( A1 => n6860, A2 => n9402, B1 => n6828, B2 => 
                           n9399, ZN => n7604);
   U7053 : AOI221_X1 port map( B1 => n9456, B2 => n7371, C1 => n9453, C2 => 
                           n7339, A => n7577, ZN => n7570);
   U7054 : OAI22_X1 port map( A1 => n7307, A2 => n9450, B1 => n7275, B2 => 
                           n9447, ZN => n7577);
   U7055 : AOI221_X1 port map( B1 => n9408, B2 => n6795, C1 => n9405, C2 => 
                           n6763, A => n7585, ZN => n7578);
   U7056 : OAI22_X1 port map( A1 => n6859, A2 => n9402, B1 => n6827, B2 => 
                           n9399, ZN => n7585);
   U7057 : AOI221_X1 port map( B1 => n9456, B2 => n7370, C1 => n9453, C2 => 
                           n7338, A => n7558, ZN => n7551);
   U7058 : OAI22_X1 port map( A1 => n7306, A2 => n9450, B1 => n7274, B2 => 
                           n9447, ZN => n7558);
   U7059 : AOI221_X1 port map( B1 => n9408, B2 => n6794, C1 => n9405, C2 => 
                           n6762, A => n7566, ZN => n7559);
   U7060 : OAI22_X1 port map( A1 => n6858, A2 => n9402, B1 => n6826, B2 => 
                           n9399, ZN => n7566);
   U7061 : AOI221_X1 port map( B1 => n9456, B2 => n7369, C1 => n9453, C2 => 
                           n7337, A => n7539, ZN => n7532);
   U7062 : OAI22_X1 port map( A1 => n7305, A2 => n9450, B1 => n7273, B2 => 
                           n9447, ZN => n7539);
   U7063 : AOI221_X1 port map( B1 => n9408, B2 => n6793, C1 => n9405, C2 => 
                           n6761, A => n7547, ZN => n7540);
   U7064 : OAI22_X1 port map( A1 => n6857, A2 => n9402, B1 => n6825, B2 => 
                           n9399, ZN => n7547);
   U7065 : AOI221_X1 port map( B1 => n9456, B2 => n7368, C1 => n9453, C2 => 
                           n7336, A => n7502, ZN => n7481);
   U7066 : OAI22_X1 port map( A1 => n7304, A2 => n9450, B1 => n7272, B2 => 
                           n9447, ZN => n7502);
   U7067 : AOI221_X1 port map( B1 => n9408, B2 => n6792, C1 => n9405, C2 => 
                           n6760, A => n7526, ZN => n7505);
   U7068 : OAI22_X1 port map( A1 => n6856, A2 => n9402, B1 => n6824, B2 => 
                           n9399, ZN => n7526);
   U7069 : AOI221_X1 port map( B1 => n9378, B2 => n7055, C1 => n9375, C2 => 
                           n7023, A => n8304, ZN => n8301);
   U7070 : OAI22_X1 port map( A1 => n7119, A2 => n9372, B1 => n7087, B2 => 
                           n9369, ZN => n8304);
   U7071 : AOI221_X1 port map( B1 => n9378, B2 => n7054, C1 => n9375, C2 => 
                           n7022, A => n8285, ZN => n8282);
   U7072 : OAI22_X1 port map( A1 => n7118, A2 => n9372, B1 => n7086, B2 => 
                           n9369, ZN => n8285);
   U7073 : AOI221_X1 port map( B1 => n9378, B2 => n7053, C1 => n9375, C2 => 
                           n7021, A => n8266, ZN => n8263);
   U7074 : OAI22_X1 port map( A1 => n7117, A2 => n9372, B1 => n7085, B2 => 
                           n9369, ZN => n8266);
   U7075 : AOI221_X1 port map( B1 => n9378, B2 => n7052, C1 => n9375, C2 => 
                           n7020, A => n8247, ZN => n8244);
   U7076 : OAI22_X1 port map( A1 => n7116, A2 => n9372, B1 => n7084, B2 => 
                           n9369, ZN => n8247);
   U7077 : AOI221_X1 port map( B1 => n9378, B2 => n7051, C1 => n9375, C2 => 
                           n7019, A => n8228, ZN => n8225);
   U7078 : OAI22_X1 port map( A1 => n7115, A2 => n9372, B1 => n7083, B2 => 
                           n9369, ZN => n8228);
   U7079 : AOI221_X1 port map( B1 => n9378, B2 => n7050, C1 => n9375, C2 => 
                           n7018, A => n8209, ZN => n8206);
   U7080 : OAI22_X1 port map( A1 => n7114, A2 => n9372, B1 => n7082, B2 => 
                           n9369, ZN => n8209);
   U7081 : AOI221_X1 port map( B1 => n9378, B2 => n7049, C1 => n9375, C2 => 
                           n7017, A => n8190, ZN => n8187);
   U7082 : OAI22_X1 port map( A1 => n7113, A2 => n9372, B1 => n7081, B2 => 
                           n9369, ZN => n8190);
   U7083 : AOI221_X1 port map( B1 => n9378, B2 => n7048, C1 => n9375, C2 => 
                           n7016, A => n8145, ZN => n8136);
   U7084 : OAI22_X1 port map( A1 => n7112, A2 => n9372, B1 => n7080, B2 => 
                           n9369, ZN => n8145);
   U7085 : AOI221_X1 port map( B1 => n9480, B2 => n7055, C1 => n9477, C2 => 
                           n7023, A => n7651, ZN => n7648);
   U7086 : OAI22_X1 port map( A1 => n7119, A2 => n9474, B1 => n7087, B2 => 
                           n9471, ZN => n7651);
   U7087 : AOI221_X1 port map( B1 => n9480, B2 => n7054, C1 => n9477, C2 => 
                           n7022, A => n7632, ZN => n7629);
   U7088 : OAI22_X1 port map( A1 => n7118, A2 => n9474, B1 => n7086, B2 => 
                           n9471, ZN => n7632);
   U7089 : AOI221_X1 port map( B1 => n9480, B2 => n7053, C1 => n9477, C2 => 
                           n7021, A => n7613, ZN => n7610);
   U7090 : OAI22_X1 port map( A1 => n7117, A2 => n9474, B1 => n7085, B2 => 
                           n9471, ZN => n7613);
   U7091 : AOI221_X1 port map( B1 => n9480, B2 => n7052, C1 => n9477, C2 => 
                           n7020, A => n7594, ZN => n7591);
   U7092 : OAI22_X1 port map( A1 => n7116, A2 => n9474, B1 => n7084, B2 => 
                           n9471, ZN => n7594);
   U7093 : AOI221_X1 port map( B1 => n9480, B2 => n7051, C1 => n9477, C2 => 
                           n7019, A => n7575, ZN => n7572);
   U7094 : OAI22_X1 port map( A1 => n7115, A2 => n9474, B1 => n7083, B2 => 
                           n9471, ZN => n7575);
   U7095 : AOI221_X1 port map( B1 => n9480, B2 => n7050, C1 => n9477, C2 => 
                           n7018, A => n7556, ZN => n7553);
   U7096 : OAI22_X1 port map( A1 => n7114, A2 => n9474, B1 => n7082, B2 => 
                           n9471, ZN => n7556);
   U7097 : AOI221_X1 port map( B1 => n9480, B2 => n7049, C1 => n9477, C2 => 
                           n7017, A => n7537, ZN => n7534);
   U7098 : OAI22_X1 port map( A1 => n7113, A2 => n9474, B1 => n7081, B2 => 
                           n9471, ZN => n7537);
   U7099 : AOI221_X1 port map( B1 => n9480, B2 => n7048, C1 => n9477, C2 => 
                           n7016, A => n7492, ZN => n7483);
   U7100 : OAI22_X1 port map( A1 => n7112, A2 => n9474, B1 => n7080, B2 => 
                           n9471, ZN => n7492);
   U7101 : OAI22_X1 port map( A1 => n9524, A2 => n9854, B1 => n7474, B2 => 
                           n7311, ZN => n2678);
   U7102 : OAI22_X1 port map( A1 => n9525, A2 => n9857, B1 => n7474, B2 => 
                           n7310, ZN => n2679);
   U7103 : OAI22_X1 port map( A1 => n9525, A2 => n9860, B1 => n7474, B2 => 
                           n7309, ZN => n2680);
   U7104 : OAI22_X1 port map( A1 => n9525, A2 => n9863, B1 => n7474, B2 => 
                           n7308, ZN => n2681);
   U7105 : OAI22_X1 port map( A1 => n9525, A2 => n9866, B1 => n7474, B2 => 
                           n7307, ZN => n2682);
   U7106 : OAI22_X1 port map( A1 => n9525, A2 => n9869, B1 => n7474, B2 => 
                           n7306, ZN => n2683);
   U7107 : OAI22_X1 port map( A1 => n9526, A2 => n9872, B1 => n7474, B2 => 
                           n7305, ZN => n2684);
   U7108 : OAI22_X1 port map( A1 => n9526, A2 => n9884, B1 => n7474, B2 => 
                           n7304, ZN => n2685);
   U7109 : OAI22_X1 port map( A1 => n9533, A2 => n9854, B1 => n7473, B2 => 
                           n7279, ZN => n2710);
   U7110 : OAI22_X1 port map( A1 => n9534, A2 => n9857, B1 => n7473, B2 => 
                           n7278, ZN => n2711);
   U7111 : OAI22_X1 port map( A1 => n9534, A2 => n9860, B1 => n7473, B2 => 
                           n7277, ZN => n2712);
   U7112 : OAI22_X1 port map( A1 => n9534, A2 => n9863, B1 => n7473, B2 => 
                           n7276, ZN => n2713);
   U7113 : OAI22_X1 port map( A1 => n9534, A2 => n9866, B1 => n7473, B2 => 
                           n7275, ZN => n2714);
   U7114 : OAI22_X1 port map( A1 => n9534, A2 => n9869, B1 => n7473, B2 => 
                           n7274, ZN => n2715);
   U7115 : OAI22_X1 port map( A1 => n9535, A2 => n9872, B1 => n7473, B2 => 
                           n7273, ZN => n2716);
   U7116 : OAI22_X1 port map( A1 => n9535, A2 => n9884, B1 => n7473, B2 => 
                           n7272, ZN => n2717);
   U7117 : OAI22_X1 port map( A1 => n9560, A2 => n9854, B1 => n7470, B2 => 
                           n7183, ZN => n2806);
   U7118 : OAI22_X1 port map( A1 => n9561, A2 => n9857, B1 => n7470, B2 => 
                           n7182, ZN => n2807);
   U7119 : OAI22_X1 port map( A1 => n9561, A2 => n9860, B1 => n7470, B2 => 
                           n7181, ZN => n2808);
   U7120 : OAI22_X1 port map( A1 => n9561, A2 => n9863, B1 => n7470, B2 => 
                           n7180, ZN => n2809);
   U7121 : OAI22_X1 port map( A1 => n9561, A2 => n9866, B1 => n7470, B2 => 
                           n7179, ZN => n2810);
   U7122 : OAI22_X1 port map( A1 => n9561, A2 => n9869, B1 => n7470, B2 => 
                           n7178, ZN => n2811);
   U7123 : OAI22_X1 port map( A1 => n9562, A2 => n9872, B1 => n7470, B2 => 
                           n7177, ZN => n2812);
   U7124 : OAI22_X1 port map( A1 => n9562, A2 => n9884, B1 => n7470, B2 => 
                           n7176, ZN => n2813);
   U7125 : OAI22_X1 port map( A1 => n9569, A2 => n9854, B1 => n7468, B2 => 
                           n7151, ZN => n2838);
   U7126 : OAI22_X1 port map( A1 => n9570, A2 => n9857, B1 => n7468, B2 => 
                           n7150, ZN => n2839);
   U7127 : OAI22_X1 port map( A1 => n9570, A2 => n9860, B1 => n7468, B2 => 
                           n7149, ZN => n2840);
   U7128 : OAI22_X1 port map( A1 => n9570, A2 => n9863, B1 => n7468, B2 => 
                           n7148, ZN => n2841);
   U7129 : OAI22_X1 port map( A1 => n9570, A2 => n9866, B1 => n7468, B2 => 
                           n7147, ZN => n2842);
   U7130 : OAI22_X1 port map( A1 => n9570, A2 => n9869, B1 => n7468, B2 => 
                           n7146, ZN => n2843);
   U7131 : OAI22_X1 port map( A1 => n9571, A2 => n9872, B1 => n7468, B2 => 
                           n7145, ZN => n2844);
   U7132 : OAI22_X1 port map( A1 => n9571, A2 => n9884, B1 => n7468, B2 => 
                           n7144, ZN => n2845);
   U7133 : OAI22_X1 port map( A1 => n9578, A2 => n9853, B1 => n7467, B2 => 
                           n7119, ZN => n2870);
   U7134 : OAI22_X1 port map( A1 => n9579, A2 => n9856, B1 => n7467, B2 => 
                           n7118, ZN => n2871);
   U7135 : OAI22_X1 port map( A1 => n9579, A2 => n9859, B1 => n7467, B2 => 
                           n7117, ZN => n2872);
   U7136 : OAI22_X1 port map( A1 => n9579, A2 => n9862, B1 => n7467, B2 => 
                           n7116, ZN => n2873);
   U7137 : OAI22_X1 port map( A1 => n9579, A2 => n9865, B1 => n7467, B2 => 
                           n7115, ZN => n2874);
   U7138 : OAI22_X1 port map( A1 => n9579, A2 => n9868, B1 => n7467, B2 => 
                           n7114, ZN => n2875);
   U7139 : OAI22_X1 port map( A1 => n9580, A2 => n9871, B1 => n7467, B2 => 
                           n7113, ZN => n2876);
   U7140 : OAI22_X1 port map( A1 => n9580, A2 => n9883, B1 => n7467, B2 => 
                           n7112, ZN => n2877);
   U7141 : OAI22_X1 port map( A1 => n9587, A2 => n9853, B1 => n7466, B2 => 
                           n7087, ZN => n2902);
   U7142 : OAI22_X1 port map( A1 => n9588, A2 => n9856, B1 => n7466, B2 => 
                           n7086, ZN => n2903);
   U7143 : OAI22_X1 port map( A1 => n9588, A2 => n9859, B1 => n7466, B2 => 
                           n7085, ZN => n2904);
   U7144 : OAI22_X1 port map( A1 => n9588, A2 => n9862, B1 => n7466, B2 => 
                           n7084, ZN => n2905);
   U7145 : OAI22_X1 port map( A1 => n9588, A2 => n9865, B1 => n7466, B2 => 
                           n7083, ZN => n2906);
   U7146 : OAI22_X1 port map( A1 => n9588, A2 => n9868, B1 => n7466, B2 => 
                           n7082, ZN => n2907);
   U7147 : OAI22_X1 port map( A1 => n9589, A2 => n9871, B1 => n7466, B2 => 
                           n7081, ZN => n2908);
   U7148 : OAI22_X1 port map( A1 => n9589, A2 => n9883, B1 => n7466, B2 => 
                           n7080, ZN => n2909);
   U7149 : OAI22_X1 port map( A1 => n9614, A2 => n9853, B1 => n7463, B2 => 
                           n6991, ZN => n2998);
   U7150 : OAI22_X1 port map( A1 => n9615, A2 => n9856, B1 => n7463, B2 => 
                           n6990, ZN => n2999);
   U7151 : OAI22_X1 port map( A1 => n9615, A2 => n9859, B1 => n7463, B2 => 
                           n6989, ZN => n3000);
   U7152 : OAI22_X1 port map( A1 => n9615, A2 => n9862, B1 => n7463, B2 => 
                           n6988, ZN => n3001);
   U7153 : OAI22_X1 port map( A1 => n9615, A2 => n9865, B1 => n7463, B2 => 
                           n6987, ZN => n3002);
   U7154 : OAI22_X1 port map( A1 => n9615, A2 => n9868, B1 => n7463, B2 => 
                           n6986, ZN => n3003);
   U7155 : OAI22_X1 port map( A1 => n9616, A2 => n9871, B1 => n7463, B2 => 
                           n6985, ZN => n3004);
   U7156 : OAI22_X1 port map( A1 => n9616, A2 => n9883, B1 => n7463, B2 => 
                           n6984, ZN => n3005);
   U7157 : OAI22_X1 port map( A1 => n9623, A2 => n9853, B1 => n7462, B2 => 
                           n6959, ZN => n3030);
   U7158 : OAI22_X1 port map( A1 => n9624, A2 => n9856, B1 => n7462, B2 => 
                           n6958, ZN => n3031);
   U7159 : OAI22_X1 port map( A1 => n9624, A2 => n9859, B1 => n7462, B2 => 
                           n6957, ZN => n3032);
   U7160 : OAI22_X1 port map( A1 => n9624, A2 => n9862, B1 => n7462, B2 => 
                           n6956, ZN => n3033);
   U7161 : OAI22_X1 port map( A1 => n9624, A2 => n9865, B1 => n7462, B2 => 
                           n6955, ZN => n3034);
   U7162 : OAI22_X1 port map( A1 => n9624, A2 => n9868, B1 => n7462, B2 => 
                           n6954, ZN => n3035);
   U7163 : OAI22_X1 port map( A1 => n9625, A2 => n9871, B1 => n7462, B2 => 
                           n6953, ZN => n3036);
   U7164 : OAI22_X1 port map( A1 => n9625, A2 => n9883, B1 => n7462, B2 => 
                           n6952, ZN => n3037);
   U7165 : OAI22_X1 port map( A1 => n9650, A2 => n9853, B1 => n7458, B2 => 
                           n6863, ZN => n3126);
   U7166 : OAI22_X1 port map( A1 => n9651, A2 => n9856, B1 => n7458, B2 => 
                           n6862, ZN => n3127);
   U7167 : OAI22_X1 port map( A1 => n9651, A2 => n9859, B1 => n7458, B2 => 
                           n6861, ZN => n3128);
   U7168 : OAI22_X1 port map( A1 => n9651, A2 => n9862, B1 => n7458, B2 => 
                           n6860, ZN => n3129);
   U7169 : OAI22_X1 port map( A1 => n9651, A2 => n9865, B1 => n7458, B2 => 
                           n6859, ZN => n3130);
   U7170 : OAI22_X1 port map( A1 => n9651, A2 => n9868, B1 => n7458, B2 => 
                           n6858, ZN => n3131);
   U7171 : OAI22_X1 port map( A1 => n9652, A2 => n9871, B1 => n7458, B2 => 
                           n6857, ZN => n3132);
   U7172 : OAI22_X1 port map( A1 => n9652, A2 => n9883, B1 => n7458, B2 => 
                           n6856, ZN => n3133);
   U7173 : OAI22_X1 port map( A1 => n9659, A2 => n9853, B1 => n7457, B2 => 
                           n6831, ZN => n3158);
   U7174 : OAI22_X1 port map( A1 => n9660, A2 => n9856, B1 => n7457, B2 => 
                           n6830, ZN => n3159);
   U7175 : OAI22_X1 port map( A1 => n9660, A2 => n9859, B1 => n7457, B2 => 
                           n6829, ZN => n3160);
   U7176 : OAI22_X1 port map( A1 => n9660, A2 => n9862, B1 => n7457, B2 => 
                           n6828, ZN => n3161);
   U7177 : OAI22_X1 port map( A1 => n9660, A2 => n9865, B1 => n7457, B2 => 
                           n6827, ZN => n3162);
   U7178 : OAI22_X1 port map( A1 => n9660, A2 => n9868, B1 => n7457, B2 => 
                           n6826, ZN => n3163);
   U7179 : OAI22_X1 port map( A1 => n9661, A2 => n9871, B1 => n7457, B2 => 
                           n6825, ZN => n3164);
   U7180 : OAI22_X1 port map( A1 => n9661, A2 => n9883, B1 => n7457, B2 => 
                           n6824, ZN => n3165);
   U7181 : OAI22_X1 port map( A1 => n9686, A2 => n9852, B1 => n7454, B2 => 
                           n6735, ZN => n3254);
   U7182 : OAI22_X1 port map( A1 => n9687, A2 => n9855, B1 => n7454, B2 => 
                           n6734, ZN => n3255);
   U7183 : OAI22_X1 port map( A1 => n9687, A2 => n9858, B1 => n7454, B2 => 
                           n6733, ZN => n3256);
   U7184 : OAI22_X1 port map( A1 => n9687, A2 => n9861, B1 => n7454, B2 => 
                           n6732, ZN => n3257);
   U7185 : OAI22_X1 port map( A1 => n9687, A2 => n9864, B1 => n7454, B2 => 
                           n6731, ZN => n3258);
   U7186 : OAI22_X1 port map( A1 => n9687, A2 => n9867, B1 => n7454, B2 => 
                           n6730, ZN => n3259);
   U7187 : OAI22_X1 port map( A1 => n9688, A2 => n9870, B1 => n7454, B2 => 
                           n6729, ZN => n3260);
   U7188 : OAI22_X1 port map( A1 => n9688, A2 => n9882, B1 => n7454, B2 => 
                           n6728, ZN => n3261);
   U7189 : OAI22_X1 port map( A1 => n9695, A2 => n9852, B1 => n7453, B2 => 
                           n6703, ZN => n3286);
   U7190 : OAI22_X1 port map( A1 => n9696, A2 => n9855, B1 => n7453, B2 => 
                           n6702, ZN => n3287);
   U7191 : OAI22_X1 port map( A1 => n9696, A2 => n9858, B1 => n7453, B2 => 
                           n6701, ZN => n3288);
   U7192 : OAI22_X1 port map( A1 => n9696, A2 => n9861, B1 => n7453, B2 => 
                           n6700, ZN => n3289);
   U7193 : OAI22_X1 port map( A1 => n9696, A2 => n9864, B1 => n7453, B2 => 
                           n6699, ZN => n3290);
   U7194 : OAI22_X1 port map( A1 => n9696, A2 => n9867, B1 => n7453, B2 => 
                           n6698, ZN => n3291);
   U7195 : OAI22_X1 port map( A1 => n9697, A2 => n9870, B1 => n7453, B2 => 
                           n6697, ZN => n3292);
   U7196 : OAI22_X1 port map( A1 => n9697, A2 => n9882, B1 => n7453, B2 => 
                           n6696, ZN => n3293);
   U7197 : OAI22_X1 port map( A1 => n9704, A2 => n9852, B1 => n7452, B2 => 
                           n6671, ZN => n3318);
   U7198 : OAI22_X1 port map( A1 => n9705, A2 => n9855, B1 => n7452, B2 => 
                           n6670, ZN => n3319);
   U7199 : OAI22_X1 port map( A1 => n9705, A2 => n9858, B1 => n7452, B2 => 
                           n6669, ZN => n3320);
   U7200 : OAI22_X1 port map( A1 => n9705, A2 => n9861, B1 => n7452, B2 => 
                           n6668, ZN => n3321);
   U7201 : OAI22_X1 port map( A1 => n9705, A2 => n9864, B1 => n7452, B2 => 
                           n6667, ZN => n3322);
   U7202 : OAI22_X1 port map( A1 => n9705, A2 => n9867, B1 => n7452, B2 => 
                           n6666, ZN => n3323);
   U7203 : OAI22_X1 port map( A1 => n9706, A2 => n9870, B1 => n7452, B2 => 
                           n6665, ZN => n3324);
   U7204 : OAI22_X1 port map( A1 => n9706, A2 => n9882, B1 => n7452, B2 => 
                           n6664, ZN => n3325);
   U7205 : OAI22_X1 port map( A1 => n9713, A2 => n9852, B1 => n7450, B2 => 
                           n6639, ZN => n3350);
   U7206 : OAI22_X1 port map( A1 => n9714, A2 => n9855, B1 => n7450, B2 => 
                           n6638, ZN => n3351);
   U7207 : OAI22_X1 port map( A1 => n9714, A2 => n9858, B1 => n7450, B2 => 
                           n6637, ZN => n3352);
   U7208 : OAI22_X1 port map( A1 => n9714, A2 => n9861, B1 => n7450, B2 => 
                           n6636, ZN => n3353);
   U7209 : OAI22_X1 port map( A1 => n9714, A2 => n9864, B1 => n7450, B2 => 
                           n6635, ZN => n3354);
   U7210 : OAI22_X1 port map( A1 => n9714, A2 => n9867, B1 => n7450, B2 => 
                           n6634, ZN => n3355);
   U7211 : OAI22_X1 port map( A1 => n9715, A2 => n9870, B1 => n7450, B2 => 
                           n6633, ZN => n3356);
   U7212 : OAI22_X1 port map( A1 => n9715, A2 => n9882, B1 => n7450, B2 => 
                           n6632, ZN => n3357);
   U7213 : OAI22_X1 port map( A1 => n9776, A2 => n9852, B1 => n7435, B2 => 
                           n6499, ZN => n3574);
   U7214 : OAI22_X1 port map( A1 => n9777, A2 => n9855, B1 => n7435, B2 => 
                           n6498, ZN => n3575);
   U7215 : OAI22_X1 port map( A1 => n9777, A2 => n9858, B1 => n7435, B2 => 
                           n6497, ZN => n3576);
   U7216 : OAI22_X1 port map( A1 => n9777, A2 => n9861, B1 => n7435, B2 => 
                           n6496, ZN => n3577);
   U7217 : OAI22_X1 port map( A1 => n9777, A2 => n9864, B1 => n7435, B2 => 
                           n6495, ZN => n3578);
   U7218 : OAI22_X1 port map( A1 => n9777, A2 => n9867, B1 => n7435, B2 => 
                           n6494, ZN => n3579);
   U7219 : OAI22_X1 port map( A1 => n9778, A2 => n9870, B1 => n7435, B2 => 
                           n6493, ZN => n3580);
   U7220 : OAI22_X1 port map( A1 => n9778, A2 => n9882, B1 => n7435, B2 => 
                           n6492, ZN => n3581);
   U7221 : OAI22_X1 port map( A1 => n9874, A2 => n9783, B1 => n7401, B2 => 
                           n6490, ZN => n3583);
   U7222 : OAI22_X1 port map( A1 => n9874, A2 => n9786, B1 => n7401, B2 => 
                           n6489, ZN => n3584);
   U7223 : OAI22_X1 port map( A1 => n9874, A2 => n9789, B1 => n7401, B2 => 
                           n6488, ZN => n3585);
   U7224 : OAI22_X1 port map( A1 => n9874, A2 => n9792, B1 => n7401, B2 => 
                           n6487, ZN => n3586);
   U7225 : OAI22_X1 port map( A1 => n9875, A2 => n9795, B1 => n7401, B2 => 
                           n6486, ZN => n3587);
   U7226 : OAI22_X1 port map( A1 => n9875, A2 => n9798, B1 => n7401, B2 => 
                           n6485, ZN => n3588);
   U7227 : OAI22_X1 port map( A1 => n9875, A2 => n9801, B1 => n7401, B2 => 
                           n6484, ZN => n3589);
   U7228 : OAI22_X1 port map( A1 => n9874, A2 => n9782, B1 => n9873, B2 => 
                           n6491, ZN => n3582);
   U7229 : OAI22_X1 port map( A1 => n9875, A2 => n9804, B1 => n9873, B2 => 
                           n6483, ZN => n3590);
   U7230 : OAI22_X1 port map( A1 => n9875, A2 => n9807, B1 => n9873, B2 => 
                           n6482, ZN => n3591);
   U7231 : OAI22_X1 port map( A1 => n9876, A2 => n9810, B1 => n9873, B2 => 
                           n6481, ZN => n3592);
   U7232 : OAI22_X1 port map( A1 => n9876, A2 => n9813, B1 => n9873, B2 => 
                           n6480, ZN => n3593);
   U7233 : OAI22_X1 port map( A1 => n9876, A2 => n9816, B1 => n9873, B2 => 
                           n6479, ZN => n3594);
   U7234 : OAI22_X1 port map( A1 => n9876, A2 => n9819, B1 => n9873, B2 => 
                           n6478, ZN => n3595);
   U7235 : OAI22_X1 port map( A1 => n9876, A2 => n9822, B1 => n9873, B2 => 
                           n6477, ZN => n3596);
   U7236 : OAI22_X1 port map( A1 => n9877, A2 => n9825, B1 => n9873, B2 => 
                           n6476, ZN => n3597);
   U7237 : OAI22_X1 port map( A1 => n9877, A2 => n9828, B1 => n9873, B2 => 
                           n6475, ZN => n3598);
   U7238 : OAI22_X1 port map( A1 => n9877, A2 => n9831, B1 => n9873, B2 => 
                           n6474, ZN => n3599);
   U7239 : OAI22_X1 port map( A1 => n9877, A2 => n9834, B1 => n9873, B2 => 
                           n6473, ZN => n3600);
   U7240 : OAI22_X1 port map( A1 => n9877, A2 => n9837, B1 => n9873, B2 => 
                           n6472, ZN => n3601);
   U7241 : OAI22_X1 port map( A1 => n9776, A2 => n9840, B1 => n9771, B2 => 
                           n6503, ZN => n3570);
   U7242 : OAI22_X1 port map( A1 => n9776, A2 => n9843, B1 => n9771, B2 => 
                           n6502, ZN => n3571);
   U7243 : OAI22_X1 port map( A1 => n9776, A2 => n9846, B1 => n9771, B2 => 
                           n6501, ZN => n3572);
   U7244 : OAI22_X1 port map( A1 => n9776, A2 => n9849, B1 => n9771, B2 => 
                           n6500, ZN => n3573);
   U7245 : OAI22_X1 port map( A1 => n9878, A2 => n9840, B1 => n7401, B2 => 
                           n6471, ZN => n3602);
   U7246 : OAI22_X1 port map( A1 => n9878, A2 => n9843, B1 => n7401, B2 => 
                           n6470, ZN => n3603);
   U7247 : OAI22_X1 port map( A1 => n9878, A2 => n9846, B1 => n7401, B2 => 
                           n6469, ZN => n3604);
   U7248 : OAI22_X1 port map( A1 => n9879, A2 => n9864, B1 => n7401, B2 => 
                           n6468, ZN => n3610);
   U7249 : OAI22_X1 port map( A1 => n9879, A2 => n9867, B1 => n9873, B2 => 
                           n6467, ZN => n3611);
   U7250 : OAI22_X1 port map( A1 => n9880, A2 => n9870, B1 => n9873, B2 => 
                           n6466, ZN => n3612);
   U7251 : OAI22_X1 port map( A1 => n9880, A2 => n9882, B1 => n9873, B2 => 
                           n6465, ZN => n3613);
   U7252 : OAI22_X1 port map( A1 => n9520, A2 => n9780, B1 => n9519, B2 => 
                           n7335, ZN => n2654);
   U7253 : OAI22_X1 port map( A1 => n9520, A2 => n9785, B1 => n9519, B2 => 
                           n7334, ZN => n2655);
   U7254 : OAI22_X1 port map( A1 => n9520, A2 => n9788, B1 => n9519, B2 => 
                           n7333, ZN => n2656);
   U7255 : OAI22_X1 port map( A1 => n9520, A2 => n9791, B1 => n9519, B2 => 
                           n7332, ZN => n2657);
   U7256 : OAI22_X1 port map( A1 => n9520, A2 => n9794, B1 => n9519, B2 => 
                           n7331, ZN => n2658);
   U7257 : OAI22_X1 port map( A1 => n9521, A2 => n9797, B1 => n9519, B2 => 
                           n7330, ZN => n2659);
   U7258 : OAI22_X1 port map( A1 => n9521, A2 => n9800, B1 => n9519, B2 => 
                           n7329, ZN => n2660);
   U7259 : OAI22_X1 port map( A1 => n9521, A2 => n9803, B1 => n9519, B2 => 
                           n7328, ZN => n2661);
   U7260 : OAI22_X1 port map( A1 => n9521, A2 => n9806, B1 => n9519, B2 => 
                           n7327, ZN => n2662);
   U7261 : OAI22_X1 port map( A1 => n9521, A2 => n9809, B1 => n9519, B2 => 
                           n7326, ZN => n2663);
   U7262 : OAI22_X1 port map( A1 => n9522, A2 => n9812, B1 => n9519, B2 => 
                           n7325, ZN => n2664);
   U7263 : OAI22_X1 port map( A1 => n9522, A2 => n9815, B1 => n9519, B2 => 
                           n7324, ZN => n2665);
   U7264 : OAI22_X1 port map( A1 => n9522, A2 => n9818, B1 => n7474, B2 => 
                           n7323, ZN => n2666);
   U7265 : OAI22_X1 port map( A1 => n9522, A2 => n9821, B1 => n7474, B2 => 
                           n7322, ZN => n2667);
   U7266 : OAI22_X1 port map( A1 => n9522, A2 => n9824, B1 => n7474, B2 => 
                           n7321, ZN => n2668);
   U7267 : OAI22_X1 port map( A1 => n9523, A2 => n9827, B1 => n9519, B2 => 
                           n7320, ZN => n2669);
   U7268 : OAI22_X1 port map( A1 => n9523, A2 => n9830, B1 => n9519, B2 => 
                           n7319, ZN => n2670);
   U7269 : OAI22_X1 port map( A1 => n9523, A2 => n9833, B1 => n9519, B2 => 
                           n7318, ZN => n2671);
   U7270 : OAI22_X1 port map( A1 => n9523, A2 => n9836, B1 => n9519, B2 => 
                           n7317, ZN => n2672);
   U7271 : OAI22_X1 port map( A1 => n9523, A2 => n9839, B1 => n9519, B2 => 
                           n7316, ZN => n2673);
   U7272 : OAI22_X1 port map( A1 => n9524, A2 => n9842, B1 => n9519, B2 => 
                           n7315, ZN => n2674);
   U7273 : OAI22_X1 port map( A1 => n9524, A2 => n9845, B1 => n9519, B2 => 
                           n7314, ZN => n2675);
   U7274 : OAI22_X1 port map( A1 => n9524, A2 => n9848, B1 => n9519, B2 => 
                           n7313, ZN => n2676);
   U7275 : OAI22_X1 port map( A1 => n9524, A2 => n9851, B1 => n9519, B2 => 
                           n7312, ZN => n2677);
   U7276 : OAI22_X1 port map( A1 => n9529, A2 => n9780, B1 => n9528, B2 => 
                           n7303, ZN => n2686);
   U7277 : OAI22_X1 port map( A1 => n9529, A2 => n9785, B1 => n9528, B2 => 
                           n7302, ZN => n2687);
   U7278 : OAI22_X1 port map( A1 => n9529, A2 => n9788, B1 => n9528, B2 => 
                           n7301, ZN => n2688);
   U7279 : OAI22_X1 port map( A1 => n9529, A2 => n9791, B1 => n9528, B2 => 
                           n7300, ZN => n2689);
   U7280 : OAI22_X1 port map( A1 => n9529, A2 => n9794, B1 => n9528, B2 => 
                           n7299, ZN => n2690);
   U7281 : OAI22_X1 port map( A1 => n9530, A2 => n9797, B1 => n9528, B2 => 
                           n7298, ZN => n2691);
   U7282 : OAI22_X1 port map( A1 => n9530, A2 => n9800, B1 => n9528, B2 => 
                           n7297, ZN => n2692);
   U7283 : OAI22_X1 port map( A1 => n9530, A2 => n9803, B1 => n9528, B2 => 
                           n7296, ZN => n2693);
   U7284 : OAI22_X1 port map( A1 => n9530, A2 => n9806, B1 => n9528, B2 => 
                           n7295, ZN => n2694);
   U7285 : OAI22_X1 port map( A1 => n9530, A2 => n9809, B1 => n9528, B2 => 
                           n7294, ZN => n2695);
   U7286 : OAI22_X1 port map( A1 => n9531, A2 => n9812, B1 => n9528, B2 => 
                           n7293, ZN => n2696);
   U7287 : OAI22_X1 port map( A1 => n9531, A2 => n9815, B1 => n9528, B2 => 
                           n7292, ZN => n2697);
   U7288 : OAI22_X1 port map( A1 => n9531, A2 => n9818, B1 => n7473, B2 => 
                           n7291, ZN => n2698);
   U7289 : OAI22_X1 port map( A1 => n9531, A2 => n9821, B1 => n7473, B2 => 
                           n7290, ZN => n2699);
   U7290 : OAI22_X1 port map( A1 => n9531, A2 => n9824, B1 => n7473, B2 => 
                           n7289, ZN => n2700);
   U7291 : OAI22_X1 port map( A1 => n9532, A2 => n9827, B1 => n9528, B2 => 
                           n7288, ZN => n2701);
   U7292 : OAI22_X1 port map( A1 => n9532, A2 => n9830, B1 => n9528, B2 => 
                           n7287, ZN => n2702);
   U7293 : OAI22_X1 port map( A1 => n9532, A2 => n9833, B1 => n9528, B2 => 
                           n7286, ZN => n2703);
   U7294 : OAI22_X1 port map( A1 => n9532, A2 => n9836, B1 => n9528, B2 => 
                           n7285, ZN => n2704);
   U7295 : OAI22_X1 port map( A1 => n9532, A2 => n9839, B1 => n9528, B2 => 
                           n7284, ZN => n2705);
   U7296 : OAI22_X1 port map( A1 => n9533, A2 => n9842, B1 => n9528, B2 => 
                           n7283, ZN => n2706);
   U7297 : OAI22_X1 port map( A1 => n9533, A2 => n9845, B1 => n9528, B2 => 
                           n7282, ZN => n2707);
   U7298 : OAI22_X1 port map( A1 => n9533, A2 => n9848, B1 => n9528, B2 => 
                           n7281, ZN => n2708);
   U7299 : OAI22_X1 port map( A1 => n9533, A2 => n9851, B1 => n9528, B2 => 
                           n7280, ZN => n2709);
   U7300 : OAI22_X1 port map( A1 => n9556, A2 => n9780, B1 => n9555, B2 => 
                           n7207, ZN => n2782);
   U7301 : OAI22_X1 port map( A1 => n9556, A2 => n9785, B1 => n9555, B2 => 
                           n7206, ZN => n2783);
   U7302 : OAI22_X1 port map( A1 => n9556, A2 => n9788, B1 => n9555, B2 => 
                           n7205, ZN => n2784);
   U7303 : OAI22_X1 port map( A1 => n9556, A2 => n9791, B1 => n9555, B2 => 
                           n7204, ZN => n2785);
   U7304 : OAI22_X1 port map( A1 => n9556, A2 => n9794, B1 => n9555, B2 => 
                           n7203, ZN => n2786);
   U7305 : OAI22_X1 port map( A1 => n9557, A2 => n9797, B1 => n9555, B2 => 
                           n7202, ZN => n2787);
   U7306 : OAI22_X1 port map( A1 => n9557, A2 => n9800, B1 => n9555, B2 => 
                           n7201, ZN => n2788);
   U7307 : OAI22_X1 port map( A1 => n9557, A2 => n9803, B1 => n9555, B2 => 
                           n7200, ZN => n2789);
   U7308 : OAI22_X1 port map( A1 => n9557, A2 => n9806, B1 => n9555, B2 => 
                           n7199, ZN => n2790);
   U7309 : OAI22_X1 port map( A1 => n9557, A2 => n9809, B1 => n9555, B2 => 
                           n7198, ZN => n2791);
   U7310 : OAI22_X1 port map( A1 => n9558, A2 => n9812, B1 => n9555, B2 => 
                           n7197, ZN => n2792);
   U7311 : OAI22_X1 port map( A1 => n9558, A2 => n9815, B1 => n9555, B2 => 
                           n7196, ZN => n2793);
   U7312 : OAI22_X1 port map( A1 => n9558, A2 => n9818, B1 => n7470, B2 => 
                           n7195, ZN => n2794);
   U7313 : OAI22_X1 port map( A1 => n9558, A2 => n9821, B1 => n7470, B2 => 
                           n7194, ZN => n2795);
   U7314 : OAI22_X1 port map( A1 => n9558, A2 => n9824, B1 => n7470, B2 => 
                           n7193, ZN => n2796);
   U7315 : OAI22_X1 port map( A1 => n9559, A2 => n9827, B1 => n9555, B2 => 
                           n7192, ZN => n2797);
   U7316 : OAI22_X1 port map( A1 => n9559, A2 => n9830, B1 => n9555, B2 => 
                           n7191, ZN => n2798);
   U7317 : OAI22_X1 port map( A1 => n9559, A2 => n9833, B1 => n9555, B2 => 
                           n7190, ZN => n2799);
   U7318 : OAI22_X1 port map( A1 => n9559, A2 => n9836, B1 => n9555, B2 => 
                           n7189, ZN => n2800);
   U7319 : OAI22_X1 port map( A1 => n9559, A2 => n9839, B1 => n9555, B2 => 
                           n7188, ZN => n2801);
   U7320 : OAI22_X1 port map( A1 => n9560, A2 => n9842, B1 => n9555, B2 => 
                           n7187, ZN => n2802);
   U7321 : OAI22_X1 port map( A1 => n9560, A2 => n9845, B1 => n9555, B2 => 
                           n7186, ZN => n2803);
   U7322 : OAI22_X1 port map( A1 => n9560, A2 => n9848, B1 => n9555, B2 => 
                           n7185, ZN => n2804);
   U7323 : OAI22_X1 port map( A1 => n9560, A2 => n9851, B1 => n9555, B2 => 
                           n7184, ZN => n2805);
   U7324 : OAI22_X1 port map( A1 => n9565, A2 => n9780, B1 => n9564, B2 => 
                           n7175, ZN => n2814);
   U7325 : OAI22_X1 port map( A1 => n9565, A2 => n9785, B1 => n9564, B2 => 
                           n7174, ZN => n2815);
   U7326 : OAI22_X1 port map( A1 => n9565, A2 => n9788, B1 => n9564, B2 => 
                           n7173, ZN => n2816);
   U7327 : OAI22_X1 port map( A1 => n9565, A2 => n9791, B1 => n9564, B2 => 
                           n7172, ZN => n2817);
   U7328 : OAI22_X1 port map( A1 => n9565, A2 => n9794, B1 => n9564, B2 => 
                           n7171, ZN => n2818);
   U7329 : OAI22_X1 port map( A1 => n9566, A2 => n9797, B1 => n9564, B2 => 
                           n7170, ZN => n2819);
   U7330 : OAI22_X1 port map( A1 => n9566, A2 => n9800, B1 => n9564, B2 => 
                           n7169, ZN => n2820);
   U7331 : OAI22_X1 port map( A1 => n9566, A2 => n9803, B1 => n9564, B2 => 
                           n7168, ZN => n2821);
   U7332 : OAI22_X1 port map( A1 => n9566, A2 => n9806, B1 => n9564, B2 => 
                           n7167, ZN => n2822);
   U7333 : OAI22_X1 port map( A1 => n9566, A2 => n9809, B1 => n9564, B2 => 
                           n7166, ZN => n2823);
   U7334 : OAI22_X1 port map( A1 => n9567, A2 => n9812, B1 => n9564, B2 => 
                           n7165, ZN => n2824);
   U7335 : OAI22_X1 port map( A1 => n9567, A2 => n9815, B1 => n9564, B2 => 
                           n7164, ZN => n2825);
   U7336 : OAI22_X1 port map( A1 => n9567, A2 => n9818, B1 => n7468, B2 => 
                           n7163, ZN => n2826);
   U7337 : OAI22_X1 port map( A1 => n9567, A2 => n9821, B1 => n7468, B2 => 
                           n7162, ZN => n2827);
   U7338 : OAI22_X1 port map( A1 => n9567, A2 => n9824, B1 => n7468, B2 => 
                           n7161, ZN => n2828);
   U7339 : OAI22_X1 port map( A1 => n9568, A2 => n9827, B1 => n9564, B2 => 
                           n7160, ZN => n2829);
   U7340 : OAI22_X1 port map( A1 => n9568, A2 => n9830, B1 => n9564, B2 => 
                           n7159, ZN => n2830);
   U7341 : OAI22_X1 port map( A1 => n9568, A2 => n9833, B1 => n9564, B2 => 
                           n7158, ZN => n2831);
   U7342 : OAI22_X1 port map( A1 => n9568, A2 => n9836, B1 => n9564, B2 => 
                           n7157, ZN => n2832);
   U7343 : OAI22_X1 port map( A1 => n9568, A2 => n9839, B1 => n9564, B2 => 
                           n7156, ZN => n2833);
   U7344 : OAI22_X1 port map( A1 => n9569, A2 => n9842, B1 => n9564, B2 => 
                           n7155, ZN => n2834);
   U7345 : OAI22_X1 port map( A1 => n9569, A2 => n9845, B1 => n9564, B2 => 
                           n7154, ZN => n2835);
   U7346 : OAI22_X1 port map( A1 => n9569, A2 => n9848, B1 => n9564, B2 => 
                           n7153, ZN => n2836);
   U7347 : OAI22_X1 port map( A1 => n9569, A2 => n9851, B1 => n9564, B2 => 
                           n7152, ZN => n2837);
   U7348 : OAI22_X1 port map( A1 => n9574, A2 => n9780, B1 => n9573, B2 => 
                           n7143, ZN => n2846);
   U7349 : OAI22_X1 port map( A1 => n9574, A2 => n9784, B1 => n9573, B2 => 
                           n7142, ZN => n2847);
   U7350 : OAI22_X1 port map( A1 => n9574, A2 => n9787, B1 => n9573, B2 => 
                           n7141, ZN => n2848);
   U7351 : OAI22_X1 port map( A1 => n9574, A2 => n9790, B1 => n9573, B2 => 
                           n7140, ZN => n2849);
   U7352 : OAI22_X1 port map( A1 => n9574, A2 => n9793, B1 => n9573, B2 => 
                           n7139, ZN => n2850);
   U7353 : OAI22_X1 port map( A1 => n9575, A2 => n9796, B1 => n9573, B2 => 
                           n7138, ZN => n2851);
   U7354 : OAI22_X1 port map( A1 => n9575, A2 => n9799, B1 => n9573, B2 => 
                           n7137, ZN => n2852);
   U7355 : OAI22_X1 port map( A1 => n9575, A2 => n9802, B1 => n9573, B2 => 
                           n7136, ZN => n2853);
   U7356 : OAI22_X1 port map( A1 => n9575, A2 => n9805, B1 => n9573, B2 => 
                           n7135, ZN => n2854);
   U7357 : OAI22_X1 port map( A1 => n9575, A2 => n9808, B1 => n9573, B2 => 
                           n7134, ZN => n2855);
   U7358 : OAI22_X1 port map( A1 => n9576, A2 => n9811, B1 => n9573, B2 => 
                           n7133, ZN => n2856);
   U7359 : OAI22_X1 port map( A1 => n9576, A2 => n9814, B1 => n9573, B2 => 
                           n7132, ZN => n2857);
   U7360 : OAI22_X1 port map( A1 => n9576, A2 => n9817, B1 => n7467, B2 => 
                           n7131, ZN => n2858);
   U7361 : OAI22_X1 port map( A1 => n9576, A2 => n9820, B1 => n7467, B2 => 
                           n7130, ZN => n2859);
   U7362 : OAI22_X1 port map( A1 => n9576, A2 => n9823, B1 => n7467, B2 => 
                           n7129, ZN => n2860);
   U7363 : OAI22_X1 port map( A1 => n9577, A2 => n9826, B1 => n9573, B2 => 
                           n7128, ZN => n2861);
   U7364 : OAI22_X1 port map( A1 => n9577, A2 => n9829, B1 => n9573, B2 => 
                           n7127, ZN => n2862);
   U7365 : OAI22_X1 port map( A1 => n9577, A2 => n9832, B1 => n9573, B2 => 
                           n7126, ZN => n2863);
   U7366 : OAI22_X1 port map( A1 => n9577, A2 => n9835, B1 => n9573, B2 => 
                           n7125, ZN => n2864);
   U7367 : OAI22_X1 port map( A1 => n9577, A2 => n9838, B1 => n9573, B2 => 
                           n7124, ZN => n2865);
   U7368 : OAI22_X1 port map( A1 => n9578, A2 => n9841, B1 => n9573, B2 => 
                           n7123, ZN => n2866);
   U7369 : OAI22_X1 port map( A1 => n9578, A2 => n9844, B1 => n9573, B2 => 
                           n7122, ZN => n2867);
   U7370 : OAI22_X1 port map( A1 => n9578, A2 => n9847, B1 => n9573, B2 => 
                           n7121, ZN => n2868);
   U7371 : OAI22_X1 port map( A1 => n9578, A2 => n9850, B1 => n9573, B2 => 
                           n7120, ZN => n2869);
   U7372 : OAI22_X1 port map( A1 => n9583, A2 => n9780, B1 => n9582, B2 => 
                           n7111, ZN => n2878);
   U7373 : OAI22_X1 port map( A1 => n9583, A2 => n9784, B1 => n9582, B2 => 
                           n7110, ZN => n2879);
   U7374 : OAI22_X1 port map( A1 => n9583, A2 => n9787, B1 => n9582, B2 => 
                           n7109, ZN => n2880);
   U7375 : OAI22_X1 port map( A1 => n9583, A2 => n9790, B1 => n9582, B2 => 
                           n7108, ZN => n2881);
   U7376 : OAI22_X1 port map( A1 => n9583, A2 => n9793, B1 => n9582, B2 => 
                           n7107, ZN => n2882);
   U7377 : OAI22_X1 port map( A1 => n9584, A2 => n9796, B1 => n9582, B2 => 
                           n7106, ZN => n2883);
   U7378 : OAI22_X1 port map( A1 => n9584, A2 => n9799, B1 => n9582, B2 => 
                           n7105, ZN => n2884);
   U7379 : OAI22_X1 port map( A1 => n9584, A2 => n9802, B1 => n9582, B2 => 
                           n7104, ZN => n2885);
   U7380 : OAI22_X1 port map( A1 => n9584, A2 => n9805, B1 => n9582, B2 => 
                           n7103, ZN => n2886);
   U7381 : OAI22_X1 port map( A1 => n9584, A2 => n9808, B1 => n9582, B2 => 
                           n7102, ZN => n2887);
   U7382 : OAI22_X1 port map( A1 => n9585, A2 => n9811, B1 => n9582, B2 => 
                           n7101, ZN => n2888);
   U7383 : OAI22_X1 port map( A1 => n9585, A2 => n9814, B1 => n9582, B2 => 
                           n7100, ZN => n2889);
   U7384 : OAI22_X1 port map( A1 => n9585, A2 => n9817, B1 => n7466, B2 => 
                           n7099, ZN => n2890);
   U7385 : OAI22_X1 port map( A1 => n9585, A2 => n9820, B1 => n7466, B2 => 
                           n7098, ZN => n2891);
   U7386 : OAI22_X1 port map( A1 => n9585, A2 => n9823, B1 => n7466, B2 => 
                           n7097, ZN => n2892);
   U7387 : OAI22_X1 port map( A1 => n9586, A2 => n9826, B1 => n9582, B2 => 
                           n7096, ZN => n2893);
   U7388 : OAI22_X1 port map( A1 => n9586, A2 => n9829, B1 => n9582, B2 => 
                           n7095, ZN => n2894);
   U7389 : OAI22_X1 port map( A1 => n9586, A2 => n9832, B1 => n9582, B2 => 
                           n7094, ZN => n2895);
   U7390 : OAI22_X1 port map( A1 => n9586, A2 => n9835, B1 => n9582, B2 => 
                           n7093, ZN => n2896);
   U7391 : OAI22_X1 port map( A1 => n9586, A2 => n9838, B1 => n9582, B2 => 
                           n7092, ZN => n2897);
   U7392 : OAI22_X1 port map( A1 => n9587, A2 => n9841, B1 => n9582, B2 => 
                           n7091, ZN => n2898);
   U7393 : OAI22_X1 port map( A1 => n9587, A2 => n9844, B1 => n9582, B2 => 
                           n7090, ZN => n2899);
   U7394 : OAI22_X1 port map( A1 => n9587, A2 => n9847, B1 => n9582, B2 => 
                           n7089, ZN => n2900);
   U7395 : OAI22_X1 port map( A1 => n9587, A2 => n9850, B1 => n9582, B2 => 
                           n7088, ZN => n2901);
   U7396 : OAI22_X1 port map( A1 => n9610, A2 => n9781, B1 => n9609, B2 => 
                           n7015, ZN => n2974);
   U7397 : OAI22_X1 port map( A1 => n9610, A2 => n9784, B1 => n9609, B2 => 
                           n7014, ZN => n2975);
   U7398 : OAI22_X1 port map( A1 => n9610, A2 => n9787, B1 => n9609, B2 => 
                           n7013, ZN => n2976);
   U7399 : OAI22_X1 port map( A1 => n9610, A2 => n9790, B1 => n9609, B2 => 
                           n7012, ZN => n2977);
   U7400 : OAI22_X1 port map( A1 => n9610, A2 => n9793, B1 => n9609, B2 => 
                           n7011, ZN => n2978);
   U7401 : OAI22_X1 port map( A1 => n9611, A2 => n9796, B1 => n9609, B2 => 
                           n7010, ZN => n2979);
   U7402 : OAI22_X1 port map( A1 => n9611, A2 => n9799, B1 => n9609, B2 => 
                           n7009, ZN => n2980);
   U7403 : OAI22_X1 port map( A1 => n9611, A2 => n9802, B1 => n9609, B2 => 
                           n7008, ZN => n2981);
   U7404 : OAI22_X1 port map( A1 => n9611, A2 => n9805, B1 => n9609, B2 => 
                           n7007, ZN => n2982);
   U7405 : OAI22_X1 port map( A1 => n9611, A2 => n9808, B1 => n9609, B2 => 
                           n7006, ZN => n2983);
   U7406 : OAI22_X1 port map( A1 => n9612, A2 => n9811, B1 => n9609, B2 => 
                           n7005, ZN => n2984);
   U7407 : OAI22_X1 port map( A1 => n9612, A2 => n9814, B1 => n9609, B2 => 
                           n7004, ZN => n2985);
   U7408 : OAI22_X1 port map( A1 => n9612, A2 => n9817, B1 => n7463, B2 => 
                           n7003, ZN => n2986);
   U7409 : OAI22_X1 port map( A1 => n9612, A2 => n9820, B1 => n7463, B2 => 
                           n7002, ZN => n2987);
   U7410 : OAI22_X1 port map( A1 => n9612, A2 => n9823, B1 => n7463, B2 => 
                           n7001, ZN => n2988);
   U7411 : OAI22_X1 port map( A1 => n9613, A2 => n9826, B1 => n9609, B2 => 
                           n7000, ZN => n2989);
   U7412 : OAI22_X1 port map( A1 => n9613, A2 => n9829, B1 => n9609, B2 => 
                           n6999, ZN => n2990);
   U7413 : OAI22_X1 port map( A1 => n9613, A2 => n9832, B1 => n9609, B2 => 
                           n6998, ZN => n2991);
   U7414 : OAI22_X1 port map( A1 => n9613, A2 => n9835, B1 => n9609, B2 => 
                           n6997, ZN => n2992);
   U7415 : OAI22_X1 port map( A1 => n9613, A2 => n9838, B1 => n9609, B2 => 
                           n6996, ZN => n2993);
   U7416 : OAI22_X1 port map( A1 => n9614, A2 => n9841, B1 => n9609, B2 => 
                           n6995, ZN => n2994);
   U7417 : OAI22_X1 port map( A1 => n9614, A2 => n9844, B1 => n9609, B2 => 
                           n6994, ZN => n2995);
   U7418 : OAI22_X1 port map( A1 => n9614, A2 => n9847, B1 => n9609, B2 => 
                           n6993, ZN => n2996);
   U7419 : OAI22_X1 port map( A1 => n9614, A2 => n9850, B1 => n9609, B2 => 
                           n6992, ZN => n2997);
   U7420 : OAI22_X1 port map( A1 => n9619, A2 => n9781, B1 => n9618, B2 => 
                           n6983, ZN => n3006);
   U7421 : OAI22_X1 port map( A1 => n9619, A2 => n9784, B1 => n9618, B2 => 
                           n6982, ZN => n3007);
   U7422 : OAI22_X1 port map( A1 => n9619, A2 => n9787, B1 => n9618, B2 => 
                           n6981, ZN => n3008);
   U7423 : OAI22_X1 port map( A1 => n9619, A2 => n9790, B1 => n9618, B2 => 
                           n6980, ZN => n3009);
   U7424 : OAI22_X1 port map( A1 => n9619, A2 => n9793, B1 => n9618, B2 => 
                           n6979, ZN => n3010);
   U7425 : OAI22_X1 port map( A1 => n9620, A2 => n9796, B1 => n9618, B2 => 
                           n6978, ZN => n3011);
   U7426 : OAI22_X1 port map( A1 => n9620, A2 => n9799, B1 => n9618, B2 => 
                           n6977, ZN => n3012);
   U7427 : OAI22_X1 port map( A1 => n9620, A2 => n9802, B1 => n9618, B2 => 
                           n6976, ZN => n3013);
   U7428 : OAI22_X1 port map( A1 => n9620, A2 => n9805, B1 => n9618, B2 => 
                           n6975, ZN => n3014);
   U7429 : OAI22_X1 port map( A1 => n9620, A2 => n9808, B1 => n9618, B2 => 
                           n6974, ZN => n3015);
   U7430 : OAI22_X1 port map( A1 => n9621, A2 => n9811, B1 => n9618, B2 => 
                           n6973, ZN => n3016);
   U7431 : OAI22_X1 port map( A1 => n9621, A2 => n9814, B1 => n9618, B2 => 
                           n6972, ZN => n3017);
   U7432 : OAI22_X1 port map( A1 => n9621, A2 => n9817, B1 => n7462, B2 => 
                           n6971, ZN => n3018);
   U7433 : OAI22_X1 port map( A1 => n9621, A2 => n9820, B1 => n7462, B2 => 
                           n6970, ZN => n3019);
   U7434 : OAI22_X1 port map( A1 => n9621, A2 => n9823, B1 => n7462, B2 => 
                           n6969, ZN => n3020);
   U7435 : OAI22_X1 port map( A1 => n9622, A2 => n9826, B1 => n9618, B2 => 
                           n6968, ZN => n3021);
   U7436 : OAI22_X1 port map( A1 => n9622, A2 => n9829, B1 => n9618, B2 => 
                           n6967, ZN => n3022);
   U7437 : OAI22_X1 port map( A1 => n9622, A2 => n9832, B1 => n9618, B2 => 
                           n6966, ZN => n3023);
   U7438 : OAI22_X1 port map( A1 => n9622, A2 => n9835, B1 => n9618, B2 => 
                           n6965, ZN => n3024);
   U7439 : OAI22_X1 port map( A1 => n9622, A2 => n9838, B1 => n9618, B2 => 
                           n6964, ZN => n3025);
   U7440 : OAI22_X1 port map( A1 => n9623, A2 => n9841, B1 => n9618, B2 => 
                           n6963, ZN => n3026);
   U7441 : OAI22_X1 port map( A1 => n9623, A2 => n9844, B1 => n9618, B2 => 
                           n6962, ZN => n3027);
   U7442 : OAI22_X1 port map( A1 => n9623, A2 => n9847, B1 => n9618, B2 => 
                           n6961, ZN => n3028);
   U7443 : OAI22_X1 port map( A1 => n9623, A2 => n9850, B1 => n9618, B2 => 
                           n6960, ZN => n3029);
   U7444 : OAI22_X1 port map( A1 => n9646, A2 => n9781, B1 => n9645, B2 => 
                           n6887, ZN => n3102);
   U7445 : OAI22_X1 port map( A1 => n9646, A2 => n9784, B1 => n9645, B2 => 
                           n6886, ZN => n3103);
   U7446 : OAI22_X1 port map( A1 => n9646, A2 => n9787, B1 => n9645, B2 => 
                           n6885, ZN => n3104);
   U7447 : OAI22_X1 port map( A1 => n9646, A2 => n9790, B1 => n9645, B2 => 
                           n6884, ZN => n3105);
   U7448 : OAI22_X1 port map( A1 => n9646, A2 => n9793, B1 => n9645, B2 => 
                           n6883, ZN => n3106);
   U7449 : OAI22_X1 port map( A1 => n9647, A2 => n9796, B1 => n9645, B2 => 
                           n6882, ZN => n3107);
   U7450 : OAI22_X1 port map( A1 => n9647, A2 => n9799, B1 => n9645, B2 => 
                           n6881, ZN => n3108);
   U7451 : OAI22_X1 port map( A1 => n9647, A2 => n9802, B1 => n9645, B2 => 
                           n6880, ZN => n3109);
   U7452 : OAI22_X1 port map( A1 => n9647, A2 => n9805, B1 => n9645, B2 => 
                           n6879, ZN => n3110);
   U7453 : OAI22_X1 port map( A1 => n9647, A2 => n9808, B1 => n9645, B2 => 
                           n6878, ZN => n3111);
   U7454 : OAI22_X1 port map( A1 => n9648, A2 => n9811, B1 => n9645, B2 => 
                           n6877, ZN => n3112);
   U7455 : OAI22_X1 port map( A1 => n9648, A2 => n9814, B1 => n9645, B2 => 
                           n6876, ZN => n3113);
   U7456 : OAI22_X1 port map( A1 => n9648, A2 => n9817, B1 => n7458, B2 => 
                           n6875, ZN => n3114);
   U7457 : OAI22_X1 port map( A1 => n9648, A2 => n9820, B1 => n7458, B2 => 
                           n6874, ZN => n3115);
   U7458 : OAI22_X1 port map( A1 => n9648, A2 => n9823, B1 => n7458, B2 => 
                           n6873, ZN => n3116);
   U7459 : OAI22_X1 port map( A1 => n9649, A2 => n9826, B1 => n9645, B2 => 
                           n6872, ZN => n3117);
   U7460 : OAI22_X1 port map( A1 => n9649, A2 => n9829, B1 => n9645, B2 => 
                           n6871, ZN => n3118);
   U7461 : OAI22_X1 port map( A1 => n9649, A2 => n9832, B1 => n9645, B2 => 
                           n6870, ZN => n3119);
   U7462 : OAI22_X1 port map( A1 => n9649, A2 => n9835, B1 => n9645, B2 => 
                           n6869, ZN => n3120);
   U7463 : OAI22_X1 port map( A1 => n9649, A2 => n9838, B1 => n9645, B2 => 
                           n6868, ZN => n3121);
   U7464 : OAI22_X1 port map( A1 => n9650, A2 => n9841, B1 => n9645, B2 => 
                           n6867, ZN => n3122);
   U7465 : OAI22_X1 port map( A1 => n9650, A2 => n9844, B1 => n9645, B2 => 
                           n6866, ZN => n3123);
   U7466 : OAI22_X1 port map( A1 => n9650, A2 => n9847, B1 => n9645, B2 => 
                           n6865, ZN => n3124);
   U7467 : OAI22_X1 port map( A1 => n9650, A2 => n9850, B1 => n9645, B2 => 
                           n6864, ZN => n3125);
   U7468 : OAI22_X1 port map( A1 => n9655, A2 => n9781, B1 => n9654, B2 => 
                           n6855, ZN => n3134);
   U7469 : OAI22_X1 port map( A1 => n9655, A2 => n9784, B1 => n9654, B2 => 
                           n6854, ZN => n3135);
   U7470 : OAI22_X1 port map( A1 => n9655, A2 => n9787, B1 => n9654, B2 => 
                           n6853, ZN => n3136);
   U7471 : OAI22_X1 port map( A1 => n9655, A2 => n9790, B1 => n9654, B2 => 
                           n6852, ZN => n3137);
   U7472 : OAI22_X1 port map( A1 => n9655, A2 => n9793, B1 => n9654, B2 => 
                           n6851, ZN => n3138);
   U7473 : OAI22_X1 port map( A1 => n9656, A2 => n9796, B1 => n9654, B2 => 
                           n6850, ZN => n3139);
   U7474 : OAI22_X1 port map( A1 => n9656, A2 => n9799, B1 => n9654, B2 => 
                           n6849, ZN => n3140);
   U7475 : OAI22_X1 port map( A1 => n9656, A2 => n9802, B1 => n9654, B2 => 
                           n6848, ZN => n3141);
   U7476 : OAI22_X1 port map( A1 => n9656, A2 => n9805, B1 => n9654, B2 => 
                           n6847, ZN => n3142);
   U7477 : OAI22_X1 port map( A1 => n9656, A2 => n9808, B1 => n9654, B2 => 
                           n6846, ZN => n3143);
   U7478 : OAI22_X1 port map( A1 => n9657, A2 => n9811, B1 => n9654, B2 => 
                           n6845, ZN => n3144);
   U7479 : OAI22_X1 port map( A1 => n9657, A2 => n9814, B1 => n9654, B2 => 
                           n6844, ZN => n3145);
   U7480 : OAI22_X1 port map( A1 => n9657, A2 => n9817, B1 => n7457, B2 => 
                           n6843, ZN => n3146);
   U7481 : OAI22_X1 port map( A1 => n9657, A2 => n9820, B1 => n7457, B2 => 
                           n6842, ZN => n3147);
   U7482 : OAI22_X1 port map( A1 => n9657, A2 => n9823, B1 => n7457, B2 => 
                           n6841, ZN => n3148);
   U7483 : OAI22_X1 port map( A1 => n9658, A2 => n9826, B1 => n9654, B2 => 
                           n6840, ZN => n3149);
   U7484 : OAI22_X1 port map( A1 => n9658, A2 => n9829, B1 => n9654, B2 => 
                           n6839, ZN => n3150);
   U7485 : OAI22_X1 port map( A1 => n9658, A2 => n9832, B1 => n9654, B2 => 
                           n6838, ZN => n3151);
   U7486 : OAI22_X1 port map( A1 => n9658, A2 => n9835, B1 => n9654, B2 => 
                           n6837, ZN => n3152);
   U7487 : OAI22_X1 port map( A1 => n9658, A2 => n9838, B1 => n9654, B2 => 
                           n6836, ZN => n3153);
   U7488 : OAI22_X1 port map( A1 => n9659, A2 => n9841, B1 => n9654, B2 => 
                           n6835, ZN => n3154);
   U7489 : OAI22_X1 port map( A1 => n9659, A2 => n9844, B1 => n9654, B2 => 
                           n6834, ZN => n3155);
   U7490 : OAI22_X1 port map( A1 => n9659, A2 => n9847, B1 => n9654, B2 => 
                           n6833, ZN => n3156);
   U7491 : OAI22_X1 port map( A1 => n9659, A2 => n9850, B1 => n9654, B2 => 
                           n6832, ZN => n3157);
   U7492 : OAI22_X1 port map( A1 => n9682, A2 => n9781, B1 => n9681, B2 => 
                           n6759, ZN => n3230);
   U7493 : OAI22_X1 port map( A1 => n9682, A2 => n9783, B1 => n9681, B2 => 
                           n6758, ZN => n3231);
   U7494 : OAI22_X1 port map( A1 => n9682, A2 => n9786, B1 => n9681, B2 => 
                           n6757, ZN => n3232);
   U7495 : OAI22_X1 port map( A1 => n9682, A2 => n9789, B1 => n9681, B2 => 
                           n6756, ZN => n3233);
   U7496 : OAI22_X1 port map( A1 => n9682, A2 => n9792, B1 => n9681, B2 => 
                           n6755, ZN => n3234);
   U7497 : OAI22_X1 port map( A1 => n9683, A2 => n9795, B1 => n9681, B2 => 
                           n6754, ZN => n3235);
   U7498 : OAI22_X1 port map( A1 => n9683, A2 => n9798, B1 => n9681, B2 => 
                           n6753, ZN => n3236);
   U7499 : OAI22_X1 port map( A1 => n9683, A2 => n9801, B1 => n9681, B2 => 
                           n6752, ZN => n3237);
   U7500 : OAI22_X1 port map( A1 => n9683, A2 => n9804, B1 => n9681, B2 => 
                           n6751, ZN => n3238);
   U7501 : OAI22_X1 port map( A1 => n9683, A2 => n9807, B1 => n9681, B2 => 
                           n6750, ZN => n3239);
   U7502 : OAI22_X1 port map( A1 => n9684, A2 => n9810, B1 => n9681, B2 => 
                           n6749, ZN => n3240);
   U7503 : OAI22_X1 port map( A1 => n9684, A2 => n9813, B1 => n9681, B2 => 
                           n6748, ZN => n3241);
   U7504 : OAI22_X1 port map( A1 => n9684, A2 => n9816, B1 => n7454, B2 => 
                           n6747, ZN => n3242);
   U7505 : OAI22_X1 port map( A1 => n9684, A2 => n9819, B1 => n7454, B2 => 
                           n6746, ZN => n3243);
   U7506 : OAI22_X1 port map( A1 => n9684, A2 => n9822, B1 => n7454, B2 => 
                           n6745, ZN => n3244);
   U7507 : OAI22_X1 port map( A1 => n9685, A2 => n9825, B1 => n9681, B2 => 
                           n6744, ZN => n3245);
   U7508 : OAI22_X1 port map( A1 => n9685, A2 => n9828, B1 => n9681, B2 => 
                           n6743, ZN => n3246);
   U7509 : OAI22_X1 port map( A1 => n9685, A2 => n9831, B1 => n9681, B2 => 
                           n6742, ZN => n3247);
   U7510 : OAI22_X1 port map( A1 => n9685, A2 => n9834, B1 => n9681, B2 => 
                           n6741, ZN => n3248);
   U7511 : OAI22_X1 port map( A1 => n9685, A2 => n9837, B1 => n9681, B2 => 
                           n6740, ZN => n3249);
   U7512 : OAI22_X1 port map( A1 => n9686, A2 => n9840, B1 => n9681, B2 => 
                           n6739, ZN => n3250);
   U7513 : OAI22_X1 port map( A1 => n9686, A2 => n9843, B1 => n9681, B2 => 
                           n6738, ZN => n3251);
   U7514 : OAI22_X1 port map( A1 => n9686, A2 => n9846, B1 => n9681, B2 => 
                           n6737, ZN => n3252);
   U7515 : OAI22_X1 port map( A1 => n9686, A2 => n9849, B1 => n9681, B2 => 
                           n6736, ZN => n3253);
   U7516 : OAI22_X1 port map( A1 => n9691, A2 => n9781, B1 => n9690, B2 => 
                           n6727, ZN => n3262);
   U7517 : OAI22_X1 port map( A1 => n9691, A2 => n9783, B1 => n9690, B2 => 
                           n6726, ZN => n3263);
   U7518 : OAI22_X1 port map( A1 => n9691, A2 => n9786, B1 => n9690, B2 => 
                           n6725, ZN => n3264);
   U7519 : OAI22_X1 port map( A1 => n9691, A2 => n9789, B1 => n9690, B2 => 
                           n6724, ZN => n3265);
   U7520 : OAI22_X1 port map( A1 => n9691, A2 => n9792, B1 => n9690, B2 => 
                           n6723, ZN => n3266);
   U7521 : OAI22_X1 port map( A1 => n9692, A2 => n9795, B1 => n9690, B2 => 
                           n6722, ZN => n3267);
   U7522 : OAI22_X1 port map( A1 => n9692, A2 => n9798, B1 => n9690, B2 => 
                           n6721, ZN => n3268);
   U7523 : OAI22_X1 port map( A1 => n9692, A2 => n9801, B1 => n9690, B2 => 
                           n6720, ZN => n3269);
   U7524 : OAI22_X1 port map( A1 => n9692, A2 => n9804, B1 => n9690, B2 => 
                           n6719, ZN => n3270);
   U7525 : OAI22_X1 port map( A1 => n9692, A2 => n9807, B1 => n9690, B2 => 
                           n6718, ZN => n3271);
   U7526 : OAI22_X1 port map( A1 => n9693, A2 => n9810, B1 => n9690, B2 => 
                           n6717, ZN => n3272);
   U7527 : OAI22_X1 port map( A1 => n9693, A2 => n9813, B1 => n9690, B2 => 
                           n6716, ZN => n3273);
   U7528 : OAI22_X1 port map( A1 => n9693, A2 => n9816, B1 => n7453, B2 => 
                           n6715, ZN => n3274);
   U7529 : OAI22_X1 port map( A1 => n9693, A2 => n9819, B1 => n7453, B2 => 
                           n6714, ZN => n3275);
   U7530 : OAI22_X1 port map( A1 => n9693, A2 => n9822, B1 => n7453, B2 => 
                           n6713, ZN => n3276);
   U7531 : OAI22_X1 port map( A1 => n9694, A2 => n9825, B1 => n9690, B2 => 
                           n6712, ZN => n3277);
   U7532 : OAI22_X1 port map( A1 => n9694, A2 => n9828, B1 => n9690, B2 => 
                           n6711, ZN => n3278);
   U7533 : OAI22_X1 port map( A1 => n9694, A2 => n9831, B1 => n9690, B2 => 
                           n6710, ZN => n3279);
   U7534 : OAI22_X1 port map( A1 => n9694, A2 => n9834, B1 => n9690, B2 => 
                           n6709, ZN => n3280);
   U7535 : OAI22_X1 port map( A1 => n9694, A2 => n9837, B1 => n9690, B2 => 
                           n6708, ZN => n3281);
   U7536 : OAI22_X1 port map( A1 => n9695, A2 => n9840, B1 => n9690, B2 => 
                           n6707, ZN => n3282);
   U7537 : OAI22_X1 port map( A1 => n9695, A2 => n9843, B1 => n9690, B2 => 
                           n6706, ZN => n3283);
   U7538 : OAI22_X1 port map( A1 => n9695, A2 => n9846, B1 => n9690, B2 => 
                           n6705, ZN => n3284);
   U7539 : OAI22_X1 port map( A1 => n9695, A2 => n9849, B1 => n9690, B2 => 
                           n6704, ZN => n3285);
   U7540 : OAI22_X1 port map( A1 => n9700, A2 => n9781, B1 => n9699, B2 => 
                           n6695, ZN => n3294);
   U7541 : OAI22_X1 port map( A1 => n9700, A2 => n9783, B1 => n9699, B2 => 
                           n6694, ZN => n3295);
   U7542 : OAI22_X1 port map( A1 => n9700, A2 => n9786, B1 => n9699, B2 => 
                           n6693, ZN => n3296);
   U7543 : OAI22_X1 port map( A1 => n9700, A2 => n9789, B1 => n9699, B2 => 
                           n6692, ZN => n3297);
   U7544 : OAI22_X1 port map( A1 => n9700, A2 => n9792, B1 => n9699, B2 => 
                           n6691, ZN => n3298);
   U7545 : OAI22_X1 port map( A1 => n9701, A2 => n9795, B1 => n9699, B2 => 
                           n6690, ZN => n3299);
   U7546 : OAI22_X1 port map( A1 => n9701, A2 => n9798, B1 => n9699, B2 => 
                           n6689, ZN => n3300);
   U7547 : OAI22_X1 port map( A1 => n9701, A2 => n9801, B1 => n9699, B2 => 
                           n6688, ZN => n3301);
   U7548 : OAI22_X1 port map( A1 => n9701, A2 => n9804, B1 => n9699, B2 => 
                           n6687, ZN => n3302);
   U7549 : OAI22_X1 port map( A1 => n9701, A2 => n9807, B1 => n9699, B2 => 
                           n6686, ZN => n3303);
   U7550 : OAI22_X1 port map( A1 => n9702, A2 => n9810, B1 => n9699, B2 => 
                           n6685, ZN => n3304);
   U7551 : OAI22_X1 port map( A1 => n9702, A2 => n9813, B1 => n9699, B2 => 
                           n6684, ZN => n3305);
   U7552 : OAI22_X1 port map( A1 => n9702, A2 => n9816, B1 => n7452, B2 => 
                           n6683, ZN => n3306);
   U7553 : OAI22_X1 port map( A1 => n9702, A2 => n9819, B1 => n7452, B2 => 
                           n6682, ZN => n3307);
   U7554 : OAI22_X1 port map( A1 => n9702, A2 => n9822, B1 => n7452, B2 => 
                           n6681, ZN => n3308);
   U7555 : OAI22_X1 port map( A1 => n9703, A2 => n9825, B1 => n9699, B2 => 
                           n6680, ZN => n3309);
   U7556 : OAI22_X1 port map( A1 => n9703, A2 => n9828, B1 => n9699, B2 => 
                           n6679, ZN => n3310);
   U7557 : OAI22_X1 port map( A1 => n9703, A2 => n9831, B1 => n9699, B2 => 
                           n6678, ZN => n3311);
   U7558 : OAI22_X1 port map( A1 => n9703, A2 => n9834, B1 => n9699, B2 => 
                           n6677, ZN => n3312);
   U7559 : OAI22_X1 port map( A1 => n9703, A2 => n9837, B1 => n9699, B2 => 
                           n6676, ZN => n3313);
   U7560 : OAI22_X1 port map( A1 => n9704, A2 => n9840, B1 => n9699, B2 => 
                           n6675, ZN => n3314);
   U7561 : OAI22_X1 port map( A1 => n9704, A2 => n9843, B1 => n9699, B2 => 
                           n6674, ZN => n3315);
   U7562 : OAI22_X1 port map( A1 => n9704, A2 => n9846, B1 => n9699, B2 => 
                           n6673, ZN => n3316);
   U7563 : OAI22_X1 port map( A1 => n9704, A2 => n9849, B1 => n9699, B2 => 
                           n6672, ZN => n3317);
   U7564 : OAI22_X1 port map( A1 => n9709, A2 => n9781, B1 => n9708, B2 => 
                           n6663, ZN => n3326);
   U7565 : OAI22_X1 port map( A1 => n9709, A2 => n9783, B1 => n9708, B2 => 
                           n6662, ZN => n3327);
   U7566 : OAI22_X1 port map( A1 => n9709, A2 => n9786, B1 => n9708, B2 => 
                           n6661, ZN => n3328);
   U7567 : OAI22_X1 port map( A1 => n9709, A2 => n9789, B1 => n9708, B2 => 
                           n6660, ZN => n3329);
   U7568 : OAI22_X1 port map( A1 => n9709, A2 => n9792, B1 => n9708, B2 => 
                           n6659, ZN => n3330);
   U7569 : OAI22_X1 port map( A1 => n9710, A2 => n9795, B1 => n9708, B2 => 
                           n6658, ZN => n3331);
   U7570 : OAI22_X1 port map( A1 => n9710, A2 => n9798, B1 => n9708, B2 => 
                           n6657, ZN => n3332);
   U7571 : OAI22_X1 port map( A1 => n9710, A2 => n9801, B1 => n9708, B2 => 
                           n6656, ZN => n3333);
   U7572 : OAI22_X1 port map( A1 => n9710, A2 => n9804, B1 => n9708, B2 => 
                           n6655, ZN => n3334);
   U7573 : OAI22_X1 port map( A1 => n9710, A2 => n9807, B1 => n9708, B2 => 
                           n6654, ZN => n3335);
   U7574 : OAI22_X1 port map( A1 => n9711, A2 => n9810, B1 => n9708, B2 => 
                           n6653, ZN => n3336);
   U7575 : OAI22_X1 port map( A1 => n9711, A2 => n9813, B1 => n9708, B2 => 
                           n6652, ZN => n3337);
   U7576 : OAI22_X1 port map( A1 => n9711, A2 => n9816, B1 => n7450, B2 => 
                           n6651, ZN => n3338);
   U7577 : OAI22_X1 port map( A1 => n9711, A2 => n9819, B1 => n7450, B2 => 
                           n6650, ZN => n3339);
   U7578 : OAI22_X1 port map( A1 => n9711, A2 => n9822, B1 => n7450, B2 => 
                           n6649, ZN => n3340);
   U7579 : OAI22_X1 port map( A1 => n9712, A2 => n9825, B1 => n9708, B2 => 
                           n6648, ZN => n3341);
   U7580 : OAI22_X1 port map( A1 => n9712, A2 => n9828, B1 => n9708, B2 => 
                           n6647, ZN => n3342);
   U7581 : OAI22_X1 port map( A1 => n9712, A2 => n9831, B1 => n9708, B2 => 
                           n6646, ZN => n3343);
   U7582 : OAI22_X1 port map( A1 => n9712, A2 => n9834, B1 => n9708, B2 => 
                           n6645, ZN => n3344);
   U7583 : OAI22_X1 port map( A1 => n9712, A2 => n9837, B1 => n9708, B2 => 
                           n6644, ZN => n3345);
   U7584 : OAI22_X1 port map( A1 => n9713, A2 => n9840, B1 => n9708, B2 => 
                           n6643, ZN => n3346);
   U7585 : OAI22_X1 port map( A1 => n9713, A2 => n9843, B1 => n9708, B2 => 
                           n6642, ZN => n3347);
   U7586 : OAI22_X1 port map( A1 => n9713, A2 => n9846, B1 => n9708, B2 => 
                           n6641, ZN => n3348);
   U7587 : OAI22_X1 port map( A1 => n9713, A2 => n9849, B1 => n9708, B2 => 
                           n6640, ZN => n3349);
   U7588 : NOR2_X1 port map( A1 => n6458, A2 => n6459, ZN => n8765);
   U7589 : NOR2_X1 port map( A1 => n6462, A2 => n6463, ZN => n8112);
   U7590 : BUF_X1 port map( A => n8130, Z => n9393);
   U7591 : BUF_X1 port map( A => n7477, Z => n9495);
   U7592 : BUF_X1 port map( A => n8130, Z => n9394);
   U7593 : BUF_X1 port map( A => n8130, Z => n9395);
   U7594 : BUF_X1 port map( A => n7477, Z => n9496);
   U7595 : BUF_X1 port map( A => n7477, Z => n9497);
   U7596 : BUF_X1 port map( A => n6451, Z => n9888);
   U7597 : BUF_X1 port map( A => n6451, Z => n9889);
   U7598 : BUF_X1 port map( A => n6451, Z => n9886);
   U7599 : BUF_X1 port map( A => n6451, Z => n9885);
   U7600 : BUF_X1 port map( A => n7432, Z => n9780);
   U7601 : BUF_X1 port map( A => n7431, Z => n9784);
   U7602 : BUF_X1 port map( A => n7430, Z => n9787);
   U7603 : BUF_X1 port map( A => n7429, Z => n9790);
   U7604 : BUF_X1 port map( A => n7428, Z => n9793);
   U7605 : BUF_X1 port map( A => n7427, Z => n9796);
   U7606 : BUF_X1 port map( A => n7426, Z => n9799);
   U7607 : BUF_X1 port map( A => n7425, Z => n9802);
   U7608 : BUF_X1 port map( A => n7424, Z => n9805);
   U7609 : BUF_X1 port map( A => n7423, Z => n9808);
   U7610 : BUF_X1 port map( A => n7422, Z => n9811);
   U7611 : BUF_X1 port map( A => n7421, Z => n9814);
   U7612 : BUF_X1 port map( A => n7420, Z => n9817);
   U7613 : BUF_X1 port map( A => n7419, Z => n9820);
   U7614 : BUF_X1 port map( A => n7418, Z => n9823);
   U7615 : BUF_X1 port map( A => n7417, Z => n9826);
   U7616 : BUF_X1 port map( A => n7416, Z => n9829);
   U7617 : BUF_X1 port map( A => n7415, Z => n9832);
   U7618 : BUF_X1 port map( A => n7414, Z => n9835);
   U7619 : BUF_X1 port map( A => n7413, Z => n9838);
   U7620 : BUF_X1 port map( A => n7412, Z => n9841);
   U7621 : BUF_X1 port map( A => n7411, Z => n9844);
   U7622 : BUF_X1 port map( A => n7410, Z => n9847);
   U7623 : BUF_X1 port map( A => n7409, Z => n9850);
   U7624 : BUF_X1 port map( A => n7408, Z => n9853);
   U7625 : BUF_X1 port map( A => n7407, Z => n9856);
   U7626 : BUF_X1 port map( A => n7406, Z => n9859);
   U7627 : BUF_X1 port map( A => n7405, Z => n9862);
   U7628 : BUF_X1 port map( A => n7404, Z => n9865);
   U7629 : BUF_X1 port map( A => n7403, Z => n9868);
   U7630 : BUF_X1 port map( A => n7402, Z => n9871);
   U7631 : BUF_X1 port map( A => n7400, Z => n9883);
   U7632 : BUF_X1 port map( A => n7432, Z => n9781);
   U7633 : BUF_X1 port map( A => n7431, Z => n9783);
   U7634 : BUF_X1 port map( A => n7430, Z => n9786);
   U7635 : BUF_X1 port map( A => n7429, Z => n9789);
   U7636 : BUF_X1 port map( A => n7428, Z => n9792);
   U7637 : BUF_X1 port map( A => n7427, Z => n9795);
   U7638 : BUF_X1 port map( A => n7426, Z => n9798);
   U7639 : BUF_X1 port map( A => n7425, Z => n9801);
   U7640 : BUF_X1 port map( A => n7424, Z => n9804);
   U7641 : BUF_X1 port map( A => n7423, Z => n9807);
   U7642 : BUF_X1 port map( A => n7422, Z => n9810);
   U7643 : BUF_X1 port map( A => n7421, Z => n9813);
   U7644 : BUF_X1 port map( A => n7420, Z => n9816);
   U7645 : BUF_X1 port map( A => n7419, Z => n9819);
   U7646 : BUF_X1 port map( A => n7418, Z => n9822);
   U7647 : BUF_X1 port map( A => n7417, Z => n9825);
   U7648 : BUF_X1 port map( A => n7416, Z => n9828);
   U7649 : BUF_X1 port map( A => n7415, Z => n9831);
   U7650 : BUF_X1 port map( A => n7414, Z => n9834);
   U7651 : BUF_X1 port map( A => n7413, Z => n9837);
   U7652 : BUF_X1 port map( A => n7412, Z => n9840);
   U7653 : BUF_X1 port map( A => n7411, Z => n9843);
   U7654 : BUF_X1 port map( A => n7410, Z => n9846);
   U7655 : BUF_X1 port map( A => n7409, Z => n9849);
   U7656 : BUF_X1 port map( A => n7408, Z => n9852);
   U7657 : BUF_X1 port map( A => n7407, Z => n9855);
   U7658 : BUF_X1 port map( A => n7406, Z => n9858);
   U7659 : BUF_X1 port map( A => n7405, Z => n9861);
   U7660 : BUF_X1 port map( A => n7404, Z => n9864);
   U7661 : BUF_X1 port map( A => n7403, Z => n9867);
   U7662 : BUF_X1 port map( A => n7402, Z => n9870);
   U7663 : BUF_X1 port map( A => n7400, Z => n9882);
   U7664 : BUF_X1 port map( A => n6451, Z => n9887);
   U7665 : BUF_X1 port map( A => n8130, Z => n9391);
   U7666 : BUF_X1 port map( A => n8130, Z => n9392);
   U7667 : BUF_X1 port map( A => n7477, Z => n9493);
   U7668 : BUF_X1 port map( A => n7477, Z => n9494);
   U7669 : BUF_X1 port map( A => n7432, Z => n9782);
   U7670 : BUF_X1 port map( A => n7431, Z => n9785);
   U7671 : BUF_X1 port map( A => n7430, Z => n9788);
   U7672 : BUF_X1 port map( A => n7429, Z => n9791);
   U7673 : BUF_X1 port map( A => n7428, Z => n9794);
   U7674 : BUF_X1 port map( A => n7427, Z => n9797);
   U7675 : BUF_X1 port map( A => n7426, Z => n9800);
   U7676 : BUF_X1 port map( A => n7425, Z => n9803);
   U7677 : BUF_X1 port map( A => n7424, Z => n9806);
   U7678 : BUF_X1 port map( A => n7423, Z => n9809);
   U7679 : BUF_X1 port map( A => n7422, Z => n9812);
   U7680 : BUF_X1 port map( A => n7421, Z => n9815);
   U7681 : BUF_X1 port map( A => n7420, Z => n9818);
   U7682 : BUF_X1 port map( A => n7419, Z => n9821);
   U7683 : BUF_X1 port map( A => n7418, Z => n9824);
   U7684 : BUF_X1 port map( A => n7417, Z => n9827);
   U7685 : BUF_X1 port map( A => n7416, Z => n9830);
   U7686 : BUF_X1 port map( A => n7415, Z => n9833);
   U7687 : BUF_X1 port map( A => n7414, Z => n9836);
   U7688 : BUF_X1 port map( A => n7413, Z => n9839);
   U7689 : BUF_X1 port map( A => n7412, Z => n9842);
   U7690 : BUF_X1 port map( A => n7411, Z => n9845);
   U7691 : BUF_X1 port map( A => n7410, Z => n9848);
   U7692 : BUF_X1 port map( A => n7409, Z => n9851);
   U7693 : BUF_X1 port map( A => n7408, Z => n9854);
   U7694 : BUF_X1 port map( A => n7407, Z => n9857);
   U7695 : BUF_X1 port map( A => n7406, Z => n9860);
   U7696 : BUF_X1 port map( A => n7405, Z => n9863);
   U7697 : BUF_X1 port map( A => n7404, Z => n9866);
   U7698 : BUF_X1 port map( A => n7403, Z => n9869);
   U7699 : BUF_X1 port map( A => n7402, Z => n9872);
   U7700 : BUF_X1 port map( A => n7400, Z => n9884);
   U7701 : NAND2_X1 port map( A1 => n8763, A2 => n8777, ZN => n8165);
   U7702 : NAND2_X1 port map( A1 => n8763, A2 => n8776, ZN => n8166);
   U7703 : NAND2_X1 port map( A1 => n8765, A2 => n8776, ZN => n8170);
   U7704 : NAND2_X1 port map( A1 => n8765, A2 => n8777, ZN => n8171);
   U7705 : NAND2_X1 port map( A1 => n8112, A2 => n8123, ZN => n7517);
   U7706 : NAND2_X1 port map( A1 => n8112, A2 => n8124, ZN => n7518);
   U7707 : NAND2_X1 port map( A1 => n8110, A2 => n8124, ZN => n7512);
   U7708 : NAND2_X1 port map( A1 => n8110, A2 => n8123, ZN => n7513);
   U7709 : NAND2_X1 port map( A1 => n8781, A2 => n8763, ZN => n8175);
   U7710 : NAND2_X1 port map( A1 => n8781, A2 => n8765, ZN => n8180);
   U7711 : NAND2_X1 port map( A1 => n8128, A2 => n8108, ZN => n7522);
   U7712 : NAND2_X1 port map( A1 => n8128, A2 => n8112, ZN => n7527);
   U7713 : NAND2_X1 port map( A1 => n8780, A2 => n8763, ZN => n8176);
   U7714 : NAND2_X1 port map( A1 => n8780, A2 => n8765, ZN => n8181);
   U7715 : NAND2_X1 port map( A1 => n8127, A2 => n8108, ZN => n7523);
   U7716 : NAND2_X1 port map( A1 => n8127, A2 => n8112, ZN => n7528);
   U7717 : NAND2_X1 port map( A1 => n8769, A2 => n8763, ZN => n8151);
   U7718 : NAND2_X1 port map( A1 => n8768, A2 => n8763, ZN => n8152);
   U7719 : NAND2_X1 port map( A1 => n8762, A2 => n8765, ZN => n8146);
   U7720 : NAND2_X1 port map( A1 => n8760, A2 => n8765, ZN => n8147);
   U7721 : NAND2_X1 port map( A1 => n8109, A2 => n8112, ZN => n7493);
   U7722 : NAND2_X1 port map( A1 => n8107, A2 => n8112, ZN => n7494);
   U7723 : NAND2_X1 port map( A1 => n8109, A2 => n8108, ZN => n7488);
   U7724 : NAND2_X1 port map( A1 => n8107, A2 => n8108, ZN => n7489);
   U7725 : NAND2_X1 port map( A1 => n8116, A2 => n8110, ZN => n7498);
   U7726 : NAND2_X1 port map( A1 => n8115, A2 => n8110, ZN => n7499);
   U7727 : NAND2_X1 port map( A1 => n8762, A2 => n8761, ZN => n8141);
   U7728 : NAND2_X1 port map( A1 => n8760, A2 => n8761, ZN => n8142);
   U7729 : NAND2_X1 port map( A1 => n8769, A2 => n8766, ZN => n8156);
   U7730 : NAND2_X1 port map( A1 => n8768, A2 => n8766, ZN => n8157);
   U7731 : NAND2_X1 port map( A1 => n8116, A2 => n8113, ZN => n7503);
   U7732 : NAND2_X1 port map( A1 => n8115, A2 => n8113, ZN => n7504);
   U7733 : AND2_X1 port map( A1 => n8108, A2 => n8124, ZN => n7509);
   U7734 : AND2_X1 port map( A1 => n8776, A2 => n8761, ZN => n8163);
   U7735 : AND2_X1 port map( A1 => n8123, A2 => n8108, ZN => n7510);
   U7736 : AND2_X1 port map( A1 => n8761, A2 => n8777, ZN => n8162);
   U7737 : AND2_X1 port map( A1 => n8766, A2 => n8776, ZN => n8167);
   U7738 : AND2_X1 port map( A1 => n8766, A2 => n8777, ZN => n8168);
   U7739 : AND2_X1 port map( A1 => n8113, A2 => n8123, ZN => n7514);
   U7740 : AND2_X1 port map( A1 => n8113, A2 => n8124, ZN => n7515);
   U7741 : AND2_X1 port map( A1 => n8762, A2 => n8763, ZN => n8138);
   U7742 : AND2_X1 port map( A1 => n8760, A2 => n8763, ZN => n8139);
   U7743 : AND2_X1 port map( A1 => n8769, A2 => n8765, ZN => n8153);
   U7744 : AND2_X1 port map( A1 => n8768, A2 => n8765, ZN => n8154);
   U7745 : AND2_X1 port map( A1 => n8116, A2 => n8112, ZN => n7500);
   U7746 : AND2_X1 port map( A1 => n8115, A2 => n8112, ZN => n7501);
   U7747 : AND2_X1 port map( A1 => n8781, A2 => n8761, ZN => n8172);
   U7748 : AND2_X1 port map( A1 => n8780, A2 => n8761, ZN => n8173);
   U7749 : AND2_X1 port map( A1 => n8781, A2 => n8766, ZN => n8177);
   U7750 : AND2_X1 port map( A1 => n8780, A2 => n8766, ZN => n8178);
   U7751 : AND2_X1 port map( A1 => n8128, A2 => n8110, ZN => n7519);
   U7752 : AND2_X1 port map( A1 => n8127, A2 => n8110, ZN => n7520);
   U7753 : AND2_X1 port map( A1 => n8128, A2 => n8113, ZN => n7524);
   U7754 : AND2_X1 port map( A1 => n8127, A2 => n8113, ZN => n7525);
   U7755 : AND2_X1 port map( A1 => n8116, A2 => n8108, ZN => n7495);
   U7756 : AND2_X1 port map( A1 => n8115, A2 => n8108, ZN => n7496);
   U7757 : AND2_X1 port map( A1 => n8109, A2 => n8110, ZN => n7485);
   U7758 : AND2_X1 port map( A1 => n8107, A2 => n8110, ZN => n7486);
   U7759 : AND2_X1 port map( A1 => n8769, A2 => n8761, ZN => n8148);
   U7760 : AND2_X1 port map( A1 => n8768, A2 => n8761, ZN => n8149);
   U7761 : AND2_X1 port map( A1 => n8762, A2 => n8766, ZN => n8143);
   U7762 : AND2_X1 port map( A1 => n8760, A2 => n8766, ZN => n8144);
   U7763 : AND2_X1 port map( A1 => n8109, A2 => n8113, ZN => n7490);
   U7764 : AND2_X1 port map( A1 => n8107, A2 => n8113, ZN => n7491);
   U7765 : BUF_X1 port map( A => n7476, Z => n9499);
   U7766 : OAI21_X1 port map( B1 => n7448, B2 => n7469, A => n9887, ZN => n7476
                           );
   U7767 : INV_X1 port map( A => n7475, ZN => n9518);
   U7768 : OAI21_X1 port map( B1 => n7446, B2 => n7469, A => n9887, ZN => n7475
                           );
   U7769 : INV_X1 port map( A => n7474, ZN => n9527);
   U7770 : OAI21_X1 port map( B1 => n7444, B2 => n7469, A => n9887, ZN => n7474
                           );
   U7771 : INV_X1 port map( A => n7473, ZN => n9536);
   U7772 : OAI21_X1 port map( B1 => n7442, B2 => n7469, A => n9888, ZN => n7473
                           );
   U7773 : INV_X1 port map( A => n7472, ZN => n9545);
   U7774 : OAI21_X1 port map( B1 => n7440, B2 => n7469, A => n9888, ZN => n7472
                           );
   U7775 : INV_X1 port map( A => n7471, ZN => n9554);
   U7776 : OAI21_X1 port map( B1 => n7438, B2 => n7469, A => n9888, ZN => n7471
                           );
   U7777 : INV_X1 port map( A => n7470, ZN => n9563);
   U7778 : OAI21_X1 port map( B1 => n7436, B2 => n7469, A => n9888, ZN => n7470
                           );
   U7779 : INV_X1 port map( A => n7468, ZN => n9572);
   U7780 : OAI21_X1 port map( B1 => n7434, B2 => n7469, A => n9888, ZN => n7468
                           );
   U7781 : INV_X1 port map( A => n7467, ZN => n9581);
   U7782 : OAI21_X1 port map( B1 => n7448, B2 => n7460, A => n9888, ZN => n7467
                           );
   U7783 : INV_X1 port map( A => n7466, ZN => n9590);
   U7784 : OAI21_X1 port map( B1 => n7446, B2 => n7460, A => n9888, ZN => n7466
                           );
   U7785 : INV_X1 port map( A => n7465, ZN => n9599);
   U7786 : OAI21_X1 port map( B1 => n7444, B2 => n7460, A => n9888, ZN => n7465
                           );
   U7787 : INV_X1 port map( A => n7464, ZN => n9608);
   U7788 : OAI21_X1 port map( B1 => n7442, B2 => n7460, A => n9888, ZN => n7464
                           );
   U7789 : INV_X1 port map( A => n7463, ZN => n9617);
   U7790 : OAI21_X1 port map( B1 => n7440, B2 => n7460, A => n9888, ZN => n7463
                           );
   U7791 : INV_X1 port map( A => n7462, ZN => n9626);
   U7792 : OAI21_X1 port map( B1 => n7438, B2 => n7460, A => n9888, ZN => n7462
                           );
   U7793 : INV_X1 port map( A => n7461, ZN => n9635);
   U7794 : OAI21_X1 port map( B1 => n7436, B2 => n7460, A => n9888, ZN => n7461
                           );
   U7795 : INV_X1 port map( A => n7459, ZN => n9644);
   U7796 : OAI21_X1 port map( B1 => n7434, B2 => n7460, A => n9888, ZN => n7459
                           );
   U7797 : INV_X1 port map( A => n7458, ZN => n9653);
   U7798 : OAI21_X1 port map( B1 => n7448, B2 => n7451, A => n9889, ZN => n7458
                           );
   U7799 : INV_X1 port map( A => n7457, ZN => n9662);
   U7800 : OAI21_X1 port map( B1 => n7446, B2 => n7451, A => n9889, ZN => n7457
                           );
   U7801 : INV_X1 port map( A => n7456, ZN => n9671);
   U7802 : OAI21_X1 port map( B1 => n7444, B2 => n7451, A => n9889, ZN => n7456
                           );
   U7803 : INV_X1 port map( A => n7455, ZN => n9680);
   U7804 : OAI21_X1 port map( B1 => n7442, B2 => n7451, A => n9889, ZN => n7455
                           );
   U7805 : INV_X1 port map( A => n7454, ZN => n9689);
   U7806 : OAI21_X1 port map( B1 => n7440, B2 => n7451, A => n9889, ZN => n7454
                           );
   U7807 : INV_X1 port map( A => n7453, ZN => n9698);
   U7808 : OAI21_X1 port map( B1 => n7438, B2 => n7451, A => n9889, ZN => n7453
                           );
   U7809 : INV_X1 port map( A => n7452, ZN => n9707);
   U7810 : OAI21_X1 port map( B1 => n7436, B2 => n7451, A => n9889, ZN => n7452
                           );
   U7811 : INV_X1 port map( A => n7450, ZN => n9716);
   U7812 : OAI21_X1 port map( B1 => n7434, B2 => n7451, A => n9889, ZN => n7450
                           );
   U7813 : INV_X1 port map( A => n7447, ZN => n9725);
   U7814 : OAI21_X1 port map( B1 => n7433, B2 => n7448, A => n9889, ZN => n7447
                           );
   U7815 : INV_X1 port map( A => n7445, ZN => n9734);
   U7816 : OAI21_X1 port map( B1 => n7433, B2 => n7446, A => n9889, ZN => n7445
                           );
   U7817 : INV_X1 port map( A => n7443, ZN => n9743);
   U7818 : OAI21_X1 port map( B1 => n7433, B2 => n7444, A => n9889, ZN => n7443
                           );
   U7819 : INV_X1 port map( A => n7441, ZN => n9752);
   U7820 : OAI21_X1 port map( B1 => n7433, B2 => n7442, A => n9889, ZN => n7441
                           );
   U7821 : INV_X1 port map( A => n7439, ZN => n9761);
   U7822 : OAI21_X1 port map( B1 => n7433, B2 => n7440, A => n9889, ZN => n7439
                           );
   U7823 : INV_X1 port map( A => n7437, ZN => n9770);
   U7824 : OAI21_X1 port map( B1 => n7433, B2 => n7438, A => n9890, ZN => n7437
                           );
   U7825 : INV_X1 port map( A => n7435, ZN => n9779);
   U7826 : OAI21_X1 port map( B1 => n7433, B2 => n7436, A => n9890, ZN => n7435
                           );
   U7827 : AOI221_X1 port map( B1 => n9340, B2 => n6535, C1 => n9337, C2 => 
                           n6567, A => n8775, ZN => n8774);
   U7828 : OAI22_X1 port map( A1 => n6491, A2 => n9334, B1 => n64, B2 => n9331,
                           ZN => n8775);
   U7829 : AOI221_X1 port map( B1 => n9340, B2 => n6534, C1 => n9337, C2 => 
                           n6566, A => n8748, ZN => n8747);
   U7830 : OAI22_X1 port map( A1 => n6490, A2 => n9334, B1 => n63, B2 => n9331,
                           ZN => n8748);
   U7831 : AOI221_X1 port map( B1 => n9340, B2 => n6533, C1 => n9337, C2 => 
                           n6565, A => n8729, ZN => n8728);
   U7832 : OAI22_X1 port map( A1 => n6489, A2 => n9334, B1 => n62, B2 => n9331,
                           ZN => n8729);
   U7833 : AOI221_X1 port map( B1 => n9340, B2 => n6532, C1 => n9337, C2 => 
                           n6564, A => n8710, ZN => n8709);
   U7834 : OAI22_X1 port map( A1 => n6488, A2 => n9334, B1 => n61, B2 => n9331,
                           ZN => n8710);
   U7835 : AOI221_X1 port map( B1 => n9340, B2 => n6531, C1 => n9337, C2 => 
                           n6563, A => n8691, ZN => n8690);
   U7836 : OAI22_X1 port map( A1 => n6487, A2 => n9334, B1 => n60, B2 => n9331,
                           ZN => n8691);
   U7837 : AOI221_X1 port map( B1 => n9340, B2 => n6530, C1 => n9337, C2 => 
                           n6562, A => n8672, ZN => n8671);
   U7838 : OAI22_X1 port map( A1 => n6486, A2 => n9334, B1 => n59, B2 => n9331,
                           ZN => n8672);
   U7839 : AOI221_X1 port map( B1 => n9340, B2 => n6529, C1 => n9337, C2 => 
                           n6561, A => n8653, ZN => n8652);
   U7840 : OAI22_X1 port map( A1 => n6485, A2 => n9334, B1 => n58, B2 => n9331,
                           ZN => n8653);
   U7841 : AOI221_X1 port map( B1 => n9340, B2 => n6528, C1 => n9337, C2 => 
                           n6560, A => n8634, ZN => n8633);
   U7842 : OAI22_X1 port map( A1 => n6484, A2 => n9334, B1 => n57, B2 => n9331,
                           ZN => n8634);
   U7843 : AOI221_X1 port map( B1 => n9340, B2 => n6527, C1 => n9337, C2 => 
                           n6559, A => n8615, ZN => n8614);
   U7844 : OAI22_X1 port map( A1 => n6483, A2 => n9334, B1 => n56, B2 => n9331,
                           ZN => n8615);
   U7845 : AOI221_X1 port map( B1 => n9340, B2 => n6526, C1 => n9337, C2 => 
                           n6558, A => n8596, ZN => n8595);
   U7846 : OAI22_X1 port map( A1 => n6482, A2 => n9334, B1 => n55, B2 => n9331,
                           ZN => n8596);
   U7847 : AOI221_X1 port map( B1 => n9340, B2 => n6525, C1 => n9337, C2 => 
                           n6557, A => n8577, ZN => n8576);
   U7848 : OAI22_X1 port map( A1 => n6481, A2 => n9334, B1 => n54, B2 => n9331,
                           ZN => n8577);
   U7849 : AOI221_X1 port map( B1 => n9340, B2 => n6524, C1 => n9337, C2 => 
                           n6556, A => n8558, ZN => n8557);
   U7850 : OAI22_X1 port map( A1 => n6480, A2 => n9334, B1 => n53, B2 => n9331,
                           ZN => n8558);
   U7851 : AOI221_X1 port map( B1 => n9341, B2 => n6523, C1 => n9338, C2 => 
                           n6555, A => n8539, ZN => n8538);
   U7852 : OAI22_X1 port map( A1 => n6479, A2 => n9335, B1 => n52, B2 => n9332,
                           ZN => n8539);
   U7853 : AOI221_X1 port map( B1 => n9341, B2 => n6522, C1 => n9338, C2 => 
                           n6554, A => n8520, ZN => n8519);
   U7854 : OAI22_X1 port map( A1 => n6478, A2 => n9335, B1 => n51, B2 => n9332,
                           ZN => n8520);
   U7855 : AOI221_X1 port map( B1 => n9341, B2 => n6521, C1 => n9338, C2 => 
                           n6553, A => n8501, ZN => n8500);
   U7856 : OAI22_X1 port map( A1 => n6477, A2 => n9335, B1 => n50, B2 => n9332,
                           ZN => n8501);
   U7857 : AOI221_X1 port map( B1 => n9341, B2 => n6520, C1 => n9338, C2 => 
                           n6552, A => n8482, ZN => n8481);
   U7858 : OAI22_X1 port map( A1 => n6476, A2 => n9335, B1 => n49, B2 => n9332,
                           ZN => n8482);
   U7859 : AOI221_X1 port map( B1 => n9341, B2 => n6519, C1 => n9338, C2 => 
                           n6551, A => n8463, ZN => n8462);
   U7860 : OAI22_X1 port map( A1 => n6475, A2 => n9335, B1 => n48, B2 => n9332,
                           ZN => n8463);
   U7861 : AOI221_X1 port map( B1 => n9341, B2 => n6518, C1 => n9338, C2 => 
                           n6550, A => n8444, ZN => n8443);
   U7862 : OAI22_X1 port map( A1 => n6474, A2 => n9335, B1 => n47, B2 => n9332,
                           ZN => n8444);
   U7863 : AOI221_X1 port map( B1 => n9341, B2 => n6517, C1 => n9338, C2 => 
                           n6549, A => n8425, ZN => n8424);
   U7864 : OAI22_X1 port map( A1 => n6473, A2 => n9335, B1 => n46, B2 => n9332,
                           ZN => n8425);
   U7865 : AOI221_X1 port map( B1 => n9341, B2 => n6516, C1 => n9338, C2 => 
                           n6548, A => n8406, ZN => n8405);
   U7866 : OAI22_X1 port map( A1 => n6472, A2 => n9335, B1 => n45, B2 => n9332,
                           ZN => n8406);
   U7867 : AOI221_X1 port map( B1 => n9341, B2 => n6512, C1 => n9338, C2 => 
                           n6544, A => n8330, ZN => n8329);
   U7868 : OAI22_X1 port map( A1 => n9, A2 => n9335, B1 => n6500, B2 => n9332, 
                           ZN => n8330);
   U7869 : AOI221_X1 port map( B1 => n9342, B2 => n6511, C1 => n9339, C2 => 
                           n6543, A => n8311, ZN => n8310);
   U7870 : OAI22_X1 port map( A1 => n8, A2 => n9336, B1 => n6499, B2 => n9333, 
                           ZN => n8311);
   U7871 : AOI221_X1 port map( B1 => n9342, B2 => n6510, C1 => n9339, C2 => 
                           n6542, A => n8292, ZN => n8291);
   U7872 : OAI22_X1 port map( A1 => n7, A2 => n9336, B1 => n6498, B2 => n9333, 
                           ZN => n8292);
   U7873 : AOI221_X1 port map( B1 => n9342, B2 => n6509, C1 => n9339, C2 => 
                           n6541, A => n8273, ZN => n8272);
   U7874 : OAI22_X1 port map( A1 => n6, A2 => n9336, B1 => n6497, B2 => n9333, 
                           ZN => n8273);
   U7875 : AOI221_X1 port map( B1 => n9342, B2 => n6508, C1 => n9339, C2 => 
                           n6540, A => n8254, ZN => n8253);
   U7876 : OAI22_X1 port map( A1 => n5, A2 => n9336, B1 => n6496, B2 => n9333, 
                           ZN => n8254);
   U7877 : AOI221_X1 port map( B1 => n9442, B2 => n6535, C1 => n9439, C2 => 
                           n6567, A => n8122, ZN => n8121);
   U7878 : OAI22_X1 port map( A1 => n6491, A2 => n9436, B1 => n64, B2 => n9433,
                           ZN => n8122);
   U7879 : AOI221_X1 port map( B1 => n9442, B2 => n6534, C1 => n9439, C2 => 
                           n6566, A => n8095, ZN => n8094);
   U7880 : OAI22_X1 port map( A1 => n6490, A2 => n9436, B1 => n63, B2 => n9433,
                           ZN => n8095);
   U7881 : AOI221_X1 port map( B1 => n9442, B2 => n6533, C1 => n9439, C2 => 
                           n6565, A => n8076, ZN => n8075);
   U7882 : OAI22_X1 port map( A1 => n6489, A2 => n9436, B1 => n62, B2 => n9433,
                           ZN => n8076);
   U7883 : AOI221_X1 port map( B1 => n9442, B2 => n6532, C1 => n9439, C2 => 
                           n6564, A => n8057, ZN => n8056);
   U7884 : OAI22_X1 port map( A1 => n6488, A2 => n9436, B1 => n61, B2 => n9433,
                           ZN => n8057);
   U7885 : AOI221_X1 port map( B1 => n9442, B2 => n6531, C1 => n9439, C2 => 
                           n6563, A => n8038, ZN => n8037);
   U7886 : OAI22_X1 port map( A1 => n6487, A2 => n9436, B1 => n60, B2 => n9433,
                           ZN => n8038);
   U7887 : AOI221_X1 port map( B1 => n9442, B2 => n6530, C1 => n9439, C2 => 
                           n6562, A => n8019, ZN => n8018);
   U7888 : OAI22_X1 port map( A1 => n6486, A2 => n9436, B1 => n59, B2 => n9433,
                           ZN => n8019);
   U7889 : AOI221_X1 port map( B1 => n9442, B2 => n6529, C1 => n9439, C2 => 
                           n6561, A => n8000, ZN => n7999);
   U7890 : OAI22_X1 port map( A1 => n6485, A2 => n9436, B1 => n58, B2 => n9433,
                           ZN => n8000);
   U7891 : AOI221_X1 port map( B1 => n9442, B2 => n6528, C1 => n9439, C2 => 
                           n6560, A => n7981, ZN => n7980);
   U7892 : OAI22_X1 port map( A1 => n6484, A2 => n9436, B1 => n57, B2 => n9433,
                           ZN => n7981);
   U7893 : AOI221_X1 port map( B1 => n9442, B2 => n6527, C1 => n9439, C2 => 
                           n6559, A => n7962, ZN => n7961);
   U7894 : OAI22_X1 port map( A1 => n6483, A2 => n9436, B1 => n56, B2 => n9433,
                           ZN => n7962);
   U7895 : AOI221_X1 port map( B1 => n9442, B2 => n6526, C1 => n9439, C2 => 
                           n6558, A => n7943, ZN => n7942);
   U7896 : OAI22_X1 port map( A1 => n6482, A2 => n9436, B1 => n55, B2 => n9433,
                           ZN => n7943);
   U7897 : AOI221_X1 port map( B1 => n9442, B2 => n6525, C1 => n9439, C2 => 
                           n6557, A => n7924, ZN => n7923);
   U7898 : OAI22_X1 port map( A1 => n6481, A2 => n9436, B1 => n54, B2 => n9433,
                           ZN => n7924);
   U7899 : AOI221_X1 port map( B1 => n9442, B2 => n6524, C1 => n9439, C2 => 
                           n6556, A => n7905, ZN => n7904);
   U7900 : OAI22_X1 port map( A1 => n6480, A2 => n9436, B1 => n53, B2 => n9433,
                           ZN => n7905);
   U7901 : AOI221_X1 port map( B1 => n9443, B2 => n6523, C1 => n9440, C2 => 
                           n6555, A => n7886, ZN => n7885);
   U7902 : OAI22_X1 port map( A1 => n6479, A2 => n9437, B1 => n52, B2 => n9434,
                           ZN => n7886);
   U7903 : AOI221_X1 port map( B1 => n9443, B2 => n6522, C1 => n9440, C2 => 
                           n6554, A => n7867, ZN => n7866);
   U7904 : OAI22_X1 port map( A1 => n6478, A2 => n9437, B1 => n51, B2 => n9434,
                           ZN => n7867);
   U7905 : AOI221_X1 port map( B1 => n9443, B2 => n6521, C1 => n9440, C2 => 
                           n6553, A => n7848, ZN => n7847);
   U7906 : OAI22_X1 port map( A1 => n6477, A2 => n9437, B1 => n50, B2 => n9434,
                           ZN => n7848);
   U7907 : AOI221_X1 port map( B1 => n9443, B2 => n6520, C1 => n9440, C2 => 
                           n6552, A => n7829, ZN => n7828);
   U7908 : OAI22_X1 port map( A1 => n6476, A2 => n9437, B1 => n49, B2 => n9434,
                           ZN => n7829);
   U7909 : AOI221_X1 port map( B1 => n9443, B2 => n6519, C1 => n9440, C2 => 
                           n6551, A => n7810, ZN => n7809);
   U7910 : OAI22_X1 port map( A1 => n6475, A2 => n9437, B1 => n48, B2 => n9434,
                           ZN => n7810);
   U7911 : AOI221_X1 port map( B1 => n9443, B2 => n6518, C1 => n9440, C2 => 
                           n6550, A => n7791, ZN => n7790);
   U7912 : OAI22_X1 port map( A1 => n6474, A2 => n9437, B1 => n47, B2 => n9434,
                           ZN => n7791);
   U7913 : AOI221_X1 port map( B1 => n9443, B2 => n6517, C1 => n9440, C2 => 
                           n6549, A => n7772, ZN => n7771);
   U7914 : OAI22_X1 port map( A1 => n6473, A2 => n9437, B1 => n46, B2 => n9434,
                           ZN => n7772);
   U7915 : AOI221_X1 port map( B1 => n9443, B2 => n6516, C1 => n9440, C2 => 
                           n6548, A => n7753, ZN => n7752);
   U7916 : OAI22_X1 port map( A1 => n6472, A2 => n9437, B1 => n45, B2 => n9434,
                           ZN => n7753);
   U7917 : AOI221_X1 port map( B1 => n9443, B2 => n6512, C1 => n9440, C2 => 
                           n6544, A => n7677, ZN => n7676);
   U7918 : OAI22_X1 port map( A1 => n9, A2 => n9437, B1 => n6500, B2 => n9434, 
                           ZN => n7677);
   U7919 : AOI221_X1 port map( B1 => n9444, B2 => n6511, C1 => n9441, C2 => 
                           n6543, A => n7658, ZN => n7657);
   U7920 : OAI22_X1 port map( A1 => n8, A2 => n9438, B1 => n6499, B2 => n9435, 
                           ZN => n7658);
   U7921 : AOI221_X1 port map( B1 => n9444, B2 => n6510, C1 => n9441, C2 => 
                           n6542, A => n7639, ZN => n7638);
   U7922 : OAI22_X1 port map( A1 => n7, A2 => n9438, B1 => n6498, B2 => n9435, 
                           ZN => n7639);
   U7923 : AOI221_X1 port map( B1 => n9444, B2 => n6509, C1 => n9441, C2 => 
                           n6541, A => n7620, ZN => n7619);
   U7924 : OAI22_X1 port map( A1 => n6, A2 => n9438, B1 => n6497, B2 => n9435, 
                           ZN => n7620);
   U7925 : AOI221_X1 port map( B1 => n9444, B2 => n6508, C1 => n9441, C2 => 
                           n6540, A => n7601, ZN => n7600);
   U7926 : OAI22_X1 port map( A1 => n5, A2 => n9438, B1 => n6496, B2 => n9435, 
                           ZN => n7601);
   U7927 : AOI221_X1 port map( B1 => n9328, B2 => n4509, C1 => n9325, C2 => 
                           n4445, A => n8778, ZN => n8773);
   U7928 : OAI22_X1 port map( A1 => n9284, A2 => n9322, B1 => n9283, B2 => 
                           n9319, ZN => n8778);
   U7929 : AOI221_X1 port map( B1 => n9328, B2 => n4508, C1 => n9325, C2 => 
                           n4444, A => n8749, ZN => n8746);
   U7930 : OAI22_X1 port map( A1 => n9269, A2 => n9322, B1 => n9268, B2 => 
                           n9319, ZN => n8749);
   U7931 : AOI221_X1 port map( B1 => n9328, B2 => n4507, C1 => n9325, C2 => 
                           n4443, A => n8730, ZN => n8727);
   U7932 : OAI22_X1 port map( A1 => n9254, A2 => n9322, B1 => n9253, B2 => 
                           n9319, ZN => n8730);
   U7933 : AOI221_X1 port map( B1 => n9328, B2 => n4506, C1 => n9325, C2 => 
                           n4442, A => n8711, ZN => n8708);
   U7934 : OAI22_X1 port map( A1 => n9239, A2 => n9322, B1 => n9238, B2 => 
                           n9319, ZN => n8711);
   U7935 : AOI221_X1 port map( B1 => n9328, B2 => n4505, C1 => n9325, C2 => 
                           n4441, A => n8692, ZN => n8689);
   U7936 : OAI22_X1 port map( A1 => n9224, A2 => n9322, B1 => n9223, B2 => 
                           n9319, ZN => n8692);
   U7937 : AOI221_X1 port map( B1 => n9328, B2 => n4504, C1 => n9325, C2 => 
                           n4440, A => n8673, ZN => n8670);
   U7938 : OAI22_X1 port map( A1 => n9209, A2 => n9322, B1 => n9208, B2 => 
                           n9319, ZN => n8673);
   U7939 : AOI221_X1 port map( B1 => n9328, B2 => n4503, C1 => n9325, C2 => 
                           n4439, A => n8654, ZN => n8651);
   U7940 : OAI22_X1 port map( A1 => n9194, A2 => n9322, B1 => n9193, B2 => 
                           n9319, ZN => n8654);
   U7941 : AOI221_X1 port map( B1 => n9328, B2 => n4502, C1 => n9325, C2 => 
                           n4438, A => n8635, ZN => n8632);
   U7942 : OAI22_X1 port map( A1 => n9179, A2 => n9322, B1 => n9178, B2 => 
                           n9319, ZN => n8635);
   U7943 : AOI221_X1 port map( B1 => n9328, B2 => n4501, C1 => n9325, C2 => 
                           n4437, A => n8616, ZN => n8613);
   U7944 : OAI22_X1 port map( A1 => n9164, A2 => n9322, B1 => n9163, B2 => 
                           n9319, ZN => n8616);
   U7945 : AOI221_X1 port map( B1 => n9328, B2 => n4500, C1 => n9325, C2 => 
                           n4436, A => n8597, ZN => n8594);
   U7946 : OAI22_X1 port map( A1 => n9149, A2 => n9322, B1 => n9148, B2 => 
                           n9319, ZN => n8597);
   U7947 : AOI221_X1 port map( B1 => n9328, B2 => n4499, C1 => n9325, C2 => 
                           n4435, A => n8578, ZN => n8575);
   U7948 : OAI22_X1 port map( A1 => n9134, A2 => n9322, B1 => n9133, B2 => 
                           n9319, ZN => n8578);
   U7949 : AOI221_X1 port map( B1 => n9328, B2 => n4498, C1 => n9325, C2 => 
                           n4434, A => n8559, ZN => n8556);
   U7950 : OAI22_X1 port map( A1 => n9119, A2 => n9322, B1 => n9118, B2 => 
                           n9319, ZN => n8559);
   U7951 : AOI221_X1 port map( B1 => n9329, B2 => n4497, C1 => n9326, C2 => 
                           n4433, A => n8540, ZN => n8537);
   U7952 : OAI22_X1 port map( A1 => n9104, A2 => n9323, B1 => n9103, B2 => 
                           n9320, ZN => n8540);
   U7953 : AOI221_X1 port map( B1 => n9329, B2 => n4496, C1 => n9326, C2 => 
                           n4432, A => n8521, ZN => n8518);
   U7954 : OAI22_X1 port map( A1 => n9089, A2 => n9323, B1 => n9088, B2 => 
                           n9320, ZN => n8521);
   U7955 : AOI221_X1 port map( B1 => n9329, B2 => n4495, C1 => n9326, C2 => 
                           n4431, A => n8502, ZN => n8499);
   U7956 : OAI22_X1 port map( A1 => n9074, A2 => n9323, B1 => n9073, B2 => 
                           n9320, ZN => n8502);
   U7957 : AOI221_X1 port map( B1 => n9329, B2 => n4494, C1 => n9326, C2 => 
                           n4430, A => n8483, ZN => n8480);
   U7958 : OAI22_X1 port map( A1 => n9059, A2 => n9323, B1 => n9058, B2 => 
                           n9320, ZN => n8483);
   U7959 : AOI221_X1 port map( B1 => n9329, B2 => n4493, C1 => n9326, C2 => 
                           n4429, A => n8464, ZN => n8461);
   U7960 : OAI22_X1 port map( A1 => n9044, A2 => n9323, B1 => n9043, B2 => 
                           n9320, ZN => n8464);
   U7961 : AOI221_X1 port map( B1 => n9329, B2 => n4492, C1 => n9326, C2 => 
                           n4428, A => n8445, ZN => n8442);
   U7962 : OAI22_X1 port map( A1 => n9029, A2 => n9323, B1 => n9028, B2 => 
                           n9320, ZN => n8445);
   U7963 : AOI221_X1 port map( B1 => n9329, B2 => n4491, C1 => n9326, C2 => 
                           n4427, A => n8426, ZN => n8423);
   U7964 : OAI22_X1 port map( A1 => n9014, A2 => n9323, B1 => n9013, B2 => 
                           n9320, ZN => n8426);
   U7965 : AOI221_X1 port map( B1 => n9329, B2 => n4490, C1 => n9326, C2 => 
                           n4426, A => n8407, ZN => n8404);
   U7966 : OAI22_X1 port map( A1 => n8999, A2 => n9323, B1 => n8998, B2 => 
                           n9320, ZN => n8407);
   U7967 : AOI221_X1 port map( B1 => n9329, B2 => n4489, C1 => n9326, C2 => 
                           n4425, A => n8388, ZN => n8385);
   U7968 : OAI22_X1 port map( A1 => n8984, A2 => n9323, B1 => n8983, B2 => 
                           n9320, ZN => n8388);
   U7969 : AOI221_X1 port map( B1 => n9329, B2 => n4488, C1 => n9326, C2 => 
                           n4424, A => n8369, ZN => n8366);
   U7970 : OAI22_X1 port map( A1 => n8969, A2 => n9323, B1 => n8968, B2 => 
                           n9320, ZN => n8369);
   U7971 : AOI221_X1 port map( B1 => n9329, B2 => n4487, C1 => n9326, C2 => 
                           n4423, A => n8350, ZN => n8347);
   U7972 : OAI22_X1 port map( A1 => n8954, A2 => n9323, B1 => n8953, B2 => 
                           n9320, ZN => n8350);
   U7973 : AOI221_X1 port map( B1 => n9329, B2 => n4486, C1 => n9326, C2 => 
                           n4422, A => n8331, ZN => n8328);
   U7974 : OAI22_X1 port map( A1 => n8939, A2 => n9323, B1 => n8938, B2 => 
                           n9320, ZN => n8331);
   U7975 : AOI221_X1 port map( B1 => n9330, B2 => n4485, C1 => n9327, C2 => 
                           n4421, A => n8312, ZN => n8309);
   U7976 : OAI22_X1 port map( A1 => n8924, A2 => n9324, B1 => n8923, B2 => 
                           n9321, ZN => n8312);
   U7977 : AOI221_X1 port map( B1 => n9330, B2 => n4484, C1 => n9327, C2 => 
                           n4420, A => n8293, ZN => n8290);
   U7978 : OAI22_X1 port map( A1 => n8909, A2 => n9324, B1 => n8908, B2 => 
                           n9321, ZN => n8293);
   U7979 : AOI221_X1 port map( B1 => n9330, B2 => n4483, C1 => n9327, C2 => 
                           n4419, A => n8274, ZN => n8271);
   U7980 : OAI22_X1 port map( A1 => n8894, A2 => n9324, B1 => n8893, B2 => 
                           n9321, ZN => n8274);
   U7981 : AOI221_X1 port map( B1 => n9330, B2 => n4482, C1 => n9327, C2 => 
                           n4418, A => n8255, ZN => n8252);
   U7982 : OAI22_X1 port map( A1 => n8879, A2 => n9324, B1 => n8878, B2 => 
                           n9321, ZN => n8255);
   U7983 : AOI221_X1 port map( B1 => n9330, B2 => n4481, C1 => n9327, C2 => 
                           n4417, A => n8236, ZN => n8233);
   U7984 : OAI22_X1 port map( A1 => n8864, A2 => n9324, B1 => n8863, B2 => 
                           n9321, ZN => n8236);
   U7985 : AOI221_X1 port map( B1 => n9330, B2 => n4480, C1 => n9327, C2 => 
                           n4416, A => n8217, ZN => n8214);
   U7986 : OAI22_X1 port map( A1 => n8849, A2 => n9324, B1 => n8848, B2 => 
                           n9321, ZN => n8217);
   U7987 : AOI221_X1 port map( B1 => n9330, B2 => n4479, C1 => n9327, C2 => 
                           n4415, A => n8198, ZN => n8195);
   U7988 : OAI22_X1 port map( A1 => n8834, A2 => n9324, B1 => n8833, B2 => 
                           n9321, ZN => n8198);
   U7989 : AOI221_X1 port map( B1 => n9330, B2 => n4478, C1 => n9327, C2 => 
                           n4414, A => n8169, ZN => n8160);
   U7990 : OAI22_X1 port map( A1 => n8819, A2 => n9324, B1 => n8818, B2 => 
                           n9321, ZN => n8169);
   U7991 : AOI221_X1 port map( B1 => n9430, B2 => n4509, C1 => n9427, C2 => 
                           n4445, A => n8125, ZN => n8120);
   U7992 : OAI22_X1 port map( A1 => n9284, A2 => n9424, B1 => n9283, B2 => 
                           n9421, ZN => n8125);
   U7993 : AOI221_X1 port map( B1 => n9430, B2 => n4508, C1 => n9427, C2 => 
                           n4444, A => n8096, ZN => n8093);
   U7994 : OAI22_X1 port map( A1 => n9269, A2 => n9424, B1 => n9268, B2 => 
                           n9421, ZN => n8096);
   U7995 : AOI221_X1 port map( B1 => n9430, B2 => n4507, C1 => n9427, C2 => 
                           n4443, A => n8077, ZN => n8074);
   U7996 : OAI22_X1 port map( A1 => n9254, A2 => n9424, B1 => n9253, B2 => 
                           n9421, ZN => n8077);
   U7997 : AOI221_X1 port map( B1 => n9430, B2 => n4506, C1 => n9427, C2 => 
                           n4442, A => n8058, ZN => n8055);
   U7998 : OAI22_X1 port map( A1 => n9239, A2 => n9424, B1 => n9238, B2 => 
                           n9421, ZN => n8058);
   U7999 : AOI221_X1 port map( B1 => n9430, B2 => n4505, C1 => n9427, C2 => 
                           n4441, A => n8039, ZN => n8036);
   U8000 : OAI22_X1 port map( A1 => n9224, A2 => n9424, B1 => n9223, B2 => 
                           n9421, ZN => n8039);
   U8001 : AOI221_X1 port map( B1 => n9430, B2 => n4504, C1 => n9427, C2 => 
                           n4440, A => n8020, ZN => n8017);
   U8002 : OAI22_X1 port map( A1 => n9209, A2 => n9424, B1 => n9208, B2 => 
                           n9421, ZN => n8020);
   U8003 : AOI221_X1 port map( B1 => n9430, B2 => n4503, C1 => n9427, C2 => 
                           n4439, A => n8001, ZN => n7998);
   U8004 : OAI22_X1 port map( A1 => n9194, A2 => n9424, B1 => n9193, B2 => 
                           n9421, ZN => n8001);
   U8005 : AOI221_X1 port map( B1 => n9430, B2 => n4502, C1 => n9427, C2 => 
                           n4438, A => n7982, ZN => n7979);
   U8006 : OAI22_X1 port map( A1 => n9179, A2 => n9424, B1 => n9178, B2 => 
                           n9421, ZN => n7982);
   U8007 : AOI221_X1 port map( B1 => n9430, B2 => n4501, C1 => n9427, C2 => 
                           n4437, A => n7963, ZN => n7960);
   U8008 : OAI22_X1 port map( A1 => n9164, A2 => n9424, B1 => n9163, B2 => 
                           n9421, ZN => n7963);
   U8009 : AOI221_X1 port map( B1 => n9430, B2 => n4500, C1 => n9427, C2 => 
                           n4436, A => n7944, ZN => n7941);
   U8010 : OAI22_X1 port map( A1 => n9149, A2 => n9424, B1 => n9148, B2 => 
                           n9421, ZN => n7944);
   U8011 : AOI221_X1 port map( B1 => n9430, B2 => n4499, C1 => n9427, C2 => 
                           n4435, A => n7925, ZN => n7922);
   U8012 : OAI22_X1 port map( A1 => n9134, A2 => n9424, B1 => n9133, B2 => 
                           n9421, ZN => n7925);
   U8013 : AOI221_X1 port map( B1 => n9430, B2 => n4498, C1 => n9427, C2 => 
                           n4434, A => n7906, ZN => n7903);
   U8014 : OAI22_X1 port map( A1 => n9119, A2 => n9424, B1 => n9118, B2 => 
                           n9421, ZN => n7906);
   U8015 : AOI221_X1 port map( B1 => n9431, B2 => n4497, C1 => n9428, C2 => 
                           n4433, A => n7887, ZN => n7884);
   U8016 : OAI22_X1 port map( A1 => n9104, A2 => n9425, B1 => n9103, B2 => 
                           n9422, ZN => n7887);
   U8017 : AOI221_X1 port map( B1 => n9431, B2 => n4496, C1 => n9428, C2 => 
                           n4432, A => n7868, ZN => n7865);
   U8018 : OAI22_X1 port map( A1 => n9089, A2 => n9425, B1 => n9088, B2 => 
                           n9422, ZN => n7868);
   U8019 : AOI221_X1 port map( B1 => n9431, B2 => n4495, C1 => n9428, C2 => 
                           n4431, A => n7849, ZN => n7846);
   U8020 : OAI22_X1 port map( A1 => n9074, A2 => n9425, B1 => n9073, B2 => 
                           n9422, ZN => n7849);
   U8021 : AOI221_X1 port map( B1 => n9431, B2 => n4494, C1 => n9428, C2 => 
                           n4430, A => n7830, ZN => n7827);
   U8022 : OAI22_X1 port map( A1 => n9059, A2 => n9425, B1 => n9058, B2 => 
                           n9422, ZN => n7830);
   U8023 : AOI221_X1 port map( B1 => n9431, B2 => n4493, C1 => n9428, C2 => 
                           n4429, A => n7811, ZN => n7808);
   U8024 : OAI22_X1 port map( A1 => n9044, A2 => n9425, B1 => n9043, B2 => 
                           n9422, ZN => n7811);
   U8025 : AOI221_X1 port map( B1 => n9431, B2 => n4492, C1 => n9428, C2 => 
                           n4428, A => n7792, ZN => n7789);
   U8026 : OAI22_X1 port map( A1 => n9029, A2 => n9425, B1 => n9028, B2 => 
                           n9422, ZN => n7792);
   U8027 : AOI221_X1 port map( B1 => n9431, B2 => n4491, C1 => n9428, C2 => 
                           n4427, A => n7773, ZN => n7770);
   U8028 : OAI22_X1 port map( A1 => n9014, A2 => n9425, B1 => n9013, B2 => 
                           n9422, ZN => n7773);
   U8029 : AOI221_X1 port map( B1 => n9431, B2 => n4490, C1 => n9428, C2 => 
                           n4426, A => n7754, ZN => n7751);
   U8030 : OAI22_X1 port map( A1 => n8999, A2 => n9425, B1 => n8998, B2 => 
                           n9422, ZN => n7754);
   U8031 : AOI221_X1 port map( B1 => n9431, B2 => n4489, C1 => n9428, C2 => 
                           n4425, A => n7735, ZN => n7732);
   U8032 : OAI22_X1 port map( A1 => n8984, A2 => n9425, B1 => n8983, B2 => 
                           n9422, ZN => n7735);
   U8033 : AOI221_X1 port map( B1 => n9431, B2 => n4488, C1 => n9428, C2 => 
                           n4424, A => n7716, ZN => n7713);
   U8034 : OAI22_X1 port map( A1 => n8969, A2 => n9425, B1 => n8968, B2 => 
                           n9422, ZN => n7716);
   U8035 : AOI221_X1 port map( B1 => n9431, B2 => n4487, C1 => n9428, C2 => 
                           n4423, A => n7697, ZN => n7694);
   U8036 : OAI22_X1 port map( A1 => n8954, A2 => n9425, B1 => n8953, B2 => 
                           n9422, ZN => n7697);
   U8037 : AOI221_X1 port map( B1 => n9431, B2 => n4486, C1 => n9428, C2 => 
                           n4422, A => n7678, ZN => n7675);
   U8038 : OAI22_X1 port map( A1 => n8939, A2 => n9425, B1 => n8938, B2 => 
                           n9422, ZN => n7678);
   U8039 : AOI221_X1 port map( B1 => n9432, B2 => n4485, C1 => n9429, C2 => 
                           n4421, A => n7659, ZN => n7656);
   U8040 : OAI22_X1 port map( A1 => n8924, A2 => n9426, B1 => n8923, B2 => 
                           n9423, ZN => n7659);
   U8041 : AOI221_X1 port map( B1 => n9432, B2 => n4484, C1 => n9429, C2 => 
                           n4420, A => n7640, ZN => n7637);
   U8042 : OAI22_X1 port map( A1 => n8909, A2 => n9426, B1 => n8908, B2 => 
                           n9423, ZN => n7640);
   U8043 : AOI221_X1 port map( B1 => n9432, B2 => n4483, C1 => n9429, C2 => 
                           n4419, A => n7621, ZN => n7618);
   U8044 : OAI22_X1 port map( A1 => n8894, A2 => n9426, B1 => n8893, B2 => 
                           n9423, ZN => n7621);
   U8045 : AOI221_X1 port map( B1 => n9432, B2 => n4482, C1 => n9429, C2 => 
                           n4418, A => n7602, ZN => n7599);
   U8046 : OAI22_X1 port map( A1 => n8879, A2 => n9426, B1 => n8878, B2 => 
                           n9423, ZN => n7602);
   U8047 : AOI221_X1 port map( B1 => n9432, B2 => n4481, C1 => n9429, C2 => 
                           n4417, A => n7583, ZN => n7580);
   U8048 : OAI22_X1 port map( A1 => n8864, A2 => n9426, B1 => n8863, B2 => 
                           n9423, ZN => n7583);
   U8049 : AOI221_X1 port map( B1 => n9432, B2 => n4480, C1 => n9429, C2 => 
                           n4416, A => n7564, ZN => n7561);
   U8050 : OAI22_X1 port map( A1 => n8849, A2 => n9426, B1 => n8848, B2 => 
                           n9423, ZN => n7564);
   U8051 : AOI221_X1 port map( B1 => n9432, B2 => n4479, C1 => n9429, C2 => 
                           n4415, A => n7545, ZN => n7542);
   U8052 : OAI22_X1 port map( A1 => n8834, A2 => n9426, B1 => n8833, B2 => 
                           n9423, ZN => n7545);
   U8053 : AOI221_X1 port map( B1 => n9432, B2 => n4478, C1 => n9429, C2 => 
                           n4414, A => n7516, ZN => n7507);
   U8054 : OAI22_X1 port map( A1 => n8819, A2 => n9426, B1 => n8818, B2 => 
                           n9423, ZN => n7516);
   U8055 : AOI221_X1 port map( B1 => n9316, B2 => n4381, C1 => n9313, C2 => 
                           n3997, A => n8779, ZN => n8772);
   U8056 : OAI22_X1 port map( A1 => n6695, A2 => n9310, B1 => n6663, B2 => 
                           n9307, ZN => n8779);
   U8057 : AOI221_X1 port map( B1 => n9316, B2 => n4380, C1 => n9313, C2 => 
                           n3996, A => n8750, ZN => n8745);
   U8058 : OAI22_X1 port map( A1 => n6694, A2 => n9310, B1 => n6662, B2 => 
                           n9307, ZN => n8750);
   U8059 : AOI221_X1 port map( B1 => n9316, B2 => n4379, C1 => n9313, C2 => 
                           n3995, A => n8731, ZN => n8726);
   U8060 : OAI22_X1 port map( A1 => n6693, A2 => n9310, B1 => n6661, B2 => 
                           n9307, ZN => n8731);
   U8061 : AOI221_X1 port map( B1 => n9316, B2 => n4378, C1 => n9313, C2 => 
                           n3994, A => n8712, ZN => n8707);
   U8062 : OAI22_X1 port map( A1 => n6692, A2 => n9310, B1 => n6660, B2 => 
                           n9307, ZN => n8712);
   U8063 : AOI221_X1 port map( B1 => n9316, B2 => n4377, C1 => n9313, C2 => 
                           n3993, A => n8693, ZN => n8688);
   U8064 : OAI22_X1 port map( A1 => n6691, A2 => n9310, B1 => n6659, B2 => 
                           n9307, ZN => n8693);
   U8065 : AOI221_X1 port map( B1 => n9316, B2 => n4376, C1 => n9313, C2 => 
                           n3992, A => n8674, ZN => n8669);
   U8066 : OAI22_X1 port map( A1 => n6690, A2 => n9310, B1 => n6658, B2 => 
                           n9307, ZN => n8674);
   U8067 : AOI221_X1 port map( B1 => n9316, B2 => n4375, C1 => n9313, C2 => 
                           n3991, A => n8655, ZN => n8650);
   U8068 : OAI22_X1 port map( A1 => n6689, A2 => n9310, B1 => n6657, B2 => 
                           n9307, ZN => n8655);
   U8069 : AOI221_X1 port map( B1 => n9316, B2 => n4374, C1 => n9313, C2 => 
                           n3990, A => n8636, ZN => n8631);
   U8070 : OAI22_X1 port map( A1 => n6688, A2 => n9310, B1 => n6656, B2 => 
                           n9307, ZN => n8636);
   U8071 : AOI221_X1 port map( B1 => n9316, B2 => n4373, C1 => n9313, C2 => 
                           n3989, A => n8617, ZN => n8612);
   U8072 : OAI22_X1 port map( A1 => n6687, A2 => n9310, B1 => n6655, B2 => 
                           n9307, ZN => n8617);
   U8073 : AOI221_X1 port map( B1 => n9316, B2 => n4372, C1 => n9313, C2 => 
                           n3988, A => n8598, ZN => n8593);
   U8074 : OAI22_X1 port map( A1 => n6686, A2 => n9310, B1 => n6654, B2 => 
                           n9307, ZN => n8598);
   U8075 : AOI221_X1 port map( B1 => n9316, B2 => n4371, C1 => n9313, C2 => 
                           n3987, A => n8579, ZN => n8574);
   U8076 : OAI22_X1 port map( A1 => n6685, A2 => n9310, B1 => n6653, B2 => 
                           n9307, ZN => n8579);
   U8077 : AOI221_X1 port map( B1 => n9316, B2 => n4370, C1 => n9313, C2 => 
                           n3986, A => n8560, ZN => n8555);
   U8078 : OAI22_X1 port map( A1 => n6684, A2 => n9310, B1 => n6652, B2 => 
                           n9307, ZN => n8560);
   U8079 : AOI221_X1 port map( B1 => n9317, B2 => n4369, C1 => n9314, C2 => 
                           n3985, A => n8541, ZN => n8536);
   U8080 : OAI22_X1 port map( A1 => n6683, A2 => n9311, B1 => n6651, B2 => 
                           n9308, ZN => n8541);
   U8081 : AOI221_X1 port map( B1 => n9317, B2 => n4368, C1 => n9314, C2 => 
                           n3984, A => n8522, ZN => n8517);
   U8082 : OAI22_X1 port map( A1 => n6682, A2 => n9311, B1 => n6650, B2 => 
                           n9308, ZN => n8522);
   U8083 : AOI221_X1 port map( B1 => n9317, B2 => n4367, C1 => n9314, C2 => 
                           n3983, A => n8503, ZN => n8498);
   U8084 : OAI22_X1 port map( A1 => n6681, A2 => n9311, B1 => n6649, B2 => 
                           n9308, ZN => n8503);
   U8085 : AOI221_X1 port map( B1 => n9317, B2 => n4366, C1 => n9314, C2 => 
                           n3982, A => n8484, ZN => n8479);
   U8086 : OAI22_X1 port map( A1 => n6680, A2 => n9311, B1 => n6648, B2 => 
                           n9308, ZN => n8484);
   U8087 : AOI221_X1 port map( B1 => n9317, B2 => n4365, C1 => n9314, C2 => 
                           n3981, A => n8465, ZN => n8460);
   U8088 : OAI22_X1 port map( A1 => n6679, A2 => n9311, B1 => n6647, B2 => 
                           n9308, ZN => n8465);
   U8089 : AOI221_X1 port map( B1 => n9317, B2 => n4364, C1 => n9314, C2 => 
                           n3980, A => n8446, ZN => n8441);
   U8090 : OAI22_X1 port map( A1 => n6678, A2 => n9311, B1 => n6646, B2 => 
                           n9308, ZN => n8446);
   U8091 : AOI221_X1 port map( B1 => n9317, B2 => n4363, C1 => n9314, C2 => 
                           n3979, A => n8427, ZN => n8422);
   U8092 : OAI22_X1 port map( A1 => n6677, A2 => n9311, B1 => n6645, B2 => 
                           n9308, ZN => n8427);
   U8093 : AOI221_X1 port map( B1 => n9317, B2 => n4362, C1 => n9314, C2 => 
                           n3978, A => n8408, ZN => n8403);
   U8094 : OAI22_X1 port map( A1 => n6676, A2 => n9311, B1 => n6644, B2 => 
                           n9308, ZN => n8408);
   U8095 : AOI221_X1 port map( B1 => n9317, B2 => n4361, C1 => n9314, C2 => 
                           n3977, A => n8389, ZN => n8384);
   U8096 : OAI22_X1 port map( A1 => n6675, A2 => n9311, B1 => n6643, B2 => 
                           n9308, ZN => n8389);
   U8097 : AOI221_X1 port map( B1 => n9317, B2 => n4360, C1 => n9314, C2 => 
                           n3976, A => n8370, ZN => n8365);
   U8098 : OAI22_X1 port map( A1 => n6674, A2 => n9311, B1 => n6642, B2 => 
                           n9308, ZN => n8370);
   U8099 : AOI221_X1 port map( B1 => n9317, B2 => n4359, C1 => n9314, C2 => 
                           n3975, A => n8351, ZN => n8346);
   U8100 : OAI22_X1 port map( A1 => n6673, A2 => n9311, B1 => n6641, B2 => 
                           n9308, ZN => n8351);
   U8101 : AOI221_X1 port map( B1 => n9317, B2 => n4358, C1 => n9314, C2 => 
                           n3974, A => n8332, ZN => n8327);
   U8102 : OAI22_X1 port map( A1 => n6672, A2 => n9311, B1 => n6640, B2 => 
                           n9308, ZN => n8332);
   U8103 : AOI221_X1 port map( B1 => n9318, B2 => n4357, C1 => n9315, C2 => 
                           n3973, A => n8313, ZN => n8308);
   U8104 : OAI22_X1 port map( A1 => n6671, A2 => n9312, B1 => n6639, B2 => 
                           n9309, ZN => n8313);
   U8105 : AOI221_X1 port map( B1 => n9318, B2 => n4356, C1 => n9315, C2 => 
                           n3972, A => n8294, ZN => n8289);
   U8106 : OAI22_X1 port map( A1 => n6670, A2 => n9312, B1 => n6638, B2 => 
                           n9309, ZN => n8294);
   U8107 : AOI221_X1 port map( B1 => n9318, B2 => n4355, C1 => n9315, C2 => 
                           n3971, A => n8275, ZN => n8270);
   U8108 : OAI22_X1 port map( A1 => n6669, A2 => n9312, B1 => n6637, B2 => 
                           n9309, ZN => n8275);
   U8109 : AOI221_X1 port map( B1 => n9318, B2 => n4354, C1 => n9315, C2 => 
                           n3970, A => n8256, ZN => n8251);
   U8110 : OAI22_X1 port map( A1 => n6668, A2 => n9312, B1 => n6636, B2 => 
                           n9309, ZN => n8256);
   U8111 : AOI221_X1 port map( B1 => n9318, B2 => n4353, C1 => n9315, C2 => 
                           n3969, A => n8237, ZN => n8232);
   U8112 : OAI22_X1 port map( A1 => n6667, A2 => n9312, B1 => n6635, B2 => 
                           n9309, ZN => n8237);
   U8113 : AOI221_X1 port map( B1 => n9318, B2 => n4352, C1 => n9315, C2 => 
                           n3968, A => n8218, ZN => n8213);
   U8114 : OAI22_X1 port map( A1 => n6666, A2 => n9312, B1 => n6634, B2 => 
                           n9309, ZN => n8218);
   U8115 : AOI221_X1 port map( B1 => n9318, B2 => n4351, C1 => n9315, C2 => 
                           n3967, A => n8199, ZN => n8194);
   U8116 : OAI22_X1 port map( A1 => n6665, A2 => n9312, B1 => n6633, B2 => 
                           n9309, ZN => n8199);
   U8117 : AOI221_X1 port map( B1 => n9318, B2 => n4350, C1 => n9315, C2 => 
                           n3966, A => n8174, ZN => n8159);
   U8118 : OAI22_X1 port map( A1 => n6664, A2 => n9312, B1 => n6632, B2 => 
                           n9309, ZN => n8174);
   U8119 : AOI221_X1 port map( B1 => n9418, B2 => n4349, C1 => n9415, C2 => 
                           n3965, A => n8126, ZN => n8119);
   U8120 : OAI22_X1 port map( A1 => n6759, A2 => n9412, B1 => n6727, B2 => 
                           n9409, ZN => n8126);
   U8121 : AOI221_X1 port map( B1 => n9418, B2 => n4348, C1 => n9415, C2 => 
                           n3964, A => n8097, ZN => n8092);
   U8122 : OAI22_X1 port map( A1 => n6758, A2 => n9412, B1 => n6726, B2 => 
                           n9409, ZN => n8097);
   U8123 : AOI221_X1 port map( B1 => n9418, B2 => n4347, C1 => n9415, C2 => 
                           n3963, A => n8078, ZN => n8073);
   U8124 : OAI22_X1 port map( A1 => n6757, A2 => n9412, B1 => n6725, B2 => 
                           n9409, ZN => n8078);
   U8125 : AOI221_X1 port map( B1 => n9418, B2 => n4346, C1 => n9415, C2 => 
                           n3962, A => n8059, ZN => n8054);
   U8126 : OAI22_X1 port map( A1 => n6756, A2 => n9412, B1 => n6724, B2 => 
                           n9409, ZN => n8059);
   U8127 : AOI221_X1 port map( B1 => n9418, B2 => n4345, C1 => n9415, C2 => 
                           n3961, A => n8040, ZN => n8035);
   U8128 : OAI22_X1 port map( A1 => n6755, A2 => n9412, B1 => n6723, B2 => 
                           n9409, ZN => n8040);
   U8129 : AOI221_X1 port map( B1 => n9418, B2 => n4344, C1 => n9415, C2 => 
                           n3960, A => n8021, ZN => n8016);
   U8130 : OAI22_X1 port map( A1 => n6754, A2 => n9412, B1 => n6722, B2 => 
                           n9409, ZN => n8021);
   U8131 : AOI221_X1 port map( B1 => n9418, B2 => n4343, C1 => n9415, C2 => 
                           n3959, A => n8002, ZN => n7997);
   U8132 : OAI22_X1 port map( A1 => n6753, A2 => n9412, B1 => n6721, B2 => 
                           n9409, ZN => n8002);
   U8133 : AOI221_X1 port map( B1 => n9418, B2 => n4342, C1 => n9415, C2 => 
                           n3958, A => n7983, ZN => n7978);
   U8134 : OAI22_X1 port map( A1 => n6752, A2 => n9412, B1 => n6720, B2 => 
                           n9409, ZN => n7983);
   U8135 : AOI221_X1 port map( B1 => n9418, B2 => n4341, C1 => n9415, C2 => 
                           n3957, A => n7964, ZN => n7959);
   U8136 : OAI22_X1 port map( A1 => n6751, A2 => n9412, B1 => n6719, B2 => 
                           n9409, ZN => n7964);
   U8137 : AOI221_X1 port map( B1 => n9418, B2 => n4340, C1 => n9415, C2 => 
                           n3956, A => n7945, ZN => n7940);
   U8138 : OAI22_X1 port map( A1 => n6750, A2 => n9412, B1 => n6718, B2 => 
                           n9409, ZN => n7945);
   U8139 : AOI221_X1 port map( B1 => n9418, B2 => n4339, C1 => n9415, C2 => 
                           n3955, A => n7926, ZN => n7921);
   U8140 : OAI22_X1 port map( A1 => n6749, A2 => n9412, B1 => n6717, B2 => 
                           n9409, ZN => n7926);
   U8141 : AOI221_X1 port map( B1 => n9418, B2 => n4338, C1 => n9415, C2 => 
                           n3954, A => n7907, ZN => n7902);
   U8142 : OAI22_X1 port map( A1 => n6748, A2 => n9412, B1 => n6716, B2 => 
                           n9409, ZN => n7907);
   U8143 : AOI221_X1 port map( B1 => n9419, B2 => n4337, C1 => n9416, C2 => 
                           n3953, A => n7888, ZN => n7883);
   U8144 : OAI22_X1 port map( A1 => n6747, A2 => n9413, B1 => n6715, B2 => 
                           n9410, ZN => n7888);
   U8145 : AOI221_X1 port map( B1 => n9419, B2 => n4336, C1 => n9416, C2 => 
                           n3952, A => n7869, ZN => n7864);
   U8146 : OAI22_X1 port map( A1 => n6746, A2 => n9413, B1 => n6714, B2 => 
                           n9410, ZN => n7869);
   U8147 : AOI221_X1 port map( B1 => n9419, B2 => n4335, C1 => n9416, C2 => 
                           n3951, A => n7850, ZN => n7845);
   U8148 : OAI22_X1 port map( A1 => n6745, A2 => n9413, B1 => n6713, B2 => 
                           n9410, ZN => n7850);
   U8149 : AOI221_X1 port map( B1 => n9419, B2 => n4334, C1 => n9416, C2 => 
                           n3950, A => n7831, ZN => n7826);
   U8150 : OAI22_X1 port map( A1 => n6744, A2 => n9413, B1 => n6712, B2 => 
                           n9410, ZN => n7831);
   U8151 : AOI221_X1 port map( B1 => n9419, B2 => n4333, C1 => n9416, C2 => 
                           n3949, A => n7812, ZN => n7807);
   U8152 : OAI22_X1 port map( A1 => n6743, A2 => n9413, B1 => n6711, B2 => 
                           n9410, ZN => n7812);
   U8153 : AOI221_X1 port map( B1 => n9419, B2 => n4332, C1 => n9416, C2 => 
                           n3948, A => n7793, ZN => n7788);
   U8154 : OAI22_X1 port map( A1 => n6742, A2 => n9413, B1 => n6710, B2 => 
                           n9410, ZN => n7793);
   U8155 : AOI221_X1 port map( B1 => n9419, B2 => n4331, C1 => n9416, C2 => 
                           n3947, A => n7774, ZN => n7769);
   U8156 : OAI22_X1 port map( A1 => n6741, A2 => n9413, B1 => n6709, B2 => 
                           n9410, ZN => n7774);
   U8157 : AOI221_X1 port map( B1 => n9419, B2 => n4330, C1 => n9416, C2 => 
                           n3946, A => n7755, ZN => n7750);
   U8158 : OAI22_X1 port map( A1 => n6740, A2 => n9413, B1 => n6708, B2 => 
                           n9410, ZN => n7755);
   U8159 : AOI221_X1 port map( B1 => n9419, B2 => n4329, C1 => n9416, C2 => 
                           n3945, A => n7736, ZN => n7731);
   U8160 : OAI22_X1 port map( A1 => n6739, A2 => n9413, B1 => n6707, B2 => 
                           n9410, ZN => n7736);
   U8161 : AOI221_X1 port map( B1 => n9419, B2 => n4328, C1 => n9416, C2 => 
                           n3944, A => n7717, ZN => n7712);
   U8162 : OAI22_X1 port map( A1 => n6738, A2 => n9413, B1 => n6706, B2 => 
                           n9410, ZN => n7717);
   U8163 : AOI221_X1 port map( B1 => n9419, B2 => n4327, C1 => n9416, C2 => 
                           n3943, A => n7698, ZN => n7693);
   U8164 : OAI22_X1 port map( A1 => n6737, A2 => n9413, B1 => n6705, B2 => 
                           n9410, ZN => n7698);
   U8165 : AOI221_X1 port map( B1 => n9419, B2 => n4326, C1 => n9416, C2 => 
                           n3942, A => n7679, ZN => n7674);
   U8166 : OAI22_X1 port map( A1 => n6736, A2 => n9413, B1 => n6704, B2 => 
                           n9410, ZN => n7679);
   U8167 : AOI221_X1 port map( B1 => n9420, B2 => n4325, C1 => n9417, C2 => 
                           n3941, A => n7660, ZN => n7655);
   U8168 : OAI22_X1 port map( A1 => n6735, A2 => n9414, B1 => n6703, B2 => 
                           n9411, ZN => n7660);
   U8169 : AOI221_X1 port map( B1 => n9420, B2 => n4324, C1 => n9417, C2 => 
                           n3940, A => n7641, ZN => n7636);
   U8170 : OAI22_X1 port map( A1 => n6734, A2 => n9414, B1 => n6702, B2 => 
                           n9411, ZN => n7641);
   U8171 : AOI221_X1 port map( B1 => n9420, B2 => n4323, C1 => n9417, C2 => 
                           n3939, A => n7622, ZN => n7617);
   U8172 : OAI22_X1 port map( A1 => n6733, A2 => n9414, B1 => n6701, B2 => 
                           n9411, ZN => n7622);
   U8173 : AOI221_X1 port map( B1 => n9420, B2 => n4322, C1 => n9417, C2 => 
                           n3938, A => n7603, ZN => n7598);
   U8174 : OAI22_X1 port map( A1 => n6732, A2 => n9414, B1 => n6700, B2 => 
                           n9411, ZN => n7603);
   U8175 : AOI221_X1 port map( B1 => n9420, B2 => n4321, C1 => n9417, C2 => 
                           n3937, A => n7584, ZN => n7579);
   U8176 : OAI22_X1 port map( A1 => n6731, A2 => n9414, B1 => n6699, B2 => 
                           n9411, ZN => n7584);
   U8177 : AOI221_X1 port map( B1 => n9420, B2 => n4320, C1 => n9417, C2 => 
                           n3936, A => n7565, ZN => n7560);
   U8178 : OAI22_X1 port map( A1 => n6730, A2 => n9414, B1 => n6698, B2 => 
                           n9411, ZN => n7565);
   U8179 : AOI221_X1 port map( B1 => n9420, B2 => n4319, C1 => n9417, C2 => 
                           n3935, A => n7546, ZN => n7541);
   U8180 : OAI22_X1 port map( A1 => n6729, A2 => n9414, B1 => n6697, B2 => 
                           n9411, ZN => n7546);
   U8181 : AOI221_X1 port map( B1 => n9420, B2 => n4318, C1 => n9417, C2 => 
                           n3934, A => n7521, ZN => n7506);
   U8182 : OAI22_X1 port map( A1 => n6728, A2 => n9414, B1 => n6696, B2 => 
                           n9411, ZN => n7521);
   U8183 : OAI22_X1 port map( A1 => n9749, A2 => n9852, B1 => n7441, B2 => 
                           n6575, ZN => n3478);
   U8184 : OAI22_X1 port map( A1 => n9750, A2 => n9855, B1 => n7441, B2 => 
                           n6574, ZN => n3479);
   U8185 : OAI22_X1 port map( A1 => n9750, A2 => n9858, B1 => n7441, B2 => 
                           n6573, ZN => n3480);
   U8186 : OAI22_X1 port map( A1 => n9750, A2 => n9861, B1 => n7441, B2 => 
                           n6572, ZN => n3481);
   U8187 : OAI22_X1 port map( A1 => n9750, A2 => n9864, B1 => n7441, B2 => 
                           n6571, ZN => n3482);
   U8188 : OAI22_X1 port map( A1 => n9750, A2 => n9867, B1 => n7441, B2 => 
                           n6570, ZN => n3483);
   U8189 : OAI22_X1 port map( A1 => n9751, A2 => n9870, B1 => n7441, B2 => 
                           n6569, ZN => n3484);
   U8190 : OAI22_X1 port map( A1 => n9751, A2 => n9882, B1 => n7441, B2 => 
                           n6568, ZN => n3485);
   U8191 : OAI22_X1 port map( A1 => n9507, A2 => n9780, B1 => n9293, B2 => 
                           n7476, ZN => n2590);
   U8192 : OAI22_X1 port map( A1 => n9515, A2 => n9854, B1 => n8934, B2 => 
                           n7475, ZN => n2646);
   U8193 : OAI22_X1 port map( A1 => n9516, A2 => n9857, B1 => n8919, B2 => 
                           n7475, ZN => n2647);
   U8194 : OAI22_X1 port map( A1 => n9516, A2 => n9860, B1 => n8904, B2 => 
                           n7475, ZN => n2648);
   U8195 : OAI22_X1 port map( A1 => n9516, A2 => n9863, B1 => n8889, B2 => 
                           n7475, ZN => n2649);
   U8196 : OAI22_X1 port map( A1 => n9516, A2 => n9866, B1 => n8874, B2 => 
                           n7475, ZN => n2650);
   U8197 : OAI22_X1 port map( A1 => n9516, A2 => n9869, B1 => n8859, B2 => 
                           n7475, ZN => n2651);
   U8198 : OAI22_X1 port map( A1 => n9517, A2 => n9872, B1 => n8844, B2 => 
                           n7475, ZN => n2652);
   U8199 : OAI22_X1 port map( A1 => n9517, A2 => n9884, B1 => n8829, B2 => 
                           n7475, ZN => n2653);
   U8200 : OAI22_X1 port map( A1 => n9542, A2 => n9854, B1 => n8931, B2 => 
                           n7472, ZN => n2742);
   U8201 : OAI22_X1 port map( A1 => n9543, A2 => n9857, B1 => n8916, B2 => 
                           n7472, ZN => n2743);
   U8202 : OAI22_X1 port map( A1 => n9543, A2 => n9860, B1 => n8901, B2 => 
                           n7472, ZN => n2744);
   U8203 : OAI22_X1 port map( A1 => n9543, A2 => n9863, B1 => n8886, B2 => 
                           n7472, ZN => n2745);
   U8204 : OAI22_X1 port map( A1 => n9543, A2 => n9866, B1 => n8871, B2 => 
                           n7472, ZN => n2746);
   U8205 : OAI22_X1 port map( A1 => n9543, A2 => n9869, B1 => n8856, B2 => 
                           n7472, ZN => n2747);
   U8206 : OAI22_X1 port map( A1 => n9544, A2 => n9872, B1 => n8841, B2 => 
                           n7472, ZN => n2748);
   U8207 : OAI22_X1 port map( A1 => n9544, A2 => n9884, B1 => n8826, B2 => 
                           n7472, ZN => n2749);
   U8208 : OAI22_X1 port map( A1 => n9551, A2 => n9854, B1 => n8932, B2 => 
                           n7471, ZN => n2774);
   U8209 : OAI22_X1 port map( A1 => n9552, A2 => n9857, B1 => n8917, B2 => 
                           n7471, ZN => n2775);
   U8210 : OAI22_X1 port map( A1 => n9552, A2 => n9860, B1 => n8902, B2 => 
                           n7471, ZN => n2776);
   U8211 : OAI22_X1 port map( A1 => n9552, A2 => n9863, B1 => n8887, B2 => 
                           n7471, ZN => n2777);
   U8212 : OAI22_X1 port map( A1 => n9552, A2 => n9866, B1 => n8872, B2 => 
                           n7471, ZN => n2778);
   U8213 : OAI22_X1 port map( A1 => n9552, A2 => n9869, B1 => n8857, B2 => 
                           n7471, ZN => n2779);
   U8214 : OAI22_X1 port map( A1 => n9553, A2 => n9872, B1 => n8842, B2 => 
                           n7471, ZN => n2780);
   U8215 : OAI22_X1 port map( A1 => n9553, A2 => n9884, B1 => n8827, B2 => 
                           n7471, ZN => n2781);
   U8216 : OAI22_X1 port map( A1 => n9596, A2 => n9853, B1 => n8929, B2 => 
                           n7465, ZN => n2934);
   U8217 : OAI22_X1 port map( A1 => n9597, A2 => n9856, B1 => n8914, B2 => 
                           n7465, ZN => n2935);
   U8218 : OAI22_X1 port map( A1 => n9597, A2 => n9859, B1 => n8899, B2 => 
                           n7465, ZN => n2936);
   U8219 : OAI22_X1 port map( A1 => n9597, A2 => n9862, B1 => n8884, B2 => 
                           n7465, ZN => n2937);
   U8220 : OAI22_X1 port map( A1 => n9597, A2 => n9865, B1 => n8869, B2 => 
                           n7465, ZN => n2938);
   U8221 : OAI22_X1 port map( A1 => n9597, A2 => n9868, B1 => n8854, B2 => 
                           n7465, ZN => n2939);
   U8222 : OAI22_X1 port map( A1 => n9598, A2 => n9871, B1 => n8839, B2 => 
                           n7465, ZN => n2940);
   U8223 : OAI22_X1 port map( A1 => n9598, A2 => n9883, B1 => n8824, B2 => 
                           n7465, ZN => n2941);
   U8224 : OAI22_X1 port map( A1 => n9605, A2 => n9853, B1 => n8930, B2 => 
                           n7464, ZN => n2966);
   U8225 : OAI22_X1 port map( A1 => n9606, A2 => n9856, B1 => n8915, B2 => 
                           n7464, ZN => n2967);
   U8226 : OAI22_X1 port map( A1 => n9606, A2 => n9859, B1 => n8900, B2 => 
                           n7464, ZN => n2968);
   U8227 : OAI22_X1 port map( A1 => n9606, A2 => n9862, B1 => n8885, B2 => 
                           n7464, ZN => n2969);
   U8228 : OAI22_X1 port map( A1 => n9606, A2 => n9865, B1 => n8870, B2 => 
                           n7464, ZN => n2970);
   U8229 : OAI22_X1 port map( A1 => n9606, A2 => n9868, B1 => n8855, B2 => 
                           n7464, ZN => n2971);
   U8230 : OAI22_X1 port map( A1 => n9607, A2 => n9871, B1 => n8840, B2 => 
                           n7464, ZN => n2972);
   U8231 : OAI22_X1 port map( A1 => n9607, A2 => n9883, B1 => n8825, B2 => 
                           n7464, ZN => n2973);
   U8232 : OAI22_X1 port map( A1 => n9632, A2 => n9853, B1 => n8927, B2 => 
                           n7461, ZN => n3062);
   U8233 : OAI22_X1 port map( A1 => n9633, A2 => n9856, B1 => n8912, B2 => 
                           n7461, ZN => n3063);
   U8234 : OAI22_X1 port map( A1 => n9633, A2 => n9859, B1 => n8897, B2 => 
                           n7461, ZN => n3064);
   U8235 : OAI22_X1 port map( A1 => n9633, A2 => n9862, B1 => n8882, B2 => 
                           n7461, ZN => n3065);
   U8236 : OAI22_X1 port map( A1 => n9633, A2 => n9865, B1 => n8867, B2 => 
                           n7461, ZN => n3066);
   U8237 : OAI22_X1 port map( A1 => n9633, A2 => n9868, B1 => n8852, B2 => 
                           n7461, ZN => n3067);
   U8238 : OAI22_X1 port map( A1 => n9634, A2 => n9871, B1 => n8837, B2 => 
                           n7461, ZN => n3068);
   U8239 : OAI22_X1 port map( A1 => n9634, A2 => n9883, B1 => n8822, B2 => 
                           n7461, ZN => n3069);
   U8240 : OAI22_X1 port map( A1 => n9641, A2 => n9853, B1 => n8928, B2 => 
                           n7459, ZN => n3094);
   U8241 : OAI22_X1 port map( A1 => n9642, A2 => n9856, B1 => n8913, B2 => 
                           n7459, ZN => n3095);
   U8242 : OAI22_X1 port map( A1 => n9642, A2 => n9859, B1 => n8898, B2 => 
                           n7459, ZN => n3096);
   U8243 : OAI22_X1 port map( A1 => n9642, A2 => n9862, B1 => n8883, B2 => 
                           n7459, ZN => n3097);
   U8244 : OAI22_X1 port map( A1 => n9642, A2 => n9865, B1 => n8868, B2 => 
                           n7459, ZN => n3098);
   U8245 : OAI22_X1 port map( A1 => n9642, A2 => n9868, B1 => n8853, B2 => 
                           n7459, ZN => n3099);
   U8246 : OAI22_X1 port map( A1 => n9643, A2 => n9871, B1 => n8838, B2 => 
                           n7459, ZN => n3100);
   U8247 : OAI22_X1 port map( A1 => n9643, A2 => n9883, B1 => n8823, B2 => 
                           n7459, ZN => n3101);
   U8248 : OAI22_X1 port map( A1 => n9668, A2 => n9853, B1 => n8925, B2 => 
                           n7456, ZN => n3190);
   U8249 : OAI22_X1 port map( A1 => n9669, A2 => n9856, B1 => n8910, B2 => 
                           n7456, ZN => n3191);
   U8250 : OAI22_X1 port map( A1 => n9669, A2 => n9859, B1 => n8895, B2 => 
                           n7456, ZN => n3192);
   U8251 : OAI22_X1 port map( A1 => n9669, A2 => n9862, B1 => n8880, B2 => 
                           n7456, ZN => n3193);
   U8252 : OAI22_X1 port map( A1 => n9669, A2 => n9865, B1 => n8865, B2 => 
                           n7456, ZN => n3194);
   U8253 : OAI22_X1 port map( A1 => n9669, A2 => n9868, B1 => n8850, B2 => 
                           n7456, ZN => n3195);
   U8254 : OAI22_X1 port map( A1 => n9670, A2 => n9871, B1 => n8835, B2 => 
                           n7456, ZN => n3196);
   U8255 : OAI22_X1 port map( A1 => n9670, A2 => n9883, B1 => n8820, B2 => 
                           n7456, ZN => n3197);
   U8256 : OAI22_X1 port map( A1 => n9677, A2 => n9853, B1 => n8926, B2 => 
                           n7455, ZN => n3222);
   U8257 : OAI22_X1 port map( A1 => n9678, A2 => n9856, B1 => n8911, B2 => 
                           n7455, ZN => n3223);
   U8258 : OAI22_X1 port map( A1 => n9678, A2 => n9859, B1 => n8896, B2 => 
                           n7455, ZN => n3224);
   U8259 : OAI22_X1 port map( A1 => n9678, A2 => n9862, B1 => n8881, B2 => 
                           n7455, ZN => n3225);
   U8260 : OAI22_X1 port map( A1 => n9678, A2 => n9865, B1 => n8866, B2 => 
                           n7455, ZN => n3226);
   U8261 : OAI22_X1 port map( A1 => n9678, A2 => n9868, B1 => n8851, B2 => 
                           n7455, ZN => n3227);
   U8262 : OAI22_X1 port map( A1 => n9679, A2 => n9871, B1 => n8836, B2 => 
                           n7455, ZN => n3228);
   U8263 : OAI22_X1 port map( A1 => n9679, A2 => n9883, B1 => n8821, B2 => 
                           n7455, ZN => n3229);
   U8264 : OAI22_X1 port map( A1 => n9722, A2 => n9852, B1 => n8924, B2 => 
                           n7447, ZN => n3382);
   U8265 : OAI22_X1 port map( A1 => n9723, A2 => n9855, B1 => n8909, B2 => 
                           n7447, ZN => n3383);
   U8266 : OAI22_X1 port map( A1 => n9723, A2 => n9858, B1 => n8894, B2 => 
                           n7447, ZN => n3384);
   U8267 : OAI22_X1 port map( A1 => n9723, A2 => n9861, B1 => n8879, B2 => 
                           n7447, ZN => n3385);
   U8268 : OAI22_X1 port map( A1 => n9723, A2 => n9864, B1 => n8864, B2 => 
                           n7447, ZN => n3386);
   U8269 : OAI22_X1 port map( A1 => n9723, A2 => n9867, B1 => n8849, B2 => 
                           n7447, ZN => n3387);
   U8270 : OAI22_X1 port map( A1 => n9724, A2 => n9870, B1 => n8834, B2 => 
                           n7447, ZN => n3388);
   U8271 : OAI22_X1 port map( A1 => n9724, A2 => n9882, B1 => n8819, B2 => 
                           n7447, ZN => n3389);
   U8272 : OAI22_X1 port map( A1 => n9731, A2 => n9852, B1 => n8923, B2 => 
                           n7445, ZN => n3414);
   U8273 : OAI22_X1 port map( A1 => n9732, A2 => n9855, B1 => n8908, B2 => 
                           n7445, ZN => n3415);
   U8274 : OAI22_X1 port map( A1 => n9732, A2 => n9858, B1 => n8893, B2 => 
                           n7445, ZN => n3416);
   U8275 : OAI22_X1 port map( A1 => n9732, A2 => n9861, B1 => n8878, B2 => 
                           n7445, ZN => n3417);
   U8276 : OAI22_X1 port map( A1 => n9732, A2 => n9864, B1 => n8863, B2 => 
                           n7445, ZN => n3418);
   U8277 : OAI22_X1 port map( A1 => n9732, A2 => n9867, B1 => n8848, B2 => 
                           n7445, ZN => n3419);
   U8278 : OAI22_X1 port map( A1 => n9733, A2 => n9870, B1 => n8833, B2 => 
                           n7445, ZN => n3420);
   U8279 : OAI22_X1 port map( A1 => n9733, A2 => n9882, B1 => n8818, B2 => 
                           n7445, ZN => n3421);
   U8280 : OAI22_X1 port map( A1 => n9758, A2 => n9852, B1 => n8922, B2 => 
                           n7439, ZN => n3510);
   U8281 : OAI22_X1 port map( A1 => n9759, A2 => n9855, B1 => n8907, B2 => 
                           n7439, ZN => n3511);
   U8282 : OAI22_X1 port map( A1 => n9759, A2 => n9858, B1 => n8892, B2 => 
                           n7439, ZN => n3512);
   U8283 : OAI22_X1 port map( A1 => n9759, A2 => n9861, B1 => n8877, B2 => 
                           n7439, ZN => n3513);
   U8284 : OAI22_X1 port map( A1 => n9759, A2 => n9864, B1 => n8862, B2 => 
                           n7439, ZN => n3514);
   U8285 : OAI22_X1 port map( A1 => n9759, A2 => n9867, B1 => n8847, B2 => 
                           n7439, ZN => n3515);
   U8286 : OAI22_X1 port map( A1 => n9760, A2 => n9870, B1 => n8832, B2 => 
                           n7439, ZN => n3516);
   U8287 : OAI22_X1 port map( A1 => n9760, A2 => n9882, B1 => n8817, B2 => 
                           n7439, ZN => n3517);
   U8288 : OAI22_X1 port map( A1 => n9767, A2 => n9852, B1 => n8921, B2 => 
                           n7437, ZN => n3542);
   U8289 : OAI22_X1 port map( A1 => n9768, A2 => n9855, B1 => n8906, B2 => 
                           n7437, ZN => n3543);
   U8290 : OAI22_X1 port map( A1 => n9768, A2 => n9858, B1 => n8891, B2 => 
                           n7437, ZN => n3544);
   U8291 : OAI22_X1 port map( A1 => n9768, A2 => n9861, B1 => n8876, B2 => 
                           n7437, ZN => n3545);
   U8292 : OAI22_X1 port map( A1 => n9768, A2 => n9864, B1 => n8861, B2 => 
                           n7437, ZN => n3546);
   U8293 : OAI22_X1 port map( A1 => n9768, A2 => n9867, B1 => n8846, B2 => 
                           n7437, ZN => n3547);
   U8294 : OAI22_X1 port map( A1 => n9769, A2 => n9870, B1 => n8831, B2 => 
                           n7437, ZN => n3548);
   U8295 : OAI22_X1 port map( A1 => n9769, A2 => n9882, B1 => n8816, B2 => 
                           n7437, ZN => n3549);
   U8296 : OAI22_X1 port map( A1 => n9745, A2 => n9782, B1 => n9744, B2 => 
                           n6599, ZN => n3454);
   U8297 : OAI22_X1 port map( A1 => n9745, A2 => n9783, B1 => n9744, B2 => 
                           n6598, ZN => n3455);
   U8298 : OAI22_X1 port map( A1 => n9745, A2 => n9786, B1 => n9744, B2 => 
                           n6597, ZN => n3456);
   U8299 : OAI22_X1 port map( A1 => n9745, A2 => n9789, B1 => n9744, B2 => 
                           n6596, ZN => n3457);
   U8300 : OAI22_X1 port map( A1 => n9745, A2 => n9792, B1 => n9744, B2 => 
                           n6595, ZN => n3458);
   U8301 : OAI22_X1 port map( A1 => n9746, A2 => n9795, B1 => n9744, B2 => 
                           n6594, ZN => n3459);
   U8302 : OAI22_X1 port map( A1 => n9746, A2 => n9798, B1 => n9744, B2 => 
                           n6593, ZN => n3460);
   U8303 : OAI22_X1 port map( A1 => n9746, A2 => n9801, B1 => n9744, B2 => 
                           n6592, ZN => n3461);
   U8304 : OAI22_X1 port map( A1 => n9746, A2 => n9804, B1 => n9744, B2 => 
                           n6591, ZN => n3462);
   U8305 : OAI22_X1 port map( A1 => n9746, A2 => n9807, B1 => n9744, B2 => 
                           n6590, ZN => n3463);
   U8306 : OAI22_X1 port map( A1 => n9747, A2 => n9810, B1 => n9744, B2 => 
                           n6589, ZN => n3464);
   U8307 : OAI22_X1 port map( A1 => n9747, A2 => n9813, B1 => n9744, B2 => 
                           n6588, ZN => n3465);
   U8308 : OAI22_X1 port map( A1 => n9747, A2 => n9816, B1 => n7441, B2 => 
                           n6587, ZN => n3466);
   U8309 : OAI22_X1 port map( A1 => n9747, A2 => n9819, B1 => n7441, B2 => 
                           n6586, ZN => n3467);
   U8310 : OAI22_X1 port map( A1 => n9747, A2 => n9822, B1 => n7441, B2 => 
                           n6585, ZN => n3468);
   U8311 : OAI22_X1 port map( A1 => n9748, A2 => n9825, B1 => n9744, B2 => 
                           n6584, ZN => n3469);
   U8312 : OAI22_X1 port map( A1 => n9748, A2 => n9828, B1 => n9744, B2 => 
                           n6583, ZN => n3470);
   U8313 : OAI22_X1 port map( A1 => n9748, A2 => n9831, B1 => n9744, B2 => 
                           n6582, ZN => n3471);
   U8314 : OAI22_X1 port map( A1 => n9748, A2 => n9834, B1 => n9744, B2 => 
                           n6581, ZN => n3472);
   U8315 : OAI22_X1 port map( A1 => n9748, A2 => n9837, B1 => n9744, B2 => 
                           n6580, ZN => n3473);
   U8316 : OAI22_X1 port map( A1 => n9749, A2 => n9840, B1 => n9744, B2 => 
                           n6579, ZN => n3474);
   U8317 : OAI22_X1 port map( A1 => n9749, A2 => n9843, B1 => n9744, B2 => 
                           n6578, ZN => n3475);
   U8318 : OAI22_X1 port map( A1 => n9749, A2 => n9846, B1 => n9744, B2 => 
                           n6577, ZN => n3476);
   U8319 : OAI22_X1 port map( A1 => n9749, A2 => n9849, B1 => n9744, B2 => 
                           n6576, ZN => n3477);
   U8320 : OAI22_X1 port map( A1 => n9278, A2 => n9499, B1 => n9507, B2 => 
                           n9785, ZN => n2591);
   U8321 : OAI22_X1 port map( A1 => n9263, A2 => n7476, B1 => n9507, B2 => 
                           n9788, ZN => n2592);
   U8322 : OAI22_X1 port map( A1 => n9248, A2 => n9499, B1 => n9507, B2 => 
                           n9791, ZN => n2593);
   U8323 : OAI22_X1 port map( A1 => n9233, A2 => n7476, B1 => n9506, B2 => 
                           n9794, ZN => n2594);
   U8324 : OAI22_X1 port map( A1 => n9218, A2 => n9499, B1 => n9506, B2 => 
                           n9797, ZN => n2595);
   U8325 : OAI22_X1 port map( A1 => n9203, A2 => n7476, B1 => n9506, B2 => 
                           n9800, ZN => n2596);
   U8326 : OAI22_X1 port map( A1 => n9188, A2 => n9499, B1 => n9506, B2 => 
                           n9803, ZN => n2597);
   U8327 : OAI22_X1 port map( A1 => n9173, A2 => n7476, B1 => n9505, B2 => 
                           n9806, ZN => n2598);
   U8328 : OAI22_X1 port map( A1 => n9158, A2 => n9499, B1 => n9505, B2 => 
                           n9809, ZN => n2599);
   U8329 : OAI22_X1 port map( A1 => n9143, A2 => n9499, B1 => n9505, B2 => 
                           n9812, ZN => n2600);
   U8330 : OAI22_X1 port map( A1 => n9128, A2 => n9499, B1 => n9505, B2 => 
                           n9815, ZN => n2601);
   U8331 : OAI22_X1 port map( A1 => n9113, A2 => n9499, B1 => n9504, B2 => 
                           n9818, ZN => n2602);
   U8332 : OAI22_X1 port map( A1 => n9098, A2 => n9499, B1 => n9504, B2 => 
                           n9821, ZN => n2603);
   U8333 : OAI22_X1 port map( A1 => n9083, A2 => n9499, B1 => n9504, B2 => 
                           n9824, ZN => n2604);
   U8334 : OAI22_X1 port map( A1 => n9068, A2 => n9499, B1 => n9504, B2 => 
                           n9827, ZN => n2605);
   U8335 : OAI22_X1 port map( A1 => n9053, A2 => n9499, B1 => n9503, B2 => 
                           n9830, ZN => n2606);
   U8336 : OAI22_X1 port map( A1 => n9038, A2 => n9499, B1 => n9503, B2 => 
                           n9833, ZN => n2607);
   U8337 : OAI22_X1 port map( A1 => n9023, A2 => n9499, B1 => n9503, B2 => 
                           n9836, ZN => n2608);
   U8338 : OAI22_X1 port map( A1 => n9008, A2 => n9499, B1 => n9503, B2 => 
                           n9839, ZN => n2609);
   U8339 : OAI22_X1 port map( A1 => n8993, A2 => n7476, B1 => n9502, B2 => 
                           n9842, ZN => n2610);
   U8340 : OAI22_X1 port map( A1 => n8978, A2 => n9499, B1 => n9502, B2 => 
                           n9845, ZN => n2611);
   U8341 : OAI22_X1 port map( A1 => n8963, A2 => n7476, B1 => n9502, B2 => 
                           n9848, ZN => n2612);
   U8342 : OAI22_X1 port map( A1 => n8948, A2 => n9499, B1 => n9502, B2 => 
                           n9851, ZN => n2613);
   U8343 : OAI22_X1 port map( A1 => n8933, A2 => n7476, B1 => n9501, B2 => 
                           n9854, ZN => n2614);
   U8344 : OAI22_X1 port map( A1 => n8918, A2 => n9499, B1 => n9501, B2 => 
                           n9857, ZN => n2615);
   U8345 : OAI22_X1 port map( A1 => n8903, A2 => n7476, B1 => n9501, B2 => 
                           n9860, ZN => n2616);
   U8346 : OAI22_X1 port map( A1 => n8888, A2 => n9499, B1 => n9501, B2 => 
                           n9863, ZN => n2617);
   U8347 : OAI22_X1 port map( A1 => n8873, A2 => n7476, B1 => n9500, B2 => 
                           n9866, ZN => n2618);
   U8348 : OAI22_X1 port map( A1 => n8858, A2 => n9499, B1 => n9500, B2 => 
                           n9869, ZN => n2619);
   U8349 : OAI22_X1 port map( A1 => n8843, A2 => n7476, B1 => n9500, B2 => 
                           n9872, ZN => n2620);
   U8350 : OAI22_X1 port map( A1 => n8828, A2 => n9499, B1 => n9500, B2 => 
                           n9884, ZN => n2621);
   U8351 : OAI22_X1 port map( A1 => n9511, A2 => n9780, B1 => n9294, B2 => 
                           n9510, ZN => n2622);
   U8352 : OAI22_X1 port map( A1 => n9511, A2 => n9785, B1 => n9279, B2 => 
                           n9510, ZN => n2623);
   U8353 : OAI22_X1 port map( A1 => n9511, A2 => n9788, B1 => n9264, B2 => 
                           n9510, ZN => n2624);
   U8354 : OAI22_X1 port map( A1 => n9511, A2 => n9791, B1 => n9249, B2 => 
                           n9510, ZN => n2625);
   U8355 : OAI22_X1 port map( A1 => n9511, A2 => n9794, B1 => n9234, B2 => 
                           n9510, ZN => n2626);
   U8356 : OAI22_X1 port map( A1 => n9512, A2 => n9797, B1 => n9219, B2 => 
                           n9510, ZN => n2627);
   U8357 : OAI22_X1 port map( A1 => n9512, A2 => n9800, B1 => n9204, B2 => 
                           n9510, ZN => n2628);
   U8358 : OAI22_X1 port map( A1 => n9512, A2 => n9803, B1 => n9189, B2 => 
                           n9510, ZN => n2629);
   U8359 : OAI22_X1 port map( A1 => n9512, A2 => n9806, B1 => n9174, B2 => 
                           n9510, ZN => n2630);
   U8360 : OAI22_X1 port map( A1 => n9512, A2 => n9809, B1 => n9159, B2 => 
                           n9510, ZN => n2631);
   U8361 : OAI22_X1 port map( A1 => n9513, A2 => n9812, B1 => n9144, B2 => 
                           n9510, ZN => n2632);
   U8362 : OAI22_X1 port map( A1 => n9513, A2 => n9815, B1 => n9129, B2 => 
                           n9510, ZN => n2633);
   U8363 : OAI22_X1 port map( A1 => n9513, A2 => n9818, B1 => n9114, B2 => 
                           n7475, ZN => n2634);
   U8364 : OAI22_X1 port map( A1 => n9513, A2 => n9821, B1 => n9099, B2 => 
                           n7475, ZN => n2635);
   U8365 : OAI22_X1 port map( A1 => n9513, A2 => n9824, B1 => n9084, B2 => 
                           n7475, ZN => n2636);
   U8366 : OAI22_X1 port map( A1 => n9514, A2 => n9827, B1 => n9069, B2 => 
                           n9510, ZN => n2637);
   U8367 : OAI22_X1 port map( A1 => n9514, A2 => n9830, B1 => n9054, B2 => 
                           n9510, ZN => n2638);
   U8368 : OAI22_X1 port map( A1 => n9514, A2 => n9833, B1 => n9039, B2 => 
                           n9510, ZN => n2639);
   U8369 : OAI22_X1 port map( A1 => n9514, A2 => n9836, B1 => n9024, B2 => 
                           n9510, ZN => n2640);
   U8370 : OAI22_X1 port map( A1 => n9514, A2 => n9839, B1 => n9009, B2 => 
                           n9510, ZN => n2641);
   U8371 : OAI22_X1 port map( A1 => n9515, A2 => n9842, B1 => n8994, B2 => 
                           n9510, ZN => n2642);
   U8372 : OAI22_X1 port map( A1 => n9515, A2 => n9845, B1 => n8979, B2 => 
                           n9510, ZN => n2643);
   U8373 : OAI22_X1 port map( A1 => n9515, A2 => n9848, B1 => n8964, B2 => 
                           n9510, ZN => n2644);
   U8374 : OAI22_X1 port map( A1 => n9515, A2 => n9851, B1 => n8949, B2 => 
                           n9510, ZN => n2645);
   U8375 : OAI22_X1 port map( A1 => n9538, A2 => n9780, B1 => n9291, B2 => 
                           n9537, ZN => n2718);
   U8376 : OAI22_X1 port map( A1 => n9538, A2 => n9785, B1 => n9276, B2 => 
                           n9537, ZN => n2719);
   U8377 : OAI22_X1 port map( A1 => n9538, A2 => n9788, B1 => n9261, B2 => 
                           n9537, ZN => n2720);
   U8378 : OAI22_X1 port map( A1 => n9538, A2 => n9791, B1 => n9246, B2 => 
                           n9537, ZN => n2721);
   U8379 : OAI22_X1 port map( A1 => n9538, A2 => n9794, B1 => n9231, B2 => 
                           n9537, ZN => n2722);
   U8380 : OAI22_X1 port map( A1 => n9539, A2 => n9797, B1 => n9216, B2 => 
                           n9537, ZN => n2723);
   U8381 : OAI22_X1 port map( A1 => n9539, A2 => n9800, B1 => n9201, B2 => 
                           n9537, ZN => n2724);
   U8382 : OAI22_X1 port map( A1 => n9539, A2 => n9803, B1 => n9186, B2 => 
                           n9537, ZN => n2725);
   U8383 : OAI22_X1 port map( A1 => n9539, A2 => n9806, B1 => n9171, B2 => 
                           n9537, ZN => n2726);
   U8384 : OAI22_X1 port map( A1 => n9539, A2 => n9809, B1 => n9156, B2 => 
                           n9537, ZN => n2727);
   U8385 : OAI22_X1 port map( A1 => n9540, A2 => n9812, B1 => n9141, B2 => 
                           n9537, ZN => n2728);
   U8386 : OAI22_X1 port map( A1 => n9540, A2 => n9815, B1 => n9126, B2 => 
                           n9537, ZN => n2729);
   U8387 : OAI22_X1 port map( A1 => n9540, A2 => n9818, B1 => n9111, B2 => 
                           n7472, ZN => n2730);
   U8388 : OAI22_X1 port map( A1 => n9540, A2 => n9821, B1 => n9096, B2 => 
                           n7472, ZN => n2731);
   U8389 : OAI22_X1 port map( A1 => n9540, A2 => n9824, B1 => n9081, B2 => 
                           n7472, ZN => n2732);
   U8390 : OAI22_X1 port map( A1 => n9541, A2 => n9827, B1 => n9066, B2 => 
                           n9537, ZN => n2733);
   U8391 : OAI22_X1 port map( A1 => n9541, A2 => n9830, B1 => n9051, B2 => 
                           n9537, ZN => n2734);
   U8392 : OAI22_X1 port map( A1 => n9541, A2 => n9833, B1 => n9036, B2 => 
                           n9537, ZN => n2735);
   U8393 : OAI22_X1 port map( A1 => n9541, A2 => n9836, B1 => n9021, B2 => 
                           n9537, ZN => n2736);
   U8394 : OAI22_X1 port map( A1 => n9541, A2 => n9839, B1 => n9006, B2 => 
                           n9537, ZN => n2737);
   U8395 : OAI22_X1 port map( A1 => n9542, A2 => n9842, B1 => n8991, B2 => 
                           n9537, ZN => n2738);
   U8396 : OAI22_X1 port map( A1 => n9542, A2 => n9845, B1 => n8976, B2 => 
                           n9537, ZN => n2739);
   U8397 : OAI22_X1 port map( A1 => n9542, A2 => n9848, B1 => n8961, B2 => 
                           n9537, ZN => n2740);
   U8398 : OAI22_X1 port map( A1 => n9542, A2 => n9851, B1 => n8946, B2 => 
                           n9537, ZN => n2741);
   U8399 : OAI22_X1 port map( A1 => n9547, A2 => n9780, B1 => n9292, B2 => 
                           n9546, ZN => n2750);
   U8400 : OAI22_X1 port map( A1 => n9547, A2 => n9785, B1 => n9277, B2 => 
                           n9546, ZN => n2751);
   U8401 : OAI22_X1 port map( A1 => n9547, A2 => n9788, B1 => n9262, B2 => 
                           n9546, ZN => n2752);
   U8402 : OAI22_X1 port map( A1 => n9547, A2 => n9791, B1 => n9247, B2 => 
                           n9546, ZN => n2753);
   U8403 : OAI22_X1 port map( A1 => n9547, A2 => n9794, B1 => n9232, B2 => 
                           n9546, ZN => n2754);
   U8404 : OAI22_X1 port map( A1 => n9548, A2 => n9797, B1 => n9217, B2 => 
                           n9546, ZN => n2755);
   U8405 : OAI22_X1 port map( A1 => n9548, A2 => n9800, B1 => n9202, B2 => 
                           n9546, ZN => n2756);
   U8406 : OAI22_X1 port map( A1 => n9548, A2 => n9803, B1 => n9187, B2 => 
                           n9546, ZN => n2757);
   U8407 : OAI22_X1 port map( A1 => n9548, A2 => n9806, B1 => n9172, B2 => 
                           n9546, ZN => n2758);
   U8408 : OAI22_X1 port map( A1 => n9548, A2 => n9809, B1 => n9157, B2 => 
                           n9546, ZN => n2759);
   U8409 : OAI22_X1 port map( A1 => n9549, A2 => n9812, B1 => n9142, B2 => 
                           n9546, ZN => n2760);
   U8410 : OAI22_X1 port map( A1 => n9549, A2 => n9815, B1 => n9127, B2 => 
                           n9546, ZN => n2761);
   U8411 : OAI22_X1 port map( A1 => n9549, A2 => n9818, B1 => n9112, B2 => 
                           n7471, ZN => n2762);
   U8412 : OAI22_X1 port map( A1 => n9549, A2 => n9821, B1 => n9097, B2 => 
                           n7471, ZN => n2763);
   U8413 : OAI22_X1 port map( A1 => n9549, A2 => n9824, B1 => n9082, B2 => 
                           n7471, ZN => n2764);
   U8414 : OAI22_X1 port map( A1 => n9550, A2 => n9827, B1 => n9067, B2 => 
                           n9546, ZN => n2765);
   U8415 : OAI22_X1 port map( A1 => n9550, A2 => n9830, B1 => n9052, B2 => 
                           n9546, ZN => n2766);
   U8416 : OAI22_X1 port map( A1 => n9550, A2 => n9833, B1 => n9037, B2 => 
                           n9546, ZN => n2767);
   U8417 : OAI22_X1 port map( A1 => n9550, A2 => n9836, B1 => n9022, B2 => 
                           n9546, ZN => n2768);
   U8418 : OAI22_X1 port map( A1 => n9550, A2 => n9839, B1 => n9007, B2 => 
                           n9546, ZN => n2769);
   U8419 : OAI22_X1 port map( A1 => n9551, A2 => n9842, B1 => n8992, B2 => 
                           n9546, ZN => n2770);
   U8420 : OAI22_X1 port map( A1 => n9551, A2 => n9845, B1 => n8977, B2 => 
                           n9546, ZN => n2771);
   U8421 : OAI22_X1 port map( A1 => n9551, A2 => n9848, B1 => n8962, B2 => 
                           n9546, ZN => n2772);
   U8422 : OAI22_X1 port map( A1 => n9551, A2 => n9851, B1 => n8947, B2 => 
                           n9546, ZN => n2773);
   U8423 : OAI22_X1 port map( A1 => n9592, A2 => n9780, B1 => n9289, B2 => 
                           n9591, ZN => n2910);
   U8424 : OAI22_X1 port map( A1 => n9592, A2 => n9784, B1 => n9274, B2 => 
                           n9591, ZN => n2911);
   U8425 : OAI22_X1 port map( A1 => n9592, A2 => n9787, B1 => n9259, B2 => 
                           n9591, ZN => n2912);
   U8426 : OAI22_X1 port map( A1 => n9592, A2 => n9790, B1 => n9244, B2 => 
                           n9591, ZN => n2913);
   U8427 : OAI22_X1 port map( A1 => n9592, A2 => n9793, B1 => n9229, B2 => 
                           n9591, ZN => n2914);
   U8428 : OAI22_X1 port map( A1 => n9593, A2 => n9796, B1 => n9214, B2 => 
                           n9591, ZN => n2915);
   U8429 : OAI22_X1 port map( A1 => n9593, A2 => n9799, B1 => n9199, B2 => 
                           n9591, ZN => n2916);
   U8430 : OAI22_X1 port map( A1 => n9593, A2 => n9802, B1 => n9184, B2 => 
                           n9591, ZN => n2917);
   U8431 : OAI22_X1 port map( A1 => n9593, A2 => n9805, B1 => n9169, B2 => 
                           n9591, ZN => n2918);
   U8432 : OAI22_X1 port map( A1 => n9593, A2 => n9808, B1 => n9154, B2 => 
                           n9591, ZN => n2919);
   U8433 : OAI22_X1 port map( A1 => n9594, A2 => n9811, B1 => n9139, B2 => 
                           n9591, ZN => n2920);
   U8434 : OAI22_X1 port map( A1 => n9594, A2 => n9814, B1 => n9124, B2 => 
                           n9591, ZN => n2921);
   U8435 : OAI22_X1 port map( A1 => n9594, A2 => n9817, B1 => n9109, B2 => 
                           n7465, ZN => n2922);
   U8436 : OAI22_X1 port map( A1 => n9594, A2 => n9820, B1 => n9094, B2 => 
                           n7465, ZN => n2923);
   U8437 : OAI22_X1 port map( A1 => n9594, A2 => n9823, B1 => n9079, B2 => 
                           n7465, ZN => n2924);
   U8438 : OAI22_X1 port map( A1 => n9595, A2 => n9826, B1 => n9064, B2 => 
                           n9591, ZN => n2925);
   U8439 : OAI22_X1 port map( A1 => n9595, A2 => n9829, B1 => n9049, B2 => 
                           n9591, ZN => n2926);
   U8440 : OAI22_X1 port map( A1 => n9595, A2 => n9832, B1 => n9034, B2 => 
                           n9591, ZN => n2927);
   U8441 : OAI22_X1 port map( A1 => n9595, A2 => n9835, B1 => n9019, B2 => 
                           n9591, ZN => n2928);
   U8442 : OAI22_X1 port map( A1 => n9595, A2 => n9838, B1 => n9004, B2 => 
                           n9591, ZN => n2929);
   U8443 : OAI22_X1 port map( A1 => n9596, A2 => n9841, B1 => n8989, B2 => 
                           n9591, ZN => n2930);
   U8444 : OAI22_X1 port map( A1 => n9596, A2 => n9844, B1 => n8974, B2 => 
                           n9591, ZN => n2931);
   U8445 : OAI22_X1 port map( A1 => n9596, A2 => n9847, B1 => n8959, B2 => 
                           n9591, ZN => n2932);
   U8446 : OAI22_X1 port map( A1 => n9596, A2 => n9850, B1 => n8944, B2 => 
                           n9591, ZN => n2933);
   U8447 : OAI22_X1 port map( A1 => n9601, A2 => n9780, B1 => n9290, B2 => 
                           n9600, ZN => n2942);
   U8448 : OAI22_X1 port map( A1 => n9601, A2 => n9784, B1 => n9275, B2 => 
                           n9600, ZN => n2943);
   U8449 : OAI22_X1 port map( A1 => n9601, A2 => n9787, B1 => n9260, B2 => 
                           n9600, ZN => n2944);
   U8450 : OAI22_X1 port map( A1 => n9601, A2 => n9790, B1 => n9245, B2 => 
                           n9600, ZN => n2945);
   U8451 : OAI22_X1 port map( A1 => n9601, A2 => n9793, B1 => n9230, B2 => 
                           n9600, ZN => n2946);
   U8452 : OAI22_X1 port map( A1 => n9602, A2 => n9796, B1 => n9215, B2 => 
                           n9600, ZN => n2947);
   U8453 : OAI22_X1 port map( A1 => n9602, A2 => n9799, B1 => n9200, B2 => 
                           n9600, ZN => n2948);
   U8454 : OAI22_X1 port map( A1 => n9602, A2 => n9802, B1 => n9185, B2 => 
                           n9600, ZN => n2949);
   U8455 : OAI22_X1 port map( A1 => n9602, A2 => n9805, B1 => n9170, B2 => 
                           n9600, ZN => n2950);
   U8456 : OAI22_X1 port map( A1 => n9602, A2 => n9808, B1 => n9155, B2 => 
                           n9600, ZN => n2951);
   U8457 : OAI22_X1 port map( A1 => n9603, A2 => n9811, B1 => n9140, B2 => 
                           n9600, ZN => n2952);
   U8458 : OAI22_X1 port map( A1 => n9603, A2 => n9814, B1 => n9125, B2 => 
                           n9600, ZN => n2953);
   U8459 : OAI22_X1 port map( A1 => n9603, A2 => n9817, B1 => n9110, B2 => 
                           n7464, ZN => n2954);
   U8460 : OAI22_X1 port map( A1 => n9603, A2 => n9820, B1 => n9095, B2 => 
                           n7464, ZN => n2955);
   U8461 : OAI22_X1 port map( A1 => n9603, A2 => n9823, B1 => n9080, B2 => 
                           n7464, ZN => n2956);
   U8462 : OAI22_X1 port map( A1 => n9604, A2 => n9826, B1 => n9065, B2 => 
                           n9600, ZN => n2957);
   U8463 : OAI22_X1 port map( A1 => n9604, A2 => n9829, B1 => n9050, B2 => 
                           n9600, ZN => n2958);
   U8464 : OAI22_X1 port map( A1 => n9604, A2 => n9832, B1 => n9035, B2 => 
                           n9600, ZN => n2959);
   U8465 : OAI22_X1 port map( A1 => n9604, A2 => n9835, B1 => n9020, B2 => 
                           n9600, ZN => n2960);
   U8466 : OAI22_X1 port map( A1 => n9604, A2 => n9838, B1 => n9005, B2 => 
                           n9600, ZN => n2961);
   U8467 : OAI22_X1 port map( A1 => n9605, A2 => n9841, B1 => n8990, B2 => 
                           n9600, ZN => n2962);
   U8468 : OAI22_X1 port map( A1 => n9605, A2 => n9844, B1 => n8975, B2 => 
                           n9600, ZN => n2963);
   U8469 : OAI22_X1 port map( A1 => n9605, A2 => n9847, B1 => n8960, B2 => 
                           n9600, ZN => n2964);
   U8470 : OAI22_X1 port map( A1 => n9605, A2 => n9850, B1 => n8945, B2 => 
                           n9600, ZN => n2965);
   U8471 : OAI22_X1 port map( A1 => n9628, A2 => n9781, B1 => n9287, B2 => 
                           n9627, ZN => n3038);
   U8472 : OAI22_X1 port map( A1 => n9628, A2 => n9784, B1 => n9272, B2 => 
                           n9627, ZN => n3039);
   U8473 : OAI22_X1 port map( A1 => n9628, A2 => n9787, B1 => n9257, B2 => 
                           n9627, ZN => n3040);
   U8474 : OAI22_X1 port map( A1 => n9628, A2 => n9790, B1 => n9242, B2 => 
                           n9627, ZN => n3041);
   U8475 : OAI22_X1 port map( A1 => n9628, A2 => n9793, B1 => n9227, B2 => 
                           n9627, ZN => n3042);
   U8476 : OAI22_X1 port map( A1 => n9629, A2 => n9796, B1 => n9212, B2 => 
                           n9627, ZN => n3043);
   U8477 : OAI22_X1 port map( A1 => n9629, A2 => n9799, B1 => n9197, B2 => 
                           n9627, ZN => n3044);
   U8478 : OAI22_X1 port map( A1 => n9629, A2 => n9802, B1 => n9182, B2 => 
                           n9627, ZN => n3045);
   U8479 : OAI22_X1 port map( A1 => n9629, A2 => n9805, B1 => n9167, B2 => 
                           n9627, ZN => n3046);
   U8480 : OAI22_X1 port map( A1 => n9629, A2 => n9808, B1 => n9152, B2 => 
                           n9627, ZN => n3047);
   U8481 : OAI22_X1 port map( A1 => n9630, A2 => n9811, B1 => n9137, B2 => 
                           n9627, ZN => n3048);
   U8482 : OAI22_X1 port map( A1 => n9630, A2 => n9814, B1 => n9122, B2 => 
                           n9627, ZN => n3049);
   U8483 : OAI22_X1 port map( A1 => n9630, A2 => n9817, B1 => n9107, B2 => 
                           n7461, ZN => n3050);
   U8484 : OAI22_X1 port map( A1 => n9630, A2 => n9820, B1 => n9092, B2 => 
                           n7461, ZN => n3051);
   U8485 : OAI22_X1 port map( A1 => n9630, A2 => n9823, B1 => n9077, B2 => 
                           n7461, ZN => n3052);
   U8486 : OAI22_X1 port map( A1 => n9631, A2 => n9826, B1 => n9062, B2 => 
                           n9627, ZN => n3053);
   U8487 : OAI22_X1 port map( A1 => n9631, A2 => n9829, B1 => n9047, B2 => 
                           n9627, ZN => n3054);
   U8488 : OAI22_X1 port map( A1 => n9631, A2 => n9832, B1 => n9032, B2 => 
                           n9627, ZN => n3055);
   U8489 : OAI22_X1 port map( A1 => n9631, A2 => n9835, B1 => n9017, B2 => 
                           n9627, ZN => n3056);
   U8490 : OAI22_X1 port map( A1 => n9631, A2 => n9838, B1 => n9002, B2 => 
                           n9627, ZN => n3057);
   U8491 : OAI22_X1 port map( A1 => n9632, A2 => n9841, B1 => n8987, B2 => 
                           n9627, ZN => n3058);
   U8492 : OAI22_X1 port map( A1 => n9632, A2 => n9844, B1 => n8972, B2 => 
                           n9627, ZN => n3059);
   U8493 : OAI22_X1 port map( A1 => n9632, A2 => n9847, B1 => n8957, B2 => 
                           n9627, ZN => n3060);
   U8494 : OAI22_X1 port map( A1 => n9632, A2 => n9850, B1 => n8942, B2 => 
                           n9627, ZN => n3061);
   U8495 : OAI22_X1 port map( A1 => n9637, A2 => n9781, B1 => n9288, B2 => 
                           n9636, ZN => n3070);
   U8496 : OAI22_X1 port map( A1 => n9637, A2 => n9784, B1 => n9273, B2 => 
                           n9636, ZN => n3071);
   U8497 : OAI22_X1 port map( A1 => n9637, A2 => n9787, B1 => n9258, B2 => 
                           n9636, ZN => n3072);
   U8498 : OAI22_X1 port map( A1 => n9637, A2 => n9790, B1 => n9243, B2 => 
                           n9636, ZN => n3073);
   U8499 : OAI22_X1 port map( A1 => n9637, A2 => n9793, B1 => n9228, B2 => 
                           n9636, ZN => n3074);
   U8500 : OAI22_X1 port map( A1 => n9638, A2 => n9796, B1 => n9213, B2 => 
                           n9636, ZN => n3075);
   U8501 : OAI22_X1 port map( A1 => n9638, A2 => n9799, B1 => n9198, B2 => 
                           n9636, ZN => n3076);
   U8502 : OAI22_X1 port map( A1 => n9638, A2 => n9802, B1 => n9183, B2 => 
                           n9636, ZN => n3077);
   U8503 : OAI22_X1 port map( A1 => n9638, A2 => n9805, B1 => n9168, B2 => 
                           n9636, ZN => n3078);
   U8504 : OAI22_X1 port map( A1 => n9638, A2 => n9808, B1 => n9153, B2 => 
                           n9636, ZN => n3079);
   U8505 : OAI22_X1 port map( A1 => n9639, A2 => n9811, B1 => n9138, B2 => 
                           n9636, ZN => n3080);
   U8506 : OAI22_X1 port map( A1 => n9639, A2 => n9814, B1 => n9123, B2 => 
                           n9636, ZN => n3081);
   U8507 : OAI22_X1 port map( A1 => n9639, A2 => n9817, B1 => n9108, B2 => 
                           n7459, ZN => n3082);
   U8508 : OAI22_X1 port map( A1 => n9639, A2 => n9820, B1 => n9093, B2 => 
                           n7459, ZN => n3083);
   U8509 : OAI22_X1 port map( A1 => n9639, A2 => n9823, B1 => n9078, B2 => 
                           n7459, ZN => n3084);
   U8510 : OAI22_X1 port map( A1 => n9640, A2 => n9826, B1 => n9063, B2 => 
                           n9636, ZN => n3085);
   U8511 : OAI22_X1 port map( A1 => n9640, A2 => n9829, B1 => n9048, B2 => 
                           n9636, ZN => n3086);
   U8512 : OAI22_X1 port map( A1 => n9640, A2 => n9832, B1 => n9033, B2 => 
                           n9636, ZN => n3087);
   U8513 : OAI22_X1 port map( A1 => n9640, A2 => n9835, B1 => n9018, B2 => 
                           n9636, ZN => n3088);
   U8514 : OAI22_X1 port map( A1 => n9640, A2 => n9838, B1 => n9003, B2 => 
                           n9636, ZN => n3089);
   U8515 : OAI22_X1 port map( A1 => n9641, A2 => n9841, B1 => n8988, B2 => 
                           n9636, ZN => n3090);
   U8516 : OAI22_X1 port map( A1 => n9641, A2 => n9844, B1 => n8973, B2 => 
                           n9636, ZN => n3091);
   U8517 : OAI22_X1 port map( A1 => n9641, A2 => n9847, B1 => n8958, B2 => 
                           n9636, ZN => n3092);
   U8518 : OAI22_X1 port map( A1 => n9641, A2 => n9850, B1 => n8943, B2 => 
                           n9636, ZN => n3093);
   U8519 : OAI22_X1 port map( A1 => n9664, A2 => n9781, B1 => n9285, B2 => 
                           n9663, ZN => n3166);
   U8520 : OAI22_X1 port map( A1 => n9664, A2 => n9784, B1 => n9270, B2 => 
                           n9663, ZN => n3167);
   U8521 : OAI22_X1 port map( A1 => n9664, A2 => n9787, B1 => n9255, B2 => 
                           n9663, ZN => n3168);
   U8522 : OAI22_X1 port map( A1 => n9664, A2 => n9790, B1 => n9240, B2 => 
                           n9663, ZN => n3169);
   U8523 : OAI22_X1 port map( A1 => n9664, A2 => n9793, B1 => n9225, B2 => 
                           n9663, ZN => n3170);
   U8524 : OAI22_X1 port map( A1 => n9665, A2 => n9796, B1 => n9210, B2 => 
                           n9663, ZN => n3171);
   U8525 : OAI22_X1 port map( A1 => n9665, A2 => n9799, B1 => n9195, B2 => 
                           n9663, ZN => n3172);
   U8526 : OAI22_X1 port map( A1 => n9665, A2 => n9802, B1 => n9180, B2 => 
                           n9663, ZN => n3173);
   U8527 : OAI22_X1 port map( A1 => n9665, A2 => n9805, B1 => n9165, B2 => 
                           n9663, ZN => n3174);
   U8528 : OAI22_X1 port map( A1 => n9665, A2 => n9808, B1 => n9150, B2 => 
                           n9663, ZN => n3175);
   U8529 : OAI22_X1 port map( A1 => n9666, A2 => n9811, B1 => n9135, B2 => 
                           n9663, ZN => n3176);
   U8530 : OAI22_X1 port map( A1 => n9666, A2 => n9814, B1 => n9120, B2 => 
                           n9663, ZN => n3177);
   U8531 : OAI22_X1 port map( A1 => n9666, A2 => n9817, B1 => n9105, B2 => 
                           n7456, ZN => n3178);
   U8532 : OAI22_X1 port map( A1 => n9666, A2 => n9820, B1 => n9090, B2 => 
                           n7456, ZN => n3179);
   U8533 : OAI22_X1 port map( A1 => n9666, A2 => n9823, B1 => n9075, B2 => 
                           n7456, ZN => n3180);
   U8534 : OAI22_X1 port map( A1 => n9667, A2 => n9826, B1 => n9060, B2 => 
                           n9663, ZN => n3181);
   U8535 : OAI22_X1 port map( A1 => n9667, A2 => n9829, B1 => n9045, B2 => 
                           n9663, ZN => n3182);
   U8536 : OAI22_X1 port map( A1 => n9667, A2 => n9832, B1 => n9030, B2 => 
                           n9663, ZN => n3183);
   U8537 : OAI22_X1 port map( A1 => n9667, A2 => n9835, B1 => n9015, B2 => 
                           n9663, ZN => n3184);
   U8538 : OAI22_X1 port map( A1 => n9667, A2 => n9838, B1 => n9000, B2 => 
                           n9663, ZN => n3185);
   U8539 : OAI22_X1 port map( A1 => n9668, A2 => n9841, B1 => n8985, B2 => 
                           n9663, ZN => n3186);
   U8540 : OAI22_X1 port map( A1 => n9668, A2 => n9844, B1 => n8970, B2 => 
                           n9663, ZN => n3187);
   U8541 : OAI22_X1 port map( A1 => n9668, A2 => n9847, B1 => n8955, B2 => 
                           n9663, ZN => n3188);
   U8542 : OAI22_X1 port map( A1 => n9668, A2 => n9850, B1 => n8940, B2 => 
                           n9663, ZN => n3189);
   U8543 : OAI22_X1 port map( A1 => n9673, A2 => n9781, B1 => n9286, B2 => 
                           n9672, ZN => n3198);
   U8544 : OAI22_X1 port map( A1 => n9673, A2 => n9784, B1 => n9271, B2 => 
                           n9672, ZN => n3199);
   U8545 : OAI22_X1 port map( A1 => n9673, A2 => n9787, B1 => n9256, B2 => 
                           n9672, ZN => n3200);
   U8546 : OAI22_X1 port map( A1 => n9673, A2 => n9790, B1 => n9241, B2 => 
                           n9672, ZN => n3201);
   U8547 : OAI22_X1 port map( A1 => n9673, A2 => n9793, B1 => n9226, B2 => 
                           n9672, ZN => n3202);
   U8548 : OAI22_X1 port map( A1 => n9674, A2 => n9796, B1 => n9211, B2 => 
                           n9672, ZN => n3203);
   U8549 : OAI22_X1 port map( A1 => n9674, A2 => n9799, B1 => n9196, B2 => 
                           n9672, ZN => n3204);
   U8550 : OAI22_X1 port map( A1 => n9674, A2 => n9802, B1 => n9181, B2 => 
                           n9672, ZN => n3205);
   U8551 : OAI22_X1 port map( A1 => n9674, A2 => n9805, B1 => n9166, B2 => 
                           n9672, ZN => n3206);
   U8552 : OAI22_X1 port map( A1 => n9674, A2 => n9808, B1 => n9151, B2 => 
                           n9672, ZN => n3207);
   U8553 : OAI22_X1 port map( A1 => n9675, A2 => n9811, B1 => n9136, B2 => 
                           n9672, ZN => n3208);
   U8554 : OAI22_X1 port map( A1 => n9675, A2 => n9814, B1 => n9121, B2 => 
                           n9672, ZN => n3209);
   U8555 : OAI22_X1 port map( A1 => n9675, A2 => n9817, B1 => n9106, B2 => 
                           n7455, ZN => n3210);
   U8556 : OAI22_X1 port map( A1 => n9675, A2 => n9820, B1 => n9091, B2 => 
                           n7455, ZN => n3211);
   U8557 : OAI22_X1 port map( A1 => n9675, A2 => n9823, B1 => n9076, B2 => 
                           n7455, ZN => n3212);
   U8558 : OAI22_X1 port map( A1 => n9676, A2 => n9826, B1 => n9061, B2 => 
                           n9672, ZN => n3213);
   U8559 : OAI22_X1 port map( A1 => n9676, A2 => n9829, B1 => n9046, B2 => 
                           n9672, ZN => n3214);
   U8560 : OAI22_X1 port map( A1 => n9676, A2 => n9832, B1 => n9031, B2 => 
                           n9672, ZN => n3215);
   U8561 : OAI22_X1 port map( A1 => n9676, A2 => n9835, B1 => n9016, B2 => 
                           n9672, ZN => n3216);
   U8562 : OAI22_X1 port map( A1 => n9676, A2 => n9838, B1 => n9001, B2 => 
                           n9672, ZN => n3217);
   U8563 : OAI22_X1 port map( A1 => n9677, A2 => n9841, B1 => n8986, B2 => 
                           n9672, ZN => n3218);
   U8564 : OAI22_X1 port map( A1 => n9677, A2 => n9844, B1 => n8971, B2 => 
                           n9672, ZN => n3219);
   U8565 : OAI22_X1 port map( A1 => n9677, A2 => n9847, B1 => n8956, B2 => 
                           n9672, ZN => n3220);
   U8566 : OAI22_X1 port map( A1 => n9677, A2 => n9850, B1 => n8941, B2 => 
                           n9672, ZN => n3221);
   U8567 : OAI22_X1 port map( A1 => n9718, A2 => n9782, B1 => n9284, B2 => 
                           n9717, ZN => n3358);
   U8568 : OAI22_X1 port map( A1 => n9718, A2 => n9783, B1 => n9269, B2 => 
                           n9717, ZN => n3359);
   U8569 : OAI22_X1 port map( A1 => n9718, A2 => n9786, B1 => n9254, B2 => 
                           n9717, ZN => n3360);
   U8570 : OAI22_X1 port map( A1 => n9718, A2 => n9789, B1 => n9239, B2 => 
                           n9717, ZN => n3361);
   U8571 : OAI22_X1 port map( A1 => n9718, A2 => n9792, B1 => n9224, B2 => 
                           n9717, ZN => n3362);
   U8572 : OAI22_X1 port map( A1 => n9719, A2 => n9795, B1 => n9209, B2 => 
                           n9717, ZN => n3363);
   U8573 : OAI22_X1 port map( A1 => n9719, A2 => n9798, B1 => n9194, B2 => 
                           n9717, ZN => n3364);
   U8574 : OAI22_X1 port map( A1 => n9719, A2 => n9801, B1 => n9179, B2 => 
                           n9717, ZN => n3365);
   U8575 : OAI22_X1 port map( A1 => n9719, A2 => n9804, B1 => n9164, B2 => 
                           n9717, ZN => n3366);
   U8576 : OAI22_X1 port map( A1 => n9719, A2 => n9807, B1 => n9149, B2 => 
                           n9717, ZN => n3367);
   U8577 : OAI22_X1 port map( A1 => n9720, A2 => n9810, B1 => n9134, B2 => 
                           n9717, ZN => n3368);
   U8578 : OAI22_X1 port map( A1 => n9720, A2 => n9813, B1 => n9119, B2 => 
                           n9717, ZN => n3369);
   U8579 : OAI22_X1 port map( A1 => n9720, A2 => n9816, B1 => n9104, B2 => 
                           n7447, ZN => n3370);
   U8580 : OAI22_X1 port map( A1 => n9720, A2 => n9819, B1 => n9089, B2 => 
                           n7447, ZN => n3371);
   U8581 : OAI22_X1 port map( A1 => n9720, A2 => n9822, B1 => n9074, B2 => 
                           n7447, ZN => n3372);
   U8582 : OAI22_X1 port map( A1 => n9721, A2 => n9825, B1 => n9059, B2 => 
                           n9717, ZN => n3373);
   U8583 : OAI22_X1 port map( A1 => n9721, A2 => n9828, B1 => n9044, B2 => 
                           n9717, ZN => n3374);
   U8584 : OAI22_X1 port map( A1 => n9721, A2 => n9831, B1 => n9029, B2 => 
                           n9717, ZN => n3375);
   U8585 : OAI22_X1 port map( A1 => n9721, A2 => n9834, B1 => n9014, B2 => 
                           n9717, ZN => n3376);
   U8586 : OAI22_X1 port map( A1 => n9721, A2 => n9837, B1 => n8999, B2 => 
                           n9717, ZN => n3377);
   U8587 : OAI22_X1 port map( A1 => n9722, A2 => n9840, B1 => n8984, B2 => 
                           n9717, ZN => n3378);
   U8588 : OAI22_X1 port map( A1 => n9722, A2 => n9843, B1 => n8969, B2 => 
                           n9717, ZN => n3379);
   U8589 : OAI22_X1 port map( A1 => n9722, A2 => n9846, B1 => n8954, B2 => 
                           n9717, ZN => n3380);
   U8590 : OAI22_X1 port map( A1 => n9722, A2 => n9849, B1 => n8939, B2 => 
                           n9717, ZN => n3381);
   U8591 : OAI22_X1 port map( A1 => n9727, A2 => n9782, B1 => n9283, B2 => 
                           n9726, ZN => n3390);
   U8592 : OAI22_X1 port map( A1 => n9727, A2 => n9783, B1 => n9268, B2 => 
                           n9726, ZN => n3391);
   U8593 : OAI22_X1 port map( A1 => n9727, A2 => n9786, B1 => n9253, B2 => 
                           n9726, ZN => n3392);
   U8594 : OAI22_X1 port map( A1 => n9727, A2 => n9789, B1 => n9238, B2 => 
                           n9726, ZN => n3393);
   U8595 : OAI22_X1 port map( A1 => n9727, A2 => n9792, B1 => n9223, B2 => 
                           n9726, ZN => n3394);
   U8596 : OAI22_X1 port map( A1 => n9728, A2 => n9795, B1 => n9208, B2 => 
                           n9726, ZN => n3395);
   U8597 : OAI22_X1 port map( A1 => n9728, A2 => n9798, B1 => n9193, B2 => 
                           n9726, ZN => n3396);
   U8598 : OAI22_X1 port map( A1 => n9728, A2 => n9801, B1 => n9178, B2 => 
                           n9726, ZN => n3397);
   U8599 : OAI22_X1 port map( A1 => n9728, A2 => n9804, B1 => n9163, B2 => 
                           n9726, ZN => n3398);
   U8600 : OAI22_X1 port map( A1 => n9728, A2 => n9807, B1 => n9148, B2 => 
                           n9726, ZN => n3399);
   U8601 : OAI22_X1 port map( A1 => n9729, A2 => n9810, B1 => n9133, B2 => 
                           n9726, ZN => n3400);
   U8602 : OAI22_X1 port map( A1 => n9729, A2 => n9813, B1 => n9118, B2 => 
                           n9726, ZN => n3401);
   U8603 : OAI22_X1 port map( A1 => n9729, A2 => n9816, B1 => n9103, B2 => 
                           n7445, ZN => n3402);
   U8604 : OAI22_X1 port map( A1 => n9729, A2 => n9819, B1 => n9088, B2 => 
                           n7445, ZN => n3403);
   U8605 : OAI22_X1 port map( A1 => n9729, A2 => n9822, B1 => n9073, B2 => 
                           n7445, ZN => n3404);
   U8606 : OAI22_X1 port map( A1 => n9730, A2 => n9825, B1 => n9058, B2 => 
                           n9726, ZN => n3405);
   U8607 : OAI22_X1 port map( A1 => n9730, A2 => n9828, B1 => n9043, B2 => 
                           n9726, ZN => n3406);
   U8608 : OAI22_X1 port map( A1 => n9730, A2 => n9831, B1 => n9028, B2 => 
                           n9726, ZN => n3407);
   U8609 : OAI22_X1 port map( A1 => n9730, A2 => n9834, B1 => n9013, B2 => 
                           n9726, ZN => n3408);
   U8610 : OAI22_X1 port map( A1 => n9730, A2 => n9837, B1 => n8998, B2 => 
                           n9726, ZN => n3409);
   U8611 : OAI22_X1 port map( A1 => n9731, A2 => n9840, B1 => n8983, B2 => 
                           n9726, ZN => n3410);
   U8612 : OAI22_X1 port map( A1 => n9731, A2 => n9843, B1 => n8968, B2 => 
                           n9726, ZN => n3411);
   U8613 : OAI22_X1 port map( A1 => n9731, A2 => n9846, B1 => n8953, B2 => 
                           n9726, ZN => n3412);
   U8614 : OAI22_X1 port map( A1 => n9731, A2 => n9849, B1 => n8938, B2 => 
                           n9726, ZN => n3413);
   U8615 : OAI22_X1 port map( A1 => n9754, A2 => n9782, B1 => n9282, B2 => 
                           n9753, ZN => n3486);
   U8616 : OAI22_X1 port map( A1 => n9754, A2 => n9783, B1 => n9267, B2 => 
                           n9753, ZN => n3487);
   U8617 : OAI22_X1 port map( A1 => n9754, A2 => n9786, B1 => n9252, B2 => 
                           n9753, ZN => n3488);
   U8618 : OAI22_X1 port map( A1 => n9754, A2 => n9789, B1 => n9237, B2 => 
                           n9753, ZN => n3489);
   U8619 : OAI22_X1 port map( A1 => n9754, A2 => n9792, B1 => n9222, B2 => 
                           n9753, ZN => n3490);
   U8620 : OAI22_X1 port map( A1 => n9755, A2 => n9795, B1 => n9207, B2 => 
                           n9753, ZN => n3491);
   U8621 : OAI22_X1 port map( A1 => n9755, A2 => n9798, B1 => n9192, B2 => 
                           n9753, ZN => n3492);
   U8622 : OAI22_X1 port map( A1 => n9755, A2 => n9801, B1 => n9177, B2 => 
                           n9753, ZN => n3493);
   U8623 : OAI22_X1 port map( A1 => n9755, A2 => n9804, B1 => n9162, B2 => 
                           n9753, ZN => n3494);
   U8624 : OAI22_X1 port map( A1 => n9755, A2 => n9807, B1 => n9147, B2 => 
                           n9753, ZN => n3495);
   U8625 : OAI22_X1 port map( A1 => n9756, A2 => n9810, B1 => n9132, B2 => 
                           n9753, ZN => n3496);
   U8626 : OAI22_X1 port map( A1 => n9756, A2 => n9813, B1 => n9117, B2 => 
                           n9753, ZN => n3497);
   U8627 : OAI22_X1 port map( A1 => n9756, A2 => n9816, B1 => n9102, B2 => 
                           n7439, ZN => n3498);
   U8628 : OAI22_X1 port map( A1 => n9756, A2 => n9819, B1 => n9087, B2 => 
                           n7439, ZN => n3499);
   U8629 : OAI22_X1 port map( A1 => n9756, A2 => n9822, B1 => n9072, B2 => 
                           n7439, ZN => n3500);
   U8630 : OAI22_X1 port map( A1 => n9757, A2 => n9825, B1 => n9057, B2 => 
                           n9753, ZN => n3501);
   U8631 : OAI22_X1 port map( A1 => n9757, A2 => n9828, B1 => n9042, B2 => 
                           n9753, ZN => n3502);
   U8632 : OAI22_X1 port map( A1 => n9757, A2 => n9831, B1 => n9027, B2 => 
                           n9753, ZN => n3503);
   U8633 : OAI22_X1 port map( A1 => n9757, A2 => n9834, B1 => n9012, B2 => 
                           n9753, ZN => n3504);
   U8634 : OAI22_X1 port map( A1 => n9757, A2 => n9837, B1 => n8997, B2 => 
                           n9753, ZN => n3505);
   U8635 : OAI22_X1 port map( A1 => n9758, A2 => n9840, B1 => n8982, B2 => 
                           n9753, ZN => n3506);
   U8636 : OAI22_X1 port map( A1 => n9758, A2 => n9843, B1 => n8967, B2 => 
                           n9753, ZN => n3507);
   U8637 : OAI22_X1 port map( A1 => n9758, A2 => n9846, B1 => n8952, B2 => 
                           n9753, ZN => n3508);
   U8638 : OAI22_X1 port map( A1 => n9758, A2 => n9849, B1 => n8937, B2 => 
                           n9753, ZN => n3509);
   U8639 : OAI22_X1 port map( A1 => n9763, A2 => n9782, B1 => n9281, B2 => 
                           n9762, ZN => n3518);
   U8640 : OAI22_X1 port map( A1 => n9763, A2 => n9783, B1 => n9266, B2 => 
                           n9762, ZN => n3519);
   U8641 : OAI22_X1 port map( A1 => n9763, A2 => n9786, B1 => n9251, B2 => 
                           n9762, ZN => n3520);
   U8642 : OAI22_X1 port map( A1 => n9763, A2 => n9789, B1 => n9236, B2 => 
                           n9762, ZN => n3521);
   U8643 : OAI22_X1 port map( A1 => n9763, A2 => n9792, B1 => n9221, B2 => 
                           n9762, ZN => n3522);
   U8644 : OAI22_X1 port map( A1 => n9764, A2 => n9795, B1 => n9206, B2 => 
                           n9762, ZN => n3523);
   U8645 : OAI22_X1 port map( A1 => n9764, A2 => n9798, B1 => n9191, B2 => 
                           n9762, ZN => n3524);
   U8646 : OAI22_X1 port map( A1 => n9764, A2 => n9801, B1 => n9176, B2 => 
                           n9762, ZN => n3525);
   U8647 : OAI22_X1 port map( A1 => n9764, A2 => n9804, B1 => n9161, B2 => 
                           n9762, ZN => n3526);
   U8648 : OAI22_X1 port map( A1 => n9764, A2 => n9807, B1 => n9146, B2 => 
                           n9762, ZN => n3527);
   U8649 : OAI22_X1 port map( A1 => n9765, A2 => n9810, B1 => n9131, B2 => 
                           n9762, ZN => n3528);
   U8650 : OAI22_X1 port map( A1 => n9765, A2 => n9813, B1 => n9116, B2 => 
                           n9762, ZN => n3529);
   U8651 : OAI22_X1 port map( A1 => n9765, A2 => n9816, B1 => n9101, B2 => 
                           n7437, ZN => n3530);
   U8652 : OAI22_X1 port map( A1 => n9765, A2 => n9819, B1 => n9086, B2 => 
                           n7437, ZN => n3531);
   U8653 : OAI22_X1 port map( A1 => n9765, A2 => n9822, B1 => n9071, B2 => 
                           n7437, ZN => n3532);
   U8654 : OAI22_X1 port map( A1 => n9766, A2 => n9825, B1 => n9056, B2 => 
                           n9762, ZN => n3533);
   U8655 : OAI22_X1 port map( A1 => n9766, A2 => n9828, B1 => n9041, B2 => 
                           n9762, ZN => n3534);
   U8656 : OAI22_X1 port map( A1 => n9766, A2 => n9831, B1 => n9026, B2 => 
                           n9762, ZN => n3535);
   U8657 : OAI22_X1 port map( A1 => n9766, A2 => n9834, B1 => n9011, B2 => 
                           n9762, ZN => n3536);
   U8658 : OAI22_X1 port map( A1 => n9766, A2 => n9837, B1 => n8996, B2 => 
                           n9762, ZN => n3537);
   U8659 : OAI22_X1 port map( A1 => n9767, A2 => n9840, B1 => n8981, B2 => 
                           n9762, ZN => n3538);
   U8660 : OAI22_X1 port map( A1 => n9767, A2 => n9843, B1 => n8966, B2 => 
                           n9762, ZN => n3539);
   U8661 : OAI22_X1 port map( A1 => n9767, A2 => n9846, B1 => n8951, B2 => 
                           n9762, ZN => n3540);
   U8662 : OAI22_X1 port map( A1 => n9767, A2 => n9849, B1 => n8936, B2 => 
                           n9762, ZN => n3541);
   U8663 : OAI22_X1 port map( A1 => n9772, A2 => n9782, B1 => n64, B2 => n7435,
                           ZN => n3550);
   U8664 : OAI22_X1 port map( A1 => n9772, A2 => n9783, B1 => n63, B2 => n7435,
                           ZN => n3551);
   U8665 : OAI22_X1 port map( A1 => n9772, A2 => n9786, B1 => n62, B2 => n7435,
                           ZN => n3552);
   U8666 : OAI22_X1 port map( A1 => n9772, A2 => n9789, B1 => n61, B2 => n9771,
                           ZN => n3553);
   U8667 : OAI22_X1 port map( A1 => n9772, A2 => n9792, B1 => n60, B2 => n9771,
                           ZN => n3554);
   U8668 : OAI22_X1 port map( A1 => n9773, A2 => n9795, B1 => n59, B2 => n9771,
                           ZN => n3555);
   U8669 : OAI22_X1 port map( A1 => n9773, A2 => n9798, B1 => n58, B2 => n9771,
                           ZN => n3556);
   U8670 : OAI22_X1 port map( A1 => n9773, A2 => n9801, B1 => n57, B2 => n9771,
                           ZN => n3557);
   U8671 : OAI22_X1 port map( A1 => n9773, A2 => n9804, B1 => n56, B2 => n9771,
                           ZN => n3558);
   U8672 : OAI22_X1 port map( A1 => n9773, A2 => n9807, B1 => n55, B2 => n9771,
                           ZN => n3559);
   U8673 : OAI22_X1 port map( A1 => n9774, A2 => n9810, B1 => n54, B2 => n9771,
                           ZN => n3560);
   U8674 : OAI22_X1 port map( A1 => n9774, A2 => n9813, B1 => n53, B2 => n9771,
                           ZN => n3561);
   U8675 : OAI22_X1 port map( A1 => n9774, A2 => n9816, B1 => n52, B2 => n9771,
                           ZN => n3562);
   U8676 : OAI22_X1 port map( A1 => n9774, A2 => n9819, B1 => n51, B2 => n9771,
                           ZN => n3563);
   U8677 : OAI22_X1 port map( A1 => n9774, A2 => n9822, B1 => n50, B2 => n9771,
                           ZN => n3564);
   U8678 : OAI22_X1 port map( A1 => n9775, A2 => n9825, B1 => n49, B2 => n9771,
                           ZN => n3565);
   U8679 : OAI22_X1 port map( A1 => n9775, A2 => n9828, B1 => n48, B2 => n9771,
                           ZN => n3566);
   U8680 : OAI22_X1 port map( A1 => n9775, A2 => n9831, B1 => n47, B2 => n9771,
                           ZN => n3567);
   U8681 : OAI22_X1 port map( A1 => n9775, A2 => n9834, B1 => n46, B2 => n9771,
                           ZN => n3568);
   U8682 : OAI22_X1 port map( A1 => n9775, A2 => n9837, B1 => n45, B2 => n9771,
                           ZN => n3569);
   U8683 : OAI22_X1 port map( A1 => n9878, A2 => n9849, B1 => n9, B2 => n9873, 
                           ZN => n3605);
   U8684 : OAI22_X1 port map( A1 => n9878, A2 => n9852, B1 => n8, B2 => n9873, 
                           ZN => n3606);
   U8685 : OAI22_X1 port map( A1 => n9879, A2 => n9855, B1 => n7, B2 => n9873, 
                           ZN => n3607);
   U8686 : OAI22_X1 port map( A1 => n9879, A2 => n9858, B1 => n6, B2 => n9873, 
                           ZN => n3608);
   U8687 : OAI22_X1 port map( A1 => n9879, A2 => n9861, B1 => n5, B2 => n9873, 
                           ZN => n3609);
   U8688 : OAI21_X1 port map( B1 => n9280, B2 => n9393, A => n8752, ZN => n2526
                           );
   U8689 : OAI21_X1 port map( B1 => n8753, B2 => n8754, A => n9396, ZN => n8752
                           );
   U8690 : NAND4_X1 port map( A1 => n8771, A2 => n8772, A3 => n8773, A4 => 
                           n8774, ZN => n8753);
   U8691 : NAND4_X1 port map( A1 => n8755, A2 => n8756, A3 => n8757, A4 => 
                           n8758, ZN => n8754);
   U8692 : OAI21_X1 port map( B1 => n9265, B2 => n9393, A => n8733, ZN => n2527
                           );
   U8693 : OAI21_X1 port map( B1 => n8734, B2 => n8735, A => n9396, ZN => n8733
                           );
   U8694 : NAND4_X1 port map( A1 => n8744, A2 => n8745, A3 => n8746, A4 => 
                           n8747, ZN => n8734);
   U8695 : NAND4_X1 port map( A1 => n8736, A2 => n8737, A3 => n8738, A4 => 
                           n8739, ZN => n8735);
   U8696 : OAI21_X1 port map( B1 => n9250, B2 => n9393, A => n8714, ZN => n2528
                           );
   U8697 : OAI21_X1 port map( B1 => n8715, B2 => n8716, A => n9395, ZN => n8714
                           );
   U8698 : NAND4_X1 port map( A1 => n8725, A2 => n8726, A3 => n8727, A4 => 
                           n8728, ZN => n8715);
   U8699 : NAND4_X1 port map( A1 => n8717, A2 => n8718, A3 => n8719, A4 => 
                           n8720, ZN => n8716);
   U8700 : OAI21_X1 port map( B1 => n9235, B2 => n9393, A => n8695, ZN => n2529
                           );
   U8701 : OAI21_X1 port map( B1 => n8696, B2 => n8697, A => n9395, ZN => n8695
                           );
   U8702 : NAND4_X1 port map( A1 => n8706, A2 => n8707, A3 => n8708, A4 => 
                           n8709, ZN => n8696);
   U8703 : NAND4_X1 port map( A1 => n8698, A2 => n8699, A3 => n8700, A4 => 
                           n8701, ZN => n8697);
   U8704 : OAI21_X1 port map( B1 => n9220, B2 => n9393, A => n8676, ZN => n2530
                           );
   U8705 : OAI21_X1 port map( B1 => n8677, B2 => n8678, A => n9395, ZN => n8676
                           );
   U8706 : NAND4_X1 port map( A1 => n8687, A2 => n8688, A3 => n8689, A4 => 
                           n8690, ZN => n8677);
   U8707 : NAND4_X1 port map( A1 => n8679, A2 => n8680, A3 => n8681, A4 => 
                           n8682, ZN => n8678);
   U8708 : OAI21_X1 port map( B1 => n9205, B2 => n9393, A => n8657, ZN => n2531
                           );
   U8709 : OAI21_X1 port map( B1 => n8658, B2 => n8659, A => n9394, ZN => n8657
                           );
   U8710 : NAND4_X1 port map( A1 => n8668, A2 => n8669, A3 => n8670, A4 => 
                           n8671, ZN => n8658);
   U8711 : NAND4_X1 port map( A1 => n8660, A2 => n8661, A3 => n8662, A4 => 
                           n8663, ZN => n8659);
   U8712 : OAI21_X1 port map( B1 => n9190, B2 => n9393, A => n8638, ZN => n2532
                           );
   U8713 : OAI21_X1 port map( B1 => n8639, B2 => n8640, A => n9395, ZN => n8638
                           );
   U8714 : NAND4_X1 port map( A1 => n8649, A2 => n8650, A3 => n8651, A4 => 
                           n8652, ZN => n8639);
   U8715 : NAND4_X1 port map( A1 => n8641, A2 => n8642, A3 => n8643, A4 => 
                           n8644, ZN => n8640);
   U8716 : OAI21_X1 port map( B1 => n9160, B2 => n9393, A => n8600, ZN => n2534
                           );
   U8717 : OAI21_X1 port map( B1 => n8601, B2 => n8602, A => n9394, ZN => n8600
                           );
   U8718 : NAND4_X1 port map( A1 => n8611, A2 => n8612, A3 => n8613, A4 => 
                           n8614, ZN => n8601);
   U8719 : NAND4_X1 port map( A1 => n8603, A2 => n8604, A3 => n8605, A4 => 
                           n8606, ZN => n8602);
   U8720 : OAI21_X1 port map( B1 => n8814, B2 => n9495, A => n8099, ZN => n2558
                           );
   U8721 : OAI21_X1 port map( B1 => n8100, B2 => n8101, A => n9498, ZN => n8099
                           );
   U8722 : NAND4_X1 port map( A1 => n8118, A2 => n8119, A3 => n8120, A4 => 
                           n8121, ZN => n8100);
   U8723 : NAND4_X1 port map( A1 => n8102, A2 => n8103, A3 => n8104, A4 => 
                           n8105, ZN => n8101);
   U8724 : OAI21_X1 port map( B1 => n8813, B2 => n9495, A => n8080, ZN => n2559
                           );
   U8725 : OAI21_X1 port map( B1 => n8081, B2 => n8082, A => n9498, ZN => n8080
                           );
   U8726 : NAND4_X1 port map( A1 => n8091, A2 => n8092, A3 => n8093, A4 => 
                           n8094, ZN => n8081);
   U8727 : NAND4_X1 port map( A1 => n8083, A2 => n8084, A3 => n8085, A4 => 
                           n8086, ZN => n8082);
   U8728 : OAI21_X1 port map( B1 => n8812, B2 => n9495, A => n8061, ZN => n2560
                           );
   U8729 : OAI21_X1 port map( B1 => n8062, B2 => n8063, A => n9497, ZN => n8061
                           );
   U8730 : NAND4_X1 port map( A1 => n8072, A2 => n8073, A3 => n8074, A4 => 
                           n8075, ZN => n8062);
   U8731 : NAND4_X1 port map( A1 => n8064, A2 => n8065, A3 => n8066, A4 => 
                           n8067, ZN => n8063);
   U8732 : OAI21_X1 port map( B1 => n8811, B2 => n9495, A => n8042, ZN => n2561
                           );
   U8733 : OAI21_X1 port map( B1 => n8043, B2 => n8044, A => n9497, ZN => n8042
                           );
   U8734 : NAND4_X1 port map( A1 => n8053, A2 => n8054, A3 => n8055, A4 => 
                           n8056, ZN => n8043);
   U8735 : NAND4_X1 port map( A1 => n8045, A2 => n8046, A3 => n8047, A4 => 
                           n8048, ZN => n8044);
   U8736 : OAI21_X1 port map( B1 => n8810, B2 => n9495, A => n8023, ZN => n2562
                           );
   U8737 : OAI21_X1 port map( B1 => n8024, B2 => n8025, A => n9497, ZN => n8023
                           );
   U8738 : NAND4_X1 port map( A1 => n8034, A2 => n8035, A3 => n8036, A4 => 
                           n8037, ZN => n8024);
   U8739 : NAND4_X1 port map( A1 => n8026, A2 => n8027, A3 => n8028, A4 => 
                           n8029, ZN => n8025);
   U8740 : OAI21_X1 port map( B1 => n8809, B2 => n9495, A => n8004, ZN => n2563
                           );
   U8741 : OAI21_X1 port map( B1 => n8005, B2 => n8006, A => n9496, ZN => n8004
                           );
   U8742 : NAND4_X1 port map( A1 => n8015, A2 => n8016, A3 => n8017, A4 => 
                           n8018, ZN => n8005);
   U8743 : NAND4_X1 port map( A1 => n8007, A2 => n8008, A3 => n8009, A4 => 
                           n8010, ZN => n8006);
   U8744 : OAI21_X1 port map( B1 => n8808, B2 => n9495, A => n7985, ZN => n2564
                           );
   U8745 : OAI21_X1 port map( B1 => n7986, B2 => n7987, A => n9497, ZN => n7985
                           );
   U8746 : NAND4_X1 port map( A1 => n7996, A2 => n7997, A3 => n7998, A4 => 
                           n7999, ZN => n7986);
   U8747 : NAND4_X1 port map( A1 => n7988, A2 => n7989, A3 => n7990, A4 => 
                           n7991, ZN => n7987);
   U8748 : OAI21_X1 port map( B1 => n8806, B2 => n9495, A => n7947, ZN => n2566
                           );
   U8749 : OAI21_X1 port map( B1 => n7948, B2 => n7949, A => n9496, ZN => n7947
                           );
   U8750 : NAND4_X1 port map( A1 => n7958, A2 => n7959, A3 => n7960, A4 => 
                           n7961, ZN => n7948);
   U8751 : NAND4_X1 port map( A1 => n7950, A2 => n7951, A3 => n7952, A4 => 
                           n7953, ZN => n7949);
   U8752 : OAI21_X1 port map( B1 => n9175, B2 => n9392, A => n8619, ZN => n2533
                           );
   U8753 : OAI21_X1 port map( B1 => n8620, B2 => n8621, A => n9394, ZN => n8619
                           );
   U8754 : NAND4_X1 port map( A1 => n8630, A2 => n8631, A3 => n8632, A4 => 
                           n8633, ZN => n8620);
   U8755 : NAND4_X1 port map( A1 => n8622, A2 => n8623, A3 => n8624, A4 => 
                           n8625, ZN => n8621);
   U8756 : OAI21_X1 port map( B1 => n9145, B2 => n9392, A => n8581, ZN => n2535
                           );
   U8757 : OAI21_X1 port map( B1 => n8582, B2 => n8583, A => n9394, ZN => n8581
                           );
   U8758 : NAND4_X1 port map( A1 => n8592, A2 => n8593, A3 => n8594, A4 => 
                           n8595, ZN => n8582);
   U8759 : NAND4_X1 port map( A1 => n8584, A2 => n8585, A3 => n8586, A4 => 
                           n8587, ZN => n8583);
   U8760 : OAI21_X1 port map( B1 => n9130, B2 => n9392, A => n8562, ZN => n2536
                           );
   U8761 : OAI21_X1 port map( B1 => n8563, B2 => n8564, A => n9393, ZN => n8562
                           );
   U8762 : NAND4_X1 port map( A1 => n8573, A2 => n8574, A3 => n8575, A4 => 
                           n8576, ZN => n8563);
   U8763 : NAND4_X1 port map( A1 => n8565, A2 => n8566, A3 => n8567, A4 => 
                           n8568, ZN => n8564);
   U8764 : OAI21_X1 port map( B1 => n9115, B2 => n9392, A => n8543, ZN => n2537
                           );
   U8765 : OAI21_X1 port map( B1 => n8544, B2 => n8545, A => n9393, ZN => n8543
                           );
   U8766 : NAND4_X1 port map( A1 => n8554, A2 => n8555, A3 => n8556, A4 => 
                           n8557, ZN => n8544);
   U8767 : NAND4_X1 port map( A1 => n8546, A2 => n8547, A3 => n8548, A4 => 
                           n8549, ZN => n8545);
   U8768 : OAI21_X1 port map( B1 => n9100, B2 => n9392, A => n8524, ZN => n2538
                           );
   U8769 : OAI21_X1 port map( B1 => n8525, B2 => n8526, A => n9394, ZN => n8524
                           );
   U8770 : NAND4_X1 port map( A1 => n8535, A2 => n8536, A3 => n8537, A4 => 
                           n8538, ZN => n8525);
   U8771 : NAND4_X1 port map( A1 => n8527, A2 => n8528, A3 => n8529, A4 => 
                           n8530, ZN => n8526);
   U8772 : OAI21_X1 port map( B1 => n9085, B2 => n9392, A => n8505, ZN => n2539
                           );
   U8773 : OAI21_X1 port map( B1 => n8506, B2 => n8507, A => n9393, ZN => n8505
                           );
   U8774 : NAND4_X1 port map( A1 => n8516, A2 => n8517, A3 => n8518, A4 => 
                           n8519, ZN => n8506);
   U8775 : NAND4_X1 port map( A1 => n8508, A2 => n8509, A3 => n8510, A4 => 
                           n8511, ZN => n8507);
   U8776 : OAI21_X1 port map( B1 => n9070, B2 => n9392, A => n8486, ZN => n2540
                           );
   U8777 : OAI21_X1 port map( B1 => n8487, B2 => n8488, A => n9393, ZN => n8486
                           );
   U8778 : NAND4_X1 port map( A1 => n8497, A2 => n8498, A3 => n8499, A4 => 
                           n8500, ZN => n8487);
   U8779 : NAND4_X1 port map( A1 => n8489, A2 => n8490, A3 => n8491, A4 => 
                           n8492, ZN => n8488);
   U8780 : OAI21_X1 port map( B1 => n9055, B2 => n9392, A => n8467, ZN => n2541
                           );
   U8781 : OAI21_X1 port map( B1 => n8468, B2 => n8469, A => n9394, ZN => n8467
                           );
   U8782 : NAND4_X1 port map( A1 => n8478, A2 => n8479, A3 => n8480, A4 => 
                           n8481, ZN => n8468);
   U8783 : NAND4_X1 port map( A1 => n8470, A2 => n8471, A3 => n8472, A4 => 
                           n8473, ZN => n8469);
   U8784 : OAI21_X1 port map( B1 => n9040, B2 => n9392, A => n8448, ZN => n2542
                           );
   U8785 : OAI21_X1 port map( B1 => n8449, B2 => n8450, A => n9394, ZN => n8448
                           );
   U8786 : NAND4_X1 port map( A1 => n8459, A2 => n8460, A3 => n8461, A4 => 
                           n8462, ZN => n8449);
   U8787 : NAND4_X1 port map( A1 => n8451, A2 => n8452, A3 => n8453, A4 => 
                           n8454, ZN => n8450);
   U8788 : OAI21_X1 port map( B1 => n9025, B2 => n9392, A => n8429, ZN => n2543
                           );
   U8789 : OAI21_X1 port map( B1 => n8430, B2 => n8431, A => n9394, ZN => n8429
                           );
   U8790 : NAND4_X1 port map( A1 => n8440, A2 => n8441, A3 => n8442, A4 => 
                           n8443, ZN => n8430);
   U8791 : NAND4_X1 port map( A1 => n8432, A2 => n8433, A3 => n8434, A4 => 
                           n8435, ZN => n8431);
   U8792 : OAI21_X1 port map( B1 => n9010, B2 => n9392, A => n8410, ZN => n2544
                           );
   U8793 : OAI21_X1 port map( B1 => n8411, B2 => n8412, A => n9394, ZN => n8410
                           );
   U8794 : NAND4_X1 port map( A1 => n8421, A2 => n8422, A3 => n8423, A4 => 
                           n8424, ZN => n8411);
   U8795 : NAND4_X1 port map( A1 => n8413, A2 => n8414, A3 => n8415, A4 => 
                           n8416, ZN => n8412);
   U8796 : OAI21_X1 port map( B1 => n8995, B2 => n9391, A => n8391, ZN => n2545
                           );
   U8797 : OAI21_X1 port map( B1 => n8392, B2 => n8393, A => n9394, ZN => n8391
                           );
   U8798 : NAND4_X1 port map( A1 => n8402, A2 => n8403, A3 => n8404, A4 => 
                           n8405, ZN => n8392);
   U8799 : NAND4_X1 port map( A1 => n8394, A2 => n8395, A3 => n8396, A4 => 
                           n8397, ZN => n8393);
   U8800 : OAI21_X1 port map( B1 => n8980, B2 => n9391, A => n8372, ZN => n2546
                           );
   U8801 : OAI21_X1 port map( B1 => n8373, B2 => n8374, A => n9394, ZN => n8372
                           );
   U8802 : NAND4_X1 port map( A1 => n8383, A2 => n8384, A3 => n8385, A4 => 
                           n8386, ZN => n8373);
   U8803 : NAND4_X1 port map( A1 => n8375, A2 => n8376, A3 => n8377, A4 => 
                           n8378, ZN => n8374);
   U8804 : OAI21_X1 port map( B1 => n8965, B2 => n9391, A => n8353, ZN => n2547
                           );
   U8805 : OAI21_X1 port map( B1 => n8354, B2 => n8355, A => n9395, ZN => n8353
                           );
   U8806 : NAND4_X1 port map( A1 => n8364, A2 => n8365, A3 => n8366, A4 => 
                           n8367, ZN => n8354);
   U8807 : NAND4_X1 port map( A1 => n8356, A2 => n8357, A3 => n8358, A4 => 
                           n8359, ZN => n8355);
   U8808 : OAI21_X1 port map( B1 => n8950, B2 => n9391, A => n8334, ZN => n2548
                           );
   U8809 : OAI21_X1 port map( B1 => n8335, B2 => n8336, A => n9394, ZN => n8334
                           );
   U8810 : NAND4_X1 port map( A1 => n8345, A2 => n8346, A3 => n8347, A4 => 
                           n8348, ZN => n8335);
   U8811 : NAND4_X1 port map( A1 => n8337, A2 => n8338, A3 => n8339, A4 => 
                           n8340, ZN => n8336);
   U8812 : OAI21_X1 port map( B1 => n8935, B2 => n9391, A => n8315, ZN => n2549
                           );
   U8813 : OAI21_X1 port map( B1 => n8316, B2 => n8317, A => n9395, ZN => n8315
                           );
   U8814 : NAND4_X1 port map( A1 => n8326, A2 => n8327, A3 => n8328, A4 => 
                           n8329, ZN => n8316);
   U8815 : NAND4_X1 port map( A1 => n8318, A2 => n8319, A3 => n8320, A4 => 
                           n8321, ZN => n8317);
   U8816 : OAI21_X1 port map( B1 => n8920, B2 => n9391, A => n8296, ZN => n2550
                           );
   U8817 : OAI21_X1 port map( B1 => n8297, B2 => n8298, A => n9395, ZN => n8296
                           );
   U8818 : NAND4_X1 port map( A1 => n8307, A2 => n8308, A3 => n8309, A4 => 
                           n8310, ZN => n8297);
   U8819 : NAND4_X1 port map( A1 => n8299, A2 => n8300, A3 => n8301, A4 => 
                           n8302, ZN => n8298);
   U8820 : OAI21_X1 port map( B1 => n8905, B2 => n9391, A => n8277, ZN => n2551
                           );
   U8821 : OAI21_X1 port map( B1 => n8278, B2 => n8279, A => n9395, ZN => n8277
                           );
   U8822 : NAND4_X1 port map( A1 => n8288, A2 => n8289, A3 => n8290, A4 => 
                           n8291, ZN => n8278);
   U8823 : NAND4_X1 port map( A1 => n8280, A2 => n8281, A3 => n8282, A4 => 
                           n8283, ZN => n8279);
   U8824 : OAI21_X1 port map( B1 => n8890, B2 => n9391, A => n8258, ZN => n2552
                           );
   U8825 : OAI21_X1 port map( B1 => n8259, B2 => n8260, A => n9395, ZN => n8258
                           );
   U8826 : NAND4_X1 port map( A1 => n8269, A2 => n8270, A3 => n8271, A4 => 
                           n8272, ZN => n8259);
   U8827 : NAND4_X1 port map( A1 => n8261, A2 => n8262, A3 => n8263, A4 => 
                           n8264, ZN => n8260);
   U8828 : OAI21_X1 port map( B1 => n8875, B2 => n9391, A => n8239, ZN => n2553
                           );
   U8829 : OAI21_X1 port map( B1 => n8240, B2 => n8241, A => n9395, ZN => n8239
                           );
   U8830 : NAND4_X1 port map( A1 => n8250, A2 => n8251, A3 => n8252, A4 => 
                           n8253, ZN => n8240);
   U8831 : NAND4_X1 port map( A1 => n8242, A2 => n8243, A3 => n8244, A4 => 
                           n8245, ZN => n8241);
   U8832 : OAI21_X1 port map( B1 => n8860, B2 => n9391, A => n8220, ZN => n2554
                           );
   U8833 : OAI21_X1 port map( B1 => n8221, B2 => n8222, A => n9395, ZN => n8220
                           );
   U8834 : NAND4_X1 port map( A1 => n8231, A2 => n8232, A3 => n8233, A4 => 
                           n8234, ZN => n8221);
   U8835 : NAND4_X1 port map( A1 => n8223, A2 => n8224, A3 => n8225, A4 => 
                           n8226, ZN => n8222);
   U8836 : OAI21_X1 port map( B1 => n8845, B2 => n9391, A => n8201, ZN => n2555
                           );
   U8837 : OAI21_X1 port map( B1 => n8202, B2 => n8203, A => n9395, ZN => n8201
                           );
   U8838 : NAND4_X1 port map( A1 => n8212, A2 => n8213, A3 => n8214, A4 => 
                           n8215, ZN => n8202);
   U8839 : NAND4_X1 port map( A1 => n8204, A2 => n8205, A3 => n8206, A4 => 
                           n8207, ZN => n8203);
   U8840 : OAI21_X1 port map( B1 => n8830, B2 => n9391, A => n8182, ZN => n2556
                           );
   U8841 : OAI21_X1 port map( B1 => n8183, B2 => n8184, A => n9396, ZN => n8182
                           );
   U8842 : NAND4_X1 port map( A1 => n8193, A2 => n8194, A3 => n8195, A4 => 
                           n8196, ZN => n8183);
   U8843 : NAND4_X1 port map( A1 => n8185, A2 => n8186, A3 => n8187, A4 => 
                           n8188, ZN => n8184);
   U8844 : OAI21_X1 port map( B1 => n8815, B2 => n9392, A => n8131, ZN => n2557
                           );
   U8845 : OAI21_X1 port map( B1 => n8132, B2 => n8133, A => n9396, ZN => n8131
                           );
   U8846 : NAND4_X1 port map( A1 => n8158, A2 => n8159, A3 => n8160, A4 => 
                           n8161, ZN => n8132);
   U8847 : NAND4_X1 port map( A1 => n8134, A2 => n8135, A3 => n8136, A4 => 
                           n8137, ZN => n8133);
   U8848 : OAI21_X1 port map( B1 => n8807, B2 => n9494, A => n7966, ZN => n2565
                           );
   U8849 : OAI21_X1 port map( B1 => n7967, B2 => n7968, A => n9496, ZN => n7966
                           );
   U8850 : NAND4_X1 port map( A1 => n7977, A2 => n7978, A3 => n7979, A4 => 
                           n7980, ZN => n7967);
   U8851 : NAND4_X1 port map( A1 => n7969, A2 => n7970, A3 => n7971, A4 => 
                           n7972, ZN => n7968);
   U8852 : OAI21_X1 port map( B1 => n8805, B2 => n9494, A => n7928, ZN => n2567
                           );
   U8853 : OAI21_X1 port map( B1 => n7929, B2 => n7930, A => n9496, ZN => n7928
                           );
   U8854 : NAND4_X1 port map( A1 => n7939, A2 => n7940, A3 => n7941, A4 => 
                           n7942, ZN => n7929);
   U8855 : NAND4_X1 port map( A1 => n7931, A2 => n7932, A3 => n7933, A4 => 
                           n7934, ZN => n7930);
   U8856 : OAI21_X1 port map( B1 => n8804, B2 => n9494, A => n7909, ZN => n2568
                           );
   U8857 : OAI21_X1 port map( B1 => n7910, B2 => n7911, A => n9495, ZN => n7909
                           );
   U8858 : NAND4_X1 port map( A1 => n7920, A2 => n7921, A3 => n7922, A4 => 
                           n7923, ZN => n7910);
   U8859 : NAND4_X1 port map( A1 => n7912, A2 => n7913, A3 => n7914, A4 => 
                           n7915, ZN => n7911);
   U8860 : OAI21_X1 port map( B1 => n8803, B2 => n9494, A => n7890, ZN => n2569
                           );
   U8861 : OAI21_X1 port map( B1 => n7891, B2 => n7892, A => n9495, ZN => n7890
                           );
   U8862 : NAND4_X1 port map( A1 => n7901, A2 => n7902, A3 => n7903, A4 => 
                           n7904, ZN => n7891);
   U8863 : NAND4_X1 port map( A1 => n7893, A2 => n7894, A3 => n7895, A4 => 
                           n7896, ZN => n7892);
   U8864 : OAI21_X1 port map( B1 => n8802, B2 => n9494, A => n7871, ZN => n2570
                           );
   U8865 : OAI21_X1 port map( B1 => n7872, B2 => n7873, A => n9496, ZN => n7871
                           );
   U8866 : NAND4_X1 port map( A1 => n7882, A2 => n7883, A3 => n7884, A4 => 
                           n7885, ZN => n7872);
   U8867 : NAND4_X1 port map( A1 => n7874, A2 => n7875, A3 => n7876, A4 => 
                           n7877, ZN => n7873);
   U8868 : OAI21_X1 port map( B1 => n8801, B2 => n9494, A => n7852, ZN => n2571
                           );
   U8869 : OAI21_X1 port map( B1 => n7853, B2 => n7854, A => n9495, ZN => n7852
                           );
   U8870 : NAND4_X1 port map( A1 => n7863, A2 => n7864, A3 => n7865, A4 => 
                           n7866, ZN => n7853);
   U8871 : NAND4_X1 port map( A1 => n7855, A2 => n7856, A3 => n7857, A4 => 
                           n7858, ZN => n7854);
   U8872 : OAI21_X1 port map( B1 => n8800, B2 => n9494, A => n7833, ZN => n2572
                           );
   U8873 : OAI21_X1 port map( B1 => n7834, B2 => n7835, A => n9495, ZN => n7833
                           );
   U8874 : NAND4_X1 port map( A1 => n7844, A2 => n7845, A3 => n7846, A4 => 
                           n7847, ZN => n7834);
   U8875 : NAND4_X1 port map( A1 => n7836, A2 => n7837, A3 => n7838, A4 => 
                           n7839, ZN => n7835);
   U8876 : OAI21_X1 port map( B1 => n8799, B2 => n9494, A => n7814, ZN => n2573
                           );
   U8877 : OAI21_X1 port map( B1 => n7815, B2 => n7816, A => n9496, ZN => n7814
                           );
   U8878 : NAND4_X1 port map( A1 => n7825, A2 => n7826, A3 => n7827, A4 => 
                           n7828, ZN => n7815);
   U8879 : NAND4_X1 port map( A1 => n7817, A2 => n7818, A3 => n7819, A4 => 
                           n7820, ZN => n7816);
   U8880 : OAI21_X1 port map( B1 => n8798, B2 => n9494, A => n7795, ZN => n2574
                           );
   U8881 : OAI21_X1 port map( B1 => n7796, B2 => n7797, A => n9496, ZN => n7795
                           );
   U8882 : NAND4_X1 port map( A1 => n7806, A2 => n7807, A3 => n7808, A4 => 
                           n7809, ZN => n7796);
   U8883 : NAND4_X1 port map( A1 => n7798, A2 => n7799, A3 => n7800, A4 => 
                           n7801, ZN => n7797);
   U8884 : OAI21_X1 port map( B1 => n8797, B2 => n9494, A => n7776, ZN => n2575
                           );
   U8885 : OAI21_X1 port map( B1 => n7777, B2 => n7778, A => n9496, ZN => n7776
                           );
   U8886 : NAND4_X1 port map( A1 => n7787, A2 => n7788, A3 => n7789, A4 => 
                           n7790, ZN => n7777);
   U8887 : NAND4_X1 port map( A1 => n7779, A2 => n7780, A3 => n7781, A4 => 
                           n7782, ZN => n7778);
   U8888 : OAI21_X1 port map( B1 => n8796, B2 => n9494, A => n7757, ZN => n2576
                           );
   U8889 : OAI21_X1 port map( B1 => n7758, B2 => n7759, A => n9496, ZN => n7757
                           );
   U8890 : NAND4_X1 port map( A1 => n7768, A2 => n7769, A3 => n7770, A4 => 
                           n7771, ZN => n7758);
   U8891 : NAND4_X1 port map( A1 => n7760, A2 => n7761, A3 => n7762, A4 => 
                           n7763, ZN => n7759);
   U8892 : OAI21_X1 port map( B1 => n8795, B2 => n9493, A => n7738, ZN => n2577
                           );
   U8893 : OAI21_X1 port map( B1 => n7739, B2 => n7740, A => n9496, ZN => n7738
                           );
   U8894 : NAND4_X1 port map( A1 => n7749, A2 => n7750, A3 => n7751, A4 => 
                           n7752, ZN => n7739);
   U8895 : NAND4_X1 port map( A1 => n7741, A2 => n7742, A3 => n7743, A4 => 
                           n7744, ZN => n7740);
   U8896 : OAI21_X1 port map( B1 => n8794, B2 => n9493, A => n7719, ZN => n2578
                           );
   U8897 : OAI21_X1 port map( B1 => n7720, B2 => n7721, A => n9496, ZN => n7719
                           );
   U8898 : NAND4_X1 port map( A1 => n7730, A2 => n7731, A3 => n7732, A4 => 
                           n7733, ZN => n7720);
   U8899 : NAND4_X1 port map( A1 => n7722, A2 => n7723, A3 => n7724, A4 => 
                           n7725, ZN => n7721);
   U8900 : OAI21_X1 port map( B1 => n8793, B2 => n9493, A => n7700, ZN => n2579
                           );
   U8901 : OAI21_X1 port map( B1 => n7701, B2 => n7702, A => n9497, ZN => n7700
                           );
   U8902 : NAND4_X1 port map( A1 => n7711, A2 => n7712, A3 => n7713, A4 => 
                           n7714, ZN => n7701);
   U8903 : NAND4_X1 port map( A1 => n7703, A2 => n7704, A3 => n7705, A4 => 
                           n7706, ZN => n7702);
   U8904 : OAI21_X1 port map( B1 => n8792, B2 => n9493, A => n7681, ZN => n2580
                           );
   U8905 : OAI21_X1 port map( B1 => n7682, B2 => n7683, A => n9496, ZN => n7681
                           );
   U8906 : NAND4_X1 port map( A1 => n7692, A2 => n7693, A3 => n7694, A4 => 
                           n7695, ZN => n7682);
   U8907 : NAND4_X1 port map( A1 => n7684, A2 => n7685, A3 => n7686, A4 => 
                           n7687, ZN => n7683);
   U8908 : OAI21_X1 port map( B1 => n8791, B2 => n9493, A => n7662, ZN => n2581
                           );
   U8909 : OAI21_X1 port map( B1 => n7663, B2 => n7664, A => n9497, ZN => n7662
                           );
   U8910 : NAND4_X1 port map( A1 => n7673, A2 => n7674, A3 => n7675, A4 => 
                           n7676, ZN => n7663);
   U8911 : NAND4_X1 port map( A1 => n7665, A2 => n7666, A3 => n7667, A4 => 
                           n7668, ZN => n7664);
   U8912 : OAI21_X1 port map( B1 => n8790, B2 => n9493, A => n7643, ZN => n2582
                           );
   U8913 : OAI21_X1 port map( B1 => n7644, B2 => n7645, A => n9497, ZN => n7643
                           );
   U8914 : NAND4_X1 port map( A1 => n7654, A2 => n7655, A3 => n7656, A4 => 
                           n7657, ZN => n7644);
   U8915 : NAND4_X1 port map( A1 => n7646, A2 => n7647, A3 => n7648, A4 => 
                           n7649, ZN => n7645);
   U8916 : OAI21_X1 port map( B1 => n8789, B2 => n9493, A => n7624, ZN => n2583
                           );
   U8917 : OAI21_X1 port map( B1 => n7625, B2 => n7626, A => n9497, ZN => n7624
                           );
   U8918 : NAND4_X1 port map( A1 => n7635, A2 => n7636, A3 => n7637, A4 => 
                           n7638, ZN => n7625);
   U8919 : NAND4_X1 port map( A1 => n7627, A2 => n7628, A3 => n7629, A4 => 
                           n7630, ZN => n7626);
   U8920 : OAI21_X1 port map( B1 => n8788, B2 => n9493, A => n7605, ZN => n2584
                           );
   U8921 : OAI21_X1 port map( B1 => n7606, B2 => n7607, A => n9497, ZN => n7605
                           );
   U8922 : NAND4_X1 port map( A1 => n7616, A2 => n7617, A3 => n7618, A4 => 
                           n7619, ZN => n7606);
   U8923 : NAND4_X1 port map( A1 => n7608, A2 => n7609, A3 => n7610, A4 => 
                           n7611, ZN => n7607);
   U8924 : OAI21_X1 port map( B1 => n8787, B2 => n9493, A => n7586, ZN => n2585
                           );
   U8925 : OAI21_X1 port map( B1 => n7587, B2 => n7588, A => n9497, ZN => n7586
                           );
   U8926 : NAND4_X1 port map( A1 => n7597, A2 => n7598, A3 => n7599, A4 => 
                           n7600, ZN => n7587);
   U8927 : NAND4_X1 port map( A1 => n7589, A2 => n7590, A3 => n7591, A4 => 
                           n7592, ZN => n7588);
   U8928 : OAI21_X1 port map( B1 => n8786, B2 => n9493, A => n7567, ZN => n2586
                           );
   U8929 : OAI21_X1 port map( B1 => n7568, B2 => n7569, A => n9497, ZN => n7567
                           );
   U8930 : NAND4_X1 port map( A1 => n7578, A2 => n7579, A3 => n7580, A4 => 
                           n7581, ZN => n7568);
   U8931 : NAND4_X1 port map( A1 => n7570, A2 => n7571, A3 => n7572, A4 => 
                           n7573, ZN => n7569);
   U8932 : OAI21_X1 port map( B1 => n8785, B2 => n9493, A => n7548, ZN => n2587
                           );
   U8933 : OAI21_X1 port map( B1 => n7549, B2 => n7550, A => n9497, ZN => n7548
                           );
   U8934 : NAND4_X1 port map( A1 => n7559, A2 => n7560, A3 => n7561, A4 => 
                           n7562, ZN => n7549);
   U8935 : NAND4_X1 port map( A1 => n7551, A2 => n7552, A3 => n7553, A4 => 
                           n7554, ZN => n7550);
   U8936 : OAI21_X1 port map( B1 => n8784, B2 => n9493, A => n7529, ZN => n2588
                           );
   U8937 : OAI21_X1 port map( B1 => n7530, B2 => n7531, A => n9498, ZN => n7529
                           );
   U8938 : NAND4_X1 port map( A1 => n7540, A2 => n7541, A3 => n7542, A4 => 
                           n7543, ZN => n7530);
   U8939 : NAND4_X1 port map( A1 => n7532, A2 => n7533, A3 => n7534, A4 => 
                           n7535, ZN => n7531);
   U8940 : OAI21_X1 port map( B1 => n8783, B2 => n9494, A => n7478, ZN => n2589
                           );
   U8941 : OAI21_X1 port map( B1 => n7479, B2 => n7480, A => n9498, ZN => n7478
                           );
   U8942 : NAND4_X1 port map( A1 => n7505, A2 => n7506, A3 => n7507, A4 => 
                           n7508, ZN => n7479);
   U8943 : NAND4_X1 port map( A1 => n7481, A2 => n7482, A3 => n7483, A4 => 
                           n7484, ZN => n7480);
   U8944 : OAI22_X1 port map( A1 => n9736, A2 => n9782, B1 => n9735, B2 => 
                           n6631, ZN => n3422);
   U8945 : OAI22_X1 port map( A1 => n9736, A2 => n9783, B1 => n9735, B2 => 
                           n6630, ZN => n3423);
   U8946 : OAI22_X1 port map( A1 => n9736, A2 => n9786, B1 => n9735, B2 => 
                           n6629, ZN => n3424);
   U8947 : OAI22_X1 port map( A1 => n9736, A2 => n9789, B1 => n9735, B2 => 
                           n6628, ZN => n3425);
   U8948 : OAI22_X1 port map( A1 => n9736, A2 => n9792, B1 => n9735, B2 => 
                           n6627, ZN => n3426);
   U8949 : OAI22_X1 port map( A1 => n9737, A2 => n9795, B1 => n9735, B2 => 
                           n6626, ZN => n3427);
   U8950 : OAI22_X1 port map( A1 => n9737, A2 => n9798, B1 => n9735, B2 => 
                           n6625, ZN => n3428);
   U8951 : OAI22_X1 port map( A1 => n9737, A2 => n9801, B1 => n9735, B2 => 
                           n6624, ZN => n3429);
   U8952 : OAI22_X1 port map( A1 => n9737, A2 => n9804, B1 => n9735, B2 => 
                           n6623, ZN => n3430);
   U8953 : OAI22_X1 port map( A1 => n9737, A2 => n9807, B1 => n9735, B2 => 
                           n6622, ZN => n3431);
   U8954 : OAI22_X1 port map( A1 => n9738, A2 => n9810, B1 => n9735, B2 => 
                           n6621, ZN => n3432);
   U8955 : OAI22_X1 port map( A1 => n9738, A2 => n9813, B1 => n9735, B2 => 
                           n6620, ZN => n3433);
   U8956 : OAI22_X1 port map( A1 => n9738, A2 => n9816, B1 => n7443, B2 => 
                           n6619, ZN => n3434);
   U8957 : OAI22_X1 port map( A1 => n9738, A2 => n9819, B1 => n7443, B2 => 
                           n6618, ZN => n3435);
   U8958 : OAI22_X1 port map( A1 => n9738, A2 => n9822, B1 => n7443, B2 => 
                           n6617, ZN => n3436);
   U8959 : OAI22_X1 port map( A1 => n9739, A2 => n9825, B1 => n9735, B2 => 
                           n6616, ZN => n3437);
   U8960 : OAI22_X1 port map( A1 => n9739, A2 => n9828, B1 => n9735, B2 => 
                           n6615, ZN => n3438);
   U8961 : OAI22_X1 port map( A1 => n9739, A2 => n9831, B1 => n9735, B2 => 
                           n6614, ZN => n3439);
   U8962 : OAI22_X1 port map( A1 => n9739, A2 => n9834, B1 => n9735, B2 => 
                           n6613, ZN => n3440);
   U8963 : OAI22_X1 port map( A1 => n9739, A2 => n9837, B1 => n9735, B2 => 
                           n6612, ZN => n3441);
   U8964 : OAI22_X1 port map( A1 => n9740, A2 => n9840, B1 => n9735, B2 => 
                           n6611, ZN => n3442);
   U8965 : OAI22_X1 port map( A1 => n9740, A2 => n9843, B1 => n9735, B2 => 
                           n6610, ZN => n3443);
   U8966 : OAI22_X1 port map( A1 => n9740, A2 => n9846, B1 => n9735, B2 => 
                           n6609, ZN => n3444);
   U8967 : OAI22_X1 port map( A1 => n9740, A2 => n9849, B1 => n9735, B2 => 
                           n6608, ZN => n3445);
   U8968 : OAI22_X1 port map( A1 => n9740, A2 => n9852, B1 => n7443, B2 => 
                           n6607, ZN => n3446);
   U8969 : OAI22_X1 port map( A1 => n9741, A2 => n9855, B1 => n7443, B2 => 
                           n6606, ZN => n3447);
   U8970 : OAI22_X1 port map( A1 => n9741, A2 => n9858, B1 => n7443, B2 => 
                           n6605, ZN => n3448);
   U8971 : OAI22_X1 port map( A1 => n9741, A2 => n9861, B1 => n7443, B2 => 
                           n6604, ZN => n3449);
   U8972 : OAI22_X1 port map( A1 => n9741, A2 => n9864, B1 => n7443, B2 => 
                           n6603, ZN => n3450);
   U8973 : OAI22_X1 port map( A1 => n9741, A2 => n9867, B1 => n7443, B2 => 
                           n6602, ZN => n3451);
   U8974 : OAI22_X1 port map( A1 => n9742, A2 => n9870, B1 => n7443, B2 => 
                           n6601, ZN => n3452);
   U8975 : OAI22_X1 port map( A1 => n9742, A2 => n9882, B1 => n7443, B2 => 
                           n6600, ZN => n3453);
   U8976 : NOR2_X1 port map( A1 => n6463, A2 => ADD_RD2(2), ZN => n8108);
   U8977 : NOR2_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), ZN => n8110);
   U8978 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => 
                           ADD_RD1(0), ZN => n8777);
   U8979 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => 
                           ADD_RD2(0), ZN => n8124);
   U8980 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => n6460, 
                           ZN => n8776);
   U8981 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => n6464, 
                           ZN => n8123);
   U8982 : NOR2_X1 port map( A1 => n6459, A2 => ADD_RD1(2), ZN => n8761);
   U8983 : NOR2_X1 port map( A1 => n6458, A2 => ADD_RD1(1), ZN => n8766);
   U8984 : NOR2_X1 port map( A1 => n6462, A2 => ADD_RD2(1), ZN => n8113);
   U8985 : NOR3_X1 port map( A1 => n6460, A2 => ADD_RD1(4), A3 => n6457, ZN => 
                           n8781);
   U8986 : NOR3_X1 port map( A1 => n6464, A2 => ADD_RD2(4), A3 => n6461, ZN => 
                           n8128);
   U8987 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(4), A3 => n6457, 
                           ZN => n8780);
   U8988 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(4), A3 => n6461, 
                           ZN => n8127);
   U8989 : INV_X1 port map( A => RESET, ZN => n6451);
   U8990 : AND3_X1 port map( A1 => ENABLE, A2 => n9890, A3 => RD1, ZN => n8130)
                           ;
   U8991 : AND3_X1 port map( A1 => ENABLE, A2 => n9890, A3 => RD2, ZN => n7477)
                           ;
   U8992 : AND3_X1 port map( A1 => n6460, A2 => n6457, A3 => ADD_RD1(4), ZN => 
                           n8760);
   U8993 : AND3_X1 port map( A1 => n6464, A2 => n6461, A3 => ADD_RD2(4), ZN => 
                           n8107);
   U8994 : AND3_X1 port map( A1 => ADD_RD1(0), A2 => n6457, A3 => ADD_RD1(4), 
                           ZN => n8762);
   U8995 : AND3_X1 port map( A1 => ADD_RD1(3), A2 => n6460, A3 => ADD_RD1(4), 
                           ZN => n8768);
   U8996 : AND3_X1 port map( A1 => ADD_RD2(0), A2 => n6461, A3 => ADD_RD2(4), 
                           ZN => n8109);
   U8997 : AND3_X1 port map( A1 => ADD_RD2(3), A2 => n6464, A3 => ADD_RD2(4), 
                           ZN => n8115);
   U8998 : AND3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(0), A3 => 
                           ADD_RD1(4), ZN => n8769);
   U8999 : AND3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(0), A3 => 
                           ADD_RD2(4), ZN => n8116);
   U9000 : NAND2_X1 port map( A1 => DATAIN(8), A2 => n9886, ZN => n7424);
   U9001 : NAND2_X1 port map( A1 => DATAIN(9), A2 => n9886, ZN => n7423);
   U9002 : NAND2_X1 port map( A1 => DATAIN(10), A2 => n9886, ZN => n7422);
   U9003 : NAND2_X1 port map( A1 => DATAIN(11), A2 => n9886, ZN => n7421);
   U9004 : NAND2_X1 port map( A1 => DATAIN(12), A2 => n9886, ZN => n7420);
   U9005 : NAND2_X1 port map( A1 => DATAIN(13), A2 => n9886, ZN => n7419);
   U9006 : NAND2_X1 port map( A1 => DATAIN(14), A2 => n9886, ZN => n7418);
   U9007 : NAND2_X1 port map( A1 => DATAIN(15), A2 => n9886, ZN => n7417);
   U9008 : NAND2_X1 port map( A1 => DATAIN(16), A2 => n9886, ZN => n7416);
   U9009 : NAND2_X1 port map( A1 => DATAIN(17), A2 => n9886, ZN => n7415);
   U9010 : NAND2_X1 port map( A1 => DATAIN(18), A2 => n9886, ZN => n7414);
   U9011 : NAND2_X1 port map( A1 => DATAIN(19), A2 => n9886, ZN => n7413);
   U9012 : NAND2_X1 port map( A1 => DATAIN(20), A2 => n9885, ZN => n7412);
   U9013 : NAND2_X1 port map( A1 => DATAIN(21), A2 => n9885, ZN => n7411);
   U9014 : NAND2_X1 port map( A1 => DATAIN(22), A2 => n9885, ZN => n7410);
   U9015 : NAND2_X1 port map( A1 => DATAIN(23), A2 => n9885, ZN => n7409);
   U9016 : NAND2_X1 port map( A1 => DATAIN(24), A2 => n9885, ZN => n7408);
   U9017 : NAND2_X1 port map( A1 => DATAIN(25), A2 => n9885, ZN => n7407);
   U9018 : NAND2_X1 port map( A1 => DATAIN(26), A2 => n9885, ZN => n7406);
   U9019 : NAND2_X1 port map( A1 => DATAIN(27), A2 => n9885, ZN => n7405);
   U9020 : NAND2_X1 port map( A1 => DATAIN(28), A2 => n9885, ZN => n7404);
   U9021 : NAND2_X1 port map( A1 => DATAIN(29), A2 => n9885, ZN => n7403);
   U9022 : NAND2_X1 port map( A1 => DATAIN(30), A2 => n9885, ZN => n7402);
   U9023 : NAND2_X1 port map( A1 => DATAIN(31), A2 => n9885, ZN => n7400);
   U9024 : NAND2_X1 port map( A1 => DATAIN(0), A2 => n9887, ZN => n7432);
   U9025 : NAND2_X1 port map( A1 => DATAIN(1), A2 => n9887, ZN => n7431);
   U9026 : NAND2_X1 port map( A1 => DATAIN(2), A2 => n9887, ZN => n7430);
   U9027 : NAND2_X1 port map( A1 => DATAIN(3), A2 => n9887, ZN => n7429);
   U9028 : NAND2_X1 port map( A1 => DATAIN(4), A2 => n9887, ZN => n7428);
   U9029 : NAND2_X1 port map( A1 => DATAIN(5), A2 => n9887, ZN => n7427);
   U9030 : NAND2_X1 port map( A1 => DATAIN(6), A2 => n9887, ZN => n7426);
   U9031 : NAND2_X1 port map( A1 => DATAIN(7), A2 => n9887, ZN => n7425);
   U9032 : INV_X1 port map( A => ADD_RD1(3), ZN => n6457);
   U9033 : INV_X1 port map( A => ADD_RD2(3), ZN => n6461);
   U9034 : INV_X1 port map( A => ADD_RD1(0), ZN => n6460);
   U9035 : INV_X1 port map( A => ADD_RD2(0), ZN => n6464);
   U9036 : AND2_X1 port map( A1 => WR, A2 => ENABLE, ZN => n7449);
   U9037 : INV_X1 port map( A => ADD_WR(2), ZN => n6454);
   U9038 : INV_X1 port map( A => ADD_WR(0), ZN => n6456);
   U9039 : INV_X1 port map( A => ADD_WR(1), ZN => n6455);
   U9040 : INV_X1 port map( A => ADD_RD1(1), ZN => n6459);
   U9041 : INV_X1 port map( A => ADD_RD2(1), ZN => n6463);
   U9042 : INV_X1 port map( A => ADD_RD1(2), ZN => n6458);
   U9043 : INV_X1 port map( A => ADD_RD2(2), ZN => n6462);
   U9044 : INV_X1 port map( A => ADD_WR(4), ZN => n6452);
   U9045 : INV_X1 port map( A => ADD_WR(3), ZN => n6453);
   U9046 : CLKBUF_X1 port map( A => n8130, Z => n9396);
   U9047 : CLKBUF_X1 port map( A => n7477, Z => n9498);
   U9048 : CLKBUF_X1 port map( A => n6451, Z => n9890);

end SYN_Behavioural;
