
module BOOTHENC_NBIT34_i0 ( A_s, A_ns, B, O, A_so, A_nso );
  input [33:0] A_s;
  input [33:0] A_ns;
  input [33:0] B;
  output [33:0] O;
  output [33:0] A_so;
  output [33:0] A_nso;
  wire   \A_s[32] , \A_s[31] , \A_s[30] , \A_s[29] , \A_s[28] , \A_s[27] ,
         \A_s[26] , \A_s[25] , \A_s[24] , \A_s[23] , \A_s[22] , \A_s[21] ,
         \A_s[20] , \A_s[19] , \A_s[18] , \A_s[17] , \A_s[16] , \A_s[15] ,
         \A_s[14] , \A_s[13] , \A_s[12] , \A_s[11] , \A_s[10] , \A_s[9] ,
         \A_s[8] , \A_s[7] , \A_s[6] , \A_s[5] , \A_s[4] , \A_s[3] , \A_s[2] ,
         \A_s[1] , \A_s[0] , \A_ns[32] , \A_ns[31] , \A_ns[30] , \A_ns[29] ,
         \A_ns[28] , \A_ns[27] , \A_ns[26] , \A_ns[25] , \A_ns[24] ,
         \A_ns[23] , \A_ns[22] , \A_ns[21] , \A_ns[20] , \A_ns[19] ,
         \A_ns[18] , \A_ns[17] , \A_ns[16] , \A_ns[15] , \A_ns[14] ,
         \A_ns[13] , \A_ns[12] , \A_ns[11] , \A_ns[10] , \A_ns[9] , \A_ns[8] ,
         \A_ns[7] , \A_ns[6] , \A_ns[5] , \A_ns[4] , \A_ns[0] , n38, n39, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, net178205, net179447, net179465, net179461, net179459,
         net180847, net180845, net180844, net180842, net180839, net180838,
         net180837, net180836, net180835, net186499, net186666, net186677,
         net186799, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355;
  assign A_nso[0] = 1'b0;
  assign A_so[0] = 1'b0;
  assign A_so[33] = \A_s[32] ;
  assign \A_s[32]  = A_s[32];
  assign A_so[32] = \A_s[31] ;
  assign \A_s[31]  = A_s[31];
  assign A_so[31] = \A_s[30] ;
  assign \A_s[30]  = A_s[30];
  assign A_so[30] = \A_s[29] ;
  assign \A_s[29]  = A_s[29];
  assign A_so[29] = \A_s[28] ;
  assign \A_s[28]  = A_s[28];
  assign A_so[28] = \A_s[27] ;
  assign \A_s[27]  = A_s[27];
  assign A_so[27] = \A_s[26] ;
  assign \A_s[26]  = A_s[26];
  assign A_so[26] = \A_s[25] ;
  assign \A_s[25]  = A_s[25];
  assign A_so[25] = \A_s[24] ;
  assign \A_s[24]  = A_s[24];
  assign A_so[24] = \A_s[23] ;
  assign \A_s[23]  = A_s[23];
  assign A_so[23] = \A_s[22] ;
  assign \A_s[22]  = A_s[22];
  assign A_so[22] = \A_s[21] ;
  assign \A_s[21]  = A_s[21];
  assign A_so[21] = \A_s[20] ;
  assign \A_s[20]  = A_s[20];
  assign A_so[20] = \A_s[19] ;
  assign \A_s[19]  = A_s[19];
  assign A_so[19] = \A_s[18] ;
  assign \A_s[18]  = A_s[18];
  assign A_so[18] = \A_s[17] ;
  assign \A_s[17]  = A_s[17];
  assign A_so[17] = \A_s[16] ;
  assign \A_s[16]  = A_s[16];
  assign A_so[16] = \A_s[15] ;
  assign \A_s[15]  = A_s[15];
  assign A_so[15] = \A_s[14] ;
  assign \A_s[14]  = A_s[14];
  assign A_so[14] = \A_s[13] ;
  assign \A_s[13]  = A_s[13];
  assign A_so[13] = \A_s[12] ;
  assign \A_s[12]  = A_s[12];
  assign A_so[12] = \A_s[11] ;
  assign \A_s[11]  = A_s[11];
  assign A_so[11] = \A_s[10] ;
  assign \A_s[10]  = A_s[10];
  assign A_so[10] = \A_s[9] ;
  assign \A_s[9]  = A_s[9];
  assign A_so[9] = \A_s[8] ;
  assign \A_s[8]  = A_s[8];
  assign A_so[8] = \A_s[7] ;
  assign \A_s[7]  = A_s[7];
  assign A_so[7] = \A_s[6] ;
  assign \A_s[6]  = A_s[6];
  assign A_so[6] = \A_s[5] ;
  assign \A_s[5]  = A_s[5];
  assign A_so[5] = \A_s[4] ;
  assign \A_s[4]  = A_s[4];
  assign A_so[4] = \A_s[3] ;
  assign \A_s[3]  = A_s[3];
  assign A_so[3] = \A_s[2] ;
  assign \A_s[2]  = A_s[2];
  assign A_so[2] = \A_s[1] ;
  assign \A_s[1]  = A_s[1];
  assign A_so[1] = \A_s[0] ;
  assign \A_s[0]  = A_s[0];
  assign A_nso[33] = \A_ns[32] ;
  assign \A_ns[32]  = A_ns[32];
  assign A_nso[32] = \A_ns[31] ;
  assign \A_ns[31]  = A_ns[31];
  assign A_nso[31] = \A_ns[30] ;
  assign \A_ns[30]  = A_ns[30];
  assign A_nso[30] = \A_ns[29] ;
  assign \A_ns[29]  = A_ns[29];
  assign A_nso[29] = \A_ns[28] ;
  assign \A_ns[28]  = A_ns[28];
  assign A_nso[28] = \A_ns[27] ;
  assign \A_ns[27]  = A_ns[27];
  assign A_nso[27] = \A_ns[26] ;
  assign \A_ns[26]  = A_ns[26];
  assign A_nso[26] = \A_ns[25] ;
  assign \A_ns[25]  = A_ns[25];
  assign A_nso[25] = \A_ns[24] ;
  assign \A_ns[24]  = A_ns[24];
  assign A_nso[24] = \A_ns[23] ;
  assign \A_ns[23]  = A_ns[23];
  assign A_nso[23] = \A_ns[22] ;
  assign \A_ns[22]  = A_ns[22];
  assign A_nso[22] = \A_ns[21] ;
  assign \A_ns[21]  = A_ns[21];
  assign A_nso[21] = \A_ns[20] ;
  assign \A_ns[20]  = A_ns[20];
  assign A_nso[20] = \A_ns[19] ;
  assign \A_ns[19]  = A_ns[19];
  assign A_nso[19] = \A_ns[18] ;
  assign \A_ns[18]  = A_ns[18];
  assign A_nso[18] = \A_ns[17] ;
  assign \A_ns[17]  = A_ns[17];
  assign A_nso[17] = \A_ns[16] ;
  assign \A_ns[16]  = A_ns[16];
  assign A_nso[16] = \A_ns[15] ;
  assign \A_ns[15]  = A_ns[15];
  assign A_nso[15] = \A_ns[14] ;
  assign \A_ns[14]  = A_ns[14];
  assign A_nso[14] = \A_ns[13] ;
  assign \A_ns[13]  = A_ns[13];
  assign A_nso[13] = \A_ns[12] ;
  assign \A_ns[12]  = A_ns[12];
  assign A_nso[12] = \A_ns[11] ;
  assign \A_ns[11]  = A_ns[11];
  assign A_nso[11] = \A_ns[10] ;
  assign \A_ns[10]  = A_ns[10];
  assign A_nso[10] = \A_ns[9] ;
  assign \A_ns[9]  = A_ns[9];
  assign A_nso[9] = \A_ns[8] ;
  assign \A_ns[8]  = A_ns[8];
  assign A_nso[8] = \A_ns[7] ;
  assign \A_ns[7]  = A_ns[7];
  assign A_nso[7] = \A_ns[6] ;
  assign \A_ns[6]  = A_ns[6];
  assign A_nso[6] = \A_ns[5] ;
  assign \A_ns[5]  = A_ns[5];
  assign A_nso[5] = \A_ns[4] ;
  assign \A_ns[4]  = A_ns[4];
  assign A_nso[1] = \A_ns[0] ;
  assign \A_ns[0]  = A_ns[0];
  assign A_nso[3] = net186499;
  assign A_nso[2] = net186799;

  BUF_X1 U3 ( .A(n39), .Z(net180839) );
  BUF_X1 U4 ( .A(n39), .Z(net180838) );
  CLKBUF_X1 U5 ( .A(n39), .Z(net180835) );
  BUF_X1 U6 ( .A(net180835), .Z(net180842) );
  OAI221_X4 U7 ( .B1(net179461), .B2(n331), .C1(net186677), .C2(n330), .A(n43), 
        .ZN(O[8]) );
  NAND2_X1 U8 ( .A1(B[1]), .A2(B[0]), .ZN(n313) );
  INV_X1 U9 ( .A(A_ns[33]), .ZN(n322) );
  INV_X1 U10 ( .A(B[1]), .ZN(n321) );
  OAI221_X1 U11 ( .B1(net179459), .B2(n345), .C1(net179447), .C2(n344), .A(n60), .ZN(O[22]) );
  NAND2_X1 U12 ( .A1(net186799), .A2(n323), .ZN(n317) );
  INV_X1 U13 ( .A(net179459), .ZN(n323) );
  NOR2_X1 U14 ( .A1(net178205), .A2(n313), .ZN(n315) );
  OAI221_X1 U15 ( .B1(net179459), .B2(n347), .C1(net179447), .C2(n346), .A(n58), .ZN(O[24]) );
  NOR2_X1 U16 ( .A1(n311), .A2(n316), .ZN(n38) );
  NOR2_X1 U17 ( .A1(n322), .A2(n313), .ZN(n316) );
  OAI211_X1 U18 ( .C1(net179447), .C2(net178205), .A(n317), .B(n63), .ZN(O[1])
         );
  BUF_X1 U19 ( .A(net180835), .Z(net180844) );
  OR2_X1 U20 ( .A1(n312), .A2(n315), .ZN(O[0]) );
  INV_X1 U21 ( .A(n313), .ZN(net179465) );
  AND2_X1 U22 ( .A1(net180844), .A2(A_s[33]), .ZN(n311) );
  AND2_X1 U23 ( .A1(net180844), .A2(\A_s[0] ), .ZN(n312) );
  BUF_X1 U24 ( .A(n326), .Z(n325) );
  OAI221_X4 U25 ( .B1(net179459), .B2(n346), .C1(net186677), .C2(n345), .A(n59), .ZN(O[23]) );
  OAI221_X4 U26 ( .B1(net179459), .B2(n338), .C1(net186677), .C2(n337), .A(n68), .ZN(O[15]) );
  OAI221_X4 U27 ( .B1(net179459), .B2(n336), .C1(net186677), .C2(n335), .A(n70), .ZN(O[13]) );
  OAI221_X4 U28 ( .B1(net179459), .B2(n339), .C1(net186677), .C2(n338), .A(n67), .ZN(O[16]) );
  OAI221_X4 U29 ( .B1(net179459), .B2(n335), .C1(net186677), .C2(n334), .A(n71), .ZN(O[12]) );
  OAI221_X4 U30 ( .B1(net179459), .B2(n334), .C1(net186677), .C2(n333), .A(n72), .ZN(O[11]) );
  OAI221_X4 U31 ( .B1(net179459), .B2(n340), .C1(net186677), .C2(n339), .A(n66), .ZN(O[17]) );
  OAI221_X4 U32 ( .B1(net179461), .B2(n329), .C1(net186677), .C2(n328), .A(n45), .ZN(O[6]) );
  OAI221_X4 U33 ( .B1(net179459), .B2(n333), .C1(net186677), .C2(n332), .A(n73), .ZN(O[10]) );
  INV_X1 U34 ( .A(A_ns[1]), .ZN(n318) );
  OAI221_X4 U35 ( .B1(net179459), .B2(n343), .C1(net186677), .C2(n342), .A(n62), .ZN(O[20]) );
  BUF_X1 U36 ( .A(A_ns[2]), .Z(net186499) );
  OAI221_X4 U37 ( .B1(net179459), .B2(n341), .C1(net186677), .C2(n340), .A(n65), .ZN(O[18]) );
  INV_X1 U38 ( .A(B[0]), .ZN(n314) );
  BUF_X2 U39 ( .A(A_ns[1]), .Z(net186799) );
  NAND2_X4 U40 ( .A1(B[1]), .A2(n314), .ZN(net186677) );
  CLKBUF_X1 U41 ( .A(net186677), .Z(net179447) );
  NAND2_X1 U42 ( .A1(n39), .A2(\A_s[2] ), .ZN(n319) );
  OAI211_X1 U43 ( .C1(net186677), .C2(n318), .A(n319), .B(n320), .ZN(O[2]) );
  NAND2_X1 U44 ( .A1(A_ns[2]), .A2(net179465), .ZN(n320) );
  AND2_X2 U45 ( .A1(B[0]), .A2(n321), .ZN(n39) );
  INV_X1 U46 ( .A(n325), .ZN(A_nso[4]) );
  OAI221_X1 U47 ( .B1(n326), .B2(net179461), .C1(net186677), .C2(net186666), 
        .A(n48), .ZN(O[3]) );
  INV_X1 U48 ( .A(net186499), .ZN(net186666) );
  INV_X1 U49 ( .A(net179465), .ZN(net179459) );
  CLKBUF_X1 U50 ( .A(n39), .Z(net180837) );
  BUF_X1 U51 ( .A(n39), .Z(net180836) );
  CLKBUF_X1 U52 ( .A(net180836), .Z(net180845) );
  OAI221_X4 U53 ( .B1(net179459), .B2(n337), .C1(net186677), .C2(n336), .A(n69), .ZN(O[14]) );
  OAI221_X1 U54 ( .B1(net179459), .B2(n351), .C1(net179447), .C2(n350), .A(n54), .ZN(O[28]) );
  OAI221_X1 U55 ( .B1(net179461), .B2(n355), .C1(net179447), .C2(n354), .A(n49), .ZN(O[32]) );
  OAI221_X1 U56 ( .B1(net179461), .B2(n328), .C1(net186677), .C2(n327), .A(n46), .ZN(O[5]) );
  NAND2_X1 U57 ( .A1(\A_s[5] ), .A2(net180837), .ZN(n46) );
  NAND2_X1 U58 ( .A1(\A_s[6] ), .A2(net180838), .ZN(n45) );
  NAND2_X1 U59 ( .A1(\A_s[8] ), .A2(net180838), .ZN(n43) );
  OAI221_X1 U60 ( .B1(n327), .B2(net179461), .C1(net186677), .C2(n325), .A(n47), .ZN(O[4]) );
  NAND2_X1 U61 ( .A1(\A_s[4] ), .A2(net180837), .ZN(n47) );
  NAND2_X1 U62 ( .A1(\A_s[3] ), .A2(net180839), .ZN(n48) );
  OAI221_X1 U63 ( .B1(net179461), .B2(n330), .C1(net186677), .C2(n329), .A(n44), .ZN(O[7]) );
  NAND2_X1 U64 ( .A1(\A_s[7] ), .A2(net180839), .ZN(n44) );
  OAI221_X1 U65 ( .B1(net179461), .B2(n332), .C1(net186677), .C2(n331), .A(n42), .ZN(O[9]) );
  NAND2_X1 U66 ( .A1(\A_s[9] ), .A2(net180836), .ZN(n42) );
  OAI221_X1 U67 ( .B1(net179459), .B2(n353), .C1(net179447), .C2(n352), .A(n51), .ZN(O[30]) );
  NAND2_X1 U68 ( .A1(\A_s[30] ), .A2(net180844), .ZN(n51) );
  OAI221_X1 U69 ( .B1(net179459), .B2(n352), .C1(net179447), .C2(n351), .A(n53), .ZN(O[29]) );
  NAND2_X1 U70 ( .A1(\A_s[29] ), .A2(net180844), .ZN(n53) );
  OAI221_X1 U71 ( .B1(net179459), .B2(n344), .C1(net179447), .C2(n343), .A(n61), .ZN(O[21]) );
  NAND2_X1 U72 ( .A1(\A_s[21] ), .A2(net180844), .ZN(n61) );
  OAI221_X1 U73 ( .B1(net179459), .B2(n342), .C1(net186677), .C2(n341), .A(n64), .ZN(O[19]) );
  NAND2_X1 U74 ( .A1(\A_s[19] ), .A2(net180844), .ZN(n64) );
  NAND2_X1 U75 ( .A1(\A_s[17] ), .A2(net180844), .ZN(n66) );
  NAND2_X1 U76 ( .A1(\A_s[15] ), .A2(net180842), .ZN(n68) );
  NAND2_X1 U77 ( .A1(\A_s[14] ), .A2(net180842), .ZN(n69) );
  NAND2_X1 U78 ( .A1(\A_s[13] ), .A2(net180845), .ZN(n70) );
  NAND2_X1 U79 ( .A1(\A_s[12] ), .A2(net180847), .ZN(n71) );
  NAND2_X1 U80 ( .A1(\A_s[20] ), .A2(net180844), .ZN(n62) );
  NAND2_X1 U81 ( .A1(\A_s[18] ), .A2(net180844), .ZN(n65) );
  NAND2_X1 U82 ( .A1(\A_s[16] ), .A2(net180842), .ZN(n67) );
  NAND2_X1 U83 ( .A1(\A_s[10] ), .A2(net180835), .ZN(n73) );
  NAND2_X1 U84 ( .A1(\A_s[22] ), .A2(net180844), .ZN(n60) );
  NAND2_X1 U85 ( .A1(\A_s[24] ), .A2(net180844), .ZN(n58) );
  NAND2_X1 U86 ( .A1(\A_s[11] ), .A2(net180847), .ZN(n72) );
  OAI221_X1 U87 ( .B1(net179459), .B2(n349), .C1(net179447), .C2(n348), .A(n56), .ZN(O[26]) );
  NAND2_X1 U88 ( .A1(\A_s[26] ), .A2(net180844), .ZN(n56) );
  NAND2_X1 U89 ( .A1(\A_s[23] ), .A2(net180844), .ZN(n59) );
  OAI21_X1 U90 ( .B1(net179447), .B2(n355), .A(n38), .ZN(O[33]) );
  OAI221_X1 U91 ( .B1(net179459), .B2(n350), .C1(net179447), .C2(n349), .A(n55), .ZN(O[27]) );
  NAND2_X1 U92 ( .A1(\A_s[27] ), .A2(net180844), .ZN(n55) );
  OAI221_X1 U93 ( .B1(net179459), .B2(n348), .C1(net179447), .C2(n347), .A(n57), .ZN(O[25]) );
  NAND2_X1 U94 ( .A1(\A_s[25] ), .A2(net180844), .ZN(n57) );
  OAI221_X1 U95 ( .B1(net179459), .B2(n354), .C1(net179447), .C2(n353), .A(n50), .ZN(O[31]) );
  NAND2_X1 U96 ( .A1(\A_s[31] ), .A2(net180844), .ZN(n50) );
  NAND2_X1 U97 ( .A1(\A_s[28] ), .A2(net180844), .ZN(n54) );
  NAND2_X1 U98 ( .A1(\A_s[32] ), .A2(net180844), .ZN(n49) );
  NAND2_X1 U99 ( .A1(\A_s[1] ), .A2(net180844), .ZN(n63) );
  BUF_X1 U100 ( .A(net180836), .Z(net180847) );
  INV_X1 U101 ( .A(net179465), .ZN(net179461) );
  INV_X1 U102 ( .A(A_ns[3]), .ZN(n326) );
  INV_X1 U103 ( .A(\A_ns[4] ), .ZN(n327) );
  INV_X1 U104 ( .A(\A_ns[5] ), .ZN(n328) );
  INV_X1 U105 ( .A(\A_ns[6] ), .ZN(n329) );
  INV_X1 U106 ( .A(\A_ns[7] ), .ZN(n330) );
  INV_X1 U107 ( .A(\A_ns[8] ), .ZN(n331) );
  INV_X1 U108 ( .A(\A_ns[9] ), .ZN(n332) );
  INV_X1 U109 ( .A(\A_ns[10] ), .ZN(n333) );
  INV_X1 U110 ( .A(\A_ns[11] ), .ZN(n334) );
  INV_X1 U111 ( .A(\A_ns[12] ), .ZN(n335) );
  INV_X1 U112 ( .A(\A_ns[13] ), .ZN(n336) );
  INV_X1 U113 ( .A(\A_ns[14] ), .ZN(n337) );
  INV_X1 U114 ( .A(\A_ns[15] ), .ZN(n338) );
  INV_X1 U115 ( .A(\A_ns[16] ), .ZN(n339) );
  INV_X1 U116 ( .A(\A_ns[17] ), .ZN(n340) );
  INV_X1 U117 ( .A(\A_ns[18] ), .ZN(n341) );
  INV_X1 U118 ( .A(\A_ns[19] ), .ZN(n342) );
  INV_X1 U119 ( .A(\A_ns[20] ), .ZN(n343) );
  INV_X1 U120 ( .A(\A_ns[21] ), .ZN(n344) );
  INV_X1 U121 ( .A(\A_ns[22] ), .ZN(n345) );
  INV_X1 U122 ( .A(\A_ns[23] ), .ZN(n346) );
  INV_X1 U123 ( .A(\A_ns[24] ), .ZN(n347) );
  INV_X1 U124 ( .A(\A_ns[25] ), .ZN(n348) );
  INV_X1 U125 ( .A(\A_ns[26] ), .ZN(n349) );
  INV_X1 U126 ( .A(\A_ns[27] ), .ZN(n350) );
  INV_X1 U127 ( .A(\A_ns[28] ), .ZN(n351) );
  INV_X1 U128 ( .A(\A_ns[29] ), .ZN(n352) );
  INV_X1 U129 ( .A(\A_ns[30] ), .ZN(n353) );
  INV_X1 U130 ( .A(\A_ns[31] ), .ZN(n354) );
  INV_X1 U131 ( .A(\A_ns[32] ), .ZN(n355) );
  INV_X1 U132 ( .A(\A_ns[0] ), .ZN(net178205) );
endmodule


module BOOTHENC_NBIT36_i2 ( A_s, A_ns, B, O, A_so, A_nso );
  input [35:0] A_s;
  input [35:0] A_ns;
  input [35:0] B;
  output [35:0] O;
  output [35:0] A_so;
  output [35:0] A_nso;
  wire   \A_s[33] , \A_s[32] , \A_s[31] , \A_s[29] , \A_s[28] , \A_s[27] ,
         \A_s[26] , \A_s[25] , \A_s[24] , \A_s[23] , \A_s[22] , \A_s[21] ,
         \A_s[20] , \A_s[19] , \A_s[18] , \A_s[17] , \A_s[16] , \A_s[1] ,
         \A_s[0] , \A_ns[2] , \A_ns[0] , n74, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n91, n92, n93, n94, n95, n96,
         n97, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         net178197, net178199, net179469, net179477, net179483, net179489,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n463, n464, n466, n468, n470, n472, n474,
         n476, n478, n480, n482, n484, n486, n488, n490, n492, n494, n496,
         n498, n500, n502, n504, n506, n508, n510, n512, n514, n516, n518,
         n520, n522, n523, n525, n527, n529, n531, n533, n535, n537, n539,
         n541, n543, n545, n547, n549, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n567, n568,
         n569, n570;
  assign A_nso[0] = 1'b0;
  assign A_nso[1] = 1'b0;
  assign A_so[0] = 1'b0;
  assign A_so[1] = 1'b0;
  assign O[0] = 1'b0;
  assign A_so[35] = \A_s[33] ;
  assign \A_s[33]  = A_s[33];
  assign A_so[34] = \A_s[32] ;
  assign \A_s[32]  = A_s[32];
  assign A_so[33] = \A_s[31] ;
  assign \A_s[31]  = A_s[31];
  assign A_so[31] = \A_s[29] ;
  assign \A_s[29]  = A_s[29];
  assign A_so[30] = \A_s[28] ;
  assign \A_s[28]  = A_s[28];
  assign A_so[29] = \A_s[27] ;
  assign \A_s[27]  = A_s[27];
  assign A_so[28] = \A_s[26] ;
  assign \A_s[26]  = A_s[26];
  assign A_so[27] = \A_s[25] ;
  assign \A_s[25]  = A_s[25];
  assign A_so[26] = \A_s[24] ;
  assign \A_s[24]  = A_s[24];
  assign A_so[25] = \A_s[23] ;
  assign \A_s[23]  = A_s[23];
  assign A_so[24] = \A_s[22] ;
  assign \A_s[22]  = A_s[22];
  assign A_so[23] = \A_s[21] ;
  assign \A_s[21]  = A_s[21];
  assign A_so[22] = \A_s[20] ;
  assign \A_s[20]  = A_s[20];
  assign A_so[21] = \A_s[19] ;
  assign \A_s[19]  = A_s[19];
  assign A_so[20] = \A_s[18] ;
  assign \A_s[18]  = A_s[18];
  assign A_so[19] = \A_s[17] ;
  assign \A_s[17]  = A_s[17];
  assign A_so[18] = \A_s[16] ;
  assign \A_s[16]  = A_s[16];
  assign A_so[3] = \A_s[1] ;
  assign \A_s[1]  = A_s[1];
  assign A_so[2] = \A_s[0] ;
  assign \A_s[0]  = A_s[0];
  assign A_nso[4] = \A_ns[2] ;
  assign \A_ns[2]  = A_ns[2];
  assign A_nso[2] = \A_ns[0] ;
  assign \A_ns[0]  = A_ns[0];
  assign A_nso[3] = net178199;

  NAND2_X1 U2 ( .A1(\A_s[0] ), .A2(n441), .ZN(n450) );
  INV_X1 U3 ( .A(\A_ns[0] ), .ZN(n449) );
  INV_X1 U4 ( .A(B[2]), .ZN(n447) );
  OAI21_X1 U5 ( .B1(net179469), .B2(n449), .A(n450), .ZN(O[1]) );
  MUX2_X1 U6 ( .A(n455), .B(n459), .S(B[3]), .Z(n460) );
  NAND2_X1 U7 ( .A1(n452), .A2(B[3]), .ZN(n453) );
  NAND2_X1 U8 ( .A1(n442), .A2(n460), .ZN(O[2]) );
  BUF_X2 U9 ( .A(A_ns[4]), .Z(A_nso[6]) );
  INV_X4 U10 ( .A(n453), .ZN(net179483) );
  NAND2_X1 U11 ( .A1(n443), .A2(n436), .ZN(n437) );
  NAND2_X1 U12 ( .A1(n444), .A2(B[3]), .ZN(n438) );
  NAND2_X1 U13 ( .A1(n437), .A2(n438), .ZN(n442) );
  INV_X1 U14 ( .A(B[3]), .ZN(n436) );
  OR2_X1 U15 ( .A1(net179469), .A2(n461), .ZN(n439) );
  OR2_X1 U16 ( .A1(net179477), .A2(net178197), .ZN(n440) );
  NAND3_X1 U17 ( .A1(n439), .A2(n440), .A3(n89), .ZN(O[3]) );
  INV_X2 U18 ( .A(n454), .ZN(n441) );
  INV_X1 U19 ( .A(n454), .ZN(net179489) );
  NAND2_X1 U20 ( .A1(n445), .A2(n448), .ZN(n454) );
  OR2_X1 U21 ( .A1(n456), .A2(net178197), .ZN(n443) );
  OR3_X1 U22 ( .A1(n449), .A2(B[2]), .A3(B[1]), .ZN(n444) );
  XOR2_X1 U23 ( .A(B[2]), .B(B[1]), .Z(n445) );
  INV_X1 U24 ( .A(\A_s[1] ), .ZN(net178197) );
  NOR2_X1 U25 ( .A1(B[2]), .A2(B[1]), .ZN(n452) );
  INV_X1 U26 ( .A(B[1]), .ZN(n446) );
  OR3_X4 U27 ( .A1(B[3]), .A2(n446), .A3(n447), .ZN(net179477) );
  NAND3_X1 U28 ( .A1(B[1]), .A2(B[2]), .A3(\A_s[0] ), .ZN(n455) );
  INV_X1 U29 ( .A(A_ns[1]), .ZN(n451) );
  OR2_X4 U30 ( .A1(n457), .A2(n448), .ZN(net179469) );
  INV_X2 U31 ( .A(n451), .ZN(net178199) );
  XNOR2_X1 U32 ( .A(B[2]), .B(B[1]), .ZN(n456) );
  XNOR2_X1 U33 ( .A(B[2]), .B(B[1]), .ZN(n457) );
  XOR2_X1 U34 ( .A(B[2]), .B(B[1]), .Z(n458) );
  INV_X1 U35 ( .A(B[3]), .ZN(n448) );
  NAND2_X1 U36 ( .A1(n458), .A2(A_ns[1]), .ZN(n459) );
  AOI22_X1 U37 ( .A1(A_nso[32]), .A2(net179483), .B1(\A_s[31] ), .B2(n441), 
        .ZN(n76) );
  AOI22_X1 U38 ( .A1(A_nso[30]), .A2(net179483), .B1(\A_s[29] ), .B2(n441), 
        .ZN(n77) );
  AOI22_X1 U39 ( .A1(A_nso[28]), .A2(net179483), .B1(\A_s[27] ), .B2(n441), 
        .ZN(n78) );
  OAI221_X1 U40 ( .B1(net179469), .B2(n468), .C1(net179477), .C2(n531), .A(n92), .ZN(O[7]) );
  AOI22_X1 U41 ( .A1(A_nso[7]), .A2(net179483), .B1(A_so[8]), .B2(n441), .ZN(
        n92) );
  OAI221_X1 U42 ( .B1(net179469), .B2(n472), .C1(net179477), .C2(n535), .A(n91), .ZN(O[9]) );
  AOI22_X1 U43 ( .A1(A_nso[9]), .A2(net179483), .B1(A_so[10]), .B2(n441), .ZN(
        n91) );
  OAI221_X1 U44 ( .B1(net179469), .B2(n523), .C1(n570), .C2(net179477), .A(n95), .ZN(O[35]) );
  OAI221_X1 U45 ( .B1(net179469), .B2(n463), .C1(net179477), .C2(n525), .A(n94), .ZN(O[4]) );
  AOI22_X1 U46 ( .A1(\A_ns[2] ), .A2(net179483), .B1(A_so[5]), .B2(net179489), 
        .ZN(n94) );
  OAI221_X1 U47 ( .B1(net179469), .B2(n466), .C1(net179477), .C2(n529), .A(n88), .ZN(O[6]) );
  AOI22_X1 U48 ( .A1(A_nso[6]), .A2(net179483), .B1(A_so[7]), .B2(n441), .ZN(
        n88) );
  OAI221_X1 U49 ( .B1(net179469), .B2(n470), .C1(net179477), .C2(n533), .A(n87), .ZN(O[8]) );
  AOI22_X1 U50 ( .A1(A_nso[8]), .A2(net179483), .B1(A_so[9]), .B2(n441), .ZN(
        n87) );
  OAI221_X1 U51 ( .B1(net179469), .B2(n464), .C1(net179477), .C2(n527), .A(n93), .ZN(O[5]) );
  AOI22_X1 U52 ( .A1(A_nso[5]), .A2(net179483), .B1(A_so[6]), .B2(n441), .ZN(
        n93) );
  OAI221_X1 U53 ( .B1(net179469), .B2(n510), .C1(net179477), .C2(n562), .A(n78), .ZN(O[28]) );
  OAI221_X1 U54 ( .B1(net179469), .B2(n518), .C1(net179477), .C2(n567), .A(n76), .ZN(O[32]) );
  OAI221_X1 U55 ( .B1(net179469), .B2(n500), .C1(net179477), .C2(n557), .A(
        n102), .ZN(O[23]) );
  OAI221_X1 U56 ( .B1(net179469), .B2(n478), .C1(net179477), .C2(n541), .A(n86), .ZN(O[12]) );
  AOI22_X1 U57 ( .A1(A_nso[12]), .A2(net179483), .B1(A_so[13]), .B2(n441), 
        .ZN(n86) );
  OAI221_X1 U58 ( .B1(net179469), .B2(n482), .C1(net179477), .C2(n545), .A(n85), .ZN(O[14]) );
  AOI22_X1 U59 ( .A1(A_nso[14]), .A2(net179483), .B1(A_so[15]), .B2(n441), 
        .ZN(n85) );
  OAI221_X1 U60 ( .B1(net179469), .B2(n498), .C1(net179477), .C2(n556), .A(n81), .ZN(O[22]) );
  AOI22_X1 U61 ( .A1(A_nso[22]), .A2(net179483), .B1(\A_s[21] ), .B2(n441), 
        .ZN(n81) );
  OAI221_X1 U62 ( .B1(net179469), .B2(n502), .C1(net179477), .C2(n558), .A(n80), .ZN(O[24]) );
  AOI22_X1 U63 ( .A1(A_nso[24]), .A2(net179483), .B1(\A_s[23] ), .B2(n441), 
        .ZN(n80) );
  OAI221_X1 U64 ( .B1(net179469), .B2(n494), .C1(net179477), .C2(n554), .A(n82), .ZN(O[20]) );
  AOI22_X1 U65 ( .A1(A_nso[20]), .A2(net179483), .B1(\A_s[19] ), .B2(n441), 
        .ZN(n82) );
  OAI221_X1 U66 ( .B1(net179469), .B2(n490), .C1(net179477), .C2(n552), .A(n83), .ZN(O[18]) );
  AOI22_X1 U67 ( .A1(A_nso[18]), .A2(net179483), .B1(\A_s[17] ), .B2(n441), 
        .ZN(n83) );
  OAI221_X1 U68 ( .B1(net179469), .B2(n474), .C1(net179477), .C2(n537), .A(
        n109), .ZN(O[10]) );
  OAI221_X1 U69 ( .B1(net179469), .B2(n486), .C1(net179477), .C2(n549), .A(n84), .ZN(O[16]) );
  AOI22_X1 U70 ( .A1(A_nso[16]), .A2(net179483), .B1(A_so[17]), .B2(n441), 
        .ZN(n84) );
  OAI221_X1 U71 ( .B1(net179469), .B2(n522), .C1(net179477), .C2(n569), .A(n74), .ZN(O[34]) );
  AOI22_X1 U72 ( .A1(A_nso[34]), .A2(net179483), .B1(\A_s[33] ), .B2(n441), 
        .ZN(n74) );
  OAI221_X1 U73 ( .B1(net179469), .B2(n506), .C1(net179477), .C2(n560), .A(n79), .ZN(O[26]) );
  AOI22_X1 U74 ( .A1(A_nso[26]), .A2(net179483), .B1(\A_s[25] ), .B2(n441), 
        .ZN(n79) );
  OAI221_X1 U75 ( .B1(net179469), .B2(n516), .C1(net179477), .C2(n565), .A(n97), .ZN(O[31]) );
  AOI22_X1 U76 ( .A1(A_nso[31]), .A2(net179483), .B1(A_so[32]), .B2(n441), 
        .ZN(n97) );
  OAI221_X1 U77 ( .B1(n520), .B2(net179469), .C1(net179477), .C2(n568), .A(n96), .ZN(O[33]) );
  AOI22_X1 U78 ( .A1(A_nso[33]), .A2(net179483), .B1(\A_s[32] ), .B2(n441), 
        .ZN(n96) );
  OAI221_X1 U79 ( .B1(net179469), .B2(n508), .C1(net179477), .C2(n561), .A(
        n100), .ZN(O[27]) );
  AOI22_X1 U80 ( .A1(net178199), .A2(net179483), .B1(A_so[4]), .B2(net179489), 
        .ZN(n89) );
  OAI221_X1 U81 ( .B1(net179469), .B2(n514), .C1(net179477), .C2(n564), .A(n77), .ZN(O[30]) );
  OAI221_X1 U82 ( .B1(net179469), .B2(n512), .C1(net179477), .C2(n563), .A(n99), .ZN(O[29]) );
  AOI22_X1 U83 ( .A1(A_nso[35]), .A2(net179483), .B1(A_s[34]), .B2(n441), .ZN(
        n95) );
  OAI221_X1 U84 ( .B1(net179469), .B2(n504), .C1(net179477), .C2(n559), .A(
        n101), .ZN(O[25]) );
  OAI221_X1 U85 ( .B1(net179469), .B2(n496), .C1(net179477), .C2(n555), .A(
        n103), .ZN(O[21]) );
  OAI221_X1 U86 ( .B1(net179469), .B2(n492), .C1(net179477), .C2(n553), .A(
        n104), .ZN(O[19]) );
  OAI221_X1 U87 ( .B1(net179469), .B2(n488), .C1(net179477), .C2(n551), .A(
        n105), .ZN(O[17]) );
  OAI221_X1 U88 ( .B1(net179469), .B2(n484), .C1(net179477), .C2(n547), .A(
        n106), .ZN(O[15]) );
  OAI221_X1 U89 ( .B1(net179469), .B2(n480), .C1(net179477), .C2(n543), .A(
        n107), .ZN(O[13]) );
  OAI221_X1 U90 ( .B1(net179469), .B2(n476), .C1(net179477), .C2(n539), .A(
        n108), .ZN(O[11]) );
  AOI22_X1 U91 ( .A1(A_nso[29]), .A2(net179483), .B1(\A_s[28] ), .B2(n441), 
        .ZN(n99) );
  AOI22_X1 U92 ( .A1(A_nso[27]), .A2(net179483), .B1(\A_s[26] ), .B2(n441), 
        .ZN(n100) );
  AOI22_X1 U93 ( .A1(A_nso[25]), .A2(net179483), .B1(\A_s[24] ), .B2(n441), 
        .ZN(n101) );
  AOI22_X1 U94 ( .A1(A_nso[23]), .A2(net179483), .B1(\A_s[22] ), .B2(n441), 
        .ZN(n102) );
  AOI22_X1 U95 ( .A1(A_nso[21]), .A2(net179483), .B1(\A_s[20] ), .B2(n441), 
        .ZN(n103) );
  AOI22_X1 U96 ( .A1(A_nso[19]), .A2(net179483), .B1(\A_s[18] ), .B2(n441), 
        .ZN(n104) );
  AOI22_X1 U97 ( .A1(A_nso[17]), .A2(net179483), .B1(\A_s[16] ), .B2(n441), 
        .ZN(n105) );
  AOI22_X1 U98 ( .A1(A_nso[15]), .A2(net179483), .B1(A_so[16]), .B2(n441), 
        .ZN(n106) );
  AOI22_X1 U99 ( .A1(A_nso[13]), .A2(net179483), .B1(A_so[14]), .B2(n441), 
        .ZN(n107) );
  AOI22_X1 U100 ( .A1(A_nso[11]), .A2(net179483), .B1(A_so[12]), .B2(n441), 
        .ZN(n108) );
  AOI22_X1 U101 ( .A1(A_nso[10]), .A2(net179483), .B1(A_so[11]), .B2(n441), 
        .ZN(n109) );
  INV_X1 U102 ( .A(\A_ns[2] ), .ZN(n461) );
  INV_X1 U103 ( .A(n463), .ZN(A_nso[5]) );
  INV_X1 U104 ( .A(A_ns[3]), .ZN(n463) );
  INV_X1 U105 ( .A(A_ns[4]), .ZN(n464) );
  INV_X1 U106 ( .A(n466), .ZN(A_nso[7]) );
  INV_X1 U107 ( .A(A_ns[5]), .ZN(n466) );
  INV_X1 U108 ( .A(n468), .ZN(A_nso[8]) );
  INV_X1 U109 ( .A(A_ns[6]), .ZN(n468) );
  INV_X1 U110 ( .A(n470), .ZN(A_nso[9]) );
  INV_X1 U111 ( .A(A_ns[7]), .ZN(n470) );
  INV_X1 U112 ( .A(n472), .ZN(A_nso[10]) );
  INV_X1 U113 ( .A(A_ns[8]), .ZN(n472) );
  INV_X1 U114 ( .A(n474), .ZN(A_nso[11]) );
  INV_X1 U115 ( .A(A_ns[9]), .ZN(n474) );
  INV_X1 U116 ( .A(n476), .ZN(A_nso[12]) );
  INV_X1 U117 ( .A(A_ns[10]), .ZN(n476) );
  INV_X1 U118 ( .A(n478), .ZN(A_nso[13]) );
  INV_X1 U119 ( .A(A_ns[11]), .ZN(n478) );
  INV_X1 U120 ( .A(n480), .ZN(A_nso[14]) );
  INV_X1 U121 ( .A(A_ns[12]), .ZN(n480) );
  INV_X1 U122 ( .A(n482), .ZN(A_nso[15]) );
  INV_X1 U123 ( .A(A_ns[13]), .ZN(n482) );
  INV_X1 U124 ( .A(n484), .ZN(A_nso[16]) );
  INV_X1 U125 ( .A(A_ns[14]), .ZN(n484) );
  INV_X1 U126 ( .A(n486), .ZN(A_nso[17]) );
  INV_X1 U127 ( .A(A_ns[15]), .ZN(n486) );
  INV_X1 U128 ( .A(n488), .ZN(A_nso[18]) );
  INV_X1 U129 ( .A(A_ns[16]), .ZN(n488) );
  INV_X1 U130 ( .A(n490), .ZN(A_nso[19]) );
  INV_X1 U131 ( .A(A_ns[17]), .ZN(n490) );
  INV_X1 U132 ( .A(n492), .ZN(A_nso[20]) );
  INV_X1 U133 ( .A(A_ns[18]), .ZN(n492) );
  INV_X1 U134 ( .A(n494), .ZN(A_nso[21]) );
  INV_X1 U135 ( .A(A_ns[19]), .ZN(n494) );
  INV_X1 U136 ( .A(n496), .ZN(A_nso[22]) );
  INV_X1 U137 ( .A(A_ns[20]), .ZN(n496) );
  INV_X1 U138 ( .A(n498), .ZN(A_nso[23]) );
  INV_X1 U139 ( .A(A_ns[21]), .ZN(n498) );
  INV_X1 U140 ( .A(n500), .ZN(A_nso[24]) );
  INV_X1 U141 ( .A(A_ns[22]), .ZN(n500) );
  INV_X1 U142 ( .A(n502), .ZN(A_nso[25]) );
  INV_X1 U143 ( .A(A_ns[23]), .ZN(n502) );
  INV_X1 U144 ( .A(n504), .ZN(A_nso[26]) );
  INV_X1 U145 ( .A(A_ns[24]), .ZN(n504) );
  INV_X1 U146 ( .A(n506), .ZN(A_nso[27]) );
  INV_X1 U147 ( .A(A_ns[25]), .ZN(n506) );
  INV_X1 U148 ( .A(n508), .ZN(A_nso[28]) );
  INV_X1 U149 ( .A(A_ns[26]), .ZN(n508) );
  INV_X1 U150 ( .A(n510), .ZN(A_nso[29]) );
  INV_X1 U151 ( .A(A_ns[27]), .ZN(n510) );
  INV_X1 U152 ( .A(n512), .ZN(A_nso[30]) );
  INV_X1 U153 ( .A(A_ns[28]), .ZN(n512) );
  INV_X1 U154 ( .A(n514), .ZN(A_nso[31]) );
  INV_X1 U155 ( .A(A_ns[29]), .ZN(n514) );
  INV_X1 U156 ( .A(n516), .ZN(A_nso[32]) );
  INV_X1 U157 ( .A(A_ns[30]), .ZN(n516) );
  INV_X1 U158 ( .A(n518), .ZN(A_nso[33]) );
  INV_X1 U159 ( .A(A_ns[31]), .ZN(n518) );
  INV_X1 U160 ( .A(n520), .ZN(A_nso[34]) );
  INV_X1 U161 ( .A(A_ns[32]), .ZN(n520) );
  INV_X1 U162 ( .A(n522), .ZN(A_nso[35]) );
  INV_X1 U163 ( .A(A_ns[33]), .ZN(n522) );
  INV_X1 U164 ( .A(A_ns[34]), .ZN(n523) );
  INV_X1 U165 ( .A(n525), .ZN(A_so[4]) );
  INV_X1 U166 ( .A(A_s[2]), .ZN(n525) );
  INV_X1 U167 ( .A(n527), .ZN(A_so[5]) );
  INV_X1 U168 ( .A(A_s[3]), .ZN(n527) );
  INV_X1 U169 ( .A(n529), .ZN(A_so[6]) );
  INV_X1 U170 ( .A(A_s[4]), .ZN(n529) );
  INV_X1 U171 ( .A(n531), .ZN(A_so[7]) );
  INV_X1 U172 ( .A(A_s[5]), .ZN(n531) );
  INV_X1 U173 ( .A(n533), .ZN(A_so[8]) );
  INV_X1 U174 ( .A(A_s[6]), .ZN(n533) );
  INV_X1 U175 ( .A(n535), .ZN(A_so[9]) );
  INV_X1 U176 ( .A(A_s[7]), .ZN(n535) );
  INV_X1 U177 ( .A(n537), .ZN(A_so[10]) );
  INV_X1 U178 ( .A(A_s[8]), .ZN(n537) );
  INV_X1 U179 ( .A(n539), .ZN(A_so[11]) );
  INV_X1 U180 ( .A(A_s[9]), .ZN(n539) );
  INV_X1 U181 ( .A(n541), .ZN(A_so[12]) );
  INV_X1 U182 ( .A(A_s[10]), .ZN(n541) );
  INV_X1 U183 ( .A(n543), .ZN(A_so[13]) );
  INV_X1 U184 ( .A(A_s[11]), .ZN(n543) );
  INV_X1 U185 ( .A(n545), .ZN(A_so[14]) );
  INV_X1 U186 ( .A(A_s[12]), .ZN(n545) );
  INV_X1 U187 ( .A(n547), .ZN(A_so[15]) );
  INV_X1 U188 ( .A(A_s[13]), .ZN(n547) );
  INV_X1 U189 ( .A(n549), .ZN(A_so[16]) );
  INV_X1 U190 ( .A(A_s[14]), .ZN(n549) );
  INV_X1 U191 ( .A(n551), .ZN(A_so[17]) );
  INV_X1 U192 ( .A(A_s[15]), .ZN(n551) );
  INV_X1 U193 ( .A(\A_s[16] ), .ZN(n552) );
  INV_X1 U194 ( .A(\A_s[17] ), .ZN(n553) );
  INV_X1 U195 ( .A(\A_s[18] ), .ZN(n554) );
  INV_X1 U196 ( .A(\A_s[19] ), .ZN(n555) );
  INV_X1 U197 ( .A(\A_s[20] ), .ZN(n556) );
  INV_X1 U198 ( .A(\A_s[21] ), .ZN(n557) );
  INV_X1 U199 ( .A(\A_s[22] ), .ZN(n558) );
  INV_X1 U200 ( .A(\A_s[23] ), .ZN(n559) );
  INV_X1 U201 ( .A(\A_s[24] ), .ZN(n560) );
  INV_X1 U202 ( .A(\A_s[25] ), .ZN(n561) );
  INV_X1 U203 ( .A(\A_s[26] ), .ZN(n562) );
  INV_X1 U204 ( .A(\A_s[27] ), .ZN(n563) );
  INV_X1 U205 ( .A(\A_s[28] ), .ZN(n564) );
  INV_X1 U206 ( .A(\A_s[29] ), .ZN(n565) );
  INV_X1 U207 ( .A(n567), .ZN(A_so[32]) );
  INV_X1 U208 ( .A(A_s[30]), .ZN(n567) );
  INV_X1 U209 ( .A(\A_s[31] ), .ZN(n568) );
  INV_X1 U210 ( .A(\A_s[32] ), .ZN(n569) );
  INV_X1 U211 ( .A(\A_s[33] ), .ZN(n570) );
endmodule


module BOOTHENC_NBIT38_i4 ( A_s, A_ns, B, O, A_so, A_nso );
  input [37:0] A_s;
  input [37:0] A_ns;
  input [37:0] B;
  output [37:0] O;
  output [37:0] A_so;
  output [37:0] A_nso;
  wire   \A_s[35] , \A_s[34] , \A_s[33] , \A_s[32] , \A_s[31] , \A_s[30] ,
         \A_s[29] , \A_s[28] , \A_s[27] , \A_s[26] , \A_s[25] , \A_s[24] ,
         \A_s[23] , \A_s[22] , \A_s[21] , \A_s[20] , \A_s[19] , \A_s[18] ,
         \A_s[17] , \A_s[16] , \A_s[15] , \A_s[14] , \A_s[13] , \A_s[12] ,
         \A_s[11] , \A_s[10] , \A_s[9] , \A_s[8] , \A_s[7] , \A_s[6] ,
         \A_s[5] , \A_s[4] , \A_s[3] , \A_s[2] , \A_s[1] , \A_s[0] ,
         \A_ns[35] , \A_ns[34] , \A_ns[33] , \A_ns[32] , \A_ns[31] ,
         \A_ns[30] , \A_ns[29] , \A_ns[28] , \A_ns[27] , \A_ns[26] ,
         \A_ns[25] , \A_ns[24] , \A_ns[23] , \A_ns[22] , \A_ns[21] ,
         \A_ns[20] , \A_ns[19] , \A_ns[18] , \A_ns[17] , \A_ns[16] ,
         \A_ns[15] , \A_ns[14] , \A_ns[13] , \A_ns[12] , \A_ns[11] ,
         \A_ns[10] , \A_ns[9] , \A_ns[8] , \A_ns[7] , \A_ns[6] , \A_ns[5] ,
         \A_ns[4] , \A_ns[3] , \A_ns[2] , \A_ns[1] , \A_ns[0] , n77, n78, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n562, n564, n566, n569, n571, n573,
         n575, n577, n579, n581, n583, n585, n587, n589, n591, n593, n595,
         n597, n599, n601, n603, n605, n607, n609, n611, n613, n615, n617,
         n619, n621, n623, n625, n627, n628, n629, n630, n631, n632;
  assign A_nso[0] = 1'b0;
  assign A_nso[1] = 1'b0;
  assign A_so[0] = 1'b0;
  assign A_so[1] = 1'b0;
  assign O[0] = 1'b0;
  assign A_so[37] = \A_s[35] ;
  assign \A_s[35]  = A_s[35];
  assign A_so[36] = \A_s[34] ;
  assign \A_s[34]  = A_s[34];
  assign A_so[35] = \A_s[33] ;
  assign \A_s[33]  = A_s[33];
  assign A_so[34] = \A_s[32] ;
  assign \A_s[32]  = A_s[32];
  assign A_so[33] = \A_s[31] ;
  assign \A_s[31]  = A_s[31];
  assign A_so[32] = \A_s[30] ;
  assign \A_s[30]  = A_s[30];
  assign A_so[31] = \A_s[29] ;
  assign \A_s[29]  = A_s[29];
  assign A_so[30] = \A_s[28] ;
  assign \A_s[28]  = A_s[28];
  assign A_so[29] = \A_s[27] ;
  assign \A_s[27]  = A_s[27];
  assign A_so[28] = \A_s[26] ;
  assign \A_s[26]  = A_s[26];
  assign A_so[27] = \A_s[25] ;
  assign \A_s[25]  = A_s[25];
  assign A_so[26] = \A_s[24] ;
  assign \A_s[24]  = A_s[24];
  assign A_so[25] = \A_s[23] ;
  assign \A_s[23]  = A_s[23];
  assign A_so[24] = \A_s[22] ;
  assign \A_s[22]  = A_s[22];
  assign A_so[23] = \A_s[21] ;
  assign \A_s[21]  = A_s[21];
  assign A_so[22] = \A_s[20] ;
  assign \A_s[20]  = A_s[20];
  assign A_so[21] = \A_s[19] ;
  assign \A_s[19]  = A_s[19];
  assign A_so[20] = \A_s[18] ;
  assign \A_s[18]  = A_s[18];
  assign A_so[19] = \A_s[17] ;
  assign \A_s[17]  = A_s[17];
  assign A_so[18] = \A_s[16] ;
  assign \A_s[16]  = A_s[16];
  assign A_so[17] = \A_s[15] ;
  assign \A_s[15]  = A_s[15];
  assign A_so[16] = \A_s[14] ;
  assign \A_s[14]  = A_s[14];
  assign A_so[15] = \A_s[13] ;
  assign \A_s[13]  = A_s[13];
  assign A_so[14] = \A_s[12] ;
  assign \A_s[12]  = A_s[12];
  assign A_so[13] = \A_s[11] ;
  assign \A_s[11]  = A_s[11];
  assign A_so[12] = \A_s[10] ;
  assign \A_s[10]  = A_s[10];
  assign A_so[11] = \A_s[9] ;
  assign \A_s[9]  = A_s[9];
  assign A_so[10] = \A_s[8] ;
  assign \A_s[8]  = A_s[8];
  assign A_so[9] = \A_s[7] ;
  assign \A_s[7]  = A_s[7];
  assign A_so[8] = \A_s[6] ;
  assign \A_s[6]  = A_s[6];
  assign A_so[7] = \A_s[5] ;
  assign \A_s[5]  = A_s[5];
  assign A_so[6] = \A_s[4] ;
  assign \A_s[4]  = A_s[4];
  assign A_so[5] = \A_s[3] ;
  assign \A_s[3]  = A_s[3];
  assign A_so[4] = \A_s[2] ;
  assign \A_s[2]  = A_s[2];
  assign A_so[3] = \A_s[1] ;
  assign \A_s[1]  = A_s[1];
  assign A_so[2] = \A_s[0] ;
  assign \A_s[0]  = A_s[0];
  assign A_nso[37] = \A_ns[35] ;
  assign \A_ns[35]  = A_ns[35];
  assign A_nso[36] = \A_ns[34] ;
  assign \A_ns[34]  = A_ns[34];
  assign A_nso[35] = \A_ns[33] ;
  assign \A_ns[33]  = A_ns[33];
  assign A_nso[34] = \A_ns[32] ;
  assign \A_ns[32]  = A_ns[32];
  assign A_nso[33] = \A_ns[31] ;
  assign \A_ns[31]  = A_ns[31];
  assign A_nso[32] = \A_ns[30] ;
  assign \A_ns[30]  = A_ns[30];
  assign A_nso[31] = \A_ns[29] ;
  assign \A_ns[29]  = A_ns[29];
  assign A_nso[30] = \A_ns[28] ;
  assign \A_ns[28]  = A_ns[28];
  assign A_nso[29] = \A_ns[27] ;
  assign \A_ns[27]  = A_ns[27];
  assign A_nso[28] = \A_ns[26] ;
  assign \A_ns[26]  = A_ns[26];
  assign A_nso[27] = \A_ns[25] ;
  assign \A_ns[25]  = A_ns[25];
  assign A_nso[26] = \A_ns[24] ;
  assign \A_ns[24]  = A_ns[24];
  assign A_nso[25] = \A_ns[23] ;
  assign \A_ns[23]  = A_ns[23];
  assign A_nso[24] = \A_ns[22] ;
  assign \A_ns[22]  = A_ns[22];
  assign A_nso[23] = \A_ns[21] ;
  assign \A_ns[21]  = A_ns[21];
  assign A_nso[22] = \A_ns[20] ;
  assign \A_ns[20]  = A_ns[20];
  assign A_nso[21] = \A_ns[19] ;
  assign \A_ns[19]  = A_ns[19];
  assign A_nso[20] = \A_ns[18] ;
  assign \A_ns[18]  = A_ns[18];
  assign A_nso[19] = \A_ns[17] ;
  assign \A_ns[17]  = A_ns[17];
  assign A_nso[18] = \A_ns[16] ;
  assign \A_ns[16]  = A_ns[16];
  assign A_nso[17] = \A_ns[15] ;
  assign \A_ns[15]  = A_ns[15];
  assign A_nso[16] = \A_ns[14] ;
  assign \A_ns[14]  = A_ns[14];
  assign A_nso[15] = \A_ns[13] ;
  assign \A_ns[13]  = A_ns[13];
  assign A_nso[14] = \A_ns[12] ;
  assign \A_ns[12]  = A_ns[12];
  assign A_nso[13] = \A_ns[11] ;
  assign \A_ns[11]  = A_ns[11];
  assign A_nso[12] = \A_ns[10] ;
  assign \A_ns[10]  = A_ns[10];
  assign A_nso[11] = \A_ns[9] ;
  assign \A_ns[9]  = A_ns[9];
  assign A_nso[10] = \A_ns[8] ;
  assign \A_ns[8]  = A_ns[8];
  assign A_nso[9] = \A_ns[7] ;
  assign \A_ns[7]  = A_ns[7];
  assign A_nso[8] = \A_ns[6] ;
  assign \A_ns[6]  = A_ns[6];
  assign A_nso[7] = \A_ns[5] ;
  assign \A_ns[5]  = A_ns[5];
  assign A_nso[6] = \A_ns[4] ;
  assign \A_ns[4]  = A_ns[4];
  assign A_nso[5] = \A_ns[3] ;
  assign \A_ns[3]  = A_ns[3];
  assign A_nso[4] = \A_ns[2] ;
  assign \A_ns[2]  = A_ns[2];
  assign A_nso[3] = \A_ns[1] ;
  assign \A_ns[1]  = A_ns[1];
  assign A_nso[2] = \A_ns[0] ;
  assign \A_ns[0]  = A_ns[0];

  NAND3_X1 U154 ( .A1(B[3]), .A2(n632), .A3(B[4]), .ZN(n77) );
  XOR2_X1 U155 ( .A(B[3]), .B(B[4]), .Z(n152) );
  CLKBUF_X1 U2 ( .A(n630), .Z(n551) );
  CLKBUF_X1 U3 ( .A(n631), .Z(n554) );
  CLKBUF_X1 U4 ( .A(n630), .Z(n550) );
  CLKBUF_X1 U5 ( .A(n631), .Z(n553) );
  CLKBUF_X1 U6 ( .A(n629), .Z(n548) );
  CLKBUF_X1 U7 ( .A(n629), .Z(n549) );
  BUF_X1 U8 ( .A(n631), .Z(n555) );
  BUF_X1 U9 ( .A(n630), .Z(n552) );
  INV_X1 U10 ( .A(\A_ns[35] ), .ZN(n558) );
  BUF_X1 U11 ( .A(n629), .Z(n547) );
  INV_X1 U12 ( .A(n109), .ZN(O[22]) );
  INV_X1 U13 ( .A(n83), .ZN(O[35]) );
  AOI221_X1 U14 ( .B1(n553), .B2(\A_ns[34] ), .C1(n550), .C2(\A_s[34] ), .A(
        n569), .ZN(n83) );
  INV_X1 U15 ( .A(n87), .ZN(O[33]) );
  AOI221_X1 U16 ( .B1(n553), .B2(\A_ns[32] ), .C1(n550), .C2(\A_s[32] ), .A(
        n573), .ZN(n87) );
  INV_X1 U17 ( .A(n89), .ZN(O[32]) );
  AOI221_X1 U18 ( .B1(n553), .B2(\A_ns[31] ), .C1(n550), .C2(\A_s[31] ), .A(
        n575), .ZN(n89) );
  INV_X1 U19 ( .A(n90), .ZN(n575) );
  INV_X1 U20 ( .A(n127), .ZN(O[13]) );
  INV_X1 U21 ( .A(n81), .ZN(n630) );
  INV_X1 U22 ( .A(n80), .ZN(n631) );
  INV_X1 U23 ( .A(n141), .ZN(O[6]) );
  AOI221_X1 U24 ( .B1(n555), .B2(\A_ns[5] ), .C1(n552), .C2(\A_s[5] ), .A(n627), .ZN(n141) );
  INV_X1 U25 ( .A(n142), .ZN(n627) );
  AOI22_X1 U26 ( .A1(\A_ns[4] ), .A2(n556), .B1(\A_s[4] ), .B2(n547), .ZN(n142) );
  INV_X1 U27 ( .A(n125), .ZN(O[14]) );
  AOI221_X1 U28 ( .B1(n554), .B2(\A_ns[13] ), .C1(n551), .C2(\A_s[13] ), .A(
        n611), .ZN(n125) );
  INV_X1 U29 ( .A(n126), .ZN(n611) );
  AOI22_X1 U30 ( .A1(\A_ns[12] ), .A2(n557), .B1(\A_s[12] ), .B2(n548), .ZN(
        n126) );
  AOI221_X1 U31 ( .B1(n554), .B2(\A_ns[12] ), .C1(n551), .C2(\A_s[12] ), .A(
        n613), .ZN(n127) );
  INV_X1 U32 ( .A(n128), .ZN(n613) );
  AOI22_X1 U33 ( .A1(\A_ns[11] ), .A2(n556), .B1(\A_s[11] ), .B2(n547), .ZN(
        n128) );
  INV_X1 U34 ( .A(n119), .ZN(O[17]) );
  AOI221_X1 U35 ( .B1(n554), .B2(\A_ns[16] ), .C1(n551), .C2(\A_s[16] ), .A(
        n605), .ZN(n119) );
  INV_X1 U36 ( .A(n120), .ZN(n605) );
  AOI22_X1 U37 ( .A1(\A_ns[15] ), .A2(n557), .B1(\A_s[15] ), .B2(n548), .ZN(
        n120) );
  INV_X1 U38 ( .A(n123), .ZN(O[15]) );
  AOI221_X1 U39 ( .B1(n554), .B2(\A_ns[14] ), .C1(n551), .C2(\A_s[14] ), .A(
        n609), .ZN(n123) );
  INV_X1 U40 ( .A(n124), .ZN(n609) );
  AOI22_X1 U41 ( .A1(\A_ns[13] ), .A2(n557), .B1(\A_s[13] ), .B2(n548), .ZN(
        n124) );
  INV_X1 U42 ( .A(n139), .ZN(O[7]) );
  AOI221_X1 U43 ( .B1(n555), .B2(\A_ns[6] ), .C1(n552), .C2(\A_s[6] ), .A(n625), .ZN(n139) );
  INV_X1 U44 ( .A(n140), .ZN(n625) );
  AOI22_X1 U45 ( .A1(\A_ns[5] ), .A2(n556), .B1(\A_s[5] ), .B2(n547), .ZN(n140) );
  INV_X1 U46 ( .A(n115), .ZN(O[19]) );
  AOI221_X1 U47 ( .B1(n554), .B2(\A_ns[18] ), .C1(n551), .C2(\A_s[18] ), .A(
        n601), .ZN(n115) );
  INV_X1 U48 ( .A(n116), .ZN(n601) );
  AOI22_X1 U49 ( .A1(\A_ns[17] ), .A2(n557), .B1(\A_s[17] ), .B2(n548), .ZN(
        n116) );
  INV_X1 U50 ( .A(n117), .ZN(O[18]) );
  AOI221_X1 U51 ( .B1(n554), .B2(\A_ns[17] ), .C1(n551), .C2(\A_s[17] ), .A(
        n603), .ZN(n117) );
  INV_X1 U52 ( .A(n118), .ZN(n603) );
  AOI22_X1 U53 ( .A1(\A_ns[16] ), .A2(n557), .B1(\A_s[16] ), .B2(n548), .ZN(
        n118) );
  INV_X1 U54 ( .A(n137), .ZN(O[8]) );
  AOI221_X1 U55 ( .B1(n555), .B2(\A_ns[7] ), .C1(n552), .C2(\A_s[7] ), .A(n623), .ZN(n137) );
  INV_X1 U56 ( .A(n138), .ZN(n623) );
  AOI22_X1 U57 ( .A1(\A_ns[6] ), .A2(n556), .B1(\A_s[6] ), .B2(n547), .ZN(n138) );
  INV_X1 U58 ( .A(n133), .ZN(O[10]) );
  AOI221_X1 U59 ( .B1(n555), .B2(\A_ns[9] ), .C1(n552), .C2(\A_s[9] ), .A(n619), .ZN(n133) );
  INV_X1 U60 ( .A(n134), .ZN(n619) );
  AOI22_X1 U61 ( .A1(\A_ns[8] ), .A2(n556), .B1(\A_s[8] ), .B2(n547), .ZN(n134) );
  INV_X1 U62 ( .A(n129), .ZN(O[12]) );
  AOI221_X1 U63 ( .B1(n554), .B2(\A_ns[11] ), .C1(n552), .C2(\A_s[11] ), .A(
        n615), .ZN(n129) );
  INV_X1 U64 ( .A(n130), .ZN(n615) );
  AOI22_X1 U65 ( .A1(\A_ns[10] ), .A2(n556), .B1(\A_s[10] ), .B2(n547), .ZN(
        n130) );
  INV_X1 U66 ( .A(n113), .ZN(O[20]) );
  AOI221_X1 U67 ( .B1(n554), .B2(\A_ns[19] ), .C1(n551), .C2(\A_s[19] ), .A(
        n599), .ZN(n113) );
  INV_X1 U68 ( .A(n114), .ZN(n599) );
  AOI22_X1 U69 ( .A1(\A_ns[18] ), .A2(n557), .B1(\A_s[18] ), .B2(n548), .ZN(
        n114) );
  INV_X1 U70 ( .A(n135), .ZN(O[9]) );
  AOI221_X1 U71 ( .B1(n555), .B2(\A_ns[8] ), .C1(n552), .C2(\A_s[8] ), .A(n621), .ZN(n135) );
  INV_X1 U72 ( .A(n136), .ZN(n621) );
  AOI22_X1 U73 ( .A1(\A_ns[7] ), .A2(n556), .B1(\A_s[7] ), .B2(n547), .ZN(n136) );
  INV_X1 U74 ( .A(n131), .ZN(O[11]) );
  AOI221_X1 U75 ( .B1(n554), .B2(\A_ns[10] ), .C1(n552), .C2(\A_s[10] ), .A(
        n617), .ZN(n131) );
  INV_X1 U76 ( .A(n132), .ZN(n617) );
  AOI22_X1 U77 ( .A1(\A_ns[9] ), .A2(n556), .B1(\A_s[9] ), .B2(n547), .ZN(n132) );
  INV_X1 U78 ( .A(n121), .ZN(O[16]) );
  AOI221_X1 U79 ( .B1(n554), .B2(\A_ns[15] ), .C1(n551), .C2(\A_s[15] ), .A(
        n607), .ZN(n121) );
  INV_X1 U80 ( .A(n122), .ZN(n607) );
  AOI22_X1 U81 ( .A1(\A_ns[14] ), .A2(n557), .B1(\A_s[14] ), .B2(n548), .ZN(
        n122) );
  AOI221_X1 U82 ( .B1(n554), .B2(\A_ns[21] ), .C1(n551), .C2(\A_s[21] ), .A(
        n595), .ZN(n109) );
  INV_X1 U83 ( .A(n110), .ZN(n595) );
  AOI22_X1 U84 ( .A1(\A_ns[20] ), .A2(n557), .B1(\A_s[20] ), .B2(n548), .ZN(
        n110) );
  AOI22_X1 U85 ( .A1(\A_ns[28] ), .A2(n557), .B1(\A_s[28] ), .B2(n549), .ZN(
        n94) );
  AOI22_X1 U86 ( .A1(\A_ns[30] ), .A2(n557), .B1(\A_s[30] ), .B2(n549), .ZN(
        n90) );
  INV_X1 U87 ( .A(n107), .ZN(O[23]) );
  AOI221_X1 U88 ( .B1(n554), .B2(\A_ns[22] ), .C1(n551), .C2(\A_s[22] ), .A(
        n593), .ZN(n107) );
  INV_X1 U89 ( .A(n108), .ZN(n593) );
  AOI22_X1 U90 ( .A1(\A_ns[21] ), .A2(n557), .B1(\A_s[21] ), .B2(n548), .ZN(
        n108) );
  INV_X1 U91 ( .A(n101), .ZN(O[26]) );
  AOI221_X1 U92 ( .B1(n553), .B2(\A_ns[25] ), .C1(n550), .C2(\A_s[25] ), .A(
        n587), .ZN(n101) );
  INV_X1 U93 ( .A(n102), .ZN(n587) );
  AOI22_X1 U94 ( .A1(\A_ns[24] ), .A2(n557), .B1(\A_s[24] ), .B2(n549), .ZN(
        n102) );
  INV_X1 U95 ( .A(n103), .ZN(O[25]) );
  AOI221_X1 U96 ( .B1(n553), .B2(\A_ns[24] ), .C1(n550), .C2(\A_s[24] ), .A(
        n589), .ZN(n103) );
  INV_X1 U97 ( .A(n104), .ZN(n589) );
  AOI22_X1 U98 ( .A1(\A_ns[23] ), .A2(n557), .B1(\A_s[23] ), .B2(n548), .ZN(
        n104) );
  INV_X1 U99 ( .A(n99), .ZN(O[27]) );
  AOI221_X1 U100 ( .B1(n553), .B2(\A_ns[26] ), .C1(n550), .C2(\A_s[26] ), .A(
        n585), .ZN(n99) );
  INV_X1 U101 ( .A(n100), .ZN(n585) );
  AOI22_X1 U102 ( .A1(\A_ns[25] ), .A2(n557), .B1(\A_s[25] ), .B2(n549), .ZN(
        n100) );
  INV_X1 U103 ( .A(n105), .ZN(O[24]) );
  AOI221_X1 U104 ( .B1(n553), .B2(\A_ns[23] ), .C1(n551), .C2(\A_s[23] ), .A(
        n591), .ZN(n105) );
  INV_X1 U105 ( .A(n106), .ZN(n591) );
  AOI22_X1 U106 ( .A1(\A_ns[22] ), .A2(n557), .B1(\A_s[22] ), .B2(n548), .ZN(
        n106) );
  INV_X1 U107 ( .A(n97), .ZN(O[28]) );
  AOI221_X1 U108 ( .B1(n553), .B2(\A_ns[27] ), .C1(n551), .C2(\A_s[27] ), .A(
        n583), .ZN(n97) );
  INV_X1 U109 ( .A(n98), .ZN(n583) );
  AOI22_X1 U110 ( .A1(\A_ns[26] ), .A2(n557), .B1(\A_s[26] ), .B2(n549), .ZN(
        n98) );
  INV_X1 U111 ( .A(n92), .ZN(n577) );
  AOI22_X1 U112 ( .A1(\A_ns[29] ), .A2(n557), .B1(\A_s[29] ), .B2(n549), .ZN(
        n92) );
  INV_X1 U113 ( .A(n96), .ZN(n581) );
  AOI22_X1 U114 ( .A1(\A_ns[27] ), .A2(n557), .B1(\A_s[27] ), .B2(n549), .ZN(
        n96) );
  INV_X1 U115 ( .A(n111), .ZN(O[21]) );
  AOI221_X1 U116 ( .B1(n554), .B2(\A_ns[20] ), .C1(n551), .C2(\A_s[20] ), .A(
        n597), .ZN(n111) );
  INV_X1 U117 ( .A(n112), .ZN(n597) );
  AOI22_X1 U118 ( .A1(\A_ns[19] ), .A2(n557), .B1(\A_s[19] ), .B2(n548), .ZN(
        n112) );
  OAI221_X1 U119 ( .B1(n558), .B2(n80), .C1(n559), .C2(n81), .A(n82), .ZN(
        O[36]) );
  AOI22_X1 U120 ( .A1(\A_ns[34] ), .A2(n557), .B1(\A_s[34] ), .B2(n549), .ZN(
        n82) );
  AOI22_X1 U121 ( .A1(A_ns[36]), .A2(n553), .B1(A_s[36]), .B2(n550), .ZN(n78)
         );
  INV_X1 U122 ( .A(n85), .ZN(O[34]) );
  AOI221_X1 U123 ( .B1(n553), .B2(\A_ns[33] ), .C1(n550), .C2(\A_s[33] ), .A(
        n571), .ZN(n85) );
  INV_X1 U124 ( .A(n86), .ZN(n571) );
  AOI22_X1 U125 ( .A1(\A_ns[32] ), .A2(n557), .B1(\A_s[32] ), .B2(n549), .ZN(
        n86) );
  INV_X1 U126 ( .A(n84), .ZN(n569) );
  AOI22_X1 U127 ( .A1(\A_ns[33] ), .A2(n557), .B1(\A_s[33] ), .B2(n549), .ZN(
        n84) );
  INV_X1 U128 ( .A(n88), .ZN(n573) );
  AOI22_X1 U129 ( .A1(\A_ns[31] ), .A2(n557), .B1(\A_s[31] ), .B2(n549), .ZN(
        n88) );
  INV_X1 U130 ( .A(\A_s[35] ), .ZN(n559) );
  OAI221_X1 U131 ( .B1(n546), .B2(n558), .C1(n77), .C2(n559), .A(n78), .ZN(
        O[37]) );
  INV_X1 U132 ( .A(n546), .ZN(n556) );
  NAND2_X1 U133 ( .A1(n152), .A2(n632), .ZN(n81) );
  NAND2_X1 U134 ( .A1(n152), .A2(n81), .ZN(n80) );
  INV_X1 U135 ( .A(n77), .ZN(n629) );
  INV_X1 U136 ( .A(n91), .ZN(O[31]) );
  AOI221_X1 U137 ( .B1(n553), .B2(\A_ns[30] ), .C1(n550), .C2(\A_s[30] ), .A(
        n577), .ZN(n91) );
  INV_X1 U138 ( .A(n93), .ZN(O[30]) );
  AOI221_X1 U139 ( .B1(n553), .B2(\A_ns[29] ), .C1(n550), .C2(\A_s[29] ), .A(
        n579), .ZN(n93) );
  INV_X1 U140 ( .A(n94), .ZN(n579) );
  INV_X1 U141 ( .A(n95), .ZN(O[29]) );
  AOI221_X1 U142 ( .B1(n553), .B2(\A_ns[28] ), .C1(n550), .C2(\A_s[28] ), .A(
        n581), .ZN(n95) );
  INV_X1 U143 ( .A(n546), .ZN(n557) );
  OR3_X1 U144 ( .A1(B[3]), .A2(B[4]), .A3(n632), .ZN(n546) );
  INV_X1 U145 ( .A(n145), .ZN(O[4]) );
  AOI221_X1 U146 ( .B1(n555), .B2(\A_ns[3] ), .C1(n552), .C2(\A_s[3] ), .A(
        n566), .ZN(n145) );
  INV_X1 U147 ( .A(n146), .ZN(n566) );
  AOI22_X1 U148 ( .A1(\A_ns[2] ), .A2(n556), .B1(\A_s[2] ), .B2(n547), .ZN(
        n146) );
  INV_X1 U149 ( .A(B[5]), .ZN(n632) );
  INV_X1 U150 ( .A(n143), .ZN(O[5]) );
  AOI221_X1 U151 ( .B1(n555), .B2(\A_ns[4] ), .C1(n552), .C2(\A_s[4] ), .A(
        n628), .ZN(n143) );
  INV_X1 U152 ( .A(n144), .ZN(n628) );
  AOI22_X1 U153 ( .A1(\A_ns[3] ), .A2(n556), .B1(\A_s[3] ), .B2(n547), .ZN(
        n144) );
  INV_X1 U156 ( .A(n147), .ZN(O[3]) );
  AOI221_X1 U157 ( .B1(n555), .B2(\A_ns[2] ), .C1(n552), .C2(\A_s[2] ), .A(
        n564), .ZN(n147) );
  INV_X1 U158 ( .A(n151), .ZN(O[1]) );
  AOI22_X1 U159 ( .A1(n550), .A2(\A_s[0] ), .B1(n555), .B2(\A_ns[0] ), .ZN(
        n151) );
  INV_X1 U160 ( .A(n149), .ZN(O[2]) );
  AOI221_X1 U161 ( .B1(n555), .B2(\A_ns[1] ), .C1(n550), .C2(\A_s[1] ), .A(
        n562), .ZN(n149) );
  INV_X1 U162 ( .A(n150), .ZN(n562) );
  AOI22_X1 U163 ( .A1(\A_ns[0] ), .A2(n556), .B1(\A_s[0] ), .B2(n547), .ZN(
        n150) );
  INV_X1 U164 ( .A(n148), .ZN(n564) );
  AOI22_X1 U165 ( .A1(\A_ns[1] ), .A2(n556), .B1(\A_s[1] ), .B2(n547), .ZN(
        n148) );
endmodule


module BOOTHENC_NBIT40_i6 ( A_s, A_ns, B, O, A_so, A_nso );
  input [39:0] A_s;
  input [39:0] A_ns;
  input [39:0] B;
  output [39:0] O;
  output [39:0] A_so;
  output [39:0] A_nso;
  wire   \A_s[37] , \A_s[36] , \A_s[35] , \A_s[34] , \A_s[33] , \A_s[32] ,
         \A_s[31] , \A_s[30] , \A_s[29] , \A_s[28] , \A_s[27] , \A_s[26] ,
         \A_s[25] , \A_s[24] , \A_s[23] , \A_s[22] , \A_s[21] , \A_s[20] ,
         \A_s[19] , \A_s[18] , \A_s[17] , \A_s[16] , \A_s[15] , \A_s[14] ,
         \A_s[13] , \A_s[12] , \A_s[11] , \A_s[10] , \A_s[9] , \A_s[8] ,
         \A_s[7] , \A_s[6] , \A_s[5] , \A_s[4] , \A_s[3] , \A_s[2] , \A_s[1] ,
         \A_s[0] , \A_ns[37] , \A_ns[36] , \A_ns[35] , \A_ns[34] , \A_ns[33] ,
         \A_ns[32] , \A_ns[31] , \A_ns[30] , \A_ns[29] , \A_ns[28] ,
         \A_ns[27] , \A_ns[26] , \A_ns[25] , \A_ns[24] , \A_ns[23] ,
         \A_ns[22] , \A_ns[21] , \A_ns[20] , \A_ns[19] , \A_ns[18] ,
         \A_ns[17] , \A_ns[16] , \A_ns[15] , \A_ns[14] , \A_ns[13] ,
         \A_ns[12] , \A_ns[11] , \A_ns[10] , \A_ns[9] , \A_ns[8] , \A_ns[7] ,
         \A_ns[6] , \A_ns[5] , \A_ns[4] , \A_ns[3] , \A_ns[2] , \A_ns[1] ,
         \A_ns[0] , n81, n82, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n596, n598, n600, n602, n604, n607, n609, n611,
         n613, n615, n617, n619, n621, n623, n625, n627, n629, n631, n633,
         n635, n637, n639, n641, n643, n645, n647, n649, n651, n653, n655,
         n657, n659, n661, n663, n665, n666, n667, n668, n669, n670;
  assign A_nso[0] = 1'b0;
  assign A_nso[1] = 1'b0;
  assign A_so[0] = 1'b0;
  assign A_so[1] = 1'b0;
  assign O[0] = 1'b0;
  assign A_so[39] = \A_s[37] ;
  assign \A_s[37]  = A_s[37];
  assign A_so[38] = \A_s[36] ;
  assign \A_s[36]  = A_s[36];
  assign A_so[37] = \A_s[35] ;
  assign \A_s[35]  = A_s[35];
  assign A_so[36] = \A_s[34] ;
  assign \A_s[34]  = A_s[34];
  assign A_so[35] = \A_s[33] ;
  assign \A_s[33]  = A_s[33];
  assign A_so[34] = \A_s[32] ;
  assign \A_s[32]  = A_s[32];
  assign A_so[33] = \A_s[31] ;
  assign \A_s[31]  = A_s[31];
  assign A_so[32] = \A_s[30] ;
  assign \A_s[30]  = A_s[30];
  assign A_so[31] = \A_s[29] ;
  assign \A_s[29]  = A_s[29];
  assign A_so[30] = \A_s[28] ;
  assign \A_s[28]  = A_s[28];
  assign A_so[29] = \A_s[27] ;
  assign \A_s[27]  = A_s[27];
  assign A_so[28] = \A_s[26] ;
  assign \A_s[26]  = A_s[26];
  assign A_so[27] = \A_s[25] ;
  assign \A_s[25]  = A_s[25];
  assign A_so[26] = \A_s[24] ;
  assign \A_s[24]  = A_s[24];
  assign A_so[25] = \A_s[23] ;
  assign \A_s[23]  = A_s[23];
  assign A_so[24] = \A_s[22] ;
  assign \A_s[22]  = A_s[22];
  assign A_so[23] = \A_s[21] ;
  assign \A_s[21]  = A_s[21];
  assign A_so[22] = \A_s[20] ;
  assign \A_s[20]  = A_s[20];
  assign A_so[21] = \A_s[19] ;
  assign \A_s[19]  = A_s[19];
  assign A_so[20] = \A_s[18] ;
  assign \A_s[18]  = A_s[18];
  assign A_so[19] = \A_s[17] ;
  assign \A_s[17]  = A_s[17];
  assign A_so[18] = \A_s[16] ;
  assign \A_s[16]  = A_s[16];
  assign A_so[17] = \A_s[15] ;
  assign \A_s[15]  = A_s[15];
  assign A_so[16] = \A_s[14] ;
  assign \A_s[14]  = A_s[14];
  assign A_so[15] = \A_s[13] ;
  assign \A_s[13]  = A_s[13];
  assign A_so[14] = \A_s[12] ;
  assign \A_s[12]  = A_s[12];
  assign A_so[13] = \A_s[11] ;
  assign \A_s[11]  = A_s[11];
  assign A_so[12] = \A_s[10] ;
  assign \A_s[10]  = A_s[10];
  assign A_so[11] = \A_s[9] ;
  assign \A_s[9]  = A_s[9];
  assign A_so[10] = \A_s[8] ;
  assign \A_s[8]  = A_s[8];
  assign A_so[9] = \A_s[7] ;
  assign \A_s[7]  = A_s[7];
  assign A_so[8] = \A_s[6] ;
  assign \A_s[6]  = A_s[6];
  assign A_so[7] = \A_s[5] ;
  assign \A_s[5]  = A_s[5];
  assign A_so[6] = \A_s[4] ;
  assign \A_s[4]  = A_s[4];
  assign A_so[5] = \A_s[3] ;
  assign \A_s[3]  = A_s[3];
  assign A_so[4] = \A_s[2] ;
  assign \A_s[2]  = A_s[2];
  assign A_so[3] = \A_s[1] ;
  assign \A_s[1]  = A_s[1];
  assign A_so[2] = \A_s[0] ;
  assign \A_s[0]  = A_s[0];
  assign A_nso[39] = \A_ns[37] ;
  assign \A_ns[37]  = A_ns[37];
  assign A_nso[38] = \A_ns[36] ;
  assign \A_ns[36]  = A_ns[36];
  assign A_nso[37] = \A_ns[35] ;
  assign \A_ns[35]  = A_ns[35];
  assign A_nso[36] = \A_ns[34] ;
  assign \A_ns[34]  = A_ns[34];
  assign A_nso[35] = \A_ns[33] ;
  assign \A_ns[33]  = A_ns[33];
  assign A_nso[34] = \A_ns[32] ;
  assign \A_ns[32]  = A_ns[32];
  assign A_nso[33] = \A_ns[31] ;
  assign \A_ns[31]  = A_ns[31];
  assign A_nso[32] = \A_ns[30] ;
  assign \A_ns[30]  = A_ns[30];
  assign A_nso[31] = \A_ns[29] ;
  assign \A_ns[29]  = A_ns[29];
  assign A_nso[30] = \A_ns[28] ;
  assign \A_ns[28]  = A_ns[28];
  assign A_nso[29] = \A_ns[27] ;
  assign \A_ns[27]  = A_ns[27];
  assign A_nso[28] = \A_ns[26] ;
  assign \A_ns[26]  = A_ns[26];
  assign A_nso[27] = \A_ns[25] ;
  assign \A_ns[25]  = A_ns[25];
  assign A_nso[26] = \A_ns[24] ;
  assign \A_ns[24]  = A_ns[24];
  assign A_nso[25] = \A_ns[23] ;
  assign \A_ns[23]  = A_ns[23];
  assign A_nso[24] = \A_ns[22] ;
  assign \A_ns[22]  = A_ns[22];
  assign A_nso[23] = \A_ns[21] ;
  assign \A_ns[21]  = A_ns[21];
  assign A_nso[22] = \A_ns[20] ;
  assign \A_ns[20]  = A_ns[20];
  assign A_nso[21] = \A_ns[19] ;
  assign \A_ns[19]  = A_ns[19];
  assign A_nso[20] = \A_ns[18] ;
  assign \A_ns[18]  = A_ns[18];
  assign A_nso[19] = \A_ns[17] ;
  assign \A_ns[17]  = A_ns[17];
  assign A_nso[18] = \A_ns[16] ;
  assign \A_ns[16]  = A_ns[16];
  assign A_nso[17] = \A_ns[15] ;
  assign \A_ns[15]  = A_ns[15];
  assign A_nso[16] = \A_ns[14] ;
  assign \A_ns[14]  = A_ns[14];
  assign A_nso[15] = \A_ns[13] ;
  assign \A_ns[13]  = A_ns[13];
  assign A_nso[14] = \A_ns[12] ;
  assign \A_ns[12]  = A_ns[12];
  assign A_nso[13] = \A_ns[11] ;
  assign \A_ns[11]  = A_ns[11];
  assign A_nso[12] = \A_ns[10] ;
  assign \A_ns[10]  = A_ns[10];
  assign A_nso[11] = \A_ns[9] ;
  assign \A_ns[9]  = A_ns[9];
  assign A_nso[10] = \A_ns[8] ;
  assign \A_ns[8]  = A_ns[8];
  assign A_nso[9] = \A_ns[7] ;
  assign \A_ns[7]  = A_ns[7];
  assign A_nso[8] = \A_ns[6] ;
  assign \A_ns[6]  = A_ns[6];
  assign A_nso[7] = \A_ns[5] ;
  assign \A_ns[5]  = A_ns[5];
  assign A_nso[6] = \A_ns[4] ;
  assign \A_ns[4]  = A_ns[4];
  assign A_nso[5] = \A_ns[3] ;
  assign \A_ns[3]  = A_ns[3];
  assign A_nso[4] = \A_ns[2] ;
  assign \A_ns[2]  = A_ns[2];
  assign A_nso[3] = \A_ns[1] ;
  assign \A_ns[1]  = A_ns[1];
  assign A_nso[2] = \A_ns[0] ;
  assign \A_ns[0]  = A_ns[0];

  NAND3_X1 U162 ( .A1(B[5]), .A2(n670), .A3(B[6]), .ZN(n81) );
  XOR2_X1 U163 ( .A(B[5]), .B(B[6]), .Z(n160) );
  AOI22_X1 U2 ( .A1(A_ns[38]), .A2(n587), .B1(A_s[38]), .B2(n584), .ZN(n82) );
  OAI221_X4 U3 ( .B1(n580), .B2(n592), .C1(n81), .C2(n593), .A(n82), .ZN(O[39]) );
  CLKBUF_X1 U4 ( .A(n668), .Z(n585) );
  CLKBUF_X1 U5 ( .A(n669), .Z(n588) );
  CLKBUF_X1 U6 ( .A(n668), .Z(n584) );
  CLKBUF_X1 U7 ( .A(n669), .Z(n587) );
  CLKBUF_X1 U8 ( .A(n667), .Z(n582) );
  CLKBUF_X1 U9 ( .A(n667), .Z(n583) );
  INV_X1 U10 ( .A(\A_ns[37] ), .ZN(n592) );
  INV_X1 U11 ( .A(\A_s[37] ), .ZN(n593) );
  INV_X1 U12 ( .A(n109), .ZN(O[26]) );
  INV_X1 U13 ( .A(n123), .ZN(O[19]) );
  INV_X1 U14 ( .A(n119), .ZN(O[21]) );
  BUF_X1 U15 ( .A(n669), .Z(n589) );
  BUF_X1 U16 ( .A(n668), .Z(n586) );
  INV_X1 U17 ( .A(n97), .ZN(O[32]) );
  AOI221_X1 U18 ( .B1(n587), .B2(\A_ns[31] ), .C1(n584), .C2(\A_s[31] ), .A(
        n617), .ZN(n97) );
  INV_X1 U19 ( .A(n89), .ZN(O[36]) );
  AOI221_X1 U20 ( .B1(n587), .B2(\A_ns[35] ), .C1(n584), .C2(\A_s[35] ), .A(
        n609), .ZN(n89) );
  INV_X1 U21 ( .A(n93), .ZN(O[34]) );
  AOI221_X1 U22 ( .B1(n587), .B2(\A_ns[33] ), .C1(n584), .C2(\A_s[33] ), .A(
        n613), .ZN(n93) );
  INV_X1 U23 ( .A(n91), .ZN(O[35]) );
  AOI221_X1 U24 ( .B1(n587), .B2(\A_ns[34] ), .C1(n584), .C2(\A_s[34] ), .A(
        n611), .ZN(n91) );
  INV_X1 U25 ( .A(n92), .ZN(n611) );
  INV_X1 U26 ( .A(n103), .ZN(O[29]) );
  AOI221_X1 U27 ( .B1(n587), .B2(\A_ns[28] ), .C1(n584), .C2(\A_s[28] ), .A(
        n623), .ZN(n103) );
  INV_X1 U28 ( .A(n104), .ZN(n623) );
  INV_X1 U29 ( .A(n95), .ZN(O[33]) );
  AOI221_X1 U30 ( .B1(n587), .B2(\A_ns[32] ), .C1(n584), .C2(\A_s[32] ), .A(
        n615), .ZN(n95) );
  INV_X1 U31 ( .A(n96), .ZN(n615) );
  INV_X1 U32 ( .A(n105), .ZN(O[28]) );
  AOI221_X1 U33 ( .B1(n587), .B2(\A_ns[27] ), .C1(n584), .C2(\A_s[27] ), .A(
        n625), .ZN(n105) );
  INV_X1 U34 ( .A(n107), .ZN(O[27]) );
  AOI221_X1 U35 ( .B1(n587), .B2(\A_ns[26] ), .C1(n584), .C2(\A_s[26] ), .A(
        n627), .ZN(n107) );
  INV_X1 U36 ( .A(n87), .ZN(O[37]) );
  AOI221_X1 U37 ( .B1(n587), .B2(\A_ns[36] ), .C1(n584), .C2(\A_s[36] ), .A(
        n607), .ZN(n87) );
  INV_X1 U38 ( .A(n88), .ZN(n607) );
  INV_X1 U39 ( .A(n139), .ZN(O[11]) );
  AOI221_X1 U40 ( .B1(n589), .B2(\A_ns[10] ), .C1(n586), .C2(\A_s[10] ), .A(
        n659), .ZN(n139) );
  INV_X1 U41 ( .A(n140), .ZN(n659) );
  AOI22_X1 U42 ( .A1(\A_ns[9] ), .A2(n590), .B1(\A_s[9] ), .B2(n581), .ZN(n140) );
  INV_X1 U43 ( .A(n133), .ZN(O[14]) );
  AOI221_X1 U44 ( .B1(n588), .B2(\A_ns[13] ), .C1(n586), .C2(\A_s[13] ), .A(
        n653), .ZN(n133) );
  INV_X1 U45 ( .A(n134), .ZN(n653) );
  AOI22_X1 U46 ( .A1(\A_ns[12] ), .A2(n591), .B1(\A_s[12] ), .B2(n582), .ZN(
        n134) );
  BUF_X1 U47 ( .A(n667), .Z(n581) );
  INV_X1 U48 ( .A(n85), .ZN(n668) );
  INV_X1 U49 ( .A(n84), .ZN(n669) );
  INV_X1 U50 ( .A(n143), .ZN(O[9]) );
  AOI221_X1 U51 ( .B1(n589), .B2(\A_ns[8] ), .C1(n586), .C2(\A_s[8] ), .A(n663), .ZN(n143) );
  INV_X1 U52 ( .A(n144), .ZN(n663) );
  AOI22_X1 U53 ( .A1(\A_ns[7] ), .A2(n590), .B1(\A_s[7] ), .B2(n581), .ZN(n144) );
  INV_X1 U54 ( .A(n131), .ZN(O[15]) );
  AOI221_X1 U55 ( .B1(n588), .B2(\A_ns[14] ), .C1(n585), .C2(\A_s[14] ), .A(
        n651), .ZN(n131) );
  INV_X1 U56 ( .A(n132), .ZN(n651) );
  AOI22_X1 U57 ( .A1(\A_ns[13] ), .A2(n591), .B1(\A_s[13] ), .B2(n582), .ZN(
        n132) );
  INV_X1 U58 ( .A(n145), .ZN(O[8]) );
  AOI221_X1 U59 ( .B1(n589), .B2(\A_ns[7] ), .C1(n586), .C2(\A_s[7] ), .A(n665), .ZN(n145) );
  INV_X1 U60 ( .A(n146), .ZN(n665) );
  AOI22_X1 U61 ( .A1(\A_ns[6] ), .A2(n590), .B1(\A_s[6] ), .B2(n581), .ZN(n146) );
  INV_X1 U62 ( .A(n141), .ZN(O[10]) );
  AOI221_X1 U63 ( .B1(n589), .B2(\A_ns[9] ), .C1(n586), .C2(\A_s[9] ), .A(n661), .ZN(n141) );
  INV_X1 U64 ( .A(n142), .ZN(n661) );
  AOI22_X1 U65 ( .A1(\A_ns[8] ), .A2(n590), .B1(\A_s[8] ), .B2(n581), .ZN(n142) );
  INV_X1 U66 ( .A(n127), .ZN(O[17]) );
  AOI221_X1 U67 ( .B1(n588), .B2(\A_ns[16] ), .C1(n585), .C2(\A_s[16] ), .A(
        n647), .ZN(n127) );
  INV_X1 U68 ( .A(n128), .ZN(n647) );
  AOI22_X1 U69 ( .A1(\A_ns[15] ), .A2(n591), .B1(\A_s[15] ), .B2(n582), .ZN(
        n128) );
  INV_X1 U70 ( .A(n137), .ZN(O[12]) );
  AOI221_X1 U71 ( .B1(n589), .B2(\A_ns[11] ), .C1(n586), .C2(\A_s[11] ), .A(
        n657), .ZN(n137) );
  INV_X1 U72 ( .A(n138), .ZN(n657) );
  AOI22_X1 U73 ( .A1(\A_ns[10] ), .A2(n590), .B1(\A_s[10] ), .B2(n581), .ZN(
        n138) );
  INV_X1 U74 ( .A(n135), .ZN(O[13]) );
  AOI221_X1 U75 ( .B1(n588), .B2(\A_ns[12] ), .C1(n586), .C2(\A_s[12] ), .A(
        n655), .ZN(n135) );
  INV_X1 U76 ( .A(n136), .ZN(n655) );
  AOI22_X1 U77 ( .A1(\A_ns[11] ), .A2(n590), .B1(\A_s[11] ), .B2(n581), .ZN(
        n136) );
  INV_X1 U78 ( .A(n129), .ZN(O[16]) );
  AOI221_X1 U79 ( .B1(n588), .B2(\A_ns[15] ), .C1(n585), .C2(\A_s[15] ), .A(
        n649), .ZN(n129) );
  INV_X1 U80 ( .A(n130), .ZN(n649) );
  AOI22_X1 U81 ( .A1(\A_ns[14] ), .A2(n591), .B1(\A_s[14] ), .B2(n582), .ZN(
        n130) );
  AOI221_X1 U82 ( .B1(n587), .B2(\A_ns[25] ), .C1(n585), .C2(\A_s[25] ), .A(
        n629), .ZN(n109) );
  INV_X1 U83 ( .A(n110), .ZN(n629) );
  AOI22_X1 U84 ( .A1(\A_ns[24] ), .A2(n591), .B1(\A_s[24] ), .B2(n583), .ZN(
        n110) );
  AOI221_X1 U85 ( .B1(n588), .B2(\A_ns[20] ), .C1(n585), .C2(\A_s[20] ), .A(
        n639), .ZN(n119) );
  INV_X1 U86 ( .A(n120), .ZN(n639) );
  AOI22_X1 U87 ( .A1(\A_ns[19] ), .A2(n591), .B1(\A_s[19] ), .B2(n582), .ZN(
        n120) );
  AOI221_X1 U88 ( .B1(n588), .B2(\A_ns[18] ), .C1(n585), .C2(\A_s[18] ), .A(
        n643), .ZN(n123) );
  INV_X1 U89 ( .A(n124), .ZN(n643) );
  AOI22_X1 U90 ( .A1(\A_ns[17] ), .A2(n591), .B1(\A_s[17] ), .B2(n582), .ZN(
        n124) );
  AOI22_X1 U91 ( .A1(\A_ns[27] ), .A2(n591), .B1(\A_s[27] ), .B2(n583), .ZN(
        n104) );
  INV_X1 U92 ( .A(n117), .ZN(O[22]) );
  AOI221_X1 U93 ( .B1(n588), .B2(\A_ns[21] ), .C1(n585), .C2(\A_s[21] ), .A(
        n637), .ZN(n117) );
  INV_X1 U94 ( .A(n118), .ZN(n637) );
  AOI22_X1 U95 ( .A1(\A_ns[20] ), .A2(n591), .B1(\A_s[20] ), .B2(n582), .ZN(
        n118) );
  INV_X1 U96 ( .A(n125), .ZN(O[18]) );
  AOI221_X1 U97 ( .B1(n588), .B2(\A_ns[17] ), .C1(n585), .C2(\A_s[17] ), .A(
        n645), .ZN(n125) );
  INV_X1 U98 ( .A(n126), .ZN(n645) );
  AOI22_X1 U99 ( .A1(\A_ns[16] ), .A2(n591), .B1(\A_s[16] ), .B2(n582), .ZN(
        n126) );
  INV_X1 U100 ( .A(n111), .ZN(O[25]) );
  AOI221_X1 U101 ( .B1(n588), .B2(\A_ns[24] ), .C1(n585), .C2(\A_s[24] ), .A(
        n631), .ZN(n111) );
  INV_X1 U102 ( .A(n112), .ZN(n631) );
  AOI22_X1 U103 ( .A1(\A_ns[23] ), .A2(n591), .B1(\A_s[23] ), .B2(n582), .ZN(
        n112) );
  INV_X1 U104 ( .A(n108), .ZN(n627) );
  AOI22_X1 U105 ( .A1(\A_ns[25] ), .A2(n591), .B1(\A_s[25] ), .B2(n583), .ZN(
        n108) );
  INV_X1 U106 ( .A(n101), .ZN(O[30]) );
  AOI221_X1 U107 ( .B1(n587), .B2(\A_ns[29] ), .C1(n585), .C2(\A_s[29] ), .A(
        n621), .ZN(n101) );
  INV_X1 U108 ( .A(n102), .ZN(n621) );
  AOI22_X1 U109 ( .A1(\A_ns[28] ), .A2(n591), .B1(\A_s[28] ), .B2(n583), .ZN(
        n102) );
  INV_X1 U110 ( .A(n121), .ZN(O[20]) );
  AOI221_X1 U111 ( .B1(n588), .B2(\A_ns[19] ), .C1(n585), .C2(\A_s[19] ), .A(
        n641), .ZN(n121) );
  INV_X1 U112 ( .A(n122), .ZN(n641) );
  AOI22_X1 U113 ( .A1(\A_ns[18] ), .A2(n591), .B1(\A_s[18] ), .B2(n582), .ZN(
        n122) );
  INV_X1 U114 ( .A(n106), .ZN(n625) );
  AOI22_X1 U115 ( .A1(\A_ns[26] ), .A2(n591), .B1(\A_s[26] ), .B2(n583), .ZN(
        n106) );
  INV_X1 U116 ( .A(n115), .ZN(O[23]) );
  AOI221_X1 U117 ( .B1(n588), .B2(\A_ns[22] ), .C1(n585), .C2(\A_s[22] ), .A(
        n635), .ZN(n115) );
  INV_X1 U118 ( .A(n116), .ZN(n635) );
  AOI22_X1 U119 ( .A1(\A_ns[21] ), .A2(n591), .B1(\A_s[21] ), .B2(n582), .ZN(
        n116) );
  INV_X1 U120 ( .A(n113), .ZN(O[24]) );
  AOI221_X1 U121 ( .B1(n588), .B2(\A_ns[23] ), .C1(n585), .C2(\A_s[23] ), .A(
        n633), .ZN(n113) );
  INV_X1 U122 ( .A(n114), .ZN(n633) );
  AOI22_X1 U123 ( .A1(\A_ns[22] ), .A2(n591), .B1(\A_s[22] ), .B2(n582), .ZN(
        n114) );
  AOI22_X1 U124 ( .A1(\A_ns[35] ), .A2(n591), .B1(\A_s[35] ), .B2(n583), .ZN(
        n88) );
  AOI22_X1 U125 ( .A1(\A_ns[33] ), .A2(n591), .B1(\A_s[33] ), .B2(n583), .ZN(
        n92) );
  AOI22_X1 U126 ( .A1(\A_ns[31] ), .A2(n591), .B1(\A_s[31] ), .B2(n583), .ZN(
        n96) );
  INV_X1 U127 ( .A(n99), .ZN(O[31]) );
  AOI221_X1 U128 ( .B1(n587), .B2(\A_ns[30] ), .C1(n584), .C2(\A_s[30] ), .A(
        n619), .ZN(n99) );
  INV_X1 U129 ( .A(n100), .ZN(n619) );
  AOI22_X1 U130 ( .A1(\A_ns[29] ), .A2(n591), .B1(\A_s[29] ), .B2(n583), .ZN(
        n100) );
  INV_X1 U131 ( .A(n90), .ZN(n609) );
  AOI22_X1 U132 ( .A1(\A_ns[34] ), .A2(n591), .B1(\A_s[34] ), .B2(n583), .ZN(
        n90) );
  INV_X1 U133 ( .A(n94), .ZN(n613) );
  AOI22_X1 U134 ( .A1(\A_ns[32] ), .A2(n591), .B1(\A_s[32] ), .B2(n583), .ZN(
        n94) );
  INV_X1 U135 ( .A(n98), .ZN(n617) );
  AOI22_X1 U136 ( .A1(\A_ns[30] ), .A2(n591), .B1(\A_s[30] ), .B2(n583), .ZN(
        n98) );
  OAI221_X1 U137 ( .B1(n592), .B2(n84), .C1(n593), .C2(n85), .A(n86), .ZN(
        O[38]) );
  AOI22_X1 U138 ( .A1(\A_ns[36] ), .A2(n591), .B1(\A_s[36] ), .B2(n583), .ZN(
        n86) );
  INV_X1 U139 ( .A(n580), .ZN(n590) );
  NAND2_X1 U140 ( .A1(n160), .A2(n670), .ZN(n85) );
  INV_X1 U141 ( .A(n81), .ZN(n667) );
  NAND2_X1 U142 ( .A1(n160), .A2(n85), .ZN(n84) );
  INV_X1 U143 ( .A(n580), .ZN(n591) );
  OR3_X1 U144 ( .A1(B[5]), .A2(B[6]), .A3(n670), .ZN(n580) );
  INV_X1 U145 ( .A(n149), .ZN(O[6]) );
  AOI221_X1 U146 ( .B1(n589), .B2(\A_ns[5] ), .C1(n586), .C2(\A_s[5] ), .A(
        n604), .ZN(n149) );
  INV_X1 U147 ( .A(n150), .ZN(n604) );
  AOI22_X1 U148 ( .A1(\A_ns[4] ), .A2(n590), .B1(\A_s[4] ), .B2(n581), .ZN(
        n150) );
  INV_X1 U149 ( .A(B[7]), .ZN(n670) );
  INV_X1 U150 ( .A(n147), .ZN(O[7]) );
  AOI221_X1 U151 ( .B1(n589), .B2(\A_ns[6] ), .C1(n586), .C2(\A_s[6] ), .A(
        n666), .ZN(n147) );
  INV_X1 U152 ( .A(n148), .ZN(n666) );
  AOI22_X1 U153 ( .A1(\A_ns[5] ), .A2(n590), .B1(\A_s[5] ), .B2(n581), .ZN(
        n148) );
  INV_X1 U154 ( .A(n159), .ZN(O[1]) );
  AOI22_X1 U155 ( .A1(n584), .A2(\A_s[0] ), .B1(n589), .B2(\A_ns[0] ), .ZN(
        n159) );
  INV_X1 U156 ( .A(n151), .ZN(O[5]) );
  AOI221_X1 U157 ( .B1(n589), .B2(\A_ns[4] ), .C1(n586), .C2(\A_s[4] ), .A(
        n602), .ZN(n151) );
  INV_X1 U158 ( .A(n155), .ZN(O[3]) );
  AOI221_X1 U159 ( .B1(n589), .B2(\A_ns[2] ), .C1(n586), .C2(\A_s[2] ), .A(
        n598), .ZN(n155) );
  INV_X1 U160 ( .A(n156), .ZN(n598) );
  INV_X1 U161 ( .A(n153), .ZN(O[4]) );
  AOI221_X1 U164 ( .B1(n589), .B2(\A_ns[3] ), .C1(n586), .C2(\A_s[3] ), .A(
        n600), .ZN(n153) );
  INV_X1 U165 ( .A(n157), .ZN(O[2]) );
  AOI221_X1 U166 ( .B1(n589), .B2(\A_ns[1] ), .C1(n584), .C2(\A_s[1] ), .A(
        n596), .ZN(n157) );
  INV_X1 U167 ( .A(n158), .ZN(n596) );
  INV_X1 U168 ( .A(n154), .ZN(n600) );
  AOI22_X1 U169 ( .A1(\A_ns[2] ), .A2(n590), .B1(\A_s[2] ), .B2(n581), .ZN(
        n154) );
  INV_X1 U170 ( .A(n152), .ZN(n602) );
  AOI22_X1 U171 ( .A1(\A_ns[3] ), .A2(n590), .B1(\A_s[3] ), .B2(n581), .ZN(
        n152) );
  AOI22_X1 U172 ( .A1(\A_ns[0] ), .A2(n590), .B1(\A_s[0] ), .B2(n581), .ZN(
        n158) );
  AOI22_X1 U173 ( .A1(\A_ns[1] ), .A2(n590), .B1(\A_s[1] ), .B2(n581), .ZN(
        n156) );
endmodule


module BOOTHENC_NBIT42_i8 ( A_s, A_ns, B, O, A_so, A_nso );
  input [41:0] A_s;
  input [41:0] A_ns;
  input [41:0] B;
  output [41:0] O;
  output [41:0] A_so;
  output [41:0] A_nso;
  wire   \A_s[39] , \A_s[38] , \A_s[37] , \A_s[36] , \A_s[35] , \A_s[34] ,
         \A_s[33] , \A_s[32] , \A_s[31] , \A_s[30] , \A_s[29] , \A_s[28] ,
         \A_s[27] , \A_s[26] , \A_s[25] , \A_s[24] , \A_s[23] , \A_s[22] ,
         \A_s[21] , \A_s[20] , \A_s[19] , \A_s[18] , \A_s[17] , \A_s[16] ,
         \A_s[15] , \A_s[14] , \A_s[13] , \A_s[12] , \A_s[11] , \A_s[10] ,
         \A_s[9] , \A_s[8] , \A_s[7] , \A_s[6] , \A_s[5] , \A_s[4] , \A_s[3] ,
         \A_s[2] , \A_s[1] , \A_s[0] , \A_ns[39] , \A_ns[38] , \A_ns[37] ,
         \A_ns[36] , \A_ns[35] , \A_ns[34] , \A_ns[33] , \A_ns[32] ,
         \A_ns[31] , \A_ns[30] , \A_ns[29] , \A_ns[28] , \A_ns[27] ,
         \A_ns[26] , \A_ns[25] , \A_ns[24] , \A_ns[23] , \A_ns[22] ,
         \A_ns[21] , \A_ns[20] , \A_ns[19] , \A_ns[18] , \A_ns[17] ,
         \A_ns[16] , \A_ns[15] , \A_ns[14] , \A_ns[13] , \A_ns[12] ,
         \A_ns[11] , \A_ns[10] , \A_ns[9] , \A_ns[8] , \A_ns[7] , \A_ns[6] ,
         \A_ns[5] , \A_ns[4] , \A_ns[3] , \A_ns[2] , \A_ns[1] , \A_ns[0] , n85,
         n86, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n633, n635,
         n637, n639, n641, n643, n645, n648, n650, n652, n654, n656, n658,
         n660, n662, n664, n666, n668, n670, n672, n674, n676, n678, n680,
         n682, n684, n686, n688, n690, n692, n694, n696, n698, n700, n702,
         n704, n706, n707, n708, n709, n710, n711;
  assign A_nso[0] = 1'b0;
  assign A_nso[1] = 1'b0;
  assign A_so[0] = 1'b0;
  assign A_so[1] = 1'b0;
  assign O[0] = 1'b0;
  assign A_so[41] = \A_s[39] ;
  assign \A_s[39]  = A_s[39];
  assign A_so[40] = \A_s[38] ;
  assign \A_s[38]  = A_s[38];
  assign A_so[39] = \A_s[37] ;
  assign \A_s[37]  = A_s[37];
  assign A_so[38] = \A_s[36] ;
  assign \A_s[36]  = A_s[36];
  assign A_so[37] = \A_s[35] ;
  assign \A_s[35]  = A_s[35];
  assign A_so[36] = \A_s[34] ;
  assign \A_s[34]  = A_s[34];
  assign A_so[35] = \A_s[33] ;
  assign \A_s[33]  = A_s[33];
  assign A_so[34] = \A_s[32] ;
  assign \A_s[32]  = A_s[32];
  assign A_so[33] = \A_s[31] ;
  assign \A_s[31]  = A_s[31];
  assign A_so[32] = \A_s[30] ;
  assign \A_s[30]  = A_s[30];
  assign A_so[31] = \A_s[29] ;
  assign \A_s[29]  = A_s[29];
  assign A_so[30] = \A_s[28] ;
  assign \A_s[28]  = A_s[28];
  assign A_so[29] = \A_s[27] ;
  assign \A_s[27]  = A_s[27];
  assign A_so[28] = \A_s[26] ;
  assign \A_s[26]  = A_s[26];
  assign A_so[27] = \A_s[25] ;
  assign \A_s[25]  = A_s[25];
  assign A_so[26] = \A_s[24] ;
  assign \A_s[24]  = A_s[24];
  assign A_so[25] = \A_s[23] ;
  assign \A_s[23]  = A_s[23];
  assign A_so[24] = \A_s[22] ;
  assign \A_s[22]  = A_s[22];
  assign A_so[23] = \A_s[21] ;
  assign \A_s[21]  = A_s[21];
  assign A_so[22] = \A_s[20] ;
  assign \A_s[20]  = A_s[20];
  assign A_so[21] = \A_s[19] ;
  assign \A_s[19]  = A_s[19];
  assign A_so[20] = \A_s[18] ;
  assign \A_s[18]  = A_s[18];
  assign A_so[19] = \A_s[17] ;
  assign \A_s[17]  = A_s[17];
  assign A_so[18] = \A_s[16] ;
  assign \A_s[16]  = A_s[16];
  assign A_so[17] = \A_s[15] ;
  assign \A_s[15]  = A_s[15];
  assign A_so[16] = \A_s[14] ;
  assign \A_s[14]  = A_s[14];
  assign A_so[15] = \A_s[13] ;
  assign \A_s[13]  = A_s[13];
  assign A_so[14] = \A_s[12] ;
  assign \A_s[12]  = A_s[12];
  assign A_so[13] = \A_s[11] ;
  assign \A_s[11]  = A_s[11];
  assign A_so[12] = \A_s[10] ;
  assign \A_s[10]  = A_s[10];
  assign A_so[11] = \A_s[9] ;
  assign \A_s[9]  = A_s[9];
  assign A_so[10] = \A_s[8] ;
  assign \A_s[8]  = A_s[8];
  assign A_so[9] = \A_s[7] ;
  assign \A_s[7]  = A_s[7];
  assign A_so[8] = \A_s[6] ;
  assign \A_s[6]  = A_s[6];
  assign A_so[7] = \A_s[5] ;
  assign \A_s[5]  = A_s[5];
  assign A_so[6] = \A_s[4] ;
  assign \A_s[4]  = A_s[4];
  assign A_so[5] = \A_s[3] ;
  assign \A_s[3]  = A_s[3];
  assign A_so[4] = \A_s[2] ;
  assign \A_s[2]  = A_s[2];
  assign A_so[3] = \A_s[1] ;
  assign \A_s[1]  = A_s[1];
  assign A_so[2] = \A_s[0] ;
  assign \A_s[0]  = A_s[0];
  assign A_nso[41] = \A_ns[39] ;
  assign \A_ns[39]  = A_ns[39];
  assign A_nso[40] = \A_ns[38] ;
  assign \A_ns[38]  = A_ns[38];
  assign A_nso[39] = \A_ns[37] ;
  assign \A_ns[37]  = A_ns[37];
  assign A_nso[38] = \A_ns[36] ;
  assign \A_ns[36]  = A_ns[36];
  assign A_nso[37] = \A_ns[35] ;
  assign \A_ns[35]  = A_ns[35];
  assign A_nso[36] = \A_ns[34] ;
  assign \A_ns[34]  = A_ns[34];
  assign A_nso[35] = \A_ns[33] ;
  assign \A_ns[33]  = A_ns[33];
  assign A_nso[34] = \A_ns[32] ;
  assign \A_ns[32]  = A_ns[32];
  assign A_nso[33] = \A_ns[31] ;
  assign \A_ns[31]  = A_ns[31];
  assign A_nso[32] = \A_ns[30] ;
  assign \A_ns[30]  = A_ns[30];
  assign A_nso[31] = \A_ns[29] ;
  assign \A_ns[29]  = A_ns[29];
  assign A_nso[30] = \A_ns[28] ;
  assign \A_ns[28]  = A_ns[28];
  assign A_nso[29] = \A_ns[27] ;
  assign \A_ns[27]  = A_ns[27];
  assign A_nso[28] = \A_ns[26] ;
  assign \A_ns[26]  = A_ns[26];
  assign A_nso[27] = \A_ns[25] ;
  assign \A_ns[25]  = A_ns[25];
  assign A_nso[26] = \A_ns[24] ;
  assign \A_ns[24]  = A_ns[24];
  assign A_nso[25] = \A_ns[23] ;
  assign \A_ns[23]  = A_ns[23];
  assign A_nso[24] = \A_ns[22] ;
  assign \A_ns[22]  = A_ns[22];
  assign A_nso[23] = \A_ns[21] ;
  assign \A_ns[21]  = A_ns[21];
  assign A_nso[22] = \A_ns[20] ;
  assign \A_ns[20]  = A_ns[20];
  assign A_nso[21] = \A_ns[19] ;
  assign \A_ns[19]  = A_ns[19];
  assign A_nso[20] = \A_ns[18] ;
  assign \A_ns[18]  = A_ns[18];
  assign A_nso[19] = \A_ns[17] ;
  assign \A_ns[17]  = A_ns[17];
  assign A_nso[18] = \A_ns[16] ;
  assign \A_ns[16]  = A_ns[16];
  assign A_nso[17] = \A_ns[15] ;
  assign \A_ns[15]  = A_ns[15];
  assign A_nso[16] = \A_ns[14] ;
  assign \A_ns[14]  = A_ns[14];
  assign A_nso[15] = \A_ns[13] ;
  assign \A_ns[13]  = A_ns[13];
  assign A_nso[14] = \A_ns[12] ;
  assign \A_ns[12]  = A_ns[12];
  assign A_nso[13] = \A_ns[11] ;
  assign \A_ns[11]  = A_ns[11];
  assign A_nso[12] = \A_ns[10] ;
  assign \A_ns[10]  = A_ns[10];
  assign A_nso[11] = \A_ns[9] ;
  assign \A_ns[9]  = A_ns[9];
  assign A_nso[10] = \A_ns[8] ;
  assign \A_ns[8]  = A_ns[8];
  assign A_nso[9] = \A_ns[7] ;
  assign \A_ns[7]  = A_ns[7];
  assign A_nso[8] = \A_ns[6] ;
  assign \A_ns[6]  = A_ns[6];
  assign A_nso[7] = \A_ns[5] ;
  assign \A_ns[5]  = A_ns[5];
  assign A_nso[6] = \A_ns[4] ;
  assign \A_ns[4]  = A_ns[4];
  assign A_nso[5] = \A_ns[3] ;
  assign \A_ns[3]  = A_ns[3];
  assign A_nso[4] = \A_ns[2] ;
  assign \A_ns[2]  = A_ns[2];
  assign A_nso[3] = \A_ns[1] ;
  assign \A_ns[1]  = A_ns[1];
  assign A_nso[2] = \A_ns[0] ;
  assign \A_ns[0]  = A_ns[0];

  NAND3_X1 U170 ( .A1(B[7]), .A2(n711), .A3(B[8]), .ZN(n85) );
  XOR2_X1 U171 ( .A(B[7]), .B(B[8]), .Z(n168) );
  CLKBUF_X1 U2 ( .A(n615), .Z(n619) );
  CLKBUF_X1 U3 ( .A(n709), .Z(n621) );
  CLKBUF_X1 U4 ( .A(n710), .Z(n624) );
  CLKBUF_X1 U5 ( .A(n614), .Z(n617) );
  CLKBUF_X1 U6 ( .A(n709), .Z(n620) );
  CLKBUF_X1 U7 ( .A(n710), .Z(n623) );
  CLKBUF_X1 U8 ( .A(n708), .Z(n615) );
  INV_X1 U9 ( .A(\A_ns[39] ), .ZN(n629) );
  INV_X1 U10 ( .A(\A_s[39] ), .ZN(n630) );
  AOI22_X1 U11 ( .A1(A_ns[40]), .A2(n623), .B1(A_s[40]), .B2(n620), .ZN(n86)
         );
  INV_X1 U12 ( .A(n119), .ZN(O[25]) );
  BUF_X1 U13 ( .A(n710), .Z(n625) );
  BUF_X1 U14 ( .A(n709), .Z(n622) );
  BUF_X1 U15 ( .A(n614), .Z(n616) );
  BUF_X1 U16 ( .A(n615), .Z(n618) );
  INV_X1 U17 ( .A(n109), .ZN(O[30]) );
  AOI221_X1 U18 ( .B1(n623), .B2(\A_ns[29] ), .C1(n621), .C2(\A_s[29] ), .A(
        n666), .ZN(n109) );
  INV_X1 U19 ( .A(n99), .ZN(O[35]) );
  AOI221_X1 U20 ( .B1(n623), .B2(\A_ns[34] ), .C1(n620), .C2(\A_s[34] ), .A(
        n656), .ZN(n99) );
  INV_X1 U21 ( .A(n100), .ZN(n656) );
  INV_X1 U22 ( .A(n111), .ZN(O[29]) );
  AOI221_X1 U23 ( .B1(n623), .B2(\A_ns[28] ), .C1(n620), .C2(\A_s[28] ), .A(
        n668), .ZN(n111) );
  INV_X1 U24 ( .A(n112), .ZN(n668) );
  INV_X1 U25 ( .A(n107), .ZN(O[31]) );
  AOI221_X1 U26 ( .B1(n623), .B2(\A_ns[30] ), .C1(n620), .C2(\A_s[30] ), .A(
        n664), .ZN(n107) );
  INV_X1 U27 ( .A(n103), .ZN(O[33]) );
  AOI221_X1 U28 ( .B1(n623), .B2(\A_ns[32] ), .C1(n620), .C2(\A_s[32] ), .A(
        n660), .ZN(n103) );
  INV_X1 U29 ( .A(n95), .ZN(O[37]) );
  AOI221_X1 U30 ( .B1(n623), .B2(\A_ns[36] ), .C1(n620), .C2(\A_s[36] ), .A(
        n652), .ZN(n95) );
  INV_X1 U31 ( .A(n96), .ZN(n652) );
  INV_X1 U32 ( .A(n113), .ZN(O[28]) );
  AOI221_X1 U33 ( .B1(n623), .B2(\A_ns[27] ), .C1(n621), .C2(\A_s[27] ), .A(
        n670), .ZN(n113) );
  INV_X1 U34 ( .A(n114), .ZN(n670) );
  INV_X1 U35 ( .A(n97), .ZN(O[36]) );
  AOI221_X1 U36 ( .B1(n623), .B2(\A_ns[35] ), .C1(n620), .C2(\A_s[35] ), .A(
        n654), .ZN(n97) );
  INV_X1 U37 ( .A(n98), .ZN(n654) );
  INV_X1 U38 ( .A(n101), .ZN(O[34]) );
  AOI221_X1 U39 ( .B1(n623), .B2(\A_ns[33] ), .C1(n620), .C2(\A_s[33] ), .A(
        n658), .ZN(n101) );
  INV_X1 U40 ( .A(n102), .ZN(n658) );
  INV_X1 U41 ( .A(n115), .ZN(O[27]) );
  AOI221_X1 U42 ( .B1(n624), .B2(\A_ns[26] ), .C1(n621), .C2(\A_s[26] ), .A(
        n672), .ZN(n115) );
  INV_X1 U43 ( .A(n125), .ZN(O[22]) );
  AOI221_X1 U44 ( .B1(n624), .B2(\A_ns[21] ), .C1(n621), .C2(\A_s[21] ), .A(
        n682), .ZN(n125) );
  INV_X1 U45 ( .A(n93), .ZN(O[38]) );
  AOI221_X1 U46 ( .B1(n623), .B2(\A_ns[37] ), .C1(n620), .C2(\A_s[37] ), .A(
        n650), .ZN(n93) );
  INV_X1 U47 ( .A(n94), .ZN(n650) );
  INV_X1 U48 ( .A(n123), .ZN(O[23]) );
  AOI221_X1 U49 ( .B1(n624), .B2(\A_ns[22] ), .C1(n621), .C2(\A_s[22] ), .A(
        n680), .ZN(n123) );
  INV_X1 U50 ( .A(n127), .ZN(O[21]) );
  AOI221_X1 U51 ( .B1(n624), .B2(\A_ns[20] ), .C1(n621), .C2(\A_s[20] ), .A(
        n684), .ZN(n127) );
  INV_X1 U52 ( .A(n89), .ZN(n709) );
  INV_X1 U53 ( .A(n88), .ZN(n710) );
  INV_X1 U54 ( .A(n145), .ZN(O[12]) );
  AOI221_X1 U55 ( .B1(n625), .B2(\A_ns[11] ), .C1(n622), .C2(\A_s[11] ), .A(
        n702), .ZN(n145) );
  INV_X1 U56 ( .A(n146), .ZN(n702) );
  AOI22_X1 U57 ( .A1(\A_ns[10] ), .A2(n626), .B1(\A_s[10] ), .B2(n616), .ZN(
        n146) );
  INV_X1 U58 ( .A(n149), .ZN(O[10]) );
  AOI221_X1 U59 ( .B1(n625), .B2(\A_ns[9] ), .C1(n622), .C2(\A_s[9] ), .A(n706), .ZN(n149) );
  INV_X1 U60 ( .A(n150), .ZN(n706) );
  AOI22_X1 U61 ( .A1(\A_ns[8] ), .A2(n626), .B1(\A_s[8] ), .B2(n616), .ZN(n150) );
  INV_X1 U62 ( .A(n143), .ZN(O[13]) );
  AOI221_X1 U63 ( .B1(n625), .B2(\A_ns[12] ), .C1(n622), .C2(\A_s[12] ), .A(
        n700), .ZN(n143) );
  INV_X1 U64 ( .A(n144), .ZN(n700) );
  AOI22_X1 U65 ( .A1(\A_ns[11] ), .A2(n626), .B1(\A_s[11] ), .B2(n616), .ZN(
        n144) );
  INV_X1 U66 ( .A(n147), .ZN(O[11]) );
  AOI221_X1 U67 ( .B1(n625), .B2(\A_ns[10] ), .C1(n622), .C2(\A_s[10] ), .A(
        n704), .ZN(n147) );
  INV_X1 U68 ( .A(n148), .ZN(n704) );
  AOI22_X1 U69 ( .A1(\A_ns[9] ), .A2(n626), .B1(\A_s[9] ), .B2(n616), .ZN(n148) );
  BUF_X1 U70 ( .A(n708), .Z(n614) );
  INV_X1 U71 ( .A(n141), .ZN(O[14]) );
  AOI221_X1 U72 ( .B1(n625), .B2(\A_ns[13] ), .C1(n622), .C2(\A_s[13] ), .A(
        n698), .ZN(n141) );
  INV_X1 U73 ( .A(n142), .ZN(n698) );
  AOI22_X1 U74 ( .A1(\A_ns[12] ), .A2(n627), .B1(\A_s[12] ), .B2(n617), .ZN(
        n142) );
  AOI221_X1 U75 ( .B1(n624), .B2(\A_ns[24] ), .C1(n621), .C2(\A_s[24] ), .A(
        n676), .ZN(n119) );
  INV_X1 U76 ( .A(n120), .ZN(n676) );
  AOI22_X1 U77 ( .A1(\A_ns[23] ), .A2(n627), .B1(\A_s[23] ), .B2(n617), .ZN(
        n120) );
  INV_X1 U78 ( .A(n137), .ZN(O[16]) );
  AOI221_X1 U79 ( .B1(n624), .B2(\A_ns[15] ), .C1(n622), .C2(\A_s[15] ), .A(
        n694), .ZN(n137) );
  INV_X1 U80 ( .A(n138), .ZN(n694) );
  AOI22_X1 U81 ( .A1(\A_ns[14] ), .A2(n627), .B1(\A_s[14] ), .B2(n617), .ZN(
        n138) );
  INV_X1 U82 ( .A(n135), .ZN(O[17]) );
  AOI221_X1 U83 ( .B1(n624), .B2(\A_ns[16] ), .C1(n621), .C2(\A_s[16] ), .A(
        n692), .ZN(n135) );
  INV_X1 U84 ( .A(n136), .ZN(n692) );
  AOI22_X1 U85 ( .A1(\A_ns[15] ), .A2(n627), .B1(\A_s[15] ), .B2(n617), .ZN(
        n136) );
  INV_X1 U86 ( .A(n131), .ZN(O[19]) );
  AOI221_X1 U87 ( .B1(n624), .B2(\A_ns[18] ), .C1(n621), .C2(\A_s[18] ), .A(
        n688), .ZN(n131) );
  INV_X1 U88 ( .A(n132), .ZN(n688) );
  AOI22_X1 U89 ( .A1(\A_ns[17] ), .A2(n627), .B1(\A_s[17] ), .B2(n617), .ZN(
        n132) );
  INV_X1 U90 ( .A(n121), .ZN(O[24]) );
  AOI221_X1 U91 ( .B1(n624), .B2(\A_ns[23] ), .C1(n621), .C2(\A_s[23] ), .A(
        n678), .ZN(n121) );
  INV_X1 U92 ( .A(n122), .ZN(n678) );
  AOI22_X1 U93 ( .A1(\A_ns[22] ), .A2(n627), .B1(\A_s[22] ), .B2(n617), .ZN(
        n122) );
  INV_X1 U94 ( .A(n117), .ZN(O[26]) );
  AOI221_X1 U95 ( .B1(n624), .B2(\A_ns[25] ), .C1(n621), .C2(\A_s[25] ), .A(
        n674), .ZN(n117) );
  INV_X1 U96 ( .A(n118), .ZN(n674) );
  AOI22_X1 U97 ( .A1(\A_ns[24] ), .A2(n628), .B1(\A_s[24] ), .B2(n618), .ZN(
        n118) );
  INV_X1 U98 ( .A(n124), .ZN(n680) );
  AOI22_X1 U99 ( .A1(\A_ns[21] ), .A2(n627), .B1(\A_s[21] ), .B2(n617), .ZN(
        n124) );
  INV_X1 U100 ( .A(n128), .ZN(n684) );
  AOI22_X1 U101 ( .A1(\A_ns[19] ), .A2(n627), .B1(\A_s[19] ), .B2(n617), .ZN(
        n128) );
  INV_X1 U102 ( .A(n126), .ZN(n682) );
  AOI22_X1 U103 ( .A1(\A_ns[20] ), .A2(n627), .B1(\A_s[20] ), .B2(n617), .ZN(
        n126) );
  INV_X1 U104 ( .A(n129), .ZN(O[20]) );
  AOI221_X1 U105 ( .B1(n624), .B2(\A_ns[19] ), .C1(n621), .C2(\A_s[19] ), .A(
        n686), .ZN(n129) );
  INV_X1 U106 ( .A(n130), .ZN(n686) );
  AOI22_X1 U107 ( .A1(\A_ns[18] ), .A2(n627), .B1(\A_s[18] ), .B2(n617), .ZN(
        n130) );
  INV_X1 U108 ( .A(n139), .ZN(O[15]) );
  AOI221_X1 U109 ( .B1(n624), .B2(\A_ns[14] ), .C1(n622), .C2(\A_s[14] ), .A(
        n696), .ZN(n139) );
  INV_X1 U110 ( .A(n140), .ZN(n696) );
  AOI22_X1 U111 ( .A1(\A_ns[13] ), .A2(n627), .B1(\A_s[13] ), .B2(n617), .ZN(
        n140) );
  INV_X1 U112 ( .A(n133), .ZN(O[18]) );
  AOI221_X1 U113 ( .B1(n624), .B2(\A_ns[17] ), .C1(n621), .C2(\A_s[17] ), .A(
        n690), .ZN(n133) );
  INV_X1 U114 ( .A(n134), .ZN(n690) );
  AOI22_X1 U115 ( .A1(\A_ns[16] ), .A2(n627), .B1(\A_s[16] ), .B2(n617), .ZN(
        n134) );
  OAI221_X1 U116 ( .B1(n629), .B2(n88), .C1(n630), .C2(n89), .A(n90), .ZN(
        O[40]) );
  AOI22_X1 U117 ( .A1(\A_ns[38] ), .A2(n628), .B1(\A_s[38] ), .B2(n619), .ZN(
        n90) );
  AOI22_X1 U118 ( .A1(\A_ns[27] ), .A2(n628), .B1(\A_s[27] ), .B2(n618), .ZN(
        n112) );
  AOI22_X1 U119 ( .A1(\A_ns[33] ), .A2(n628), .B1(\A_s[33] ), .B2(n618), .ZN(
        n100) );
  AOI22_X1 U120 ( .A1(\A_ns[35] ), .A2(n628), .B1(\A_s[35] ), .B2(n618), .ZN(
        n96) );
  AOI22_X1 U121 ( .A1(\A_ns[36] ), .A2(n628), .B1(\A_s[36] ), .B2(n619), .ZN(
        n94) );
  AOI22_X1 U122 ( .A1(\A_ns[32] ), .A2(n628), .B1(\A_s[32] ), .B2(n618), .ZN(
        n102) );
  AOI22_X1 U123 ( .A1(\A_ns[34] ), .A2(n628), .B1(\A_s[34] ), .B2(n618), .ZN(
        n98) );
  AOI22_X1 U124 ( .A1(\A_ns[26] ), .A2(n628), .B1(\A_s[26] ), .B2(n618), .ZN(
        n114) );
  INV_X1 U125 ( .A(n91), .ZN(O[39]) );
  AOI221_X1 U126 ( .B1(n623), .B2(\A_ns[38] ), .C1(n620), .C2(\A_s[38] ), .A(
        n648), .ZN(n91) );
  INV_X1 U127 ( .A(n92), .ZN(n648) );
  AOI22_X1 U128 ( .A1(\A_ns[37] ), .A2(n628), .B1(\A_s[37] ), .B2(n619), .ZN(
        n92) );
  INV_X1 U129 ( .A(n108), .ZN(n664) );
  AOI22_X1 U130 ( .A1(\A_ns[29] ), .A2(n628), .B1(\A_s[29] ), .B2(n618), .ZN(
        n108) );
  INV_X1 U131 ( .A(n104), .ZN(n660) );
  AOI22_X1 U132 ( .A1(\A_ns[31] ), .A2(n628), .B1(\A_s[31] ), .B2(n618), .ZN(
        n104) );
  INV_X1 U133 ( .A(n116), .ZN(n672) );
  AOI22_X1 U134 ( .A1(\A_ns[25] ), .A2(n628), .B1(\A_s[25] ), .B2(n618), .ZN(
        n116) );
  INV_X1 U135 ( .A(n105), .ZN(O[32]) );
  AOI221_X1 U136 ( .B1(n623), .B2(\A_ns[31] ), .C1(n620), .C2(\A_s[31] ), .A(
        n662), .ZN(n105) );
  INV_X1 U137 ( .A(n106), .ZN(n662) );
  AOI22_X1 U138 ( .A1(\A_ns[30] ), .A2(n628), .B1(\A_s[30] ), .B2(n618), .ZN(
        n106) );
  INV_X1 U139 ( .A(n110), .ZN(n666) );
  AOI22_X1 U140 ( .A1(\A_ns[28] ), .A2(n628), .B1(\A_s[28] ), .B2(n618), .ZN(
        n110) );
  OAI221_X1 U141 ( .B1(n613), .B2(n629), .C1(n85), .C2(n630), .A(n86), .ZN(
        O[41]) );
  INV_X1 U142 ( .A(n613), .ZN(n626) );
  NAND2_X1 U143 ( .A1(n168), .A2(n711), .ZN(n89) );
  NAND2_X1 U144 ( .A1(n168), .A2(n89), .ZN(n88) );
  INV_X1 U145 ( .A(n85), .ZN(n708) );
  INV_X1 U146 ( .A(n613), .ZN(n627) );
  INV_X1 U147 ( .A(n613), .ZN(n628) );
  OR3_X1 U148 ( .A1(B[7]), .A2(B[8]), .A3(n711), .ZN(n613) );
  INV_X1 U149 ( .A(n153), .ZN(O[8]) );
  AOI221_X1 U150 ( .B1(n625), .B2(\A_ns[7] ), .C1(n622), .C2(\A_s[7] ), .A(
        n645), .ZN(n153) );
  INV_X1 U151 ( .A(n154), .ZN(n645) );
  AOI22_X1 U152 ( .A1(\A_ns[6] ), .A2(n626), .B1(\A_s[6] ), .B2(n616), .ZN(
        n154) );
  INV_X1 U153 ( .A(B[9]), .ZN(n711) );
  INV_X1 U154 ( .A(n151), .ZN(O[9]) );
  AOI221_X1 U155 ( .B1(n625), .B2(\A_ns[8] ), .C1(n622), .C2(\A_s[8] ), .A(
        n707), .ZN(n151) );
  INV_X1 U156 ( .A(n152), .ZN(n707) );
  AOI22_X1 U157 ( .A1(\A_ns[7] ), .A2(n626), .B1(\A_s[7] ), .B2(n616), .ZN(
        n152) );
  INV_X1 U158 ( .A(n163), .ZN(O[3]) );
  AOI221_X1 U159 ( .B1(n625), .B2(\A_ns[2] ), .C1(n620), .C2(\A_s[2] ), .A(
        n635), .ZN(n163) );
  INV_X1 U160 ( .A(n164), .ZN(n635) );
  INV_X1 U161 ( .A(n165), .ZN(O[2]) );
  AOI221_X1 U162 ( .B1(n625), .B2(\A_ns[1] ), .C1(n620), .C2(\A_s[1] ), .A(
        n633), .ZN(n165) );
  INV_X1 U163 ( .A(n166), .ZN(n633) );
  AOI22_X1 U164 ( .A1(\A_ns[0] ), .A2(n626), .B1(\A_s[0] ), .B2(n616), .ZN(
        n166) );
  INV_X1 U165 ( .A(n161), .ZN(O[4]) );
  AOI221_X1 U166 ( .B1(n625), .B2(\A_ns[3] ), .C1(n622), .C2(\A_s[3] ), .A(
        n637), .ZN(n161) );
  INV_X1 U167 ( .A(n162), .ZN(n637) );
  AOI22_X1 U168 ( .A1(\A_ns[2] ), .A2(n626), .B1(\A_s[2] ), .B2(n616), .ZN(
        n162) );
  INV_X1 U169 ( .A(n157), .ZN(O[6]) );
  AOI221_X1 U172 ( .B1(n625), .B2(\A_ns[5] ), .C1(n622), .C2(\A_s[5] ), .A(
        n641), .ZN(n157) );
  INV_X1 U173 ( .A(n158), .ZN(n641) );
  AOI22_X1 U174 ( .A1(\A_ns[4] ), .A2(n626), .B1(\A_s[4] ), .B2(n616), .ZN(
        n158) );
  INV_X1 U175 ( .A(n159), .ZN(O[5]) );
  AOI221_X1 U176 ( .B1(n625), .B2(\A_ns[4] ), .C1(n622), .C2(\A_s[4] ), .A(
        n639), .ZN(n159) );
  INV_X1 U177 ( .A(n160), .ZN(n639) );
  AOI22_X1 U178 ( .A1(\A_ns[3] ), .A2(n626), .B1(\A_s[3] ), .B2(n616), .ZN(
        n160) );
  INV_X1 U179 ( .A(n155), .ZN(O[7]) );
  AOI221_X1 U180 ( .B1(n625), .B2(\A_ns[6] ), .C1(n622), .C2(\A_s[6] ), .A(
        n643), .ZN(n155) );
  INV_X1 U181 ( .A(n156), .ZN(n643) );
  AOI22_X1 U182 ( .A1(\A_ns[5] ), .A2(n626), .B1(\A_s[5] ), .B2(n616), .ZN(
        n156) );
  INV_X1 U183 ( .A(n167), .ZN(O[1]) );
  AOI22_X1 U184 ( .A1(n620), .A2(\A_s[0] ), .B1(n623), .B2(\A_ns[0] ), .ZN(
        n167) );
  AOI22_X1 U185 ( .A1(\A_ns[1] ), .A2(n626), .B1(\A_s[1] ), .B2(n616), .ZN(
        n164) );
endmodule


module BOOTHENC_NBIT44_i10 ( A_s, A_ns, B, O, A_so, A_nso );
  input [43:0] A_s;
  input [43:0] A_ns;
  input [43:0] B;
  output [43:0] O;
  output [43:0] A_so;
  output [43:0] A_nso;
  wire   \A_s[41] , \A_s[40] , \A_s[39] , \A_s[38] , \A_s[37] , \A_s[36] ,
         \A_s[35] , \A_s[34] , \A_s[33] , \A_s[32] , \A_s[31] , \A_s[30] ,
         \A_s[29] , \A_s[28] , \A_s[27] , \A_s[26] , \A_s[25] , \A_s[24] ,
         \A_s[23] , \A_s[22] , \A_s[21] , \A_s[20] , \A_s[19] , \A_s[18] ,
         \A_s[17] , \A_s[16] , \A_s[15] , \A_s[14] , \A_s[13] , \A_s[12] ,
         \A_s[11] , \A_s[10] , \A_s[9] , \A_s[8] , \A_s[7] , \A_s[6] ,
         \A_s[5] , \A_s[4] , \A_s[3] , \A_s[2] , \A_s[1] , \A_s[0] ,
         \A_ns[40] , \A_ns[39] , \A_ns[38] , \A_ns[37] , \A_ns[36] ,
         \A_ns[35] , \A_ns[34] , \A_ns[33] , \A_ns[32] , \A_ns[31] ,
         \A_ns[30] , \A_ns[29] , \A_ns[28] , \A_ns[27] , \A_ns[26] ,
         \A_ns[25] , \A_ns[24] , \A_ns[23] , \A_ns[22] , \A_ns[21] ,
         \A_ns[20] , \A_ns[19] , \A_ns[18] , \A_ns[17] , \A_ns[16] ,
         \A_ns[15] , \A_ns[14] , \A_ns[13] , \A_ns[12] , \A_ns[11] ,
         \A_ns[10] , \A_ns[9] , \A_ns[8] , \A_ns[7] , \A_ns[6] , \A_ns[5] ,
         \A_ns[4] , \A_ns[3] , \A_ns[2] , \A_ns[1] , \A_ns[0] , n89, n90, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n663, n664, n667, n669, n671, n673, n675,
         n677, n679, n681, n683, n686, n688, n690, n692, n694, n696, n698,
         n700, n702, n704, n706, n708, n710, n712, n714, n716, n718, n720,
         n722, n724, n726, n728, n730, n732, n734, n736, n738, n740, n742,
         n744, n745, n746, n747, n748, n749;
  assign A_nso[0] = 1'b0;
  assign A_nso[1] = 1'b0;
  assign A_so[0] = 1'b0;
  assign A_so[1] = 1'b0;
  assign O[0] = 1'b0;
  assign A_so[43] = \A_s[41] ;
  assign \A_s[41]  = A_s[41];
  assign A_so[42] = \A_s[40] ;
  assign \A_s[40]  = A_s[40];
  assign A_so[41] = \A_s[39] ;
  assign \A_s[39]  = A_s[39];
  assign A_so[40] = \A_s[38] ;
  assign \A_s[38]  = A_s[38];
  assign A_so[39] = \A_s[37] ;
  assign \A_s[37]  = A_s[37];
  assign A_so[38] = \A_s[36] ;
  assign \A_s[36]  = A_s[36];
  assign A_so[37] = \A_s[35] ;
  assign \A_s[35]  = A_s[35];
  assign A_so[36] = \A_s[34] ;
  assign \A_s[34]  = A_s[34];
  assign A_so[35] = \A_s[33] ;
  assign \A_s[33]  = A_s[33];
  assign A_so[34] = \A_s[32] ;
  assign \A_s[32]  = A_s[32];
  assign A_so[33] = \A_s[31] ;
  assign \A_s[31]  = A_s[31];
  assign A_so[32] = \A_s[30] ;
  assign \A_s[30]  = A_s[30];
  assign A_so[31] = \A_s[29] ;
  assign \A_s[29]  = A_s[29];
  assign A_so[30] = \A_s[28] ;
  assign \A_s[28]  = A_s[28];
  assign A_so[29] = \A_s[27] ;
  assign \A_s[27]  = A_s[27];
  assign A_so[28] = \A_s[26] ;
  assign \A_s[26]  = A_s[26];
  assign A_so[27] = \A_s[25] ;
  assign \A_s[25]  = A_s[25];
  assign A_so[26] = \A_s[24] ;
  assign \A_s[24]  = A_s[24];
  assign A_so[25] = \A_s[23] ;
  assign \A_s[23]  = A_s[23];
  assign A_so[24] = \A_s[22] ;
  assign \A_s[22]  = A_s[22];
  assign A_so[23] = \A_s[21] ;
  assign \A_s[21]  = A_s[21];
  assign A_so[22] = \A_s[20] ;
  assign \A_s[20]  = A_s[20];
  assign A_so[21] = \A_s[19] ;
  assign \A_s[19]  = A_s[19];
  assign A_so[20] = \A_s[18] ;
  assign \A_s[18]  = A_s[18];
  assign A_so[19] = \A_s[17] ;
  assign \A_s[17]  = A_s[17];
  assign A_so[18] = \A_s[16] ;
  assign \A_s[16]  = A_s[16];
  assign A_so[17] = \A_s[15] ;
  assign \A_s[15]  = A_s[15];
  assign A_so[16] = \A_s[14] ;
  assign \A_s[14]  = A_s[14];
  assign A_so[15] = \A_s[13] ;
  assign \A_s[13]  = A_s[13];
  assign A_so[14] = \A_s[12] ;
  assign \A_s[12]  = A_s[12];
  assign A_so[13] = \A_s[11] ;
  assign \A_s[11]  = A_s[11];
  assign A_so[12] = \A_s[10] ;
  assign \A_s[10]  = A_s[10];
  assign A_so[11] = \A_s[9] ;
  assign \A_s[9]  = A_s[9];
  assign A_so[10] = \A_s[8] ;
  assign \A_s[8]  = A_s[8];
  assign A_so[9] = \A_s[7] ;
  assign \A_s[7]  = A_s[7];
  assign A_so[8] = \A_s[6] ;
  assign \A_s[6]  = A_s[6];
  assign A_so[7] = \A_s[5] ;
  assign \A_s[5]  = A_s[5];
  assign A_so[6] = \A_s[4] ;
  assign \A_s[4]  = A_s[4];
  assign A_so[5] = \A_s[3] ;
  assign \A_s[3]  = A_s[3];
  assign A_so[4] = \A_s[2] ;
  assign \A_s[2]  = A_s[2];
  assign A_so[3] = \A_s[1] ;
  assign \A_s[1]  = A_s[1];
  assign A_so[2] = \A_s[0] ;
  assign \A_s[0]  = A_s[0];
  assign A_nso[42] = \A_ns[40] ;
  assign \A_ns[40]  = A_ns[40];
  assign A_nso[41] = \A_ns[39] ;
  assign \A_ns[39]  = A_ns[39];
  assign A_nso[40] = \A_ns[38] ;
  assign \A_ns[38]  = A_ns[38];
  assign A_nso[39] = \A_ns[37] ;
  assign \A_ns[37]  = A_ns[37];
  assign A_nso[38] = \A_ns[36] ;
  assign \A_ns[36]  = A_ns[36];
  assign A_nso[37] = \A_ns[35] ;
  assign \A_ns[35]  = A_ns[35];
  assign A_nso[36] = \A_ns[34] ;
  assign \A_ns[34]  = A_ns[34];
  assign A_nso[35] = \A_ns[33] ;
  assign \A_ns[33]  = A_ns[33];
  assign A_nso[34] = \A_ns[32] ;
  assign \A_ns[32]  = A_ns[32];
  assign A_nso[33] = \A_ns[31] ;
  assign \A_ns[31]  = A_ns[31];
  assign A_nso[32] = \A_ns[30] ;
  assign \A_ns[30]  = A_ns[30];
  assign A_nso[31] = \A_ns[29] ;
  assign \A_ns[29]  = A_ns[29];
  assign A_nso[30] = \A_ns[28] ;
  assign \A_ns[28]  = A_ns[28];
  assign A_nso[29] = \A_ns[27] ;
  assign \A_ns[27]  = A_ns[27];
  assign A_nso[28] = \A_ns[26] ;
  assign \A_ns[26]  = A_ns[26];
  assign A_nso[27] = \A_ns[25] ;
  assign \A_ns[25]  = A_ns[25];
  assign A_nso[26] = \A_ns[24] ;
  assign \A_ns[24]  = A_ns[24];
  assign A_nso[25] = \A_ns[23] ;
  assign \A_ns[23]  = A_ns[23];
  assign A_nso[24] = \A_ns[22] ;
  assign \A_ns[22]  = A_ns[22];
  assign A_nso[23] = \A_ns[21] ;
  assign \A_ns[21]  = A_ns[21];
  assign A_nso[22] = \A_ns[20] ;
  assign \A_ns[20]  = A_ns[20];
  assign A_nso[21] = \A_ns[19] ;
  assign \A_ns[19]  = A_ns[19];
  assign A_nso[20] = \A_ns[18] ;
  assign \A_ns[18]  = A_ns[18];
  assign A_nso[19] = \A_ns[17] ;
  assign \A_ns[17]  = A_ns[17];
  assign A_nso[18] = \A_ns[16] ;
  assign \A_ns[16]  = A_ns[16];
  assign A_nso[17] = \A_ns[15] ;
  assign \A_ns[15]  = A_ns[15];
  assign A_nso[16] = \A_ns[14] ;
  assign \A_ns[14]  = A_ns[14];
  assign A_nso[15] = \A_ns[13] ;
  assign \A_ns[13]  = A_ns[13];
  assign A_nso[14] = \A_ns[12] ;
  assign \A_ns[12]  = A_ns[12];
  assign A_nso[13] = \A_ns[11] ;
  assign \A_ns[11]  = A_ns[11];
  assign A_nso[12] = \A_ns[10] ;
  assign \A_ns[10]  = A_ns[10];
  assign A_nso[11] = \A_ns[9] ;
  assign \A_ns[9]  = A_ns[9];
  assign A_nso[10] = \A_ns[8] ;
  assign \A_ns[8]  = A_ns[8];
  assign A_nso[9] = \A_ns[7] ;
  assign \A_ns[7]  = A_ns[7];
  assign A_nso[8] = \A_ns[6] ;
  assign \A_ns[6]  = A_ns[6];
  assign A_nso[7] = \A_ns[5] ;
  assign \A_ns[5]  = A_ns[5];
  assign A_nso[6] = \A_ns[4] ;
  assign \A_ns[4]  = A_ns[4];
  assign A_nso[5] = \A_ns[3] ;
  assign \A_ns[3]  = A_ns[3];
  assign A_nso[4] = \A_ns[2] ;
  assign \A_ns[2]  = A_ns[2];
  assign A_nso[3] = \A_ns[1] ;
  assign \A_ns[1]  = A_ns[1];
  assign A_nso[2] = \A_ns[0] ;
  assign \A_ns[0]  = A_ns[0];

  OAI221_X2 U2 ( .B1(n641), .B2(n663), .C1(n89), .C2(n664), .A(n90), .ZN(O[43]) );
  NAND3_X1 U178 ( .A1(B[10]), .A2(n749), .A3(B[9]), .ZN(n89) );
  XOR2_X1 U179 ( .A(B[10]), .B(B[9]), .Z(n176) );
  AOI22_X1 U3 ( .A1(A_ns[42]), .A2(n656), .B1(A_s[42]), .B2(n650), .ZN(n90) );
  OAI221_X1 U4 ( .B1(n663), .B2(n92), .C1(n664), .C2(n93), .A(n94), .ZN(O[42])
         );
  CLKBUF_X1 U5 ( .A(n654), .Z(n656) );
  CLKBUF_X1 U6 ( .A(n649), .Z(n653) );
  CLKBUF_X1 U7 ( .A(n655), .Z(n659) );
  CLKBUF_X1 U8 ( .A(n642), .Z(n645) );
  CLKBUF_X1 U9 ( .A(n748), .Z(n654) );
  CLKBUF_X1 U10 ( .A(n747), .Z(n648) );
  CLKBUF_X1 U11 ( .A(n746), .Z(n643) );
  INV_X1 U12 ( .A(A_ns[41]), .ZN(n663) );
  INV_X1 U13 ( .A(\A_s[41] ), .ZN(n664) );
  BUF_X1 U14 ( .A(n654), .Z(n657) );
  BUF_X1 U15 ( .A(n655), .Z(n658) );
  BUF_X1 U16 ( .A(n649), .Z(n652) );
  BUF_X1 U17 ( .A(n648), .Z(n650) );
  BUF_X1 U18 ( .A(n648), .Z(n651) );
  BUF_X1 U19 ( .A(n642), .Z(n644) );
  BUF_X1 U20 ( .A(n747), .Z(n649) );
  BUF_X1 U21 ( .A(n748), .Z(n655) );
  BUF_X1 U22 ( .A(n643), .Z(n646) );
  BUF_X1 U23 ( .A(n643), .Z(n647) );
  INV_X1 U24 ( .A(n153), .ZN(O[12]) );
  INV_X1 U25 ( .A(n151), .ZN(O[13]) );
  AOI221_X1 U26 ( .B1(n658), .B2(\A_ns[12] ), .C1(n652), .C2(\A_s[12] ), .A(
        n742), .ZN(n151) );
  AOI22_X1 U27 ( .A1(\A_ns[40] ), .A2(n661), .B1(\A_s[40] ), .B2(n647), .ZN(
        n94) );
  INV_X1 U28 ( .A(n133), .ZN(O[22]) );
  AOI221_X1 U29 ( .B1(n657), .B2(\A_ns[21] ), .C1(n651), .C2(\A_s[21] ), .A(
        n724), .ZN(n133) );
  INV_X1 U30 ( .A(n134), .ZN(n724) );
  AOI22_X1 U31 ( .A1(\A_ns[20] ), .A2(n661), .B1(\A_s[20] ), .B2(n645), .ZN(
        n134) );
  AOI221_X1 U32 ( .B1(n658), .B2(\A_ns[11] ), .C1(n652), .C2(\A_s[11] ), .A(
        n744), .ZN(n153) );
  INV_X1 U33 ( .A(n154), .ZN(n744) );
  AOI22_X1 U34 ( .A1(\A_ns[10] ), .A2(n660), .B1(\A_s[10] ), .B2(n644), .ZN(
        n154) );
  INV_X1 U35 ( .A(n135), .ZN(O[21]) );
  AOI221_X1 U36 ( .B1(n657), .B2(\A_ns[20] ), .C1(n651), .C2(\A_s[20] ), .A(
        n726), .ZN(n135) );
  INV_X1 U37 ( .A(n136), .ZN(n726) );
  AOI22_X1 U38 ( .A1(\A_ns[19] ), .A2(n661), .B1(\A_s[19] ), .B2(n645), .ZN(
        n136) );
  INV_X1 U39 ( .A(n149), .ZN(O[14]) );
  AOI221_X1 U40 ( .B1(n658), .B2(\A_ns[13] ), .C1(n652), .C2(\A_s[13] ), .A(
        n740), .ZN(n149) );
  INV_X1 U41 ( .A(n150), .ZN(n740) );
  AOI22_X1 U42 ( .A1(\A_ns[12] ), .A2(n661), .B1(\A_s[12] ), .B2(n645), .ZN(
        n150) );
  INV_X1 U43 ( .A(n139), .ZN(O[19]) );
  AOI221_X1 U44 ( .B1(n657), .B2(\A_ns[18] ), .C1(n651), .C2(\A_s[18] ), .A(
        n730), .ZN(n139) );
  INV_X1 U45 ( .A(n140), .ZN(n730) );
  AOI22_X1 U46 ( .A1(\A_ns[17] ), .A2(n661), .B1(\A_s[17] ), .B2(n645), .ZN(
        n140) );
  INV_X1 U47 ( .A(n131), .ZN(O[23]) );
  AOI221_X1 U48 ( .B1(n657), .B2(\A_ns[22] ), .C1(n651), .C2(\A_s[22] ), .A(
        n722), .ZN(n131) );
  INV_X1 U49 ( .A(n132), .ZN(n722) );
  AOI22_X1 U50 ( .A1(\A_ns[21] ), .A2(n661), .B1(\A_s[21] ), .B2(n645), .ZN(
        n132) );
  INV_X1 U51 ( .A(n143), .ZN(O[17]) );
  AOI221_X1 U52 ( .B1(n657), .B2(\A_ns[16] ), .C1(n652), .C2(\A_s[16] ), .A(
        n734), .ZN(n143) );
  INV_X1 U53 ( .A(n144), .ZN(n734) );
  AOI22_X1 U54 ( .A1(\A_ns[15] ), .A2(n661), .B1(\A_s[15] ), .B2(n645), .ZN(
        n144) );
  INV_X1 U55 ( .A(n152), .ZN(n742) );
  AOI22_X1 U56 ( .A1(\A_ns[11] ), .A2(n660), .B1(\A_s[11] ), .B2(n644), .ZN(
        n152) );
  INV_X1 U57 ( .A(n145), .ZN(O[16]) );
  AOI221_X1 U58 ( .B1(n658), .B2(\A_ns[15] ), .C1(n652), .C2(\A_s[15] ), .A(
        n736), .ZN(n145) );
  INV_X1 U59 ( .A(n146), .ZN(n736) );
  AOI22_X1 U60 ( .A1(\A_ns[14] ), .A2(n661), .B1(\A_s[14] ), .B2(n645), .ZN(
        n146) );
  INV_X1 U61 ( .A(n147), .ZN(O[15]) );
  AOI221_X1 U62 ( .B1(n658), .B2(\A_ns[14] ), .C1(n652), .C2(\A_s[14] ), .A(
        n738), .ZN(n147) );
  INV_X1 U63 ( .A(n148), .ZN(n738) );
  AOI22_X1 U64 ( .A1(\A_ns[13] ), .A2(n661), .B1(\A_s[13] ), .B2(n645), .ZN(
        n148) );
  BUF_X1 U65 ( .A(n746), .Z(n642) );
  INV_X1 U66 ( .A(n137), .ZN(O[20]) );
  AOI221_X1 U67 ( .B1(n657), .B2(\A_ns[19] ), .C1(n651), .C2(\A_s[19] ), .A(
        n728), .ZN(n137) );
  INV_X1 U68 ( .A(n138), .ZN(n728) );
  AOI22_X1 U69 ( .A1(\A_ns[18] ), .A2(n661), .B1(\A_s[18] ), .B2(n645), .ZN(
        n138) );
  INV_X1 U70 ( .A(n141), .ZN(O[18]) );
  AOI221_X1 U71 ( .B1(n657), .B2(\A_ns[17] ), .C1(n652), .C2(\A_s[17] ), .A(
        n732), .ZN(n141) );
  INV_X1 U72 ( .A(n142), .ZN(n732) );
  AOI22_X1 U73 ( .A1(\A_ns[16] ), .A2(n661), .B1(\A_s[16] ), .B2(n645), .ZN(
        n142) );
  INV_X1 U74 ( .A(n93), .ZN(n747) );
  INV_X1 U75 ( .A(n92), .ZN(n748) );
  INV_X1 U76 ( .A(n115), .ZN(O[31]) );
  AOI221_X1 U77 ( .B1(n656), .B2(\A_ns[30] ), .C1(n650), .C2(\A_s[30] ), .A(
        n706), .ZN(n115) );
  INV_X1 U78 ( .A(n116), .ZN(n706) );
  AOI22_X1 U79 ( .A1(\A_ns[29] ), .A2(n660), .B1(\A_s[29] ), .B2(n646), .ZN(
        n116) );
  INV_X1 U80 ( .A(n101), .ZN(O[38]) );
  AOI221_X1 U81 ( .B1(n656), .B2(\A_ns[37] ), .C1(n650), .C2(\A_s[37] ), .A(
        n692), .ZN(n101) );
  INV_X1 U82 ( .A(n102), .ZN(n692) );
  AOI22_X1 U83 ( .A1(\A_ns[36] ), .A2(n660), .B1(\A_s[36] ), .B2(n647), .ZN(
        n102) );
  INV_X1 U84 ( .A(n105), .ZN(O[36]) );
  AOI221_X1 U85 ( .B1(n656), .B2(\A_ns[35] ), .C1(n650), .C2(\A_s[35] ), .A(
        n696), .ZN(n105) );
  INV_X1 U86 ( .A(n106), .ZN(n696) );
  AOI22_X1 U87 ( .A1(\A_ns[34] ), .A2(n660), .B1(\A_s[34] ), .B2(n646), .ZN(
        n106) );
  INV_X1 U88 ( .A(n113), .ZN(O[32]) );
  AOI221_X1 U89 ( .B1(n656), .B2(\A_ns[31] ), .C1(n651), .C2(\A_s[31] ), .A(
        n704), .ZN(n113) );
  INV_X1 U90 ( .A(n114), .ZN(n704) );
  AOI22_X1 U91 ( .A1(\A_ns[30] ), .A2(n660), .B1(\A_s[30] ), .B2(n646), .ZN(
        n114) );
  INV_X1 U92 ( .A(n109), .ZN(O[34]) );
  AOI221_X1 U93 ( .B1(n656), .B2(\A_ns[33] ), .C1(n650), .C2(\A_s[33] ), .A(
        n700), .ZN(n109) );
  INV_X1 U94 ( .A(n110), .ZN(n700) );
  AOI22_X1 U95 ( .A1(\A_ns[32] ), .A2(n660), .B1(\A_s[32] ), .B2(n646), .ZN(
        n110) );
  INV_X1 U96 ( .A(n111), .ZN(O[33]) );
  AOI221_X1 U97 ( .B1(n656), .B2(\A_ns[32] ), .C1(n650), .C2(\A_s[32] ), .A(
        n702), .ZN(n111) );
  INV_X1 U98 ( .A(n112), .ZN(n702) );
  AOI22_X1 U99 ( .A1(\A_ns[31] ), .A2(n660), .B1(\A_s[31] ), .B2(n646), .ZN(
        n112) );
  INV_X1 U100 ( .A(n127), .ZN(O[25]) );
  AOI221_X1 U101 ( .B1(n657), .B2(\A_ns[24] ), .C1(n651), .C2(\A_s[24] ), .A(
        n718), .ZN(n127) );
  INV_X1 U102 ( .A(n128), .ZN(n718) );
  AOI22_X1 U103 ( .A1(\A_ns[23] ), .A2(n661), .B1(\A_s[23] ), .B2(n645), .ZN(
        n128) );
  INV_X1 U104 ( .A(n107), .ZN(O[35]) );
  AOI221_X1 U105 ( .B1(n656), .B2(\A_ns[34] ), .C1(n650), .C2(\A_s[34] ), .A(
        n698), .ZN(n107) );
  INV_X1 U106 ( .A(n108), .ZN(n698) );
  AOI22_X1 U107 ( .A1(\A_ns[33] ), .A2(n660), .B1(\A_s[33] ), .B2(n646), .ZN(
        n108) );
  INV_X1 U108 ( .A(n119), .ZN(O[29]) );
  AOI221_X1 U109 ( .B1(n657), .B2(\A_ns[28] ), .C1(n651), .C2(\A_s[28] ), .A(
        n710), .ZN(n119) );
  INV_X1 U110 ( .A(n120), .ZN(n710) );
  AOI22_X1 U111 ( .A1(\A_ns[27] ), .A2(n660), .B1(\A_s[27] ), .B2(n646), .ZN(
        n120) );
  INV_X1 U112 ( .A(n99), .ZN(O[39]) );
  AOI221_X1 U113 ( .B1(n656), .B2(\A_ns[38] ), .C1(n650), .C2(\A_s[38] ), .A(
        n690), .ZN(n99) );
  INV_X1 U114 ( .A(n100), .ZN(n690) );
  AOI22_X1 U115 ( .A1(\A_ns[37] ), .A2(n661), .B1(\A_s[37] ), .B2(n647), .ZN(
        n100) );
  INV_X1 U116 ( .A(n97), .ZN(O[40]) );
  AOI221_X1 U117 ( .B1(n656), .B2(\A_ns[39] ), .C1(n650), .C2(\A_s[39] ), .A(
        n688), .ZN(n97) );
  INV_X1 U118 ( .A(n98), .ZN(n688) );
  AOI22_X1 U119 ( .A1(\A_ns[38] ), .A2(n660), .B1(\A_s[38] ), .B2(n647), .ZN(
        n98) );
  INV_X1 U120 ( .A(n125), .ZN(O[26]) );
  AOI221_X1 U121 ( .B1(n657), .B2(\A_ns[25] ), .C1(n651), .C2(\A_s[25] ), .A(
        n716), .ZN(n125) );
  INV_X1 U122 ( .A(n126), .ZN(n716) );
  AOI22_X1 U123 ( .A1(\A_ns[24] ), .A2(n660), .B1(\A_s[24] ), .B2(n646), .ZN(
        n126) );
  INV_X1 U124 ( .A(n129), .ZN(O[24]) );
  AOI221_X1 U125 ( .B1(n657), .B2(\A_ns[23] ), .C1(n651), .C2(\A_s[23] ), .A(
        n720), .ZN(n129) );
  INV_X1 U126 ( .A(n130), .ZN(n720) );
  AOI22_X1 U127 ( .A1(\A_ns[22] ), .A2(n661), .B1(\A_s[22] ), .B2(n645), .ZN(
        n130) );
  INV_X1 U128 ( .A(n117), .ZN(O[30]) );
  AOI221_X1 U129 ( .B1(n656), .B2(\A_ns[29] ), .C1(n651), .C2(\A_s[29] ), .A(
        n708), .ZN(n117) );
  INV_X1 U130 ( .A(n118), .ZN(n708) );
  AOI22_X1 U131 ( .A1(\A_ns[28] ), .A2(n660), .B1(\A_s[28] ), .B2(n646), .ZN(
        n118) );
  INV_X1 U132 ( .A(n121), .ZN(O[28]) );
  AOI221_X1 U133 ( .B1(n657), .B2(\A_ns[27] ), .C1(n651), .C2(\A_s[27] ), .A(
        n712), .ZN(n121) );
  INV_X1 U134 ( .A(n122), .ZN(n712) );
  AOI22_X1 U135 ( .A1(\A_ns[26] ), .A2(n660), .B1(\A_s[26] ), .B2(n646), .ZN(
        n122) );
  INV_X1 U136 ( .A(n103), .ZN(O[37]) );
  AOI221_X1 U137 ( .B1(n656), .B2(\A_ns[36] ), .C1(n650), .C2(\A_s[36] ), .A(
        n694), .ZN(n103) );
  INV_X1 U138 ( .A(n104), .ZN(n694) );
  AOI22_X1 U139 ( .A1(\A_ns[35] ), .A2(n661), .B1(\A_s[35] ), .B2(n646), .ZN(
        n104) );
  INV_X1 U140 ( .A(n123), .ZN(O[27]) );
  AOI221_X1 U141 ( .B1(n657), .B2(\A_ns[26] ), .C1(n651), .C2(\A_s[26] ), .A(
        n714), .ZN(n123) );
  INV_X1 U142 ( .A(n124), .ZN(n714) );
  AOI22_X1 U143 ( .A1(\A_ns[25] ), .A2(n660), .B1(\A_s[25] ), .B2(n646), .ZN(
        n124) );
  INV_X1 U144 ( .A(n95), .ZN(O[41]) );
  AOI221_X1 U145 ( .B1(n656), .B2(\A_ns[40] ), .C1(n650), .C2(\A_s[40] ), .A(
        n686), .ZN(n95) );
  INV_X1 U146 ( .A(n96), .ZN(n686) );
  AOI22_X1 U147 ( .A1(\A_ns[39] ), .A2(n661), .B1(\A_s[39] ), .B2(n647), .ZN(
        n96) );
  INV_X1 U148 ( .A(n641), .ZN(n661) );
  INV_X1 U149 ( .A(n641), .ZN(n660) );
  NAND2_X1 U150 ( .A1(n176), .A2(n749), .ZN(n93) );
  NAND2_X1 U151 ( .A1(n176), .A2(n93), .ZN(n92) );
  INV_X1 U152 ( .A(n89), .ZN(n746) );
  OR3_X1 U153 ( .A1(B[10]), .A2(B[9]), .A3(n749), .ZN(n641) );
  INV_X1 U154 ( .A(n155), .ZN(O[11]) );
  AOI221_X1 U155 ( .B1(n658), .B2(\A_ns[10] ), .C1(n652), .C2(\A_s[10] ), .A(
        n745), .ZN(n155) );
  INV_X1 U156 ( .A(n156), .ZN(n745) );
  AOI22_X1 U157 ( .A1(\A_ns[9] ), .A2(n660), .B1(\A_s[9] ), .B2(n644), .ZN(
        n156) );
  INV_X1 U158 ( .A(n157), .ZN(O[10]) );
  AOI221_X1 U159 ( .B1(n658), .B2(\A_ns[9] ), .C1(n652), .C2(\A_s[9] ), .A(
        n683), .ZN(n157) );
  INV_X1 U160 ( .A(n158), .ZN(n683) );
  AOI22_X1 U161 ( .A1(\A_ns[8] ), .A2(n660), .B1(\A_s[8] ), .B2(n644), .ZN(
        n158) );
  INV_X1 U162 ( .A(B[11]), .ZN(n749) );
  INV_X1 U163 ( .A(n159), .ZN(O[9]) );
  AOI221_X1 U164 ( .B1(n658), .B2(\A_ns[8] ), .C1(n652), .C2(\A_s[8] ), .A(
        n681), .ZN(n159) );
  INV_X1 U165 ( .A(n161), .ZN(O[8]) );
  AOI221_X1 U166 ( .B1(n658), .B2(\A_ns[7] ), .C1(n652), .C2(\A_s[7] ), .A(
        n679), .ZN(n161) );
  INV_X1 U167 ( .A(n163), .ZN(O[7]) );
  AOI221_X1 U168 ( .B1(n658), .B2(\A_ns[6] ), .C1(n652), .C2(\A_s[6] ), .A(
        n677), .ZN(n163) );
  INV_X1 U169 ( .A(n175), .ZN(O[1]) );
  INV_X1 U170 ( .A(n173), .ZN(O[2]) );
  AOI221_X1 U171 ( .B1(n659), .B2(\A_ns[1] ), .C1(n650), .C2(\A_s[1] ), .A(
        n667), .ZN(n173) );
  INV_X1 U172 ( .A(n169), .ZN(O[4]) );
  AOI221_X1 U173 ( .B1(n658), .B2(\A_ns[3] ), .C1(n653), .C2(\A_s[3] ), .A(
        n671), .ZN(n169) );
  INV_X1 U174 ( .A(n167), .ZN(O[5]) );
  AOI221_X1 U175 ( .B1(n658), .B2(\A_ns[4] ), .C1(n653), .C2(\A_s[4] ), .A(
        n673), .ZN(n167) );
  INV_X1 U176 ( .A(n165), .ZN(O[6]) );
  AOI221_X1 U177 ( .B1(n658), .B2(\A_ns[5] ), .C1(n652), .C2(\A_s[5] ), .A(
        n675), .ZN(n165) );
  INV_X1 U180 ( .A(n171), .ZN(O[3]) );
  AOI221_X1 U181 ( .B1(n659), .B2(\A_ns[2] ), .C1(n653), .C2(\A_s[2] ), .A(
        n669), .ZN(n171) );
  INV_X1 U182 ( .A(n174), .ZN(n667) );
  AOI22_X1 U183 ( .A1(\A_ns[0] ), .A2(n660), .B1(\A_s[0] ), .B2(n644), .ZN(
        n174) );
  INV_X1 U184 ( .A(n172), .ZN(n669) );
  AOI22_X1 U185 ( .A1(\A_ns[1] ), .A2(n660), .B1(\A_s[1] ), .B2(n644), .ZN(
        n172) );
  INV_X1 U186 ( .A(n170), .ZN(n671) );
  AOI22_X1 U187 ( .A1(\A_ns[2] ), .A2(n660), .B1(\A_s[2] ), .B2(n644), .ZN(
        n170) );
  INV_X1 U188 ( .A(n168), .ZN(n673) );
  AOI22_X1 U189 ( .A1(\A_ns[3] ), .A2(n660), .B1(\A_s[3] ), .B2(n644), .ZN(
        n168) );
  INV_X1 U190 ( .A(n166), .ZN(n675) );
  AOI22_X1 U191 ( .A1(\A_ns[4] ), .A2(n660), .B1(\A_s[4] ), .B2(n644), .ZN(
        n166) );
  INV_X1 U192 ( .A(n164), .ZN(n677) );
  AOI22_X1 U193 ( .A1(\A_ns[5] ), .A2(n660), .B1(\A_s[5] ), .B2(n644), .ZN(
        n164) );
  INV_X1 U194 ( .A(n162), .ZN(n679) );
  AOI22_X1 U195 ( .A1(\A_ns[6] ), .A2(n660), .B1(\A_s[6] ), .B2(n644), .ZN(
        n162) );
  INV_X1 U196 ( .A(n160), .ZN(n681) );
  AOI22_X1 U197 ( .A1(\A_ns[7] ), .A2(n660), .B1(\A_s[7] ), .B2(n644), .ZN(
        n160) );
  AOI22_X1 U198 ( .A1(n650), .A2(\A_s[0] ), .B1(n659), .B2(\A_ns[0] ), .ZN(
        n175) );
  INV_X1 U199 ( .A(n663), .ZN(A_nso[43]) );
endmodule


module BOOTHENC_NBIT46_i12 ( A_s, A_ns, B, O, A_so, A_nso );
  input [45:0] A_s;
  input [45:0] A_ns;
  input [45:0] B;
  output [45:0] O;
  output [45:0] A_so;
  output [45:0] A_nso;
  wire   \A_s[43] , \A_s[42] , \A_s[41] , \A_s[40] , \A_s[39] , \A_s[38] ,
         \A_s[37] , \A_s[36] , \A_s[35] , \A_s[34] , \A_s[33] , \A_s[32] ,
         \A_s[31] , \A_s[30] , \A_s[29] , \A_s[28] , \A_s[27] , \A_s[26] ,
         \A_s[25] , \A_s[24] , \A_s[23] , \A_s[22] , \A_s[21] , \A_s[20] ,
         \A_s[19] , \A_s[18] , \A_s[17] , \A_s[16] , \A_s[15] , \A_s[14] ,
         \A_s[13] , \A_s[12] , \A_s[11] , \A_s[10] , \A_s[9] , \A_s[8] ,
         \A_s[7] , \A_s[6] , \A_s[5] , \A_s[4] , \A_s[3] , \A_s[2] , \A_s[1] ,
         \A_s[0] , \A_ns[43] , \A_ns[42] , \A_ns[41] , \A_ns[40] , \A_ns[39] ,
         \A_ns[38] , \A_ns[37] , \A_ns[36] , \A_ns[35] , \A_ns[34] ,
         \A_ns[33] , \A_ns[32] , \A_ns[31] , \A_ns[30] , \A_ns[29] ,
         \A_ns[28] , \A_ns[27] , \A_ns[26] , \A_ns[25] , \A_ns[24] ,
         \A_ns[23] , \A_ns[22] , \A_ns[21] , \A_ns[20] , \A_ns[19] ,
         \A_ns[18] , \A_ns[17] , \A_ns[16] , \A_ns[15] , \A_ns[14] ,
         \A_ns[13] , \A_ns[12] , \A_ns[11] , \A_ns[10] , \A_ns[9] , \A_ns[8] ,
         \A_ns[7] , \A_ns[6] , \A_ns[5] , \A_ns[4] , \A_ns[3] , \A_ns[2] ,
         \A_ns[1] , \A_ns[0] , n93, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n694, n696, n698, n700, n702,
         n704, n706, n708, n710, n712, n714, n716, n719, n721, n723, n725,
         n727, n729, n731, n733, n735, n737, n739, n741, n743, n745, n747,
         n749, n751, n753, n755, n757, n759, n761, n763, n765, n767, n769,
         n771, n773, n775, n776, n777, n778, n779, n780;
  assign A_nso[0] = 1'b0;
  assign A_nso[1] = 1'b0;
  assign A_so[0] = 1'b0;
  assign A_so[1] = 1'b0;
  assign O[0] = 1'b0;
  assign A_so[45] = \A_s[43] ;
  assign \A_s[43]  = A_s[43];
  assign A_so[44] = \A_s[42] ;
  assign \A_s[42]  = A_s[42];
  assign A_so[43] = \A_s[41] ;
  assign \A_s[41]  = A_s[41];
  assign A_so[42] = \A_s[40] ;
  assign \A_s[40]  = A_s[40];
  assign A_so[41] = \A_s[39] ;
  assign \A_s[39]  = A_s[39];
  assign A_so[40] = \A_s[38] ;
  assign \A_s[38]  = A_s[38];
  assign A_so[39] = \A_s[37] ;
  assign \A_s[37]  = A_s[37];
  assign A_so[38] = \A_s[36] ;
  assign \A_s[36]  = A_s[36];
  assign A_so[37] = \A_s[35] ;
  assign \A_s[35]  = A_s[35];
  assign A_so[36] = \A_s[34] ;
  assign \A_s[34]  = A_s[34];
  assign A_so[35] = \A_s[33] ;
  assign \A_s[33]  = A_s[33];
  assign A_so[34] = \A_s[32] ;
  assign \A_s[32]  = A_s[32];
  assign A_so[33] = \A_s[31] ;
  assign \A_s[31]  = A_s[31];
  assign A_so[32] = \A_s[30] ;
  assign \A_s[30]  = A_s[30];
  assign A_so[31] = \A_s[29] ;
  assign \A_s[29]  = A_s[29];
  assign A_so[30] = \A_s[28] ;
  assign \A_s[28]  = A_s[28];
  assign A_so[29] = \A_s[27] ;
  assign \A_s[27]  = A_s[27];
  assign A_so[28] = \A_s[26] ;
  assign \A_s[26]  = A_s[26];
  assign A_so[27] = \A_s[25] ;
  assign \A_s[25]  = A_s[25];
  assign A_so[26] = \A_s[24] ;
  assign \A_s[24]  = A_s[24];
  assign A_so[25] = \A_s[23] ;
  assign \A_s[23]  = A_s[23];
  assign A_so[24] = \A_s[22] ;
  assign \A_s[22]  = A_s[22];
  assign A_so[23] = \A_s[21] ;
  assign \A_s[21]  = A_s[21];
  assign A_so[22] = \A_s[20] ;
  assign \A_s[20]  = A_s[20];
  assign A_so[21] = \A_s[19] ;
  assign \A_s[19]  = A_s[19];
  assign A_so[20] = \A_s[18] ;
  assign \A_s[18]  = A_s[18];
  assign A_so[19] = \A_s[17] ;
  assign \A_s[17]  = A_s[17];
  assign A_so[18] = \A_s[16] ;
  assign \A_s[16]  = A_s[16];
  assign A_so[17] = \A_s[15] ;
  assign \A_s[15]  = A_s[15];
  assign A_so[16] = \A_s[14] ;
  assign \A_s[14]  = A_s[14];
  assign A_so[15] = \A_s[13] ;
  assign \A_s[13]  = A_s[13];
  assign A_so[14] = \A_s[12] ;
  assign \A_s[12]  = A_s[12];
  assign A_so[13] = \A_s[11] ;
  assign \A_s[11]  = A_s[11];
  assign A_so[12] = \A_s[10] ;
  assign \A_s[10]  = A_s[10];
  assign A_so[11] = \A_s[9] ;
  assign \A_s[9]  = A_s[9];
  assign A_so[10] = \A_s[8] ;
  assign \A_s[8]  = A_s[8];
  assign A_so[9] = \A_s[7] ;
  assign \A_s[7]  = A_s[7];
  assign A_so[8] = \A_s[6] ;
  assign \A_s[6]  = A_s[6];
  assign A_so[7] = \A_s[5] ;
  assign \A_s[5]  = A_s[5];
  assign A_so[6] = \A_s[4] ;
  assign \A_s[4]  = A_s[4];
  assign A_so[5] = \A_s[3] ;
  assign \A_s[3]  = A_s[3];
  assign A_so[4] = \A_s[2] ;
  assign \A_s[2]  = A_s[2];
  assign A_so[3] = \A_s[1] ;
  assign \A_s[1]  = A_s[1];
  assign A_so[2] = \A_s[0] ;
  assign \A_s[0]  = A_s[0];
  assign A_nso[45] = \A_ns[43] ;
  assign \A_ns[43]  = A_ns[43];
  assign A_nso[44] = \A_ns[42] ;
  assign \A_ns[42]  = A_ns[42];
  assign A_nso[43] = \A_ns[41] ;
  assign \A_ns[41]  = A_ns[41];
  assign A_nso[42] = \A_ns[40] ;
  assign \A_ns[40]  = A_ns[40];
  assign A_nso[41] = \A_ns[39] ;
  assign \A_ns[39]  = A_ns[39];
  assign A_nso[40] = \A_ns[38] ;
  assign \A_ns[38]  = A_ns[38];
  assign A_nso[39] = \A_ns[37] ;
  assign \A_ns[37]  = A_ns[37];
  assign A_nso[38] = \A_ns[36] ;
  assign \A_ns[36]  = A_ns[36];
  assign A_nso[37] = \A_ns[35] ;
  assign \A_ns[35]  = A_ns[35];
  assign A_nso[36] = \A_ns[34] ;
  assign \A_ns[34]  = A_ns[34];
  assign A_nso[35] = \A_ns[33] ;
  assign \A_ns[33]  = A_ns[33];
  assign A_nso[34] = \A_ns[32] ;
  assign \A_ns[32]  = A_ns[32];
  assign A_nso[33] = \A_ns[31] ;
  assign \A_ns[31]  = A_ns[31];
  assign A_nso[32] = \A_ns[30] ;
  assign \A_ns[30]  = A_ns[30];
  assign A_nso[31] = \A_ns[29] ;
  assign \A_ns[29]  = A_ns[29];
  assign A_nso[30] = \A_ns[28] ;
  assign \A_ns[28]  = A_ns[28];
  assign A_nso[29] = \A_ns[27] ;
  assign \A_ns[27]  = A_ns[27];
  assign A_nso[28] = \A_ns[26] ;
  assign \A_ns[26]  = A_ns[26];
  assign A_nso[27] = \A_ns[25] ;
  assign \A_ns[25]  = A_ns[25];
  assign A_nso[26] = \A_ns[24] ;
  assign \A_ns[24]  = A_ns[24];
  assign A_nso[25] = \A_ns[23] ;
  assign \A_ns[23]  = A_ns[23];
  assign A_nso[24] = \A_ns[22] ;
  assign \A_ns[22]  = A_ns[22];
  assign A_nso[23] = \A_ns[21] ;
  assign \A_ns[21]  = A_ns[21];
  assign A_nso[22] = \A_ns[20] ;
  assign \A_ns[20]  = A_ns[20];
  assign A_nso[21] = \A_ns[19] ;
  assign \A_ns[19]  = A_ns[19];
  assign A_nso[20] = \A_ns[18] ;
  assign \A_ns[18]  = A_ns[18];
  assign A_nso[19] = \A_ns[17] ;
  assign \A_ns[17]  = A_ns[17];
  assign A_nso[18] = \A_ns[16] ;
  assign \A_ns[16]  = A_ns[16];
  assign A_nso[17] = \A_ns[15] ;
  assign \A_ns[15]  = A_ns[15];
  assign A_nso[16] = \A_ns[14] ;
  assign \A_ns[14]  = A_ns[14];
  assign A_nso[15] = \A_ns[13] ;
  assign \A_ns[13]  = A_ns[13];
  assign A_nso[14] = \A_ns[12] ;
  assign \A_ns[12]  = A_ns[12];
  assign A_nso[13] = \A_ns[11] ;
  assign \A_ns[11]  = A_ns[11];
  assign A_nso[12] = \A_ns[10] ;
  assign \A_ns[10]  = A_ns[10];
  assign A_nso[11] = \A_ns[9] ;
  assign \A_ns[9]  = A_ns[9];
  assign A_nso[10] = \A_ns[8] ;
  assign \A_ns[8]  = A_ns[8];
  assign A_nso[9] = \A_ns[7] ;
  assign \A_ns[7]  = A_ns[7];
  assign A_nso[8] = \A_ns[6] ;
  assign \A_ns[6]  = A_ns[6];
  assign A_nso[7] = \A_ns[5] ;
  assign \A_ns[5]  = A_ns[5];
  assign A_nso[6] = \A_ns[4] ;
  assign \A_ns[4]  = A_ns[4];
  assign A_nso[5] = \A_ns[3] ;
  assign \A_ns[3]  = A_ns[3];
  assign A_nso[4] = \A_ns[2] ;
  assign \A_ns[2]  = A_ns[2];
  assign A_nso[3] = \A_ns[1] ;
  assign \A_ns[1]  = A_ns[1];
  assign A_nso[2] = \A_ns[0] ;
  assign \A_ns[0]  = A_ns[0];

  NAND3_X1 U186 ( .A1(B[11]), .A2(n780), .A3(B[12]), .ZN(n96) );
  XOR2_X1 U187 ( .A(B[11]), .B(B[12]), .Z(n184) );
  INV_X1 U2 ( .A(n101), .ZN(O[42]) );
  OAI221_X1 U3 ( .B1(n98), .B2(n690), .C1(n99), .C2(n691), .A(n100), .ZN(O[43]) );
  OAI221_X1 U4 ( .B1(n669), .B2(n690), .C1(n96), .C2(n691), .A(n97), .ZN(O[44]) );
  CLKBUF_X1 U5 ( .A(n682), .Z(n684) );
  CLKBUF_X1 U6 ( .A(n677), .Z(n681) );
  CLKBUF_X1 U7 ( .A(n683), .Z(n687) );
  CLKBUF_X1 U8 ( .A(n778), .Z(n676) );
  CLKBUF_X1 U9 ( .A(n779), .Z(n682) );
  CLKBUF_X1 U10 ( .A(n777), .Z(n671) );
  BUF_X1 U11 ( .A(n683), .Z(n686) );
  BUF_X1 U12 ( .A(n677), .Z(n680) );
  BUF_X1 U13 ( .A(n682), .Z(n685) );
  BUF_X1 U14 ( .A(n676), .Z(n678) );
  BUF_X1 U15 ( .A(n676), .Z(n679) );
  BUF_X1 U16 ( .A(n670), .Z(n673) );
  BUF_X1 U17 ( .A(n670), .Z(n672) );
  BUF_X1 U18 ( .A(n778), .Z(n677) );
  BUF_X1 U19 ( .A(n779), .Z(n683) );
  BUF_X1 U20 ( .A(n671), .Z(n674) );
  BUF_X1 U21 ( .A(n671), .Z(n675) );
  INV_X1 U22 ( .A(n93), .ZN(O[45]) );
  AOI221_X1 U23 ( .B1(n684), .B2(\A_ns[41] ), .C1(n678), .C2(\A_s[41] ), .A(
        n719), .ZN(n101) );
  INV_X1 U24 ( .A(n151), .ZN(O[17]) );
  AOI221_X1 U25 ( .B1(n686), .B2(\A_ns[16] ), .C1(n680), .C2(\A_s[16] ), .A(
        n769), .ZN(n151) );
  INV_X1 U26 ( .A(n152), .ZN(n769) );
  AOI22_X1 U27 ( .A1(\A_ns[15] ), .A2(n689), .B1(\A_s[15] ), .B2(n673), .ZN(
        n152) );
  INV_X1 U28 ( .A(n155), .ZN(O[15]) );
  AOI221_X1 U29 ( .B1(n686), .B2(\A_ns[14] ), .C1(n680), .C2(\A_s[14] ), .A(
        n773), .ZN(n155) );
  INV_X1 U30 ( .A(n156), .ZN(n773) );
  AOI22_X1 U31 ( .A1(\A_ns[13] ), .A2(n689), .B1(\A_s[13] ), .B2(n673), .ZN(
        n156) );
  INV_X1 U32 ( .A(n149), .ZN(O[18]) );
  AOI221_X1 U33 ( .B1(n685), .B2(\A_ns[17] ), .C1(n680), .C2(\A_s[17] ), .A(
        n767), .ZN(n149) );
  INV_X1 U34 ( .A(n150), .ZN(n767) );
  AOI22_X1 U35 ( .A1(\A_ns[16] ), .A2(n689), .B1(\A_s[16] ), .B2(n673), .ZN(
        n150) );
  INV_X1 U36 ( .A(n153), .ZN(O[16]) );
  AOI221_X1 U37 ( .B1(n686), .B2(\A_ns[15] ), .C1(n680), .C2(\A_s[15] ), .A(
        n771), .ZN(n153) );
  INV_X1 U38 ( .A(n154), .ZN(n771) );
  AOI22_X1 U39 ( .A1(\A_ns[14] ), .A2(n689), .B1(\A_s[14] ), .B2(n673), .ZN(
        n154) );
  INV_X1 U40 ( .A(n157), .ZN(O[14]) );
  AOI221_X1 U41 ( .B1(n686), .B2(\A_ns[13] ), .C1(n680), .C2(\A_s[13] ), .A(
        n775), .ZN(n157) );
  INV_X1 U42 ( .A(n158), .ZN(n775) );
  AOI22_X1 U43 ( .A1(\A_ns[12] ), .A2(n689), .B1(\A_s[12] ), .B2(n673), .ZN(
        n158) );
  INV_X1 U44 ( .A(n147), .ZN(O[19]) );
  AOI221_X1 U45 ( .B1(n685), .B2(\A_ns[18] ), .C1(n680), .C2(\A_s[18] ), .A(
        n765), .ZN(n147) );
  INV_X1 U46 ( .A(n148), .ZN(n765) );
  AOI22_X1 U47 ( .A1(\A_ns[17] ), .A2(n689), .B1(\A_s[17] ), .B2(n673), .ZN(
        n148) );
  BUF_X1 U48 ( .A(n777), .Z(n670) );
  INV_X1 U49 ( .A(n99), .ZN(n778) );
  INV_X1 U50 ( .A(n98), .ZN(n779) );
  AOI22_X1 U51 ( .A1(\A_ns[41] ), .A2(n689), .B1(\A_s[41] ), .B2(n675), .ZN(
        n100) );
  INV_X1 U52 ( .A(n135), .ZN(O[25]) );
  AOI221_X1 U53 ( .B1(n685), .B2(\A_ns[24] ), .C1(n679), .C2(\A_s[24] ), .A(
        n753), .ZN(n135) );
  INV_X1 U54 ( .A(n136), .ZN(n753) );
  AOI22_X1 U55 ( .A1(\A_ns[23] ), .A2(n689), .B1(\A_s[23] ), .B2(n673), .ZN(
        n136) );
  AOI221_X1 U56 ( .B1(n689), .B2(\A_ns[43] ), .C1(n675), .C2(\A_s[43] ), .A(
        n716), .ZN(n93) );
  INV_X1 U57 ( .A(n95), .ZN(n716) );
  AOI22_X1 U58 ( .A1(A_ns[44]), .A2(n684), .B1(A_s[44]), .B2(n678), .ZN(n95)
         );
  INV_X1 U59 ( .A(n139), .ZN(O[23]) );
  AOI221_X1 U60 ( .B1(n685), .B2(\A_ns[22] ), .C1(n679), .C2(\A_s[22] ), .A(
        n757), .ZN(n139) );
  INV_X1 U61 ( .A(n140), .ZN(n757) );
  AOI22_X1 U62 ( .A1(\A_ns[21] ), .A2(n689), .B1(\A_s[21] ), .B2(n673), .ZN(
        n140) );
  INV_X1 U63 ( .A(n127), .ZN(O[29]) );
  AOI221_X1 U64 ( .B1(n685), .B2(\A_ns[28] ), .C1(n679), .C2(\A_s[28] ), .A(
        n745), .ZN(n127) );
  INV_X1 U65 ( .A(n128), .ZN(n745) );
  AOI22_X1 U66 ( .A1(\A_ns[27] ), .A2(n688), .B1(\A_s[27] ), .B2(n674), .ZN(
        n128) );
  INV_X1 U67 ( .A(n103), .ZN(O[41]) );
  AOI221_X1 U68 ( .B1(n684), .B2(\A_ns[40] ), .C1(n678), .C2(\A_s[40] ), .A(
        n721), .ZN(n103) );
  INV_X1 U69 ( .A(n104), .ZN(n721) );
  AOI22_X1 U70 ( .A1(\A_ns[39] ), .A2(n689), .B1(\A_s[39] ), .B2(n675), .ZN(
        n104) );
  INV_X1 U71 ( .A(n102), .ZN(n719) );
  AOI22_X1 U72 ( .A1(\A_ns[40] ), .A2(n689), .B1(\A_s[40] ), .B2(n675), .ZN(
        n102) );
  INV_X1 U73 ( .A(n133), .ZN(O[26]) );
  AOI221_X1 U74 ( .B1(n685), .B2(\A_ns[25] ), .C1(n679), .C2(\A_s[25] ), .A(
        n751), .ZN(n133) );
  INV_X1 U75 ( .A(n134), .ZN(n751) );
  AOI22_X1 U76 ( .A1(\A_ns[24] ), .A2(n688), .B1(\A_s[24] ), .B2(n674), .ZN(
        n134) );
  INV_X1 U77 ( .A(n129), .ZN(O[28]) );
  AOI221_X1 U78 ( .B1(n685), .B2(\A_ns[27] ), .C1(n679), .C2(\A_s[27] ), .A(
        n747), .ZN(n129) );
  INV_X1 U79 ( .A(n130), .ZN(n747) );
  AOI22_X1 U80 ( .A1(\A_ns[26] ), .A2(n688), .B1(\A_s[26] ), .B2(n674), .ZN(
        n130) );
  INV_X1 U81 ( .A(n109), .ZN(O[38]) );
  AOI221_X1 U82 ( .B1(n684), .B2(\A_ns[37] ), .C1(n678), .C2(\A_s[37] ), .A(
        n727), .ZN(n109) );
  INV_X1 U83 ( .A(n110), .ZN(n727) );
  AOI22_X1 U84 ( .A1(\A_ns[36] ), .A2(n688), .B1(\A_s[36] ), .B2(n675), .ZN(
        n110) );
  INV_X1 U85 ( .A(n105), .ZN(O[40]) );
  AOI221_X1 U86 ( .B1(n684), .B2(\A_ns[39] ), .C1(n678), .C2(\A_s[39] ), .A(
        n723), .ZN(n105) );
  INV_X1 U87 ( .A(n106), .ZN(n723) );
  AOI22_X1 U88 ( .A1(\A_ns[38] ), .A2(n689), .B1(\A_s[38] ), .B2(n675), .ZN(
        n106) );
  INV_X1 U89 ( .A(n143), .ZN(O[21]) );
  AOI221_X1 U90 ( .B1(n685), .B2(\A_ns[20] ), .C1(n679), .C2(\A_s[20] ), .A(
        n761), .ZN(n143) );
  INV_X1 U91 ( .A(n144), .ZN(n761) );
  AOI22_X1 U92 ( .A1(\A_ns[19] ), .A2(n689), .B1(\A_s[19] ), .B2(n673), .ZN(
        n144) );
  INV_X1 U93 ( .A(n123), .ZN(O[31]) );
  AOI221_X1 U94 ( .B1(n684), .B2(\A_ns[30] ), .C1(n679), .C2(\A_s[30] ), .A(
        n741), .ZN(n123) );
  INV_X1 U95 ( .A(n124), .ZN(n741) );
  AOI22_X1 U96 ( .A1(\A_ns[29] ), .A2(n688), .B1(\A_s[29] ), .B2(n674), .ZN(
        n124) );
  INV_X1 U97 ( .A(n131), .ZN(O[27]) );
  AOI221_X1 U98 ( .B1(n685), .B2(\A_ns[26] ), .C1(n679), .C2(\A_s[26] ), .A(
        n749), .ZN(n131) );
  INV_X1 U99 ( .A(n132), .ZN(n749) );
  AOI22_X1 U100 ( .A1(\A_ns[25] ), .A2(n688), .B1(\A_s[25] ), .B2(n674), .ZN(
        n132) );
  INV_X1 U101 ( .A(n119), .ZN(O[33]) );
  AOI221_X1 U102 ( .B1(n684), .B2(\A_ns[32] ), .C1(n678), .C2(\A_s[32] ), .A(
        n737), .ZN(n119) );
  INV_X1 U103 ( .A(n120), .ZN(n737) );
  AOI22_X1 U104 ( .A1(\A_ns[31] ), .A2(n688), .B1(\A_s[31] ), .B2(n674), .ZN(
        n120) );
  INV_X1 U105 ( .A(n115), .ZN(O[35]) );
  AOI221_X1 U106 ( .B1(n684), .B2(\A_ns[34] ), .C1(n678), .C2(\A_s[34] ), .A(
        n733), .ZN(n115) );
  INV_X1 U107 ( .A(n116), .ZN(n733) );
  AOI22_X1 U108 ( .A1(\A_ns[33] ), .A2(n688), .B1(\A_s[33] ), .B2(n674), .ZN(
        n116) );
  INV_X1 U109 ( .A(n111), .ZN(O[37]) );
  AOI221_X1 U110 ( .B1(n684), .B2(\A_ns[36] ), .C1(n678), .C2(\A_s[36] ), .A(
        n729), .ZN(n111) );
  INV_X1 U111 ( .A(n112), .ZN(n729) );
  AOI22_X1 U112 ( .A1(\A_ns[35] ), .A2(n688), .B1(\A_s[35] ), .B2(n674), .ZN(
        n112) );
  INV_X1 U113 ( .A(n107), .ZN(O[39]) );
  AOI221_X1 U114 ( .B1(n684), .B2(\A_ns[38] ), .C1(n678), .C2(\A_s[38] ), .A(
        n725), .ZN(n107) );
  INV_X1 U115 ( .A(n108), .ZN(n725) );
  AOI22_X1 U116 ( .A1(\A_ns[37] ), .A2(n689), .B1(\A_s[37] ), .B2(n675), .ZN(
        n108) );
  INV_X1 U117 ( .A(n137), .ZN(O[24]) );
  AOI221_X1 U118 ( .B1(n685), .B2(\A_ns[23] ), .C1(n679), .C2(\A_s[23] ), .A(
        n755), .ZN(n137) );
  INV_X1 U119 ( .A(n138), .ZN(n755) );
  AOI22_X1 U120 ( .A1(\A_ns[22] ), .A2(n689), .B1(\A_s[22] ), .B2(n673), .ZN(
        n138) );
  INV_X1 U121 ( .A(n117), .ZN(O[34]) );
  AOI221_X1 U122 ( .B1(n685), .B2(\A_ns[33] ), .C1(n679), .C2(\A_s[33] ), .A(
        n735), .ZN(n117) );
  INV_X1 U123 ( .A(n118), .ZN(n735) );
  AOI22_X1 U124 ( .A1(\A_ns[32] ), .A2(n688), .B1(\A_s[32] ), .B2(n674), .ZN(
        n118) );
  INV_X1 U125 ( .A(n141), .ZN(O[22]) );
  AOI221_X1 U126 ( .B1(n685), .B2(\A_ns[21] ), .C1(n679), .C2(\A_s[21] ), .A(
        n759), .ZN(n141) );
  INV_X1 U127 ( .A(n142), .ZN(n759) );
  AOI22_X1 U128 ( .A1(\A_ns[20] ), .A2(n689), .B1(\A_s[20] ), .B2(n673), .ZN(
        n142) );
  INV_X1 U129 ( .A(n125), .ZN(O[30]) );
  AOI221_X1 U130 ( .B1(n684), .B2(\A_ns[29] ), .C1(n679), .C2(\A_s[29] ), .A(
        n743), .ZN(n125) );
  INV_X1 U131 ( .A(n126), .ZN(n743) );
  AOI22_X1 U132 ( .A1(\A_ns[28] ), .A2(n688), .B1(\A_s[28] ), .B2(n674), .ZN(
        n126) );
  INV_X1 U133 ( .A(n145), .ZN(O[20]) );
  AOI221_X1 U134 ( .B1(n685), .B2(\A_ns[19] ), .C1(n679), .C2(\A_s[19] ), .A(
        n763), .ZN(n145) );
  INV_X1 U135 ( .A(n146), .ZN(n763) );
  AOI22_X1 U136 ( .A1(\A_ns[18] ), .A2(n689), .B1(\A_s[18] ), .B2(n673), .ZN(
        n146) );
  INV_X1 U137 ( .A(n121), .ZN(O[32]) );
  AOI221_X1 U138 ( .B1(n684), .B2(\A_ns[31] ), .C1(n678), .C2(\A_s[31] ), .A(
        n739), .ZN(n121) );
  INV_X1 U139 ( .A(n122), .ZN(n739) );
  AOI22_X1 U140 ( .A1(\A_ns[30] ), .A2(n688), .B1(\A_s[30] ), .B2(n674), .ZN(
        n122) );
  INV_X1 U141 ( .A(n113), .ZN(O[36]) );
  AOI221_X1 U142 ( .B1(n684), .B2(\A_ns[35] ), .C1(n678), .C2(\A_s[35] ), .A(
        n731), .ZN(n113) );
  INV_X1 U143 ( .A(n114), .ZN(n731) );
  AOI22_X1 U144 ( .A1(\A_ns[34] ), .A2(n688), .B1(\A_s[34] ), .B2(n674), .ZN(
        n114) );
  INV_X1 U145 ( .A(n669), .ZN(n689) );
  INV_X1 U146 ( .A(n669), .ZN(n688) );
  NAND2_X1 U147 ( .A1(n184), .A2(n780), .ZN(n99) );
  NAND2_X1 U148 ( .A1(n184), .A2(n99), .ZN(n98) );
  INV_X1 U149 ( .A(n96), .ZN(n777) );
  AOI22_X1 U150 ( .A1(n687), .A2(\A_ns[43] ), .B1(n681), .B2(\A_s[43] ), .ZN(
        n97) );
  OR3_X1 U151 ( .A1(B[11]), .A2(B[12]), .A3(n780), .ZN(n669) );
  INV_X1 U152 ( .A(n161), .ZN(O[12]) );
  AOI221_X1 U153 ( .B1(n686), .B2(\A_ns[11] ), .C1(n680), .C2(\A_s[11] ), .A(
        n714), .ZN(n161) );
  INV_X1 U154 ( .A(n162), .ZN(n714) );
  AOI22_X1 U155 ( .A1(\A_ns[10] ), .A2(n688), .B1(\A_s[10] ), .B2(n672), .ZN(
        n162) );
  INV_X1 U156 ( .A(B[13]), .ZN(n780) );
  INV_X1 U157 ( .A(n159), .ZN(O[13]) );
  AOI221_X1 U158 ( .B1(n686), .B2(\A_ns[12] ), .C1(n680), .C2(\A_s[12] ), .A(
        n776), .ZN(n159) );
  INV_X1 U159 ( .A(n160), .ZN(n776) );
  AOI22_X1 U160 ( .A1(\A_ns[11] ), .A2(n688), .B1(\A_s[11] ), .B2(n672), .ZN(
        n160) );
  INV_X1 U161 ( .A(n163), .ZN(O[11]) );
  AOI221_X1 U162 ( .B1(n686), .B2(\A_ns[10] ), .C1(n680), .C2(\A_s[10] ), .A(
        n712), .ZN(n163) );
  INV_X1 U163 ( .A(n171), .ZN(O[7]) );
  AOI221_X1 U164 ( .B1(n686), .B2(\A_ns[6] ), .C1(n680), .C2(\A_s[6] ), .A(
        n704), .ZN(n171) );
  INV_X1 U165 ( .A(n172), .ZN(n704) );
  INV_X1 U166 ( .A(n169), .ZN(O[8]) );
  AOI221_X1 U167 ( .B1(n686), .B2(\A_ns[7] ), .C1(n680), .C2(\A_s[7] ), .A(
        n706), .ZN(n169) );
  INV_X1 U168 ( .A(n170), .ZN(n706) );
  INV_X1 U169 ( .A(n167), .ZN(O[9]) );
  AOI221_X1 U170 ( .B1(n686), .B2(\A_ns[8] ), .C1(n680), .C2(\A_s[8] ), .A(
        n708), .ZN(n167) );
  INV_X1 U171 ( .A(n168), .ZN(n708) );
  INV_X1 U172 ( .A(n165), .ZN(O[10]) );
  AOI221_X1 U173 ( .B1(n686), .B2(\A_ns[9] ), .C1(n680), .C2(\A_s[9] ), .A(
        n710), .ZN(n165) );
  INV_X1 U174 ( .A(n183), .ZN(O[1]) );
  AOI22_X1 U175 ( .A1(n678), .A2(\A_s[0] ), .B1(n687), .B2(\A_ns[0] ), .ZN(
        n183) );
  INV_X1 U176 ( .A(n181), .ZN(O[2]) );
  AOI221_X1 U177 ( .B1(n687), .B2(\A_ns[1] ), .C1(n678), .C2(\A_s[1] ), .A(
        n694), .ZN(n181) );
  INV_X1 U178 ( .A(n182), .ZN(n694) );
  INV_X1 U179 ( .A(n179), .ZN(O[3]) );
  AOI221_X1 U180 ( .B1(n687), .B2(\A_ns[2] ), .C1(n681), .C2(\A_s[2] ), .A(
        n696), .ZN(n179) );
  INV_X1 U181 ( .A(n180), .ZN(n696) );
  INV_X1 U182 ( .A(n177), .ZN(O[4]) );
  AOI221_X1 U183 ( .B1(n687), .B2(\A_ns[3] ), .C1(n681), .C2(\A_s[3] ), .A(
        n698), .ZN(n177) );
  INV_X1 U184 ( .A(n178), .ZN(n698) );
  INV_X1 U185 ( .A(n175), .ZN(O[5]) );
  AOI221_X1 U188 ( .B1(n686), .B2(\A_ns[4] ), .C1(n681), .C2(\A_s[4] ), .A(
        n700), .ZN(n175) );
  INV_X1 U189 ( .A(n176), .ZN(n700) );
  INV_X1 U190 ( .A(n173), .ZN(O[6]) );
  AOI221_X1 U191 ( .B1(n686), .B2(\A_ns[5] ), .C1(n681), .C2(\A_s[5] ), .A(
        n702), .ZN(n173) );
  INV_X1 U192 ( .A(n174), .ZN(n702) );
  INV_X1 U193 ( .A(n166), .ZN(n710) );
  AOI22_X1 U194 ( .A1(\A_ns[8] ), .A2(n688), .B1(\A_s[8] ), .B2(n672), .ZN(
        n166) );
  INV_X1 U195 ( .A(n164), .ZN(n712) );
  AOI22_X1 U196 ( .A1(\A_ns[9] ), .A2(n688), .B1(\A_s[9] ), .B2(n672), .ZN(
        n164) );
  AOI22_X1 U197 ( .A1(\A_ns[0] ), .A2(n688), .B1(\A_s[0] ), .B2(n672), .ZN(
        n182) );
  AOI22_X1 U198 ( .A1(\A_ns[1] ), .A2(n688), .B1(\A_s[1] ), .B2(n672), .ZN(
        n180) );
  AOI22_X1 U199 ( .A1(\A_ns[2] ), .A2(n688), .B1(\A_s[2] ), .B2(n672), .ZN(
        n178) );
  AOI22_X1 U200 ( .A1(\A_ns[3] ), .A2(n688), .B1(\A_s[3] ), .B2(n672), .ZN(
        n176) );
  AOI22_X1 U201 ( .A1(\A_ns[4] ), .A2(n688), .B1(\A_s[4] ), .B2(n672), .ZN(
        n174) );
  AOI22_X1 U202 ( .A1(\A_ns[5] ), .A2(n688), .B1(\A_s[5] ), .B2(n672), .ZN(
        n172) );
  AOI22_X1 U203 ( .A1(\A_ns[6] ), .A2(n688), .B1(\A_s[6] ), .B2(n672), .ZN(
        n170) );
  AOI22_X1 U204 ( .A1(\A_ns[7] ), .A2(n688), .B1(\A_s[7] ), .B2(n672), .ZN(
        n168) );
  INV_X1 U205 ( .A(\A_ns[42] ), .ZN(n690) );
  INV_X1 U206 ( .A(\A_s[42] ), .ZN(n691) );
endmodule


module BOOTHENC_NBIT48_i14 ( A_s, A_ns, B, O, A_so, A_nso );
  input [47:0] A_s;
  input [47:0] A_ns;
  input [47:0] B;
  output [47:0] O;
  output [47:0] A_so;
  output [47:0] A_nso;
  wire   \A_s[45] , \A_s[44] , \A_s[43] , \A_s[42] , \A_s[41] , \A_s[40] ,
         \A_s[39] , \A_s[38] , \A_s[37] , \A_s[36] , \A_s[35] , \A_s[34] ,
         \A_s[33] , \A_s[32] , \A_s[31] , \A_s[30] , \A_s[29] , \A_s[28] ,
         \A_s[27] , \A_s[26] , \A_s[25] , \A_s[24] , \A_s[23] , \A_s[22] ,
         \A_s[21] , \A_s[20] , \A_s[19] , \A_s[18] , \A_s[17] , \A_s[16] ,
         \A_s[15] , \A_s[14] , \A_s[13] , \A_s[12] , \A_s[11] , \A_s[10] ,
         \A_s[9] , \A_s[8] , \A_s[7] , \A_s[6] , \A_s[5] , \A_s[4] , \A_s[3] ,
         \A_s[2] , \A_s[1] , \A_s[0] , \A_ns[45] , \A_ns[44] , \A_ns[43] ,
         \A_ns[42] , \A_ns[41] , \A_ns[40] , \A_ns[39] , \A_ns[38] ,
         \A_ns[37] , \A_ns[36] , \A_ns[35] , \A_ns[34] , \A_ns[33] ,
         \A_ns[32] , \A_ns[31] , \A_ns[30] , \A_ns[29] , \A_ns[28] ,
         \A_ns[27] , \A_ns[26] , \A_ns[25] , \A_ns[24] , \A_ns[23] ,
         \A_ns[22] , \A_ns[21] , \A_ns[20] , \A_ns[19] , \A_ns[18] ,
         \A_ns[17] , \A_ns[16] , \A_ns[15] , \A_ns[14] , \A_ns[13] ,
         \A_ns[12] , \A_ns[11] , \A_ns[10] , \A_ns[9] , \A_ns[8] , \A_ns[7] ,
         \A_ns[6] , \A_ns[5] , \A_ns[4] , \A_ns[3] , \A_ns[2] , \A_ns[1] ,
         \A_ns[0] , n97, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n722, n724,
         n726, n728, n730, n732, n734, n736, n738, n740, n742, n744, n746,
         n748, n751, n753, n755, n757, n759, n761, n763, n765, n767, n769,
         n771, n773, n775, n777, n779, n781, n783, n785, n787, n789, n791,
         n793, n795, n797, n799, n801, n803, n805, n807, n808, n809, n810,
         n811, n812;
  assign A_nso[0] = 1'b0;
  assign A_nso[1] = 1'b0;
  assign A_so[0] = 1'b0;
  assign A_so[1] = 1'b0;
  assign O[0] = 1'b0;
  assign A_so[47] = \A_s[45] ;
  assign \A_s[45]  = A_s[45];
  assign A_so[46] = \A_s[44] ;
  assign \A_s[44]  = A_s[44];
  assign A_so[45] = \A_s[43] ;
  assign \A_s[43]  = A_s[43];
  assign A_so[44] = \A_s[42] ;
  assign \A_s[42]  = A_s[42];
  assign A_so[43] = \A_s[41] ;
  assign \A_s[41]  = A_s[41];
  assign A_so[42] = \A_s[40] ;
  assign \A_s[40]  = A_s[40];
  assign A_so[41] = \A_s[39] ;
  assign \A_s[39]  = A_s[39];
  assign A_so[40] = \A_s[38] ;
  assign \A_s[38]  = A_s[38];
  assign A_so[39] = \A_s[37] ;
  assign \A_s[37]  = A_s[37];
  assign A_so[38] = \A_s[36] ;
  assign \A_s[36]  = A_s[36];
  assign A_so[37] = \A_s[35] ;
  assign \A_s[35]  = A_s[35];
  assign A_so[36] = \A_s[34] ;
  assign \A_s[34]  = A_s[34];
  assign A_so[35] = \A_s[33] ;
  assign \A_s[33]  = A_s[33];
  assign A_so[34] = \A_s[32] ;
  assign \A_s[32]  = A_s[32];
  assign A_so[33] = \A_s[31] ;
  assign \A_s[31]  = A_s[31];
  assign A_so[32] = \A_s[30] ;
  assign \A_s[30]  = A_s[30];
  assign A_so[31] = \A_s[29] ;
  assign \A_s[29]  = A_s[29];
  assign A_so[30] = \A_s[28] ;
  assign \A_s[28]  = A_s[28];
  assign A_so[29] = \A_s[27] ;
  assign \A_s[27]  = A_s[27];
  assign A_so[28] = \A_s[26] ;
  assign \A_s[26]  = A_s[26];
  assign A_so[27] = \A_s[25] ;
  assign \A_s[25]  = A_s[25];
  assign A_so[26] = \A_s[24] ;
  assign \A_s[24]  = A_s[24];
  assign A_so[25] = \A_s[23] ;
  assign \A_s[23]  = A_s[23];
  assign A_so[24] = \A_s[22] ;
  assign \A_s[22]  = A_s[22];
  assign A_so[23] = \A_s[21] ;
  assign \A_s[21]  = A_s[21];
  assign A_so[22] = \A_s[20] ;
  assign \A_s[20]  = A_s[20];
  assign A_so[21] = \A_s[19] ;
  assign \A_s[19]  = A_s[19];
  assign A_so[20] = \A_s[18] ;
  assign \A_s[18]  = A_s[18];
  assign A_so[19] = \A_s[17] ;
  assign \A_s[17]  = A_s[17];
  assign A_so[18] = \A_s[16] ;
  assign \A_s[16]  = A_s[16];
  assign A_so[17] = \A_s[15] ;
  assign \A_s[15]  = A_s[15];
  assign A_so[16] = \A_s[14] ;
  assign \A_s[14]  = A_s[14];
  assign A_so[15] = \A_s[13] ;
  assign \A_s[13]  = A_s[13];
  assign A_so[14] = \A_s[12] ;
  assign \A_s[12]  = A_s[12];
  assign A_so[13] = \A_s[11] ;
  assign \A_s[11]  = A_s[11];
  assign A_so[12] = \A_s[10] ;
  assign \A_s[10]  = A_s[10];
  assign A_so[11] = \A_s[9] ;
  assign \A_s[9]  = A_s[9];
  assign A_so[10] = \A_s[8] ;
  assign \A_s[8]  = A_s[8];
  assign A_so[9] = \A_s[7] ;
  assign \A_s[7]  = A_s[7];
  assign A_so[8] = \A_s[6] ;
  assign \A_s[6]  = A_s[6];
  assign A_so[7] = \A_s[5] ;
  assign \A_s[5]  = A_s[5];
  assign A_so[6] = \A_s[4] ;
  assign \A_s[4]  = A_s[4];
  assign A_so[5] = \A_s[3] ;
  assign \A_s[3]  = A_s[3];
  assign A_so[4] = \A_s[2] ;
  assign \A_s[2]  = A_s[2];
  assign A_so[3] = \A_s[1] ;
  assign \A_s[1]  = A_s[1];
  assign A_so[2] = \A_s[0] ;
  assign \A_s[0]  = A_s[0];
  assign A_nso[47] = \A_ns[45] ;
  assign \A_ns[45]  = A_ns[45];
  assign A_nso[46] = \A_ns[44] ;
  assign \A_ns[44]  = A_ns[44];
  assign A_nso[45] = \A_ns[43] ;
  assign \A_ns[43]  = A_ns[43];
  assign A_nso[44] = \A_ns[42] ;
  assign \A_ns[42]  = A_ns[42];
  assign A_nso[43] = \A_ns[41] ;
  assign \A_ns[41]  = A_ns[41];
  assign A_nso[42] = \A_ns[40] ;
  assign \A_ns[40]  = A_ns[40];
  assign A_nso[41] = \A_ns[39] ;
  assign \A_ns[39]  = A_ns[39];
  assign A_nso[40] = \A_ns[38] ;
  assign \A_ns[38]  = A_ns[38];
  assign A_nso[39] = \A_ns[37] ;
  assign \A_ns[37]  = A_ns[37];
  assign A_nso[38] = \A_ns[36] ;
  assign \A_ns[36]  = A_ns[36];
  assign A_nso[37] = \A_ns[35] ;
  assign \A_ns[35]  = A_ns[35];
  assign A_nso[36] = \A_ns[34] ;
  assign \A_ns[34]  = A_ns[34];
  assign A_nso[35] = \A_ns[33] ;
  assign \A_ns[33]  = A_ns[33];
  assign A_nso[34] = \A_ns[32] ;
  assign \A_ns[32]  = A_ns[32];
  assign A_nso[33] = \A_ns[31] ;
  assign \A_ns[31]  = A_ns[31];
  assign A_nso[32] = \A_ns[30] ;
  assign \A_ns[30]  = A_ns[30];
  assign A_nso[31] = \A_ns[29] ;
  assign \A_ns[29]  = A_ns[29];
  assign A_nso[30] = \A_ns[28] ;
  assign \A_ns[28]  = A_ns[28];
  assign A_nso[29] = \A_ns[27] ;
  assign \A_ns[27]  = A_ns[27];
  assign A_nso[28] = \A_ns[26] ;
  assign \A_ns[26]  = A_ns[26];
  assign A_nso[27] = \A_ns[25] ;
  assign \A_ns[25]  = A_ns[25];
  assign A_nso[26] = \A_ns[24] ;
  assign \A_ns[24]  = A_ns[24];
  assign A_nso[25] = \A_ns[23] ;
  assign \A_ns[23]  = A_ns[23];
  assign A_nso[24] = \A_ns[22] ;
  assign \A_ns[22]  = A_ns[22];
  assign A_nso[23] = \A_ns[21] ;
  assign \A_ns[21]  = A_ns[21];
  assign A_nso[22] = \A_ns[20] ;
  assign \A_ns[20]  = A_ns[20];
  assign A_nso[21] = \A_ns[19] ;
  assign \A_ns[19]  = A_ns[19];
  assign A_nso[20] = \A_ns[18] ;
  assign \A_ns[18]  = A_ns[18];
  assign A_nso[19] = \A_ns[17] ;
  assign \A_ns[17]  = A_ns[17];
  assign A_nso[18] = \A_ns[16] ;
  assign \A_ns[16]  = A_ns[16];
  assign A_nso[17] = \A_ns[15] ;
  assign \A_ns[15]  = A_ns[15];
  assign A_nso[16] = \A_ns[14] ;
  assign \A_ns[14]  = A_ns[14];
  assign A_nso[15] = \A_ns[13] ;
  assign \A_ns[13]  = A_ns[13];
  assign A_nso[14] = \A_ns[12] ;
  assign \A_ns[12]  = A_ns[12];
  assign A_nso[13] = \A_ns[11] ;
  assign \A_ns[11]  = A_ns[11];
  assign A_nso[12] = \A_ns[10] ;
  assign \A_ns[10]  = A_ns[10];
  assign A_nso[11] = \A_ns[9] ;
  assign \A_ns[9]  = A_ns[9];
  assign A_nso[10] = \A_ns[8] ;
  assign \A_ns[8]  = A_ns[8];
  assign A_nso[9] = \A_ns[7] ;
  assign \A_ns[7]  = A_ns[7];
  assign A_nso[8] = \A_ns[6] ;
  assign \A_ns[6]  = A_ns[6];
  assign A_nso[7] = \A_ns[5] ;
  assign \A_ns[5]  = A_ns[5];
  assign A_nso[6] = \A_ns[4] ;
  assign \A_ns[4]  = A_ns[4];
  assign A_nso[5] = \A_ns[3] ;
  assign \A_ns[3]  = A_ns[3];
  assign A_nso[4] = \A_ns[2] ;
  assign \A_ns[2]  = A_ns[2];
  assign A_nso[3] = \A_ns[1] ;
  assign \A_ns[1]  = A_ns[1];
  assign A_nso[2] = \A_ns[0] ;
  assign \A_ns[0]  = A_ns[0];

  NAND3_X1 U194 ( .A1(B[13]), .A2(n812), .A3(B[14]), .ZN(n100) );
  XOR2_X1 U195 ( .A(B[13]), .B(B[14]), .Z(n192) );
  OAI221_X1 U2 ( .B1(n697), .B2(n718), .C1(n100), .C2(n719), .A(n101), .ZN(
        O[46]) );
  AOI221_X1 U3 ( .B1(n717), .B2(\A_ns[45] ), .C1(n703), .C2(\A_s[45] ), .A(
        n748), .ZN(n97) );
  INV_X1 U4 ( .A(n145), .ZN(O[24]) );
  INV_X1 U5 ( .A(n97), .ZN(O[47]) );
  CLKBUF_X1 U6 ( .A(n704), .Z(n706) );
  CLKBUF_X1 U7 ( .A(n705), .Z(n709) );
  CLKBUF_X1 U8 ( .A(n711), .Z(n715) );
  CLKBUF_X1 U9 ( .A(n810), .Z(n704) );
  CLKBUF_X1 U10 ( .A(n811), .Z(n710) );
  CLKBUF_X1 U11 ( .A(n698), .Z(n700) );
  CLKBUF_X1 U12 ( .A(n809), .Z(n699) );
  INV_X1 U13 ( .A(n99), .ZN(n748) );
  AOI22_X1 U14 ( .A1(A_ns[46]), .A2(n712), .B1(A_s[46]), .B2(n706), .ZN(n99)
         );
  BUF_X1 U15 ( .A(n711), .Z(n714) );
  BUF_X1 U16 ( .A(n705), .Z(n708) );
  BUF_X1 U17 ( .A(n710), .Z(n712) );
  BUF_X1 U18 ( .A(n710), .Z(n713) );
  BUF_X1 U19 ( .A(n704), .Z(n707) );
  BUF_X1 U20 ( .A(n698), .Z(n701) );
  BUF_X1 U21 ( .A(n810), .Z(n705) );
  BUF_X1 U22 ( .A(n811), .Z(n711) );
  BUF_X1 U23 ( .A(n699), .Z(n702) );
  BUF_X1 U24 ( .A(n699), .Z(n703) );
  BUF_X1 U25 ( .A(n809), .Z(n698) );
  INV_X1 U26 ( .A(n103), .ZN(n810) );
  INV_X1 U27 ( .A(n102), .ZN(n811) );
  AOI221_X1 U28 ( .B1(n713), .B2(\A_ns[23] ), .C1(n707), .C2(\A_s[23] ), .A(
        n791), .ZN(n145) );
  INV_X1 U29 ( .A(n146), .ZN(n791) );
  AOI22_X1 U30 ( .A1(\A_ns[22] ), .A2(n716), .B1(\A_s[22] ), .B2(n701), .ZN(
        n146) );
  INV_X1 U31 ( .A(n127), .ZN(O[33]) );
  AOI221_X1 U32 ( .B1(n712), .B2(\A_ns[32] ), .C1(n707), .C2(\A_s[32] ), .A(
        n773), .ZN(n127) );
  INV_X1 U33 ( .A(n128), .ZN(n773) );
  AOI22_X1 U34 ( .A1(\A_ns[31] ), .A2(n717), .B1(\A_s[31] ), .B2(n702), .ZN(
        n128) );
  INV_X1 U35 ( .A(n107), .ZN(O[43]) );
  AOI221_X1 U36 ( .B1(n712), .B2(\A_ns[42] ), .C1(n706), .C2(\A_s[42] ), .A(
        n753), .ZN(n107) );
  INV_X1 U37 ( .A(n108), .ZN(n753) );
  AOI22_X1 U38 ( .A1(\A_ns[41] ), .A2(n717), .B1(\A_s[41] ), .B2(n703), .ZN(
        n108) );
  INV_X1 U39 ( .A(n153), .ZN(O[20]) );
  AOI221_X1 U40 ( .B1(n713), .B2(\A_ns[19] ), .C1(n708), .C2(\A_s[19] ), .A(
        n799), .ZN(n153) );
  INV_X1 U41 ( .A(n154), .ZN(n799) );
  AOI22_X1 U42 ( .A1(\A_ns[18] ), .A2(n716), .B1(\A_s[18] ), .B2(n701), .ZN(
        n154) );
  INV_X1 U43 ( .A(n157), .ZN(O[18]) );
  AOI221_X1 U44 ( .B1(n714), .B2(\A_ns[17] ), .C1(n708), .C2(\A_s[17] ), .A(
        n803), .ZN(n157) );
  INV_X1 U45 ( .A(n158), .ZN(n803) );
  AOI22_X1 U46 ( .A1(\A_ns[16] ), .A2(n716), .B1(\A_s[16] ), .B2(n701), .ZN(
        n158) );
  INV_X1 U47 ( .A(n139), .ZN(O[27]) );
  AOI221_X1 U48 ( .B1(n713), .B2(\A_ns[26] ), .C1(n707), .C2(\A_s[26] ), .A(
        n785), .ZN(n139) );
  INV_X1 U49 ( .A(n140), .ZN(n785) );
  AOI22_X1 U50 ( .A1(\A_ns[25] ), .A2(n717), .B1(\A_s[25] ), .B2(n702), .ZN(
        n140) );
  INV_X1 U51 ( .A(n155), .ZN(O[19]) );
  AOI221_X1 U52 ( .B1(n714), .B2(\A_ns[18] ), .C1(n708), .C2(\A_s[18] ), .A(
        n801), .ZN(n155) );
  INV_X1 U53 ( .A(n156), .ZN(n801) );
  AOI22_X1 U54 ( .A1(\A_ns[17] ), .A2(n716), .B1(\A_s[17] ), .B2(n701), .ZN(
        n156) );
  INV_X1 U55 ( .A(n141), .ZN(O[26]) );
  AOI221_X1 U56 ( .B1(n713), .B2(\A_ns[25] ), .C1(n707), .C2(\A_s[25] ), .A(
        n787), .ZN(n141) );
  INV_X1 U57 ( .A(n142), .ZN(n787) );
  AOI22_X1 U58 ( .A1(\A_ns[24] ), .A2(n717), .B1(\A_s[24] ), .B2(n702), .ZN(
        n142) );
  INV_X1 U59 ( .A(n159), .ZN(O[17]) );
  AOI221_X1 U60 ( .B1(n714), .B2(\A_ns[16] ), .C1(n708), .C2(\A_s[16] ), .A(
        n805), .ZN(n159) );
  INV_X1 U61 ( .A(n160), .ZN(n805) );
  AOI22_X1 U62 ( .A1(\A_ns[15] ), .A2(n716), .B1(\A_s[15] ), .B2(n701), .ZN(
        n160) );
  INV_X1 U63 ( .A(n115), .ZN(O[39]) );
  AOI221_X1 U64 ( .B1(n712), .B2(\A_ns[38] ), .C1(n706), .C2(\A_s[38] ), .A(
        n761), .ZN(n115) );
  INV_X1 U65 ( .A(n116), .ZN(n761) );
  AOI22_X1 U66 ( .A1(\A_ns[37] ), .A2(n717), .B1(\A_s[37] ), .B2(n703), .ZN(
        n116) );
  INV_X1 U67 ( .A(n137), .ZN(O[28]) );
  AOI221_X1 U68 ( .B1(n713), .B2(\A_ns[27] ), .C1(n707), .C2(\A_s[27] ), .A(
        n783), .ZN(n137) );
  INV_X1 U69 ( .A(n138), .ZN(n783) );
  AOI22_X1 U70 ( .A1(\A_ns[26] ), .A2(n717), .B1(\A_s[26] ), .B2(n702), .ZN(
        n138) );
  INV_X1 U71 ( .A(n117), .ZN(O[38]) );
  AOI221_X1 U72 ( .B1(n712), .B2(\A_ns[37] ), .C1(n706), .C2(\A_s[37] ), .A(
        n763), .ZN(n117) );
  INV_X1 U73 ( .A(n118), .ZN(n763) );
  AOI22_X1 U74 ( .A1(\A_ns[36] ), .A2(n717), .B1(\A_s[36] ), .B2(n703), .ZN(
        n118) );
  INV_X1 U75 ( .A(n113), .ZN(O[40]) );
  AOI221_X1 U76 ( .B1(n712), .B2(\A_ns[39] ), .C1(n706), .C2(\A_s[39] ), .A(
        n759), .ZN(n113) );
  INV_X1 U77 ( .A(n114), .ZN(n759) );
  AOI22_X1 U78 ( .A1(\A_ns[38] ), .A2(n717), .B1(\A_s[38] ), .B2(n703), .ZN(
        n114) );
  INV_X1 U79 ( .A(n135), .ZN(O[29]) );
  AOI221_X1 U80 ( .B1(n713), .B2(\A_ns[28] ), .C1(n707), .C2(\A_s[28] ), .A(
        n781), .ZN(n135) );
  INV_X1 U81 ( .A(n136), .ZN(n781) );
  AOI22_X1 U82 ( .A1(\A_ns[27] ), .A2(n717), .B1(\A_s[27] ), .B2(n702), .ZN(
        n136) );
  INV_X1 U83 ( .A(n111), .ZN(O[41]) );
  AOI221_X1 U84 ( .B1(n712), .B2(\A_ns[40] ), .C1(n706), .C2(\A_s[40] ), .A(
        n757), .ZN(n111) );
  INV_X1 U85 ( .A(n112), .ZN(n757) );
  AOI22_X1 U86 ( .A1(\A_ns[39] ), .A2(n717), .B1(\A_s[39] ), .B2(n703), .ZN(
        n112) );
  INV_X1 U87 ( .A(n131), .ZN(O[31]) );
  AOI221_X1 U88 ( .B1(n713), .B2(\A_ns[30] ), .C1(n707), .C2(\A_s[30] ), .A(
        n777), .ZN(n131) );
  INV_X1 U89 ( .A(n132), .ZN(n777) );
  AOI22_X1 U90 ( .A1(\A_ns[29] ), .A2(n717), .B1(\A_s[29] ), .B2(n702), .ZN(
        n132) );
  INV_X1 U91 ( .A(n143), .ZN(O[25]) );
  AOI221_X1 U92 ( .B1(n713), .B2(\A_ns[24] ), .C1(n707), .C2(\A_s[24] ), .A(
        n789), .ZN(n143) );
  INV_X1 U93 ( .A(n144), .ZN(n789) );
  AOI22_X1 U94 ( .A1(\A_ns[23] ), .A2(n716), .B1(\A_s[23] ), .B2(n701), .ZN(
        n144) );
  INV_X1 U95 ( .A(n161), .ZN(O[16]) );
  AOI221_X1 U96 ( .B1(n714), .B2(\A_ns[15] ), .C1(n708), .C2(\A_s[15] ), .A(
        n807), .ZN(n161) );
  INV_X1 U97 ( .A(n162), .ZN(n807) );
  AOI22_X1 U98 ( .A1(\A_ns[14] ), .A2(n716), .B1(\A_s[14] ), .B2(n701), .ZN(
        n162) );
  INV_X1 U99 ( .A(n123), .ZN(O[35]) );
  AOI221_X1 U100 ( .B1(n712), .B2(\A_ns[34] ), .C1(n706), .C2(\A_s[34] ), .A(
        n769), .ZN(n123) );
  INV_X1 U101 ( .A(n124), .ZN(n769) );
  AOI22_X1 U102 ( .A1(\A_ns[33] ), .A2(n717), .B1(\A_s[33] ), .B2(n702), .ZN(
        n124) );
  INV_X1 U103 ( .A(n119), .ZN(O[37]) );
  AOI221_X1 U104 ( .B1(n712), .B2(\A_ns[36] ), .C1(n706), .C2(\A_s[36] ), .A(
        n765), .ZN(n119) );
  INV_X1 U105 ( .A(n120), .ZN(n765) );
  AOI22_X1 U106 ( .A1(\A_ns[35] ), .A2(n717), .B1(\A_s[35] ), .B2(n702), .ZN(
        n120) );
  INV_X1 U107 ( .A(n147), .ZN(O[23]) );
  AOI221_X1 U108 ( .B1(n713), .B2(\A_ns[22] ), .C1(n707), .C2(\A_s[22] ), .A(
        n793), .ZN(n147) );
  INV_X1 U109 ( .A(n148), .ZN(n793) );
  AOI22_X1 U110 ( .A1(\A_ns[21] ), .A2(n716), .B1(\A_s[21] ), .B2(n701), .ZN(
        n148) );
  INV_X1 U111 ( .A(n151), .ZN(O[21]) );
  AOI221_X1 U112 ( .B1(n713), .B2(\A_ns[20] ), .C1(n708), .C2(\A_s[20] ), .A(
        n797), .ZN(n151) );
  INV_X1 U113 ( .A(n152), .ZN(n797) );
  AOI22_X1 U114 ( .A1(\A_ns[19] ), .A2(n716), .B1(\A_s[19] ), .B2(n701), .ZN(
        n152) );
  INV_X1 U115 ( .A(n129), .ZN(O[32]) );
  AOI221_X1 U116 ( .B1(n712), .B2(\A_ns[31] ), .C1(n707), .C2(\A_s[31] ), .A(
        n775), .ZN(n129) );
  INV_X1 U117 ( .A(n130), .ZN(n775) );
  AOI22_X1 U118 ( .A1(\A_ns[30] ), .A2(n717), .B1(\A_s[30] ), .B2(n702), .ZN(
        n130) );
  INV_X1 U119 ( .A(n125), .ZN(O[34]) );
  AOI221_X1 U120 ( .B1(n712), .B2(\A_ns[33] ), .C1(n706), .C2(\A_s[33] ), .A(
        n771), .ZN(n125) );
  INV_X1 U121 ( .A(n126), .ZN(n771) );
  AOI22_X1 U122 ( .A1(\A_ns[32] ), .A2(n717), .B1(\A_s[32] ), .B2(n702), .ZN(
        n126) );
  INV_X1 U123 ( .A(n121), .ZN(O[36]) );
  AOI221_X1 U124 ( .B1(n713), .B2(\A_ns[35] ), .C1(n707), .C2(\A_s[35] ), .A(
        n767), .ZN(n121) );
  INV_X1 U125 ( .A(n122), .ZN(n767) );
  AOI22_X1 U126 ( .A1(\A_ns[34] ), .A2(n717), .B1(\A_s[34] ), .B2(n702), .ZN(
        n122) );
  INV_X1 U127 ( .A(n149), .ZN(O[22]) );
  AOI221_X1 U128 ( .B1(n713), .B2(\A_ns[21] ), .C1(n707), .C2(\A_s[21] ), .A(
        n795), .ZN(n149) );
  INV_X1 U129 ( .A(n150), .ZN(n795) );
  AOI22_X1 U130 ( .A1(\A_ns[20] ), .A2(n716), .B1(\A_s[20] ), .B2(n701), .ZN(
        n150) );
  INV_X1 U131 ( .A(n133), .ZN(O[30]) );
  AOI221_X1 U132 ( .B1(n713), .B2(\A_ns[29] ), .C1(n707), .C2(\A_s[29] ), .A(
        n779), .ZN(n133) );
  INV_X1 U133 ( .A(n134), .ZN(n779) );
  AOI22_X1 U134 ( .A1(\A_ns[28] ), .A2(n717), .B1(\A_s[28] ), .B2(n702), .ZN(
        n134) );
  OAI221_X1 U135 ( .B1(n102), .B2(n718), .C1(n103), .C2(n719), .A(n104), .ZN(
        O[45]) );
  AOI22_X1 U136 ( .A1(\A_ns[43] ), .A2(n717), .B1(\A_s[43] ), .B2(n703), .ZN(
        n104) );
  INV_X1 U137 ( .A(n109), .ZN(O[42]) );
  AOI221_X1 U138 ( .B1(n712), .B2(\A_ns[41] ), .C1(n706), .C2(\A_s[41] ), .A(
        n755), .ZN(n109) );
  INV_X1 U139 ( .A(n110), .ZN(n755) );
  AOI22_X1 U140 ( .A1(\A_ns[40] ), .A2(n717), .B1(\A_s[40] ), .B2(n703), .ZN(
        n110) );
  INV_X1 U141 ( .A(n105), .ZN(O[44]) );
  AOI221_X1 U142 ( .B1(n712), .B2(\A_ns[43] ), .C1(n706), .C2(\A_s[43] ), .A(
        n751), .ZN(n105) );
  INV_X1 U143 ( .A(n106), .ZN(n751) );
  AOI22_X1 U144 ( .A1(\A_ns[42] ), .A2(n717), .B1(\A_s[42] ), .B2(n703), .ZN(
        n106) );
  AOI22_X1 U145 ( .A1(n715), .A2(\A_ns[45] ), .B1(n709), .B2(\A_s[45] ), .ZN(
        n101) );
  INV_X1 U146 ( .A(n697), .ZN(n716) );
  NAND2_X1 U147 ( .A1(n192), .A2(n812), .ZN(n103) );
  NAND2_X1 U148 ( .A1(n192), .A2(n103), .ZN(n102) );
  INV_X1 U149 ( .A(n100), .ZN(n809) );
  INV_X1 U150 ( .A(n697), .ZN(n717) );
  OR3_X1 U151 ( .A1(B[13]), .A2(B[14]), .A3(n812), .ZN(n697) );
  INV_X1 U152 ( .A(n165), .ZN(O[14]) );
  AOI221_X1 U153 ( .B1(n714), .B2(\A_ns[13] ), .C1(n708), .C2(\A_s[13] ), .A(
        n746), .ZN(n165) );
  INV_X1 U154 ( .A(n166), .ZN(n746) );
  AOI22_X1 U155 ( .A1(\A_ns[12] ), .A2(n716), .B1(\A_s[12] ), .B2(n701), .ZN(
        n166) );
  INV_X1 U156 ( .A(n163), .ZN(O[15]) );
  AOI221_X1 U157 ( .B1(n714), .B2(\A_ns[14] ), .C1(n708), .C2(\A_s[14] ), .A(
        n808), .ZN(n163) );
  INV_X1 U158 ( .A(n164), .ZN(n808) );
  AOI22_X1 U159 ( .A1(\A_ns[13] ), .A2(n716), .B1(\A_s[13] ), .B2(n701), .ZN(
        n164) );
  INV_X1 U160 ( .A(B[15]), .ZN(n812) );
  INV_X1 U161 ( .A(n167), .ZN(O[13]) );
  AOI221_X1 U162 ( .B1(n714), .B2(\A_ns[12] ), .C1(n708), .C2(\A_s[12] ), .A(
        n744), .ZN(n167) );
  INV_X1 U163 ( .A(n179), .ZN(O[7]) );
  AOI221_X1 U164 ( .B1(n714), .B2(\A_ns[6] ), .C1(n709), .C2(\A_s[6] ), .A(
        n732), .ZN(n179) );
  INV_X1 U165 ( .A(n180), .ZN(n732) );
  INV_X1 U166 ( .A(n177), .ZN(O[8]) );
  AOI221_X1 U167 ( .B1(n714), .B2(\A_ns[7] ), .C1(n709), .C2(\A_s[7] ), .A(
        n734), .ZN(n177) );
  INV_X1 U168 ( .A(n178), .ZN(n734) );
  INV_X1 U169 ( .A(n175), .ZN(O[9]) );
  AOI221_X1 U170 ( .B1(n714), .B2(\A_ns[8] ), .C1(n708), .C2(\A_s[8] ), .A(
        n736), .ZN(n175) );
  INV_X1 U171 ( .A(n176), .ZN(n736) );
  INV_X1 U172 ( .A(n173), .ZN(O[10]) );
  AOI221_X1 U173 ( .B1(n714), .B2(\A_ns[9] ), .C1(n708), .C2(\A_s[9] ), .A(
        n738), .ZN(n173) );
  INV_X1 U174 ( .A(n174), .ZN(n738) );
  INV_X1 U175 ( .A(n171), .ZN(O[11]) );
  AOI221_X1 U176 ( .B1(n714), .B2(\A_ns[10] ), .C1(n708), .C2(\A_s[10] ), .A(
        n740), .ZN(n171) );
  INV_X1 U177 ( .A(n172), .ZN(n740) );
  INV_X1 U178 ( .A(n169), .ZN(O[12]) );
  AOI221_X1 U179 ( .B1(n714), .B2(\A_ns[11] ), .C1(n708), .C2(\A_s[11] ), .A(
        n742), .ZN(n169) );
  INV_X1 U180 ( .A(n191), .ZN(O[1]) );
  AOI22_X1 U181 ( .A1(n706), .A2(\A_s[0] ), .B1(n715), .B2(\A_ns[0] ), .ZN(
        n191) );
  INV_X1 U182 ( .A(n189), .ZN(O[2]) );
  AOI221_X1 U183 ( .B1(n715), .B2(\A_ns[1] ), .C1(n706), .C2(\A_s[1] ), .A(
        n722), .ZN(n189) );
  INV_X1 U184 ( .A(n190), .ZN(n722) );
  INV_X1 U185 ( .A(n187), .ZN(O[3]) );
  AOI221_X1 U186 ( .B1(n715), .B2(\A_ns[2] ), .C1(n709), .C2(\A_s[2] ), .A(
        n724), .ZN(n187) );
  INV_X1 U187 ( .A(n188), .ZN(n724) );
  INV_X1 U188 ( .A(n185), .ZN(O[4]) );
  AOI221_X1 U189 ( .B1(n715), .B2(\A_ns[3] ), .C1(n709), .C2(\A_s[3] ), .A(
        n726), .ZN(n185) );
  INV_X1 U190 ( .A(n186), .ZN(n726) );
  INV_X1 U191 ( .A(n183), .ZN(O[5]) );
  AOI221_X1 U192 ( .B1(n715), .B2(\A_ns[4] ), .C1(n709), .C2(\A_s[4] ), .A(
        n728), .ZN(n183) );
  INV_X1 U193 ( .A(n184), .ZN(n728) );
  INV_X1 U196 ( .A(n181), .ZN(O[6]) );
  AOI221_X1 U197 ( .B1(n715), .B2(\A_ns[5] ), .C1(n709), .C2(\A_s[5] ), .A(
        n730), .ZN(n181) );
  INV_X1 U198 ( .A(n182), .ZN(n730) );
  INV_X1 U199 ( .A(n170), .ZN(n742) );
  AOI22_X1 U200 ( .A1(\A_ns[10] ), .A2(n717), .B1(\A_s[10] ), .B2(n700), .ZN(
        n170) );
  INV_X1 U201 ( .A(n168), .ZN(n744) );
  AOI22_X1 U202 ( .A1(\A_ns[11] ), .A2(n717), .B1(\A_s[11] ), .B2(n700), .ZN(
        n168) );
  AOI22_X1 U203 ( .A1(\A_ns[0] ), .A2(n717), .B1(\A_s[0] ), .B2(n700), .ZN(
        n190) );
  AOI22_X1 U204 ( .A1(\A_ns[1] ), .A2(n716), .B1(\A_s[1] ), .B2(n700), .ZN(
        n188) );
  AOI22_X1 U205 ( .A1(\A_ns[2] ), .A2(n716), .B1(\A_s[2] ), .B2(n700), .ZN(
        n186) );
  AOI22_X1 U206 ( .A1(\A_ns[3] ), .A2(n716), .B1(\A_s[3] ), .B2(n700), .ZN(
        n184) );
  AOI22_X1 U207 ( .A1(\A_ns[4] ), .A2(n716), .B1(\A_s[4] ), .B2(n700), .ZN(
        n182) );
  AOI22_X1 U208 ( .A1(\A_ns[5] ), .A2(n716), .B1(\A_s[5] ), .B2(n700), .ZN(
        n180) );
  AOI22_X1 U209 ( .A1(\A_ns[6] ), .A2(n716), .B1(\A_s[6] ), .B2(n700), .ZN(
        n178) );
  AOI22_X1 U210 ( .A1(\A_ns[7] ), .A2(n716), .B1(\A_s[7] ), .B2(n700), .ZN(
        n176) );
  AOI22_X1 U211 ( .A1(\A_ns[8] ), .A2(n716), .B1(\A_s[8] ), .B2(n700), .ZN(
        n174) );
  AOI22_X1 U212 ( .A1(\A_ns[9] ), .A2(n716), .B1(\A_s[9] ), .B2(n700), .ZN(
        n172) );
  INV_X1 U213 ( .A(\A_ns[44] ), .ZN(n718) );
  INV_X1 U214 ( .A(\A_s[44] ), .ZN(n719) );
endmodule


module BOOTHENC_NBIT50_i16 ( A_s, A_ns, B, O, A_so, A_nso );
  input [49:0] A_s;
  input [49:0] A_ns;
  input [49:0] B;
  output [49:0] O;
  output [49:0] A_so;
  output [49:0] A_nso;
  wire   \A_s[47] , \A_s[46] , \A_s[44] , \A_s[43] , \A_s[42] , \A_s[41] ,
         \A_s[40] , \A_s[39] , \A_s[38] , \A_s[37] , \A_s[36] , \A_s[35] ,
         \A_s[33] , \A_s[32] , \A_s[31] , \A_s[30] , \A_s[29] , \A_s[28] ,
         \A_s[14] , \A_s[13] , \A_s[12] , \A_s[11] , \A_s[10] , \A_s[9] ,
         \A_s[8] , \A_s[7] , \A_s[6] , \A_s[5] , \A_s[4] , \A_s[3] , \A_s[2] ,
         \A_s[1] , \A_s[0] , \A_ns[47] , \A_ns[46] , \A_ns[43] , \A_ns[42] ,
         \A_ns[41] , \A_ns[14] , \A_ns[13] , \A_ns[12] , \A_ns[11] ,
         \A_ns[10] , \A_ns[9] , \A_ns[8] , \A_ns[7] , \A_ns[6] , \A_ns[5] ,
         \A_ns[4] , \A_ns[3] , \A_ns[2] , \A_ns[1] , \A_ns[0] , n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n664, n666,
         n668, n670, n672, n674, n676, n678, n680, n682, n684, n686, n688,
         n690, n692, n694, n696, n698, n700, n702, n704, n706, n708, n710,
         n712, n713, n714, n715, n717, n719, n720, n721, n723, n725, n727,
         n729, n731, n733, n735, n737, n739, n741, n743, n745, n747, n749,
         n750, n751, n752, n753, n754, n755, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804;
  assign A_nso[0] = 1'b0;
  assign A_nso[1] = 1'b0;
  assign A_so[0] = 1'b0;
  assign A_so[1] = 1'b0;
  assign O[0] = 1'b0;
  assign A_so[49] = \A_s[47] ;
  assign \A_s[47]  = A_s[47];
  assign A_so[48] = \A_s[46] ;
  assign \A_s[46]  = A_s[46];
  assign A_so[46] = \A_s[44] ;
  assign \A_s[44]  = A_s[44];
  assign A_so[45] = \A_s[43] ;
  assign \A_s[43]  = A_s[43];
  assign A_so[44] = \A_s[42] ;
  assign \A_s[42]  = A_s[42];
  assign A_so[43] = \A_s[41] ;
  assign \A_s[41]  = A_s[41];
  assign A_so[42] = \A_s[40] ;
  assign \A_s[40]  = A_s[40];
  assign A_so[41] = \A_s[39] ;
  assign \A_s[39]  = A_s[39];
  assign A_so[40] = \A_s[38] ;
  assign \A_s[38]  = A_s[38];
  assign A_so[39] = \A_s[37] ;
  assign \A_s[37]  = A_s[37];
  assign A_so[38] = \A_s[36] ;
  assign \A_s[36]  = A_s[36];
  assign A_so[37] = \A_s[35] ;
  assign \A_s[35]  = A_s[35];
  assign A_so[35] = \A_s[33] ;
  assign \A_s[33]  = A_s[33];
  assign A_so[34] = \A_s[32] ;
  assign \A_s[32]  = A_s[32];
  assign A_so[33] = \A_s[31] ;
  assign \A_s[31]  = A_s[31];
  assign A_so[32] = \A_s[30] ;
  assign \A_s[30]  = A_s[30];
  assign A_so[31] = \A_s[29] ;
  assign \A_s[29]  = A_s[29];
  assign A_so[30] = \A_s[28] ;
  assign \A_s[28]  = A_s[28];
  assign A_so[16] = \A_s[14] ;
  assign \A_s[14]  = A_s[14];
  assign A_so[15] = \A_s[13] ;
  assign \A_s[13]  = A_s[13];
  assign A_so[14] = \A_s[12] ;
  assign \A_s[12]  = A_s[12];
  assign A_so[13] = \A_s[11] ;
  assign \A_s[11]  = A_s[11];
  assign A_so[12] = \A_s[10] ;
  assign \A_s[10]  = A_s[10];
  assign A_so[11] = \A_s[9] ;
  assign \A_s[9]  = A_s[9];
  assign A_so[10] = \A_s[8] ;
  assign \A_s[8]  = A_s[8];
  assign A_so[9] = \A_s[7] ;
  assign \A_s[7]  = A_s[7];
  assign A_so[8] = \A_s[6] ;
  assign \A_s[6]  = A_s[6];
  assign A_so[7] = \A_s[5] ;
  assign \A_s[5]  = A_s[5];
  assign A_so[6] = \A_s[4] ;
  assign \A_s[4]  = A_s[4];
  assign A_so[5] = \A_s[3] ;
  assign \A_s[3]  = A_s[3];
  assign A_so[4] = \A_s[2] ;
  assign \A_s[2]  = A_s[2];
  assign A_so[3] = \A_s[1] ;
  assign \A_s[1]  = A_s[1];
  assign A_so[2] = \A_s[0] ;
  assign \A_s[0]  = A_s[0];
  assign A_nso[49] = \A_ns[47] ;
  assign \A_ns[47]  = A_ns[47];
  assign A_nso[48] = \A_ns[46] ;
  assign \A_ns[46]  = A_ns[46];
  assign A_nso[45] = \A_ns[43] ;
  assign \A_ns[43]  = A_ns[43];
  assign A_nso[44] = \A_ns[42] ;
  assign \A_ns[42]  = A_ns[42];
  assign A_nso[43] = \A_ns[41] ;
  assign \A_ns[41]  = A_ns[41];
  assign A_nso[16] = \A_ns[14] ;
  assign \A_ns[14]  = A_ns[14];
  assign A_nso[15] = \A_ns[13] ;
  assign \A_ns[13]  = A_ns[13];
  assign A_nso[14] = \A_ns[12] ;
  assign \A_ns[12]  = A_ns[12];
  assign A_nso[13] = \A_ns[11] ;
  assign \A_ns[11]  = A_ns[11];
  assign A_nso[12] = \A_ns[10] ;
  assign \A_ns[10]  = A_ns[10];
  assign A_nso[11] = \A_ns[9] ;
  assign \A_ns[9]  = A_ns[9];
  assign A_nso[10] = \A_ns[8] ;
  assign \A_ns[8]  = A_ns[8];
  assign A_nso[9] = \A_ns[7] ;
  assign \A_ns[7]  = A_ns[7];
  assign A_nso[8] = \A_ns[6] ;
  assign \A_ns[6]  = A_ns[6];
  assign A_nso[7] = \A_ns[5] ;
  assign \A_ns[5]  = A_ns[5];
  assign A_nso[6] = \A_ns[4] ;
  assign \A_ns[4]  = A_ns[4];
  assign A_nso[5] = \A_ns[3] ;
  assign \A_ns[3]  = A_ns[3];
  assign A_nso[4] = \A_ns[2] ;
  assign \A_ns[2]  = A_ns[2];
  assign A_nso[3] = \A_ns[1] ;
  assign \A_ns[1]  = A_ns[1];
  assign A_nso[2] = \A_ns[0] ;
  assign \A_ns[0]  = A_ns[0];

  XOR2_X1 U201 ( .A(B[15]), .B(B[16]), .Z(n152) );
  NAND3_X1 U202 ( .A1(B[16]), .A2(n804), .A3(B[15]), .ZN(n103) );
  OAI221_X1 U2 ( .B1(n659), .B2(n702), .C1(n654), .C2(n758), .A(n123), .ZN(
        O[37]) );
  CLKBUF_X1 U3 ( .A(n645), .Z(n648) );
  CLKBUF_X1 U4 ( .A(n639), .Z(n642) );
  CLKBUF_X1 U5 ( .A(n802), .Z(n640) );
  CLKBUF_X1 U6 ( .A(n803), .Z(n646) );
  CLKBUF_X1 U7 ( .A(n652), .Z(n655) );
  CLKBUF_X1 U8 ( .A(n662), .Z(n658) );
  CLKBUF_X1 U9 ( .A(n102), .Z(n661) );
  AOI22_X1 U10 ( .A1(A_ns[48]), .A2(n650), .B1(A_s[48]), .B2(n644), .ZN(n110)
         );
  BUF_X1 U11 ( .A(n645), .Z(n647) );
  BUF_X1 U12 ( .A(n639), .Z(n641) );
  BUF_X1 U13 ( .A(n646), .Z(n649) );
  BUF_X1 U14 ( .A(n640), .Z(n643) );
  AOI22_X1 U15 ( .A1(A_nso[42]), .A2(n649), .B1(\A_s[40] ), .B2(n643), .ZN(
        n118) );
  BUF_X1 U16 ( .A(n646), .Z(n650) );
  BUF_X1 U17 ( .A(n640), .Z(n644) );
  OAI221_X1 U18 ( .B1(n660), .B2(n721), .C1(n653), .C2(n771), .A(n110), .ZN(
        O[49]) );
  OAI221_X1 U19 ( .B1(n659), .B2(n712), .C1(n654), .C2(n763), .A(n117), .ZN(
        O[42]) );
  AOI22_X1 U20 ( .A1(\A_ns[41] ), .A2(n649), .B1(\A_s[41] ), .B2(n643), .ZN(
        n117) );
  OAI221_X1 U21 ( .B1(n660), .B2(n713), .C1(n654), .C2(n764), .A(n116), .ZN(
        O[43]) );
  AOI22_X1 U22 ( .A1(\A_ns[42] ), .A2(n649), .B1(\A_s[42] ), .B2(n643), .ZN(
        n116) );
  OAI221_X1 U23 ( .B1(n659), .B2(n710), .C1(n654), .C2(n762), .A(n118), .ZN(
        O[41]) );
  OAI221_X1 U24 ( .B1(n659), .B2(n714), .C1(n654), .C2(n765), .A(n115), .ZN(
        O[44]) );
  AOI22_X1 U25 ( .A1(\A_ns[43] ), .A2(n650), .B1(\A_s[43] ), .B2(n644), .ZN(
        n115) );
  AOI22_X1 U26 ( .A1(A_nso[38]), .A2(n649), .B1(\A_s[36] ), .B2(n643), .ZN(
        n123) );
  OAI221_X1 U27 ( .B1(n657), .B2(n666), .C1(n656), .C2(n729), .A(n142), .ZN(
        O[19]) );
  AOI22_X1 U28 ( .A1(A_nso[20]), .A2(n647), .B1(A_so[20]), .B2(n641), .ZN(n142) );
  OAI221_X1 U29 ( .B1(n657), .B2(n664), .C1(n656), .C2(n727), .A(n143), .ZN(
        O[18]) );
  AOI22_X1 U30 ( .A1(A_nso[19]), .A2(n647), .B1(A_so[19]), .B2(n641), .ZN(n143) );
  OAI221_X1 U31 ( .B1(n658), .B2(n678), .C1(n655), .C2(n741), .A(n136), .ZN(
        O[25]) );
  AOI22_X1 U32 ( .A1(A_nso[26]), .A2(n648), .B1(A_so[26]), .B2(n642), .ZN(n136) );
  OAI221_X1 U33 ( .B1(n658), .B2(n686), .C1(n655), .C2(n749), .A(n132), .ZN(
        O[29]) );
  AOI22_X1 U34 ( .A1(A_nso[30]), .A2(n648), .B1(\A_s[28] ), .B2(n642), .ZN(
        n132) );
  OAI221_X1 U35 ( .B1(n658), .B2(n690), .C1(n655), .C2(n751), .A(n129), .ZN(
        O[31]) );
  AOI22_X1 U36 ( .A1(A_nso[32]), .A2(n648), .B1(\A_s[30] ), .B2(n642), .ZN(
        n129) );
  OAI221_X1 U37 ( .B1(n659), .B2(n698), .C1(n654), .C2(n755), .A(n125), .ZN(
        O[35]) );
  AOI22_X1 U38 ( .A1(A_nso[36]), .A2(n649), .B1(A_so[36]), .B2(n643), .ZN(n125) );
  OAI221_X1 U39 ( .B1(n658), .B2(n680), .C1(n655), .C2(n743), .A(n135), .ZN(
        O[26]) );
  AOI22_X1 U40 ( .A1(A_nso[27]), .A2(n648), .B1(A_so[27]), .B2(n642), .ZN(n135) );
  OAI221_X1 U41 ( .B1(n658), .B2(n684), .C1(n655), .C2(n747), .A(n133), .ZN(
        O[28]) );
  AOI22_X1 U42 ( .A1(A_nso[29]), .A2(n648), .B1(A_so[29]), .B2(n642), .ZN(n133) );
  OAI221_X1 U43 ( .B1(n658), .B2(n672), .C1(n655), .C2(n735), .A(n139), .ZN(
        O[22]) );
  AOI22_X1 U44 ( .A1(A_nso[23]), .A2(n648), .B1(A_so[23]), .B2(n642), .ZN(n139) );
  OAI221_X1 U45 ( .B1(n658), .B2(n688), .C1(n655), .C2(n750), .A(n130), .ZN(
        O[30]) );
  AOI22_X1 U46 ( .A1(A_nso[31]), .A2(n648), .B1(\A_s[29] ), .B2(n642), .ZN(
        n130) );
  OAI221_X1 U47 ( .B1(n658), .B2(n692), .C1(n655), .C2(n752), .A(n128), .ZN(
        O[32]) );
  AOI22_X1 U48 ( .A1(A_nso[33]), .A2(n648), .B1(\A_s[31] ), .B2(n642), .ZN(
        n128) );
  OAI221_X1 U49 ( .B1(n659), .B2(n696), .C1(n654), .C2(n754), .A(n126), .ZN(
        O[34]) );
  AOI22_X1 U50 ( .A1(A_nso[35]), .A2(n649), .B1(\A_s[33] ), .B2(n643), .ZN(
        n126) );
  OAI221_X1 U51 ( .B1(n659), .B2(n700), .C1(n654), .C2(n757), .A(n124), .ZN(
        O[36]) );
  AOI22_X1 U52 ( .A1(A_nso[37]), .A2(n649), .B1(\A_s[35] ), .B2(n643), .ZN(
        n124) );
  OAI221_X1 U53 ( .B1(n659), .B2(n704), .C1(n654), .C2(n759), .A(n122), .ZN(
        O[38]) );
  AOI22_X1 U54 ( .A1(A_nso[39]), .A2(n649), .B1(\A_s[37] ), .B2(n643), .ZN(
        n122) );
  OAI221_X1 U55 ( .B1(n658), .B2(n676), .C1(n655), .C2(n739), .A(n137), .ZN(
        O[24]) );
  AOI22_X1 U56 ( .A1(A_nso[25]), .A2(n648), .B1(A_so[25]), .B2(n642), .ZN(n137) );
  OAI221_X1 U57 ( .B1(n658), .B2(n694), .C1(n655), .C2(n753), .A(n127), .ZN(
        O[33]) );
  AOI22_X1 U58 ( .A1(A_nso[34]), .A2(n649), .B1(\A_s[32] ), .B2(n643), .ZN(
        n127) );
  OAI221_X1 U59 ( .B1(n658), .B2(n682), .C1(n655), .C2(n745), .A(n134), .ZN(
        O[27]) );
  AOI22_X1 U60 ( .A1(A_nso[28]), .A2(n648), .B1(A_so[28]), .B2(n642), .ZN(n134) );
  OAI221_X1 U61 ( .B1(n657), .B2(n668), .C1(n656), .C2(n731), .A(n141), .ZN(
        O[20]) );
  AOI22_X1 U62 ( .A1(A_nso[21]), .A2(n647), .B1(A_so[21]), .B2(n641), .ZN(n141) );
  OAI221_X1 U63 ( .B1(n658), .B2(n674), .C1(n655), .C2(n737), .A(n138), .ZN(
        O[23]) );
  AOI22_X1 U64 ( .A1(A_nso[24]), .A2(n648), .B1(A_so[24]), .B2(n642), .ZN(n138) );
  OAI221_X1 U65 ( .B1(n657), .B2(n670), .C1(n655), .C2(n733), .A(n140), .ZN(
        O[21]) );
  AOI22_X1 U66 ( .A1(A_nso[22]), .A2(n647), .B1(A_so[22]), .B2(n641), .ZN(n140) );
  BUF_X1 U67 ( .A(n802), .Z(n639) );
  BUF_X1 U68 ( .A(n803), .Z(n645) );
  OAI221_X1 U69 ( .B1(n660), .B2(n715), .C1(n653), .C2(n766), .A(n114), .ZN(
        O[45]) );
  AOI22_X1 U70 ( .A1(A_nso[46]), .A2(n650), .B1(\A_s[44] ), .B2(n644), .ZN(
        n114) );
  OAI221_X1 U71 ( .B1(n659), .B2(n717), .C1(n653), .C2(n767), .A(n113), .ZN(
        O[46]) );
  AOI22_X1 U72 ( .A1(A_nso[47]), .A2(n650), .B1(A_so[47]), .B2(n644), .ZN(n113) );
  OAI221_X1 U73 ( .B1(n659), .B2(n706), .C1(n654), .C2(n760), .A(n121), .ZN(
        O[39]) );
  AOI22_X1 U74 ( .A1(A_nso[40]), .A2(n649), .B1(\A_s[38] ), .B2(n643), .ZN(
        n121) );
  OAI221_X1 U75 ( .B1(n660), .B2(n719), .C1(n653), .C2(n769), .A(n112), .ZN(
        O[47]) );
  AOI22_X1 U76 ( .A1(\A_ns[46] ), .A2(n650), .B1(\A_s[46] ), .B2(n644), .ZN(
        n112) );
  OAI221_X1 U77 ( .B1(n659), .B2(n708), .C1(n654), .C2(n761), .A(n119), .ZN(
        O[40]) );
  AOI22_X1 U78 ( .A1(A_nso[41]), .A2(n649), .B1(\A_s[39] ), .B2(n643), .ZN(
        n119) );
  OAI221_X1 U79 ( .B1(n660), .B2(n720), .C1(n653), .C2(n770), .A(n111), .ZN(
        O[48]) );
  AOI22_X1 U80 ( .A1(\A_ns[47] ), .A2(n650), .B1(\A_s[47] ), .B2(n644), .ZN(
        n111) );
  BUF_X1 U81 ( .A(n662), .Z(n657) );
  BUF_X1 U82 ( .A(n652), .Z(n656) );
  INV_X1 U83 ( .A(n100), .ZN(n802) );
  INV_X1 U84 ( .A(n101), .ZN(n803) );
  BUF_X1 U85 ( .A(n661), .Z(n659) );
  BUF_X1 U86 ( .A(n651), .Z(n654) );
  BUF_X1 U87 ( .A(n661), .Z(n660) );
  BUF_X1 U88 ( .A(n651), .Z(n653) );
  OAI221_X1 U89 ( .B1(n657), .B2(n723), .C1(n656), .C2(n725), .A(n144), .ZN(
        O[17]) );
  AOI22_X1 U90 ( .A1(A_nso[18]), .A2(n647), .B1(A_so[18]), .B2(n641), .ZN(n144) );
  NAND2_X1 U91 ( .A1(n152), .A2(n804), .ZN(n100) );
  NAND2_X1 U92 ( .A1(n152), .A2(n100), .ZN(n101) );
  BUF_X1 U93 ( .A(n103), .Z(n652) );
  BUF_X1 U94 ( .A(n102), .Z(n662) );
  CLKBUF_X1 U95 ( .A(n103), .Z(n651) );
  OAI221_X1 U96 ( .B1(n657), .B2(n800), .C1(n656), .C2(n801), .A(n145), .ZN(
        O[16]) );
  INV_X1 U97 ( .A(\A_ns[14] ), .ZN(n800) );
  INV_X1 U98 ( .A(\A_s[14] ), .ZN(n801) );
  AOI22_X1 U99 ( .A1(A_nso[17]), .A2(n647), .B1(A_so[17]), .B2(n641), .ZN(n145) );
  INV_X1 U100 ( .A(B[17]), .ZN(n804) );
  OR3_X1 U101 ( .A1(B[15]), .A2(B[16]), .A3(n804), .ZN(n102) );
  OAI221_X1 U102 ( .B1(n657), .B2(n797), .C1(n656), .C2(n799), .A(n146), .ZN(
        O[15]) );
  INV_X1 U103 ( .A(\A_ns[13] ), .ZN(n797) );
  OAI221_X1 U104 ( .B1(n660), .B2(n781), .C1(n653), .C2(n783), .A(n106), .ZN(
        O[7]) );
  INV_X1 U105 ( .A(\A_ns[5] ), .ZN(n781) );
  INV_X1 U106 ( .A(\A_s[5] ), .ZN(n783) );
  OAI221_X1 U107 ( .B1(n660), .B2(n784), .C1(n653), .C2(n786), .A(n105), .ZN(
        O[8]) );
  INV_X1 U108 ( .A(\A_ns[6] ), .ZN(n784) );
  INV_X1 U109 ( .A(\A_s[6] ), .ZN(n786) );
  OAI221_X1 U110 ( .B1(n657), .B2(n785), .C1(n654), .C2(n787), .A(n104), .ZN(
        O[9]) );
  INV_X1 U111 ( .A(\A_ns[7] ), .ZN(n785) );
  INV_X1 U112 ( .A(\A_s[7] ), .ZN(n787) );
  OAI221_X1 U113 ( .B1(n788), .B2(n660), .C1(n790), .C2(n653), .A(n151), .ZN(
        O[10]) );
  INV_X1 U114 ( .A(\A_s[8] ), .ZN(n790) );
  INV_X1 U115 ( .A(\A_ns[8] ), .ZN(n788) );
  OAI221_X1 U116 ( .B1(n657), .B2(n789), .C1(n653), .C2(n791), .A(n150), .ZN(
        O[11]) );
  INV_X1 U117 ( .A(\A_ns[9] ), .ZN(n789) );
  INV_X1 U118 ( .A(\A_s[9] ), .ZN(n791) );
  OAI221_X1 U119 ( .B1(n657), .B2(n792), .C1(n656), .C2(n794), .A(n149), .ZN(
        O[12]) );
  INV_X1 U120 ( .A(\A_ns[10] ), .ZN(n792) );
  INV_X1 U121 ( .A(\A_s[10] ), .ZN(n794) );
  OAI221_X1 U122 ( .B1(n657), .B2(n793), .C1(n656), .C2(n795), .A(n148), .ZN(
        O[13]) );
  INV_X1 U123 ( .A(\A_ns[11] ), .ZN(n793) );
  INV_X1 U124 ( .A(\A_s[11] ), .ZN(n795) );
  OAI221_X1 U125 ( .B1(n657), .B2(n796), .C1(n656), .C2(n798), .A(n147), .ZN(
        O[14]) );
  INV_X1 U126 ( .A(\A_ns[12] ), .ZN(n796) );
  OAI22_X1 U127 ( .A1(n100), .A2(n774), .B1(n101), .B2(n772), .ZN(O[1]) );
  OAI221_X1 U128 ( .B1(n772), .B2(n660), .C1(n774), .C2(n653), .A(n131), .ZN(
        O[2]) );
  AOI22_X1 U129 ( .A1(\A_ns[1] ), .A2(n648), .B1(\A_s[1] ), .B2(n642), .ZN(
        n131) );
  OAI221_X1 U130 ( .B1(n659), .B2(n773), .C1(n654), .C2(n775), .A(n120), .ZN(
        O[3]) );
  INV_X1 U131 ( .A(\A_ns[1] ), .ZN(n773) );
  INV_X1 U132 ( .A(\A_s[1] ), .ZN(n775) );
  OAI221_X1 U133 ( .B1(n660), .B2(n776), .C1(n653), .C2(n778), .A(n109), .ZN(
        O[4]) );
  INV_X1 U134 ( .A(\A_ns[2] ), .ZN(n776) );
  INV_X1 U135 ( .A(\A_s[2] ), .ZN(n778) );
  OAI221_X1 U136 ( .B1(n660), .B2(n777), .C1(n653), .C2(n779), .A(n108), .ZN(
        O[5]) );
  INV_X1 U137 ( .A(\A_ns[3] ), .ZN(n777) );
  INV_X1 U138 ( .A(\A_s[3] ), .ZN(n779) );
  OAI221_X1 U139 ( .B1(n660), .B2(n780), .C1(n653), .C2(n782), .A(n107), .ZN(
        O[6]) );
  INV_X1 U140 ( .A(\A_ns[4] ), .ZN(n780) );
  INV_X1 U141 ( .A(\A_s[4] ), .ZN(n782) );
  INV_X1 U142 ( .A(\A_ns[0] ), .ZN(n772) );
  INV_X1 U143 ( .A(\A_s[0] ), .ZN(n774) );
  AOI22_X1 U144 ( .A1(\A_ns[2] ), .A2(n649), .B1(\A_s[2] ), .B2(n643), .ZN(
        n120) );
  AOI22_X1 U145 ( .A1(\A_ns[3] ), .A2(n650), .B1(\A_s[3] ), .B2(n644), .ZN(
        n109) );
  AOI22_X1 U146 ( .A1(\A_ns[4] ), .A2(n650), .B1(\A_s[4] ), .B2(n644), .ZN(
        n108) );
  AOI22_X1 U147 ( .A1(\A_ns[5] ), .A2(n650), .B1(\A_s[5] ), .B2(n644), .ZN(
        n107) );
  AOI22_X1 U148 ( .A1(\A_ns[6] ), .A2(n650), .B1(\A_s[6] ), .B2(n644), .ZN(
        n106) );
  AOI22_X1 U149 ( .A1(\A_ns[7] ), .A2(n650), .B1(\A_s[7] ), .B2(n644), .ZN(
        n105) );
  AOI22_X1 U150 ( .A1(\A_ns[8] ), .A2(n650), .B1(\A_s[8] ), .B2(n644), .ZN(
        n104) );
  AOI22_X1 U151 ( .A1(\A_ns[9] ), .A2(n647), .B1(\A_s[9] ), .B2(n641), .ZN(
        n151) );
  AOI22_X1 U152 ( .A1(\A_ns[10] ), .A2(n647), .B1(\A_s[10] ), .B2(n641), .ZN(
        n150) );
  AOI22_X1 U153 ( .A1(\A_ns[11] ), .A2(n647), .B1(\A_s[11] ), .B2(n641), .ZN(
        n149) );
  AOI22_X1 U154 ( .A1(\A_ns[12] ), .A2(n647), .B1(\A_s[12] ), .B2(n641), .ZN(
        n148) );
  AOI22_X1 U155 ( .A1(\A_ns[13] ), .A2(n647), .B1(\A_s[13] ), .B2(n641), .ZN(
        n147) );
  AOI22_X1 U156 ( .A1(\A_ns[14] ), .A2(n647), .B1(\A_s[14] ), .B2(n641), .ZN(
        n146) );
  INV_X1 U157 ( .A(\A_s[12] ), .ZN(n798) );
  INV_X1 U158 ( .A(\A_s[13] ), .ZN(n799) );
  INV_X1 U159 ( .A(n664), .ZN(A_nso[18]) );
  INV_X1 U160 ( .A(A_ns[16]), .ZN(n664) );
  INV_X1 U161 ( .A(n666), .ZN(A_nso[19]) );
  INV_X1 U162 ( .A(A_ns[17]), .ZN(n666) );
  INV_X1 U163 ( .A(n668), .ZN(A_nso[20]) );
  INV_X1 U164 ( .A(A_ns[18]), .ZN(n668) );
  INV_X1 U165 ( .A(n670), .ZN(A_nso[21]) );
  INV_X1 U166 ( .A(A_ns[19]), .ZN(n670) );
  INV_X1 U167 ( .A(n672), .ZN(A_nso[22]) );
  INV_X1 U168 ( .A(A_ns[20]), .ZN(n672) );
  INV_X1 U169 ( .A(n674), .ZN(A_nso[23]) );
  INV_X1 U170 ( .A(A_ns[21]), .ZN(n674) );
  INV_X1 U171 ( .A(n676), .ZN(A_nso[24]) );
  INV_X1 U172 ( .A(A_ns[22]), .ZN(n676) );
  INV_X1 U173 ( .A(n678), .ZN(A_nso[25]) );
  INV_X1 U174 ( .A(A_ns[23]), .ZN(n678) );
  INV_X1 U175 ( .A(n680), .ZN(A_nso[26]) );
  INV_X1 U176 ( .A(A_ns[24]), .ZN(n680) );
  INV_X1 U177 ( .A(n682), .ZN(A_nso[27]) );
  INV_X1 U178 ( .A(A_ns[25]), .ZN(n682) );
  INV_X1 U179 ( .A(n684), .ZN(A_nso[28]) );
  INV_X1 U180 ( .A(A_ns[26]), .ZN(n684) );
  INV_X1 U181 ( .A(n686), .ZN(A_nso[29]) );
  INV_X1 U182 ( .A(A_ns[27]), .ZN(n686) );
  INV_X1 U183 ( .A(n688), .ZN(A_nso[30]) );
  INV_X1 U184 ( .A(A_ns[28]), .ZN(n688) );
  INV_X1 U185 ( .A(n690), .ZN(A_nso[31]) );
  INV_X1 U186 ( .A(A_ns[29]), .ZN(n690) );
  INV_X1 U187 ( .A(n692), .ZN(A_nso[32]) );
  INV_X1 U188 ( .A(A_ns[30]), .ZN(n692) );
  INV_X1 U189 ( .A(n694), .ZN(A_nso[33]) );
  INV_X1 U190 ( .A(A_ns[31]), .ZN(n694) );
  INV_X1 U191 ( .A(n696), .ZN(A_nso[34]) );
  INV_X1 U192 ( .A(A_ns[32]), .ZN(n696) );
  INV_X1 U193 ( .A(n698), .ZN(A_nso[35]) );
  INV_X1 U194 ( .A(A_ns[33]), .ZN(n698) );
  INV_X1 U195 ( .A(n700), .ZN(A_nso[36]) );
  INV_X1 U196 ( .A(A_ns[34]), .ZN(n700) );
  INV_X1 U197 ( .A(n702), .ZN(A_nso[37]) );
  INV_X1 U198 ( .A(A_ns[35]), .ZN(n702) );
  INV_X1 U199 ( .A(n704), .ZN(A_nso[38]) );
  INV_X1 U200 ( .A(A_ns[36]), .ZN(n704) );
  INV_X1 U203 ( .A(n706), .ZN(A_nso[39]) );
  INV_X1 U204 ( .A(A_ns[37]), .ZN(n706) );
  INV_X1 U205 ( .A(n708), .ZN(A_nso[40]) );
  INV_X1 U206 ( .A(A_ns[38]), .ZN(n708) );
  INV_X1 U207 ( .A(n710), .ZN(A_nso[41]) );
  INV_X1 U208 ( .A(A_ns[39]), .ZN(n710) );
  INV_X1 U209 ( .A(n712), .ZN(A_nso[42]) );
  INV_X1 U210 ( .A(A_ns[40]), .ZN(n712) );
  INV_X1 U211 ( .A(\A_ns[41] ), .ZN(n713) );
  INV_X1 U212 ( .A(\A_ns[42] ), .ZN(n714) );
  INV_X1 U213 ( .A(\A_ns[43] ), .ZN(n715) );
  INV_X1 U214 ( .A(n717), .ZN(A_nso[46]) );
  INV_X1 U215 ( .A(A_ns[44]), .ZN(n717) );
  INV_X1 U216 ( .A(n719), .ZN(A_nso[47]) );
  INV_X1 U217 ( .A(A_ns[45]), .ZN(n719) );
  INV_X1 U218 ( .A(\A_ns[46] ), .ZN(n720) );
  INV_X1 U219 ( .A(\A_ns[47] ), .ZN(n721) );
  INV_X1 U220 ( .A(n723), .ZN(A_nso[17]) );
  INV_X1 U221 ( .A(A_ns[15]), .ZN(n723) );
  INV_X1 U222 ( .A(n725), .ZN(A_so[17]) );
  INV_X1 U223 ( .A(A_s[15]), .ZN(n725) );
  INV_X1 U224 ( .A(n727), .ZN(A_so[18]) );
  INV_X1 U225 ( .A(A_s[16]), .ZN(n727) );
  INV_X1 U226 ( .A(n729), .ZN(A_so[19]) );
  INV_X1 U227 ( .A(A_s[17]), .ZN(n729) );
  INV_X1 U228 ( .A(n731), .ZN(A_so[20]) );
  INV_X1 U229 ( .A(A_s[18]), .ZN(n731) );
  INV_X1 U230 ( .A(n733), .ZN(A_so[21]) );
  INV_X1 U231 ( .A(A_s[19]), .ZN(n733) );
  INV_X1 U232 ( .A(n735), .ZN(A_so[22]) );
  INV_X1 U233 ( .A(A_s[20]), .ZN(n735) );
  INV_X1 U234 ( .A(n737), .ZN(A_so[23]) );
  INV_X1 U235 ( .A(A_s[21]), .ZN(n737) );
  INV_X1 U236 ( .A(n739), .ZN(A_so[24]) );
  INV_X1 U237 ( .A(A_s[22]), .ZN(n739) );
  INV_X1 U238 ( .A(n741), .ZN(A_so[25]) );
  INV_X1 U239 ( .A(A_s[23]), .ZN(n741) );
  INV_X1 U240 ( .A(n743), .ZN(A_so[26]) );
  INV_X1 U241 ( .A(A_s[24]), .ZN(n743) );
  INV_X1 U242 ( .A(n745), .ZN(A_so[27]) );
  INV_X1 U243 ( .A(A_s[25]), .ZN(n745) );
  INV_X1 U244 ( .A(n747), .ZN(A_so[28]) );
  INV_X1 U245 ( .A(A_s[26]), .ZN(n747) );
  INV_X1 U246 ( .A(n749), .ZN(A_so[29]) );
  INV_X1 U247 ( .A(A_s[27]), .ZN(n749) );
  INV_X1 U248 ( .A(\A_s[28] ), .ZN(n750) );
  INV_X1 U249 ( .A(\A_s[29] ), .ZN(n751) );
  INV_X1 U250 ( .A(\A_s[30] ), .ZN(n752) );
  INV_X1 U251 ( .A(\A_s[31] ), .ZN(n753) );
  INV_X1 U252 ( .A(\A_s[32] ), .ZN(n754) );
  INV_X1 U253 ( .A(\A_s[33] ), .ZN(n755) );
  INV_X1 U254 ( .A(n757), .ZN(A_so[36]) );
  INV_X1 U255 ( .A(A_s[34]), .ZN(n757) );
  INV_X1 U256 ( .A(\A_s[35] ), .ZN(n758) );
  INV_X1 U257 ( .A(\A_s[36] ), .ZN(n759) );
  INV_X1 U258 ( .A(\A_s[37] ), .ZN(n760) );
  INV_X1 U259 ( .A(\A_s[38] ), .ZN(n761) );
  INV_X1 U260 ( .A(\A_s[39] ), .ZN(n762) );
  INV_X1 U261 ( .A(\A_s[40] ), .ZN(n763) );
  INV_X1 U262 ( .A(\A_s[41] ), .ZN(n764) );
  INV_X1 U263 ( .A(\A_s[42] ), .ZN(n765) );
  INV_X1 U264 ( .A(\A_s[43] ), .ZN(n766) );
  INV_X1 U265 ( .A(\A_s[44] ), .ZN(n767) );
  INV_X1 U266 ( .A(n769), .ZN(A_so[47]) );
  INV_X1 U267 ( .A(A_s[45]), .ZN(n769) );
  INV_X1 U268 ( .A(\A_s[46] ), .ZN(n770) );
  INV_X1 U269 ( .A(\A_s[47] ), .ZN(n771) );
endmodule


module BOOTHENC_NBIT52_i18 ( A_s, A_ns, B, O, A_so, A_nso );
  input [51:0] A_s;
  input [51:0] A_ns;
  input [51:0] B;
  output [51:0] O;
  output [51:0] A_so;
  output [51:0] A_nso;
  wire   \A_s[49] , \A_s[48] , \A_s[47] , \A_s[46] , \A_s[45] , \A_s[44] ,
         \A_s[43] , \A_s[42] , \A_s[41] , \A_s[40] , \A_s[39] , \A_s[37] ,
         \A_s[36] , \A_s[35] , \A_s[34] , \A_s[33] , \A_s[32] , \A_s[31] ,
         \A_s[30] , \A_s[29] , \A_s[28] , \A_s[27] , \A_s[26] , \A_s[25] ,
         \A_s[24] , \A_s[23] , \A_s[22] , \A_s[21] , \A_s[20] , \A_s[19] ,
         \A_s[18] , \A_s[17] , \A_s[16] , \A_s[15] , \A_s[14] , \A_s[13] ,
         \A_s[12] , \A_s[11] , \A_s[10] , \A_s[9] , \A_s[8] , \A_s[7] ,
         \A_s[6] , \A_s[5] , \A_s[4] , \A_s[3] , \A_s[2] , \A_s[1] , \A_s[0] ,
         \A_ns[49] , \A_ns[48] , \A_ns[47] , \A_ns[46] , \A_ns[42] ,
         \A_ns[41] , \A_ns[40] , \A_ns[39] , \A_ns[38] , \A_ns[37] ,
         \A_ns[36] , \A_ns[35] , \A_ns[34] , \A_ns[33] , \A_ns[32] ,
         \A_ns[31] , \A_ns[30] , \A_ns[29] , \A_ns[28] , \A_ns[27] ,
         \A_ns[26] , \A_ns[25] , \A_ns[24] , \A_ns[23] , \A_ns[22] ,
         \A_ns[21] , \A_ns[20] , \A_ns[19] , \A_ns[18] , \A_ns[17] ,
         \A_ns[16] , \A_ns[15] , \A_ns[14] , \A_ns[13] , \A_ns[12] ,
         \A_ns[11] , \A_ns[10] , \A_ns[9] , \A_ns[8] , \A_ns[7] , \A_ns[6] ,
         \A_ns[5] , \A_ns[4] , \A_ns[3] , \A_ns[2] , \A_ns[1] , \A_ns[0] ,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n708, n710, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788;
  assign A_nso[0] = 1'b0;
  assign A_nso[1] = 1'b0;
  assign A_so[0] = 1'b0;
  assign A_so[1] = 1'b0;
  assign O[0] = 1'b0;
  assign A_so[51] = \A_s[49] ;
  assign \A_s[49]  = A_s[49];
  assign A_so[50] = \A_s[48] ;
  assign \A_s[48]  = A_s[48];
  assign A_so[49] = \A_s[47] ;
  assign \A_s[47]  = A_s[47];
  assign A_so[48] = \A_s[46] ;
  assign \A_s[46]  = A_s[46];
  assign A_so[47] = \A_s[45] ;
  assign \A_s[45]  = A_s[45];
  assign A_so[46] = \A_s[44] ;
  assign \A_s[44]  = A_s[44];
  assign A_so[45] = \A_s[43] ;
  assign \A_s[43]  = A_s[43];
  assign A_so[44] = \A_s[42] ;
  assign \A_s[42]  = A_s[42];
  assign A_so[43] = \A_s[41] ;
  assign \A_s[41]  = A_s[41];
  assign A_so[42] = \A_s[40] ;
  assign \A_s[40]  = A_s[40];
  assign A_so[41] = \A_s[39] ;
  assign \A_s[39]  = A_s[39];
  assign A_so[39] = \A_s[37] ;
  assign \A_s[37]  = A_s[37];
  assign A_so[38] = \A_s[36] ;
  assign \A_s[36]  = A_s[36];
  assign A_so[37] = \A_s[35] ;
  assign \A_s[35]  = A_s[35];
  assign A_so[36] = \A_s[34] ;
  assign \A_s[34]  = A_s[34];
  assign A_so[35] = \A_s[33] ;
  assign \A_s[33]  = A_s[33];
  assign A_so[34] = \A_s[32] ;
  assign \A_s[32]  = A_s[32];
  assign A_so[33] = \A_s[31] ;
  assign \A_s[31]  = A_s[31];
  assign A_so[32] = \A_s[30] ;
  assign \A_s[30]  = A_s[30];
  assign A_so[31] = \A_s[29] ;
  assign \A_s[29]  = A_s[29];
  assign A_so[30] = \A_s[28] ;
  assign \A_s[28]  = A_s[28];
  assign A_so[29] = \A_s[27] ;
  assign \A_s[27]  = A_s[27];
  assign A_so[28] = \A_s[26] ;
  assign \A_s[26]  = A_s[26];
  assign A_so[27] = \A_s[25] ;
  assign \A_s[25]  = A_s[25];
  assign A_so[26] = \A_s[24] ;
  assign \A_s[24]  = A_s[24];
  assign A_so[25] = \A_s[23] ;
  assign \A_s[23]  = A_s[23];
  assign A_so[24] = \A_s[22] ;
  assign \A_s[22]  = A_s[22];
  assign A_so[23] = \A_s[21] ;
  assign \A_s[21]  = A_s[21];
  assign A_so[22] = \A_s[20] ;
  assign \A_s[20]  = A_s[20];
  assign A_so[21] = \A_s[19] ;
  assign \A_s[19]  = A_s[19];
  assign A_so[20] = \A_s[18] ;
  assign \A_s[18]  = A_s[18];
  assign A_so[19] = \A_s[17] ;
  assign \A_s[17]  = A_s[17];
  assign A_so[18] = \A_s[16] ;
  assign \A_s[16]  = A_s[16];
  assign A_so[17] = \A_s[15] ;
  assign \A_s[15]  = A_s[15];
  assign A_so[16] = \A_s[14] ;
  assign \A_s[14]  = A_s[14];
  assign A_so[15] = \A_s[13] ;
  assign \A_s[13]  = A_s[13];
  assign A_so[14] = \A_s[12] ;
  assign \A_s[12]  = A_s[12];
  assign A_so[13] = \A_s[11] ;
  assign \A_s[11]  = A_s[11];
  assign A_so[12] = \A_s[10] ;
  assign \A_s[10]  = A_s[10];
  assign A_so[11] = \A_s[9] ;
  assign \A_s[9]  = A_s[9];
  assign A_so[10] = \A_s[8] ;
  assign \A_s[8]  = A_s[8];
  assign A_so[9] = \A_s[7] ;
  assign \A_s[7]  = A_s[7];
  assign A_so[8] = \A_s[6] ;
  assign \A_s[6]  = A_s[6];
  assign A_so[7] = \A_s[5] ;
  assign \A_s[5]  = A_s[5];
  assign A_so[6] = \A_s[4] ;
  assign \A_s[4]  = A_s[4];
  assign A_so[5] = \A_s[3] ;
  assign \A_s[3]  = A_s[3];
  assign A_so[4] = \A_s[2] ;
  assign \A_s[2]  = A_s[2];
  assign A_so[3] = \A_s[1] ;
  assign \A_s[1]  = A_s[1];
  assign A_so[2] = \A_s[0] ;
  assign \A_s[0]  = A_s[0];
  assign A_nso[51] = \A_ns[49] ;
  assign \A_ns[49]  = A_ns[49];
  assign A_nso[50] = \A_ns[48] ;
  assign \A_ns[48]  = A_ns[48];
  assign A_nso[49] = \A_ns[47] ;
  assign \A_ns[47]  = A_ns[47];
  assign A_nso[48] = \A_ns[46] ;
  assign \A_ns[46]  = A_ns[46];
  assign A_nso[44] = \A_ns[42] ;
  assign \A_ns[42]  = A_ns[42];
  assign A_nso[43] = \A_ns[41] ;
  assign \A_ns[41]  = A_ns[41];
  assign A_nso[42] = \A_ns[40] ;
  assign \A_ns[40]  = A_ns[40];
  assign A_nso[41] = \A_ns[39] ;
  assign \A_ns[39]  = A_ns[39];
  assign A_nso[40] = \A_ns[38] ;
  assign \A_ns[38]  = A_ns[38];
  assign A_nso[39] = \A_ns[37] ;
  assign \A_ns[37]  = A_ns[37];
  assign A_nso[38] = \A_ns[36] ;
  assign \A_ns[36]  = A_ns[36];
  assign A_nso[37] = \A_ns[35] ;
  assign \A_ns[35]  = A_ns[35];
  assign A_nso[36] = \A_ns[34] ;
  assign \A_ns[34]  = A_ns[34];
  assign A_nso[35] = \A_ns[33] ;
  assign \A_ns[33]  = A_ns[33];
  assign A_nso[34] = \A_ns[32] ;
  assign \A_ns[32]  = A_ns[32];
  assign A_nso[33] = \A_ns[31] ;
  assign \A_ns[31]  = A_ns[31];
  assign A_nso[32] = \A_ns[30] ;
  assign \A_ns[30]  = A_ns[30];
  assign A_nso[31] = \A_ns[29] ;
  assign \A_ns[29]  = A_ns[29];
  assign A_nso[30] = \A_ns[28] ;
  assign \A_ns[28]  = A_ns[28];
  assign A_nso[29] = \A_ns[27] ;
  assign \A_ns[27]  = A_ns[27];
  assign A_nso[28] = \A_ns[26] ;
  assign \A_ns[26]  = A_ns[26];
  assign A_nso[27] = \A_ns[25] ;
  assign \A_ns[25]  = A_ns[25];
  assign A_nso[26] = \A_ns[24] ;
  assign \A_ns[24]  = A_ns[24];
  assign A_nso[25] = \A_ns[23] ;
  assign \A_ns[23]  = A_ns[23];
  assign A_nso[24] = \A_ns[22] ;
  assign \A_ns[22]  = A_ns[22];
  assign A_nso[23] = \A_ns[21] ;
  assign \A_ns[21]  = A_ns[21];
  assign A_nso[22] = \A_ns[20] ;
  assign \A_ns[20]  = A_ns[20];
  assign A_nso[21] = \A_ns[19] ;
  assign \A_ns[19]  = A_ns[19];
  assign A_nso[20] = \A_ns[18] ;
  assign \A_ns[18]  = A_ns[18];
  assign A_nso[19] = \A_ns[17] ;
  assign \A_ns[17]  = A_ns[17];
  assign A_nso[18] = \A_ns[16] ;
  assign \A_ns[16]  = A_ns[16];
  assign A_nso[17] = \A_ns[15] ;
  assign \A_ns[15]  = A_ns[15];
  assign A_nso[16] = \A_ns[14] ;
  assign \A_ns[14]  = A_ns[14];
  assign A_nso[15] = \A_ns[13] ;
  assign \A_ns[13]  = A_ns[13];
  assign A_nso[14] = \A_ns[12] ;
  assign \A_ns[12]  = A_ns[12];
  assign A_nso[13] = \A_ns[11] ;
  assign \A_ns[11]  = A_ns[11];
  assign A_nso[12] = \A_ns[10] ;
  assign \A_ns[10]  = A_ns[10];
  assign A_nso[11] = \A_ns[9] ;
  assign \A_ns[9]  = A_ns[9];
  assign A_nso[10] = \A_ns[8] ;
  assign \A_ns[8]  = A_ns[8];
  assign A_nso[9] = \A_ns[7] ;
  assign \A_ns[7]  = A_ns[7];
  assign A_nso[8] = \A_ns[6] ;
  assign \A_ns[6]  = A_ns[6];
  assign A_nso[7] = \A_ns[5] ;
  assign \A_ns[5]  = A_ns[5];
  assign A_nso[6] = \A_ns[4] ;
  assign \A_ns[4]  = A_ns[4];
  assign A_nso[5] = \A_ns[3] ;
  assign \A_ns[3]  = A_ns[3];
  assign A_nso[4] = \A_ns[2] ;
  assign \A_ns[2]  = A_ns[2];
  assign A_nso[3] = \A_ns[1] ;
  assign \A_ns[1]  = A_ns[1];
  assign A_nso[2] = \A_ns[0] ;
  assign \A_ns[0]  = A_ns[0];

  OAI221_X2 U13 ( .B1(n678), .B2(n716), .C1(n671), .C2(n751), .A(n113), .ZN(
        O[51]) );
  XOR2_X1 U209 ( .A(B[17]), .B(B[18]), .Z(n158) );
  NAND3_X1 U210 ( .A1(B[18]), .A2(n788), .A3(B[17]), .ZN(n107) );
  OAI221_X1 U2 ( .B1(n677), .B2(n699), .C1(n672), .C2(n736), .A(n129), .ZN(
        O[37]) );
  AOI22_X1 U3 ( .A1(A_ns[50]), .A2(n667), .B1(A_s[50]), .B2(n660), .ZN(n113)
         );
  OAI221_X1 U4 ( .B1(n678), .B2(n715), .C1(n671), .C2(n750), .A(n114), .ZN(
        O[50]) );
  OAI221_X1 U5 ( .B1(n676), .B2(n686), .C1(n673), .C2(n723), .A(n143), .ZN(
        O[24]) );
  OAI221_X4 U6 ( .B1(n678), .B2(n714), .C1(n671), .C2(n749), .A(n116), .ZN(
        O[49]) );
  OAI221_X4 U7 ( .B1(n678), .B2(n713), .C1(n672), .C2(n748), .A(n117), .ZN(
        O[48]) );
  CLKBUF_X1 U8 ( .A(n662), .Z(n666) );
  CLKBUF_X1 U9 ( .A(n655), .Z(n659) );
  CLKBUF_X1 U10 ( .A(n662), .Z(n665) );
  CLKBUF_X1 U11 ( .A(n655), .Z(n658) );
  CLKBUF_X1 U12 ( .A(n786), .Z(n656) );
  CLKBUF_X1 U14 ( .A(n787), .Z(n663) );
  AOI22_X1 U15 ( .A1(\A_ns[47] ), .A2(n667), .B1(\A_s[47] ), .B2(n660), .ZN(
        n117) );
  BUF_X1 U16 ( .A(n662), .Z(n664) );
  BUF_X1 U17 ( .A(n655), .Z(n657) );
  BUF_X1 U18 ( .A(n663), .Z(n667) );
  BUF_X1 U19 ( .A(n656), .Z(n660) );
  BUF_X1 U20 ( .A(n663), .Z(n668) );
  BUF_X1 U21 ( .A(n656), .Z(n661) );
  AOI22_X1 U22 ( .A1(\A_ns[49] ), .A2(n667), .B1(\A_s[49] ), .B2(n660), .ZN(
        n114) );
  AOI22_X1 U23 ( .A1(\A_ns[36] ), .A2(n666), .B1(\A_s[36] ), .B2(n659), .ZN(
        n129) );
  AOI22_X1 U24 ( .A1(\A_ns[23] ), .A2(n665), .B1(\A_s[23] ), .B2(n658), .ZN(
        n143) );
  OAI221_X1 U25 ( .B1(n675), .B2(n682), .C1(n674), .C2(n719), .A(n147), .ZN(
        O[20]) );
  AOI22_X1 U26 ( .A1(\A_ns[19] ), .A2(n664), .B1(\A_s[19] ), .B2(n657), .ZN(
        n147) );
  OAI221_X1 U27 ( .B1(n676), .B2(n687), .C1(n673), .C2(n724), .A(n142), .ZN(
        O[25]) );
  AOI22_X1 U28 ( .A1(\A_ns[24] ), .A2(n665), .B1(\A_s[24] ), .B2(n658), .ZN(
        n142) );
  OAI221_X1 U29 ( .B1(n675), .B2(n683), .C1(n674), .C2(n720), .A(n146), .ZN(
        O[21]) );
  AOI22_X1 U30 ( .A1(\A_ns[20] ), .A2(n664), .B1(\A_s[20] ), .B2(n657), .ZN(
        n146) );
  OAI221_X1 U31 ( .B1(n676), .B2(n685), .C1(n673), .C2(n722), .A(n144), .ZN(
        O[23]) );
  AOI22_X1 U32 ( .A1(\A_ns[22] ), .A2(n665), .B1(\A_s[22] ), .B2(n658), .ZN(
        n144) );
  OAI221_X1 U33 ( .B1(n676), .B2(n689), .C1(n673), .C2(n726), .A(n140), .ZN(
        O[27]) );
  AOI22_X1 U34 ( .A1(\A_ns[26] ), .A2(n665), .B1(\A_s[26] ), .B2(n658), .ZN(
        n140) );
  OAI221_X1 U35 ( .B1(n676), .B2(n693), .C1(n673), .C2(n730), .A(n135), .ZN(
        O[31]) );
  AOI22_X1 U36 ( .A1(\A_ns[30] ), .A2(n665), .B1(\A_s[30] ), .B2(n658), .ZN(
        n135) );
  OAI221_X1 U37 ( .B1(n676), .B2(n695), .C1(n673), .C2(n732), .A(n133), .ZN(
        O[33]) );
  AOI22_X1 U38 ( .A1(\A_ns[32] ), .A2(n666), .B1(\A_s[32] ), .B2(n659), .ZN(
        n133) );
  OAI221_X1 U39 ( .B1(n677), .B2(n684), .C1(n674), .C2(n721), .A(n145), .ZN(
        O[22]) );
  AOI22_X1 U40 ( .A1(\A_ns[21] ), .A2(n665), .B1(\A_s[21] ), .B2(n658), .ZN(
        n145) );
  OAI221_X1 U41 ( .B1(n676), .B2(n692), .C1(n673), .C2(n729), .A(n136), .ZN(
        O[30]) );
  AOI22_X1 U42 ( .A1(\A_ns[29] ), .A2(n665), .B1(\A_s[29] ), .B2(n658), .ZN(
        n136) );
  OAI221_X1 U43 ( .B1(n676), .B2(n694), .C1(n673), .C2(n731), .A(n134), .ZN(
        O[32]) );
  AOI22_X1 U44 ( .A1(\A_ns[31] ), .A2(n665), .B1(\A_s[31] ), .B2(n658), .ZN(
        n134) );
  OAI221_X1 U45 ( .B1(n676), .B2(n696), .C1(n673), .C2(n733), .A(n132), .ZN(
        O[34]) );
  AOI22_X1 U46 ( .A1(\A_ns[33] ), .A2(n666), .B1(\A_s[33] ), .B2(n659), .ZN(
        n132) );
  OAI221_X1 U47 ( .B1(n677), .B2(n697), .C1(n672), .C2(n734), .A(n131), .ZN(
        O[35]) );
  AOI22_X1 U48 ( .A1(\A_ns[34] ), .A2(n666), .B1(\A_s[34] ), .B2(n659), .ZN(
        n131) );
  OAI221_X1 U49 ( .B1(n676), .B2(n688), .C1(n673), .C2(n725), .A(n141), .ZN(
        O[26]) );
  AOI22_X1 U50 ( .A1(\A_ns[25] ), .A2(n665), .B1(\A_s[25] ), .B2(n658), .ZN(
        n141) );
  OAI221_X1 U51 ( .B1(n675), .B2(n717), .C1(n674), .C2(n718), .A(n148), .ZN(
        O[19]) );
  AOI22_X1 U52 ( .A1(\A_ns[18] ), .A2(n664), .B1(\A_s[18] ), .B2(n657), .ZN(
        n148) );
  OAI221_X1 U53 ( .B1(n676), .B2(n690), .C1(n673), .C2(n727), .A(n139), .ZN(
        O[28]) );
  AOI22_X1 U54 ( .A1(\A_ns[27] ), .A2(n665), .B1(\A_s[27] ), .B2(n658), .ZN(
        n139) );
  OAI221_X1 U55 ( .B1(n676), .B2(n691), .C1(n673), .C2(n728), .A(n138), .ZN(
        O[29]) );
  AOI22_X1 U56 ( .A1(\A_ns[28] ), .A2(n665), .B1(\A_s[28] ), .B2(n658), .ZN(
        n138) );
  BUF_X1 U57 ( .A(n786), .Z(n655) );
  BUF_X1 U58 ( .A(n787), .Z(n662) );
  OAI221_X1 U59 ( .B1(n678), .B2(n708), .C1(n672), .C2(n745), .A(n120), .ZN(
        O[45]) );
  AOI22_X1 U60 ( .A1(A_nso[46]), .A2(n667), .B1(\A_s[44] ), .B2(n660), .ZN(
        n120) );
  OAI221_X1 U61 ( .B1(n677), .B2(n705), .C1(n672), .C2(n743), .A(n122), .ZN(
        O[43]) );
  AOI22_X1 U62 ( .A1(\A_ns[42] ), .A2(n666), .B1(\A_s[42] ), .B2(n659), .ZN(
        n122) );
  AOI22_X1 U63 ( .A1(\A_ns[48] ), .A2(n667), .B1(\A_s[48] ), .B2(n660), .ZN(
        n116) );
  OAI221_X1 U64 ( .B1(n677), .B2(n704), .C1(n672), .C2(n742), .A(n123), .ZN(
        O[42]) );
  AOI22_X1 U65 ( .A1(\A_ns[41] ), .A2(n666), .B1(\A_s[41] ), .B2(n659), .ZN(
        n123) );
  OAI221_X1 U66 ( .B1(n677), .B2(n701), .C1(n672), .C2(n738), .A(n127), .ZN(
        O[39]) );
  AOI22_X1 U67 ( .A1(\A_ns[38] ), .A2(n666), .B1(A_so[40]), .B2(n659), .ZN(
        n127) );
  OAI221_X1 U68 ( .B1(n677), .B2(n703), .C1(n672), .C2(n741), .A(n124), .ZN(
        O[41]) );
  AOI22_X1 U69 ( .A1(\A_ns[40] ), .A2(n666), .B1(\A_s[40] ), .B2(n659), .ZN(
        n124) );
  OAI221_X1 U70 ( .B1(n677), .B2(n698), .C1(n672), .C2(n735), .A(n130), .ZN(
        O[36]) );
  AOI22_X1 U71 ( .A1(\A_ns[35] ), .A2(n666), .B1(\A_s[35] ), .B2(n659), .ZN(
        n130) );
  OAI221_X1 U72 ( .B1(n677), .B2(n700), .C1(n672), .C2(n737), .A(n128), .ZN(
        O[38]) );
  AOI22_X1 U73 ( .A1(\A_ns[37] ), .A2(n666), .B1(\A_s[37] ), .B2(n659), .ZN(
        n128) );
  OAI221_X1 U74 ( .B1(n677), .B2(n702), .C1(n672), .C2(n740), .A(n125), .ZN(
        O[40]) );
  AOI22_X1 U75 ( .A1(\A_ns[39] ), .A2(n666), .B1(\A_s[39] ), .B2(n659), .ZN(
        n125) );
  OAI221_X1 U76 ( .B1(n678), .B2(n706), .C1(n672), .C2(n744), .A(n121), .ZN(
        O[44]) );
  AOI22_X1 U77 ( .A1(A_nso[45]), .A2(n667), .B1(\A_s[43] ), .B2(n660), .ZN(
        n121) );
  OAI221_X1 U78 ( .B1(n677), .B2(n710), .C1(n671), .C2(n746), .A(n119), .ZN(
        O[46]) );
  AOI22_X1 U79 ( .A1(A_nso[47]), .A2(n667), .B1(\A_s[45] ), .B2(n660), .ZN(
        n119) );
  OAI221_X1 U80 ( .B1(n678), .B2(n712), .C1(n671), .C2(n747), .A(n118), .ZN(
        O[47]) );
  AOI22_X1 U81 ( .A1(\A_ns[46] ), .A2(n667), .B1(\A_s[46] ), .B2(n660), .ZN(
        n118) );
  BUF_X1 U82 ( .A(n681), .Z(n676) );
  BUF_X1 U83 ( .A(n681), .Z(n675) );
  BUF_X1 U84 ( .A(n680), .Z(n677) );
  BUF_X1 U85 ( .A(n670), .Z(n673) );
  BUF_X1 U86 ( .A(n670), .Z(n674) );
  INV_X1 U87 ( .A(n104), .ZN(n786) );
  INV_X1 U88 ( .A(n105), .ZN(n787) );
  BUF_X1 U89 ( .A(n669), .Z(n672) );
  BUF_X1 U90 ( .A(n680), .Z(n678) );
  BUF_X1 U91 ( .A(n669), .Z(n671) );
  BUF_X1 U92 ( .A(n680), .Z(n679) );
  NAND2_X1 U93 ( .A1(n158), .A2(n788), .ZN(n104) );
  NAND2_X1 U94 ( .A1(n158), .A2(n104), .ZN(n105) );
  BUF_X1 U95 ( .A(n107), .Z(n670) );
  BUF_X1 U96 ( .A(n106), .Z(n680) );
  BUF_X1 U97 ( .A(n106), .Z(n681) );
  BUF_X1 U98 ( .A(n107), .Z(n669) );
  OAI221_X1 U99 ( .B1(n675), .B2(n784), .C1(n674), .C2(n785), .A(n149), .ZN(
        O[18]) );
  INV_X1 U100 ( .A(\A_ns[16] ), .ZN(n784) );
  INV_X1 U101 ( .A(\A_s[16] ), .ZN(n785) );
  AOI22_X1 U102 ( .A1(\A_ns[17] ), .A2(n664), .B1(\A_s[17] ), .B2(n657), .ZN(
        n149) );
  INV_X1 U103 ( .A(B[19]), .ZN(n788) );
  OR3_X1 U104 ( .A1(B[17]), .A2(B[18]), .A3(n788), .ZN(n106) );
  OAI221_X1 U105 ( .B1(n675), .B2(n780), .C1(n674), .C2(n782), .A(n151), .ZN(
        O[16]) );
  INV_X1 U106 ( .A(\A_ns[14] ), .ZN(n780) );
  OAI221_X1 U107 ( .B1(n675), .B2(n781), .C1(n674), .C2(n783), .A(n150), .ZN(
        O[17]) );
  INV_X1 U108 ( .A(\A_ns[15] ), .ZN(n781) );
  OAI221_X1 U109 ( .B1(n675), .B2(n777), .C1(n674), .C2(n779), .A(n152), .ZN(
        O[15]) );
  INV_X1 U110 ( .A(\A_ns[13] ), .ZN(n777) );
  INV_X1 U111 ( .A(\A_s[13] ), .ZN(n779) );
  OAI221_X1 U112 ( .B1(n678), .B2(n761), .C1(n671), .C2(n763), .A(n110), .ZN(
        O[7]) );
  INV_X1 U113 ( .A(\A_ns[5] ), .ZN(n761) );
  INV_X1 U114 ( .A(\A_s[5] ), .ZN(n763) );
  OAI221_X1 U115 ( .B1(n678), .B2(n764), .C1(n671), .C2(n766), .A(n109), .ZN(
        O[8]) );
  INV_X1 U116 ( .A(\A_ns[6] ), .ZN(n764) );
  INV_X1 U117 ( .A(\A_s[6] ), .ZN(n766) );
  OAI221_X1 U118 ( .B1(n675), .B2(n765), .C1(n673), .C2(n767), .A(n108), .ZN(
        O[9]) );
  INV_X1 U119 ( .A(\A_ns[7] ), .ZN(n765) );
  INV_X1 U120 ( .A(\A_s[7] ), .ZN(n767) );
  OAI221_X1 U121 ( .B1(n768), .B2(n679), .C1(n770), .C2(n671), .A(n157), .ZN(
        O[10]) );
  INV_X1 U122 ( .A(\A_s[8] ), .ZN(n770) );
  INV_X1 U123 ( .A(\A_ns[8] ), .ZN(n768) );
  OAI221_X1 U124 ( .B1(n675), .B2(n769), .C1(n671), .C2(n771), .A(n156), .ZN(
        O[11]) );
  INV_X1 U125 ( .A(\A_ns[9] ), .ZN(n769) );
  INV_X1 U126 ( .A(\A_s[9] ), .ZN(n771) );
  OAI221_X1 U127 ( .B1(n675), .B2(n772), .C1(n674), .C2(n774), .A(n155), .ZN(
        O[12]) );
  INV_X1 U128 ( .A(\A_ns[10] ), .ZN(n772) );
  INV_X1 U129 ( .A(\A_s[10] ), .ZN(n774) );
  OAI221_X1 U130 ( .B1(n675), .B2(n773), .C1(n674), .C2(n775), .A(n154), .ZN(
        O[13]) );
  INV_X1 U131 ( .A(\A_ns[11] ), .ZN(n773) );
  INV_X1 U132 ( .A(\A_s[11] ), .ZN(n775) );
  OAI221_X1 U133 ( .B1(n675), .B2(n776), .C1(n674), .C2(n778), .A(n153), .ZN(
        O[14]) );
  INV_X1 U134 ( .A(\A_ns[12] ), .ZN(n776) );
  INV_X1 U135 ( .A(\A_s[12] ), .ZN(n778) );
  OAI22_X1 U136 ( .A1(n104), .A2(n754), .B1(n105), .B2(n752), .ZN(O[1]) );
  OAI221_X1 U137 ( .B1(n752), .B2(n679), .C1(n754), .C2(n671), .A(n137), .ZN(
        O[2]) );
  AOI22_X1 U138 ( .A1(\A_ns[1] ), .A2(n665), .B1(\A_s[1] ), .B2(n658), .ZN(
        n137) );
  OAI221_X1 U139 ( .B1(n677), .B2(n753), .C1(n672), .C2(n755), .A(n126), .ZN(
        O[3]) );
  INV_X1 U140 ( .A(\A_ns[1] ), .ZN(n753) );
  INV_X1 U141 ( .A(\A_s[1] ), .ZN(n755) );
  OAI221_X1 U142 ( .B1(n678), .B2(n756), .C1(n671), .C2(n758), .A(n115), .ZN(
        O[4]) );
  INV_X1 U143 ( .A(\A_ns[2] ), .ZN(n756) );
  INV_X1 U144 ( .A(\A_s[2] ), .ZN(n758) );
  OAI221_X1 U145 ( .B1(n678), .B2(n757), .C1(n671), .C2(n759), .A(n112), .ZN(
        O[5]) );
  INV_X1 U146 ( .A(\A_ns[3] ), .ZN(n757) );
  INV_X1 U147 ( .A(\A_s[3] ), .ZN(n759) );
  OAI221_X1 U148 ( .B1(n678), .B2(n760), .C1(n671), .C2(n762), .A(n111), .ZN(
        O[6]) );
  INV_X1 U149 ( .A(\A_ns[4] ), .ZN(n760) );
  INV_X1 U150 ( .A(\A_s[4] ), .ZN(n762) );
  INV_X1 U151 ( .A(\A_ns[0] ), .ZN(n752) );
  INV_X1 U152 ( .A(\A_s[0] ), .ZN(n754) );
  AOI22_X1 U153 ( .A1(\A_ns[16] ), .A2(n664), .B1(\A_s[16] ), .B2(n657), .ZN(
        n150) );
  AOI22_X1 U154 ( .A1(\A_ns[2] ), .A2(n666), .B1(\A_s[2] ), .B2(n659), .ZN(
        n126) );
  AOI22_X1 U155 ( .A1(\A_ns[3] ), .A2(n667), .B1(\A_s[3] ), .B2(n660), .ZN(
        n115) );
  AOI22_X1 U156 ( .A1(\A_ns[4] ), .A2(n667), .B1(\A_s[4] ), .B2(n660), .ZN(
        n112) );
  AOI22_X1 U157 ( .A1(\A_ns[5] ), .A2(n667), .B1(\A_s[5] ), .B2(n660), .ZN(
        n111) );
  AOI22_X1 U158 ( .A1(\A_ns[6] ), .A2(n667), .B1(\A_s[6] ), .B2(n660), .ZN(
        n110) );
  AOI22_X1 U159 ( .A1(\A_ns[7] ), .A2(n668), .B1(\A_s[7] ), .B2(n661), .ZN(
        n109) );
  AOI22_X1 U160 ( .A1(\A_ns[8] ), .A2(n668), .B1(\A_s[8] ), .B2(n661), .ZN(
        n108) );
  AOI22_X1 U161 ( .A1(\A_ns[9] ), .A2(n664), .B1(\A_s[9] ), .B2(n657), .ZN(
        n157) );
  AOI22_X1 U162 ( .A1(\A_ns[10] ), .A2(n664), .B1(\A_s[10] ), .B2(n657), .ZN(
        n156) );
  AOI22_X1 U163 ( .A1(\A_ns[11] ), .A2(n664), .B1(\A_s[11] ), .B2(n657), .ZN(
        n155) );
  AOI22_X1 U164 ( .A1(\A_ns[12] ), .A2(n664), .B1(\A_s[12] ), .B2(n657), .ZN(
        n154) );
  AOI22_X1 U165 ( .A1(\A_ns[13] ), .A2(n664), .B1(\A_s[13] ), .B2(n657), .ZN(
        n153) );
  AOI22_X1 U166 ( .A1(\A_ns[14] ), .A2(n664), .B1(\A_s[14] ), .B2(n657), .ZN(
        n152) );
  AOI22_X1 U167 ( .A1(\A_ns[15] ), .A2(n664), .B1(\A_s[15] ), .B2(n657), .ZN(
        n151) );
  INV_X1 U168 ( .A(\A_s[15] ), .ZN(n783) );
  INV_X1 U169 ( .A(\A_s[14] ), .ZN(n782) );
  INV_X1 U170 ( .A(\A_ns[18] ), .ZN(n682) );
  INV_X1 U171 ( .A(\A_ns[19] ), .ZN(n683) );
  INV_X1 U172 ( .A(\A_ns[20] ), .ZN(n684) );
  INV_X1 U173 ( .A(\A_ns[21] ), .ZN(n685) );
  INV_X1 U174 ( .A(\A_ns[22] ), .ZN(n686) );
  INV_X1 U175 ( .A(\A_ns[23] ), .ZN(n687) );
  INV_X1 U176 ( .A(\A_ns[24] ), .ZN(n688) );
  INV_X1 U177 ( .A(\A_ns[25] ), .ZN(n689) );
  INV_X1 U178 ( .A(\A_ns[26] ), .ZN(n690) );
  INV_X1 U179 ( .A(\A_ns[27] ), .ZN(n691) );
  INV_X1 U180 ( .A(\A_ns[28] ), .ZN(n692) );
  INV_X1 U181 ( .A(\A_ns[29] ), .ZN(n693) );
  INV_X1 U182 ( .A(\A_ns[30] ), .ZN(n694) );
  INV_X1 U183 ( .A(\A_ns[31] ), .ZN(n695) );
  INV_X1 U184 ( .A(\A_ns[32] ), .ZN(n696) );
  INV_X1 U185 ( .A(\A_ns[33] ), .ZN(n697) );
  INV_X1 U186 ( .A(\A_ns[34] ), .ZN(n698) );
  INV_X1 U187 ( .A(\A_ns[35] ), .ZN(n699) );
  INV_X1 U188 ( .A(\A_ns[36] ), .ZN(n700) );
  INV_X1 U189 ( .A(\A_ns[37] ), .ZN(n701) );
  INV_X1 U190 ( .A(\A_ns[38] ), .ZN(n702) );
  INV_X1 U191 ( .A(\A_ns[39] ), .ZN(n703) );
  INV_X1 U192 ( .A(\A_ns[40] ), .ZN(n704) );
  INV_X1 U193 ( .A(\A_ns[41] ), .ZN(n705) );
  INV_X1 U194 ( .A(\A_ns[42] ), .ZN(n706) );
  INV_X1 U195 ( .A(n708), .ZN(A_nso[45]) );
  INV_X1 U196 ( .A(A_ns[43]), .ZN(n708) );
  INV_X1 U197 ( .A(n710), .ZN(A_nso[46]) );
  INV_X1 U198 ( .A(A_ns[44]), .ZN(n710) );
  INV_X1 U199 ( .A(n712), .ZN(A_nso[47]) );
  INV_X1 U200 ( .A(A_ns[45]), .ZN(n712) );
  INV_X1 U201 ( .A(\A_ns[46] ), .ZN(n713) );
  INV_X1 U202 ( .A(\A_ns[47] ), .ZN(n714) );
  INV_X1 U203 ( .A(\A_ns[48] ), .ZN(n715) );
  INV_X1 U204 ( .A(\A_ns[49] ), .ZN(n716) );
  INV_X1 U205 ( .A(\A_ns[17] ), .ZN(n717) );
  INV_X1 U206 ( .A(\A_s[17] ), .ZN(n718) );
  INV_X1 U207 ( .A(\A_s[18] ), .ZN(n719) );
  INV_X1 U208 ( .A(\A_s[19] ), .ZN(n720) );
  INV_X1 U211 ( .A(\A_s[20] ), .ZN(n721) );
  INV_X1 U212 ( .A(\A_s[21] ), .ZN(n722) );
  INV_X1 U213 ( .A(\A_s[22] ), .ZN(n723) );
  INV_X1 U214 ( .A(\A_s[23] ), .ZN(n724) );
  INV_X1 U215 ( .A(\A_s[24] ), .ZN(n725) );
  INV_X1 U216 ( .A(\A_s[25] ), .ZN(n726) );
  INV_X1 U217 ( .A(\A_s[26] ), .ZN(n727) );
  INV_X1 U218 ( .A(\A_s[27] ), .ZN(n728) );
  INV_X1 U219 ( .A(\A_s[28] ), .ZN(n729) );
  INV_X1 U220 ( .A(\A_s[29] ), .ZN(n730) );
  INV_X1 U221 ( .A(\A_s[30] ), .ZN(n731) );
  INV_X1 U222 ( .A(\A_s[31] ), .ZN(n732) );
  INV_X1 U223 ( .A(\A_s[32] ), .ZN(n733) );
  INV_X1 U224 ( .A(\A_s[33] ), .ZN(n734) );
  INV_X1 U225 ( .A(\A_s[34] ), .ZN(n735) );
  INV_X1 U226 ( .A(\A_s[35] ), .ZN(n736) );
  INV_X1 U227 ( .A(\A_s[36] ), .ZN(n737) );
  INV_X1 U228 ( .A(\A_s[37] ), .ZN(n738) );
  INV_X1 U229 ( .A(n740), .ZN(A_so[40]) );
  INV_X1 U230 ( .A(A_s[38]), .ZN(n740) );
  INV_X1 U231 ( .A(\A_s[39] ), .ZN(n741) );
  INV_X1 U232 ( .A(\A_s[40] ), .ZN(n742) );
  INV_X1 U233 ( .A(\A_s[41] ), .ZN(n743) );
  INV_X1 U234 ( .A(\A_s[42] ), .ZN(n744) );
  INV_X1 U235 ( .A(\A_s[43] ), .ZN(n745) );
  INV_X1 U236 ( .A(\A_s[44] ), .ZN(n746) );
  INV_X1 U237 ( .A(\A_s[45] ), .ZN(n747) );
  INV_X1 U238 ( .A(\A_s[46] ), .ZN(n748) );
  INV_X1 U239 ( .A(\A_s[47] ), .ZN(n749) );
  INV_X1 U240 ( .A(\A_s[48] ), .ZN(n750) );
  INV_X1 U241 ( .A(\A_s[49] ), .ZN(n751) );
endmodule


module BOOTHENC_NBIT54_i20 ( A_s, A_ns, B, O, A_so, A_nso );
  input [53:0] A_s;
  input [53:0] A_ns;
  input [53:0] B;
  output [53:0] O;
  output [53:0] A_so;
  output [53:0] A_nso;
  wire   \A_s[51] , \A_s[50] , \A_s[49] , \A_s[48] , \A_s[47] , \A_s[46] ,
         \A_s[45] , \A_s[44] , \A_s[43] , \A_s[42] , \A_s[41] , \A_s[40] ,
         \A_s[39] , \A_s[38] , \A_s[37] , \A_s[36] , \A_s[35] , \A_s[34] ,
         \A_s[33] , \A_s[32] , \A_s[31] , \A_s[30] , \A_s[29] , \A_s[28] ,
         \A_s[27] , \A_s[26] , \A_s[25] , \A_s[24] , \A_s[23] , \A_s[22] ,
         \A_s[21] , \A_s[20] , \A_s[19] , \A_s[18] , \A_s[17] , \A_s[16] ,
         \A_s[15] , \A_s[14] , \A_s[13] , \A_s[12] , \A_s[11] , \A_s[10] ,
         \A_s[9] , \A_s[8] , \A_s[7] , \A_s[6] , \A_s[5] , \A_s[4] , \A_s[3] ,
         \A_s[2] , \A_s[1] , \A_s[0] , \A_ns[51] , \A_ns[49] , \A_ns[48] ,
         \A_ns[47] , \A_ns[46] , \A_ns[45] , \A_ns[44] , \A_ns[43] ,
         \A_ns[42] , \A_ns[40] , \A_ns[38] , \A_ns[37] , \A_ns[36] ,
         \A_ns[35] , \A_ns[34] , \A_ns[33] , \A_ns[32] , \A_ns[31] ,
         \A_ns[30] , \A_ns[29] , \A_ns[28] , \A_ns[27] , \A_ns[26] ,
         \A_ns[25] , \A_ns[24] , \A_ns[23] , \A_ns[22] , \A_ns[21] ,
         \A_ns[20] , \A_ns[19] , \A_ns[18] , \A_ns[17] , \A_ns[16] ,
         \A_ns[15] , \A_ns[14] , \A_ns[13] , \A_ns[12] , \A_ns[11] ,
         \A_ns[10] , \A_ns[9] , \A_ns[8] , \A_ns[7] , \A_ns[6] , \A_ns[5] ,
         \A_ns[4] , \A_ns[3] , \A_ns[2] , \A_ns[1] , \A_ns[0] , n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n669, n670, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758;
  assign A_nso[0] = 1'b0;
  assign A_nso[1] = 1'b0;
  assign A_so[0] = 1'b0;
  assign A_so[1] = 1'b0;
  assign O[0] = 1'b0;
  assign A_so[53] = \A_s[51] ;
  assign \A_s[51]  = A_s[51];
  assign A_so[52] = \A_s[50] ;
  assign \A_s[50]  = A_s[50];
  assign A_so[51] = \A_s[49] ;
  assign \A_s[49]  = A_s[49];
  assign A_so[50] = \A_s[48] ;
  assign \A_s[48]  = A_s[48];
  assign A_so[49] = \A_s[47] ;
  assign \A_s[47]  = A_s[47];
  assign A_so[48] = \A_s[46] ;
  assign \A_s[46]  = A_s[46];
  assign A_so[47] = \A_s[45] ;
  assign \A_s[45]  = A_s[45];
  assign A_so[46] = \A_s[44] ;
  assign \A_s[44]  = A_s[44];
  assign A_so[45] = \A_s[43] ;
  assign \A_s[43]  = A_s[43];
  assign A_so[44] = \A_s[42] ;
  assign \A_s[42]  = A_s[42];
  assign A_so[43] = \A_s[41] ;
  assign \A_s[41]  = A_s[41];
  assign A_so[42] = \A_s[40] ;
  assign \A_s[40]  = A_s[40];
  assign A_so[41] = \A_s[39] ;
  assign \A_s[39]  = A_s[39];
  assign A_so[40] = \A_s[38] ;
  assign \A_s[38]  = A_s[38];
  assign A_so[39] = \A_s[37] ;
  assign \A_s[37]  = A_s[37];
  assign A_so[38] = \A_s[36] ;
  assign \A_s[36]  = A_s[36];
  assign A_so[37] = \A_s[35] ;
  assign \A_s[35]  = A_s[35];
  assign A_so[36] = \A_s[34] ;
  assign \A_s[34]  = A_s[34];
  assign A_so[35] = \A_s[33] ;
  assign \A_s[33]  = A_s[33];
  assign A_so[34] = \A_s[32] ;
  assign \A_s[32]  = A_s[32];
  assign A_so[33] = \A_s[31] ;
  assign \A_s[31]  = A_s[31];
  assign A_so[32] = \A_s[30] ;
  assign \A_s[30]  = A_s[30];
  assign A_so[31] = \A_s[29] ;
  assign \A_s[29]  = A_s[29];
  assign A_so[30] = \A_s[28] ;
  assign \A_s[28]  = A_s[28];
  assign A_so[29] = \A_s[27] ;
  assign \A_s[27]  = A_s[27];
  assign A_so[28] = \A_s[26] ;
  assign \A_s[26]  = A_s[26];
  assign A_so[27] = \A_s[25] ;
  assign \A_s[25]  = A_s[25];
  assign A_so[26] = \A_s[24] ;
  assign \A_s[24]  = A_s[24];
  assign A_so[25] = \A_s[23] ;
  assign \A_s[23]  = A_s[23];
  assign A_so[24] = \A_s[22] ;
  assign \A_s[22]  = A_s[22];
  assign A_so[23] = \A_s[21] ;
  assign \A_s[21]  = A_s[21];
  assign A_so[22] = \A_s[20] ;
  assign \A_s[20]  = A_s[20];
  assign A_so[21] = \A_s[19] ;
  assign \A_s[19]  = A_s[19];
  assign A_so[20] = \A_s[18] ;
  assign \A_s[18]  = A_s[18];
  assign A_so[19] = \A_s[17] ;
  assign \A_s[17]  = A_s[17];
  assign A_so[18] = \A_s[16] ;
  assign \A_s[16]  = A_s[16];
  assign A_so[17] = \A_s[15] ;
  assign \A_s[15]  = A_s[15];
  assign A_so[16] = \A_s[14] ;
  assign \A_s[14]  = A_s[14];
  assign A_so[15] = \A_s[13] ;
  assign \A_s[13]  = A_s[13];
  assign A_so[14] = \A_s[12] ;
  assign \A_s[12]  = A_s[12];
  assign A_so[13] = \A_s[11] ;
  assign \A_s[11]  = A_s[11];
  assign A_so[12] = \A_s[10] ;
  assign \A_s[10]  = A_s[10];
  assign A_so[11] = \A_s[9] ;
  assign \A_s[9]  = A_s[9];
  assign A_so[10] = \A_s[8] ;
  assign \A_s[8]  = A_s[8];
  assign A_so[9] = \A_s[7] ;
  assign \A_s[7]  = A_s[7];
  assign A_so[8] = \A_s[6] ;
  assign \A_s[6]  = A_s[6];
  assign A_so[7] = \A_s[5] ;
  assign \A_s[5]  = A_s[5];
  assign A_so[6] = \A_s[4] ;
  assign \A_s[4]  = A_s[4];
  assign A_so[5] = \A_s[3] ;
  assign \A_s[3]  = A_s[3];
  assign A_so[4] = \A_s[2] ;
  assign \A_s[2]  = A_s[2];
  assign A_so[3] = \A_s[1] ;
  assign \A_s[1]  = A_s[1];
  assign A_so[2] = \A_s[0] ;
  assign \A_s[0]  = A_s[0];
  assign A_nso[53] = \A_ns[51] ;
  assign \A_ns[51]  = A_ns[51];
  assign A_nso[51] = \A_ns[49] ;
  assign \A_ns[49]  = A_ns[49];
  assign A_nso[50] = \A_ns[48] ;
  assign \A_ns[48]  = A_ns[48];
  assign A_nso[49] = \A_ns[47] ;
  assign \A_ns[47]  = A_ns[47];
  assign A_nso[48] = \A_ns[46] ;
  assign \A_ns[46]  = A_ns[46];
  assign A_nso[47] = \A_ns[45] ;
  assign \A_ns[45]  = A_ns[45];
  assign A_nso[46] = \A_ns[44] ;
  assign \A_ns[44]  = A_ns[44];
  assign A_nso[45] = \A_ns[43] ;
  assign \A_ns[43]  = A_ns[43];
  assign A_nso[44] = \A_ns[42] ;
  assign \A_ns[42]  = A_ns[42];
  assign A_nso[42] = \A_ns[40] ;
  assign \A_ns[40]  = A_ns[40];
  assign A_nso[40] = \A_ns[38] ;
  assign \A_ns[38]  = A_ns[38];
  assign A_nso[39] = \A_ns[37] ;
  assign \A_ns[37]  = A_ns[37];
  assign A_nso[38] = \A_ns[36] ;
  assign \A_ns[36]  = A_ns[36];
  assign A_nso[37] = \A_ns[35] ;
  assign \A_ns[35]  = A_ns[35];
  assign A_nso[36] = \A_ns[34] ;
  assign \A_ns[34]  = A_ns[34];
  assign A_nso[35] = \A_ns[33] ;
  assign \A_ns[33]  = A_ns[33];
  assign A_nso[34] = \A_ns[32] ;
  assign \A_ns[32]  = A_ns[32];
  assign A_nso[33] = \A_ns[31] ;
  assign \A_ns[31]  = A_ns[31];
  assign A_nso[32] = \A_ns[30] ;
  assign \A_ns[30]  = A_ns[30];
  assign A_nso[31] = \A_ns[29] ;
  assign \A_ns[29]  = A_ns[29];
  assign A_nso[30] = \A_ns[28] ;
  assign \A_ns[28]  = A_ns[28];
  assign A_nso[29] = \A_ns[27] ;
  assign \A_ns[27]  = A_ns[27];
  assign A_nso[28] = \A_ns[26] ;
  assign \A_ns[26]  = A_ns[26];
  assign A_nso[27] = \A_ns[25] ;
  assign \A_ns[25]  = A_ns[25];
  assign A_nso[26] = \A_ns[24] ;
  assign \A_ns[24]  = A_ns[24];
  assign A_nso[25] = \A_ns[23] ;
  assign \A_ns[23]  = A_ns[23];
  assign A_nso[24] = \A_ns[22] ;
  assign \A_ns[22]  = A_ns[22];
  assign A_nso[23] = \A_ns[21] ;
  assign \A_ns[21]  = A_ns[21];
  assign A_nso[22] = \A_ns[20] ;
  assign \A_ns[20]  = A_ns[20];
  assign A_nso[21] = \A_ns[19] ;
  assign \A_ns[19]  = A_ns[19];
  assign A_nso[20] = \A_ns[18] ;
  assign \A_ns[18]  = A_ns[18];
  assign A_nso[19] = \A_ns[17] ;
  assign \A_ns[17]  = A_ns[17];
  assign A_nso[18] = \A_ns[16] ;
  assign \A_ns[16]  = A_ns[16];
  assign A_nso[17] = \A_ns[15] ;
  assign \A_ns[15]  = A_ns[15];
  assign A_nso[16] = \A_ns[14] ;
  assign \A_ns[14]  = A_ns[14];
  assign A_nso[15] = \A_ns[13] ;
  assign \A_ns[13]  = A_ns[13];
  assign A_nso[14] = \A_ns[12] ;
  assign \A_ns[12]  = A_ns[12];
  assign A_nso[13] = \A_ns[11] ;
  assign \A_ns[11]  = A_ns[11];
  assign A_nso[12] = \A_ns[10] ;
  assign \A_ns[10]  = A_ns[10];
  assign A_nso[11] = \A_ns[9] ;
  assign \A_ns[9]  = A_ns[9];
  assign A_nso[10] = \A_ns[8] ;
  assign \A_ns[8]  = A_ns[8];
  assign A_nso[9] = \A_ns[7] ;
  assign \A_ns[7]  = A_ns[7];
  assign A_nso[8] = \A_ns[6] ;
  assign \A_ns[6]  = A_ns[6];
  assign A_nso[7] = \A_ns[5] ;
  assign \A_ns[5]  = A_ns[5];
  assign A_nso[6] = \A_ns[4] ;
  assign \A_ns[4]  = A_ns[4];
  assign A_nso[5] = \A_ns[3] ;
  assign \A_ns[3]  = A_ns[3];
  assign A_nso[4] = \A_ns[2] ;
  assign \A_ns[2]  = A_ns[2];
  assign A_nso[3] = \A_ns[1] ;
  assign \A_ns[1]  = A_ns[1];
  assign A_nso[2] = \A_ns[0] ;
  assign \A_ns[0]  = A_ns[0];

  XOR2_X1 U217 ( .A(B[19]), .B(B[20]), .Z(n164) );
  NAND3_X1 U218 ( .A1(B[20]), .A2(n758), .A3(B[19]), .ZN(n111) );
  OAI221_X1 U2 ( .B1(n644), .B2(n672), .C1(n639), .C2(n707), .A(n128), .ZN(
        O[43]) );
  OAI221_X1 U3 ( .B1(n645), .B2(n675), .C1(n639), .C2(n710), .A(n125), .ZN(
        O[46]) );
  OAI221_X1 U4 ( .B1(n645), .B2(n678), .C1(n638), .C2(n713), .A(n122), .ZN(
        O[49]) );
  OAI221_X1 U5 ( .B1(n644), .B2(n662), .C1(n640), .C2(n699), .A(n137), .ZN(
        O[35]) );
  OAI221_X1 U6 ( .B1(n645), .B2(n682), .C1(n638), .C2(n716), .A(n118), .ZN(
        O[52]) );
  AOI22_X1 U7 ( .A1(\A_ns[45] ), .A2(n634), .B1(\A_s[45] ), .B2(n627), .ZN(
        n125) );
  BUF_X1 U8 ( .A(n629), .Z(n631) );
  BUF_X1 U9 ( .A(n629), .Z(n632) );
  BUF_X1 U10 ( .A(n622), .Z(n624) );
  BUF_X1 U11 ( .A(n622), .Z(n625) );
  BUF_X1 U12 ( .A(n629), .Z(n633) );
  BUF_X1 U13 ( .A(n622), .Z(n626) );
  BUF_X1 U14 ( .A(n630), .Z(n634) );
  BUF_X1 U15 ( .A(n623), .Z(n627) );
  BUF_X1 U16 ( .A(n630), .Z(n635) );
  BUF_X1 U17 ( .A(n623), .Z(n628) );
  OAI221_X1 U18 ( .B1(n645), .B2(n683), .C1(n638), .C2(n717), .A(n117), .ZN(
        O[53]) );
  AOI22_X1 U19 ( .A1(A_ns[52]), .A2(n634), .B1(A_s[52]), .B2(n627), .ZN(n117)
         );
  OAI221_X1 U20 ( .B1(n645), .B2(n679), .C1(n638), .C2(n714), .A(n120), .ZN(
        O[50]) );
  AOI22_X1 U21 ( .A1(\A_ns[49] ), .A2(n634), .B1(\A_s[49] ), .B2(n627), .ZN(
        n120) );
  OAI221_X1 U22 ( .B1(n645), .B2(n676), .C1(n639), .C2(n711), .A(n124), .ZN(
        O[47]) );
  AOI22_X1 U23 ( .A1(\A_ns[46] ), .A2(n634), .B1(\A_s[46] ), .B2(n627), .ZN(
        n124) );
  OAI221_X1 U24 ( .B1(n645), .B2(n677), .C1(n639), .C2(n712), .A(n123), .ZN(
        O[48]) );
  AOI22_X1 U25 ( .A1(\A_ns[47] ), .A2(n634), .B1(\A_s[47] ), .B2(n627), .ZN(
        n123) );
  AOI22_X1 U26 ( .A1(\A_ns[51] ), .A2(n634), .B1(\A_s[51] ), .B2(n627), .ZN(
        n118) );
  OAI221_X1 U27 ( .B1(n644), .B2(n649), .C1(n641), .C2(n686), .A(n151), .ZN(
        O[22]) );
  AOI22_X1 U28 ( .A1(\A_ns[21] ), .A2(n632), .B1(\A_s[21] ), .B2(n625), .ZN(
        n151) );
  OAI221_X1 U29 ( .B1(n643), .B2(n660), .C1(n640), .C2(n697), .A(n139), .ZN(
        O[33]) );
  AOI22_X1 U30 ( .A1(\A_ns[32] ), .A2(n633), .B1(\A_s[32] ), .B2(n626), .ZN(
        n139) );
  OAI221_X1 U31 ( .B1(n643), .B2(n650), .C1(n641), .C2(n687), .A(n150), .ZN(
        O[23]) );
  AOI22_X1 U32 ( .A1(\A_ns[22] ), .A2(n632), .B1(\A_s[22] ), .B2(n625), .ZN(
        n150) );
  OAI221_X1 U33 ( .B1(n642), .B2(n684), .C1(n641), .C2(n685), .A(n152), .ZN(
        O[21]) );
  AOI22_X1 U34 ( .A1(\A_ns[20] ), .A2(n631), .B1(\A_s[20] ), .B2(n624), .ZN(
        n152) );
  OAI221_X1 U35 ( .B1(n643), .B2(n651), .C1(n641), .C2(n688), .A(n149), .ZN(
        O[24]) );
  AOI22_X1 U36 ( .A1(\A_ns[23] ), .A2(n632), .B1(\A_s[23] ), .B2(n625), .ZN(
        n149) );
  OAI221_X1 U37 ( .B1(n643), .B2(n652), .C1(n640), .C2(n689), .A(n148), .ZN(
        O[25]) );
  AOI22_X1 U38 ( .A1(\A_ns[24] ), .A2(n632), .B1(\A_s[24] ), .B2(n625), .ZN(
        n148) );
  OAI221_X1 U39 ( .B1(n643), .B2(n653), .C1(n640), .C2(n690), .A(n147), .ZN(
        O[26]) );
  AOI22_X1 U40 ( .A1(\A_ns[25] ), .A2(n632), .B1(\A_s[25] ), .B2(n625), .ZN(
        n147) );
  OAI221_X1 U41 ( .B1(n643), .B2(n654), .C1(n640), .C2(n691), .A(n146), .ZN(
        O[27]) );
  AOI22_X1 U42 ( .A1(\A_ns[26] ), .A2(n632), .B1(\A_s[26] ), .B2(n625), .ZN(
        n146) );
  OAI221_X1 U43 ( .B1(n643), .B2(n657), .C1(n640), .C2(n694), .A(n142), .ZN(
        O[30]) );
  AOI22_X1 U44 ( .A1(\A_ns[29] ), .A2(n632), .B1(\A_s[29] ), .B2(n625), .ZN(
        n142) );
  OAI221_X1 U45 ( .B1(n643), .B2(n658), .C1(n640), .C2(n695), .A(n141), .ZN(
        O[31]) );
  AOI22_X1 U46 ( .A1(\A_ns[30] ), .A2(n632), .B1(\A_s[30] ), .B2(n625), .ZN(
        n141) );
  OAI221_X1 U47 ( .B1(n643), .B2(n659), .C1(n640), .C2(n696), .A(n140), .ZN(
        O[32]) );
  AOI22_X1 U48 ( .A1(\A_ns[31] ), .A2(n632), .B1(\A_s[31] ), .B2(n625), .ZN(
        n140) );
  OAI221_X1 U49 ( .B1(n643), .B2(n655), .C1(n640), .C2(n692), .A(n145), .ZN(
        O[28]) );
  AOI22_X1 U50 ( .A1(\A_ns[27] ), .A2(n632), .B1(\A_s[27] ), .B2(n625), .ZN(
        n145) );
  OAI221_X1 U51 ( .B1(n643), .B2(n656), .C1(n640), .C2(n693), .A(n144), .ZN(
        O[29]) );
  AOI22_X1 U52 ( .A1(\A_ns[28] ), .A2(n632), .B1(\A_s[28] ), .B2(n625), .ZN(
        n144) );
  AOI22_X1 U53 ( .A1(\A_ns[34] ), .A2(n633), .B1(\A_s[34] ), .B2(n626), .ZN(
        n137) );
  BUF_X1 U54 ( .A(n756), .Z(n622) );
  BUF_X1 U55 ( .A(n757), .Z(n629) );
  AOI22_X1 U56 ( .A1(\A_ns[42] ), .A2(n633), .B1(\A_s[42] ), .B2(n626), .ZN(
        n128) );
  OAI221_X1 U57 ( .B1(n643), .B2(n661), .C1(n640), .C2(n698), .A(n138), .ZN(
        O[34]) );
  AOI22_X1 U58 ( .A1(\A_ns[33] ), .A2(n633), .B1(\A_s[33] ), .B2(n626), .ZN(
        n138) );
  OAI221_X1 U59 ( .B1(n644), .B2(n663), .C1(n640), .C2(n700), .A(n136), .ZN(
        O[36]) );
  AOI22_X1 U60 ( .A1(\A_ns[35] ), .A2(n633), .B1(\A_s[35] ), .B2(n626), .ZN(
        n136) );
  OAI221_X1 U61 ( .B1(n644), .B2(n664), .C1(n639), .C2(n701), .A(n135), .ZN(
        O[37]) );
  AOI22_X1 U62 ( .A1(\A_ns[36] ), .A2(n633), .B1(\A_s[36] ), .B2(n626), .ZN(
        n135) );
  OAI221_X1 U63 ( .B1(n644), .B2(n665), .C1(n639), .C2(n702), .A(n134), .ZN(
        O[38]) );
  AOI22_X1 U64 ( .A1(\A_ns[37] ), .A2(n633), .B1(\A_s[37] ), .B2(n626), .ZN(
        n134) );
  OAI221_X1 U65 ( .B1(n644), .B2(n666), .C1(n639), .C2(n703), .A(n133), .ZN(
        O[39]) );
  AOI22_X1 U66 ( .A1(\A_ns[38] ), .A2(n633), .B1(\A_s[38] ), .B2(n626), .ZN(
        n133) );
  OAI221_X1 U67 ( .B1(n644), .B2(n667), .C1(n639), .C2(n704), .A(n131), .ZN(
        O[40]) );
  AOI22_X1 U68 ( .A1(A_nso[41]), .A2(n633), .B1(\A_s[39] ), .B2(n626), .ZN(
        n131) );
  OAI221_X1 U69 ( .B1(n644), .B2(n669), .C1(n639), .C2(n705), .A(n130), .ZN(
        O[41]) );
  AOI22_X1 U70 ( .A1(\A_ns[40] ), .A2(n633), .B1(\A_s[40] ), .B2(n626), .ZN(
        n130) );
  OAI221_X1 U71 ( .B1(n644), .B2(n670), .C1(n639), .C2(n706), .A(n129), .ZN(
        O[42]) );
  AOI22_X1 U72 ( .A1(A_nso[43]), .A2(n633), .B1(\A_s[41] ), .B2(n626), .ZN(
        n129) );
  OAI221_X1 U73 ( .B1(n644), .B2(n673), .C1(n639), .C2(n708), .A(n127), .ZN(
        O[44]) );
  AOI22_X1 U74 ( .A1(\A_ns[43] ), .A2(n634), .B1(\A_s[43] ), .B2(n627), .ZN(
        n127) );
  OAI221_X1 U75 ( .B1(n645), .B2(n674), .C1(n639), .C2(n709), .A(n126), .ZN(
        O[45]) );
  AOI22_X1 U76 ( .A1(\A_ns[44] ), .A2(n634), .B1(\A_s[44] ), .B2(n627), .ZN(
        n126) );
  OAI221_X1 U77 ( .B1(n645), .B2(n680), .C1(n638), .C2(n715), .A(n119), .ZN(
        O[51]) );
  AOI22_X1 U78 ( .A1(A_nso[52]), .A2(n634), .B1(\A_s[50] ), .B2(n627), .ZN(
        n119) );
  AOI22_X1 U79 ( .A1(\A_ns[48] ), .A2(n634), .B1(\A_s[48] ), .B2(n627), .ZN(
        n122) );
  BUF_X1 U80 ( .A(n756), .Z(n623) );
  BUF_X1 U81 ( .A(n757), .Z(n630) );
  BUF_X1 U82 ( .A(n648), .Z(n642) );
  BUF_X1 U83 ( .A(n648), .Z(n643) );
  BUF_X1 U84 ( .A(n647), .Z(n644) );
  BUF_X1 U85 ( .A(n637), .Z(n640) );
  BUF_X1 U86 ( .A(n637), .Z(n641) );
  INV_X1 U87 ( .A(n108), .ZN(n756) );
  INV_X1 U88 ( .A(n109), .ZN(n757) );
  BUF_X1 U89 ( .A(n636), .Z(n639) );
  BUF_X1 U90 ( .A(n647), .Z(n645) );
  BUF_X1 U91 ( .A(n636), .Z(n638) );
  BUF_X1 U92 ( .A(n647), .Z(n646) );
  NAND2_X1 U93 ( .A1(n164), .A2(n758), .ZN(n108) );
  NAND2_X1 U94 ( .A1(n164), .A2(n108), .ZN(n109) );
  BUF_X1 U95 ( .A(n111), .Z(n637) );
  BUF_X1 U96 ( .A(n110), .Z(n647) );
  BUF_X1 U97 ( .A(n110), .Z(n648) );
  BUF_X1 U98 ( .A(n111), .Z(n636) );
  OAI221_X1 U99 ( .B1(n642), .B2(n754), .C1(n641), .C2(n755), .A(n153), .ZN(
        O[20]) );
  INV_X1 U100 ( .A(\A_ns[18] ), .ZN(n754) );
  INV_X1 U101 ( .A(\A_s[18] ), .ZN(n755) );
  AOI22_X1 U102 ( .A1(\A_ns[19] ), .A2(n631), .B1(\A_s[19] ), .B2(n624), .ZN(
        n153) );
  INV_X1 U103 ( .A(B[21]), .ZN(n758) );
  OR3_X1 U104 ( .A1(B[19]), .A2(B[20]), .A3(n758), .ZN(n110) );
  OAI221_X1 U105 ( .B1(n642), .B2(n743), .C1(n641), .C2(n745), .A(n158), .ZN(
        O[15]) );
  INV_X1 U106 ( .A(\A_ns[13] ), .ZN(n743) );
  INV_X1 U107 ( .A(\A_s[13] ), .ZN(n745) );
  OAI221_X1 U108 ( .B1(n646), .B2(n727), .C1(n638), .C2(n729), .A(n114), .ZN(
        O[7]) );
  INV_X1 U109 ( .A(\A_ns[5] ), .ZN(n727) );
  INV_X1 U110 ( .A(\A_s[5] ), .ZN(n729) );
  OAI221_X1 U111 ( .B1(n645), .B2(n730), .C1(n638), .C2(n732), .A(n113), .ZN(
        O[8]) );
  INV_X1 U112 ( .A(\A_ns[6] ), .ZN(n730) );
  INV_X1 U113 ( .A(\A_s[6] ), .ZN(n732) );
  OAI221_X1 U114 ( .B1(n642), .B2(n731), .C1(n640), .C2(n733), .A(n112), .ZN(
        O[9]) );
  INV_X1 U115 ( .A(\A_ns[7] ), .ZN(n731) );
  INV_X1 U116 ( .A(\A_s[7] ), .ZN(n733) );
  OAI221_X1 U117 ( .B1(n734), .B2(n646), .C1(n736), .C2(n638), .A(n163), .ZN(
        O[10]) );
  INV_X1 U118 ( .A(\A_s[8] ), .ZN(n736) );
  INV_X1 U119 ( .A(\A_ns[8] ), .ZN(n734) );
  OAI221_X1 U120 ( .B1(n642), .B2(n735), .C1(n638), .C2(n737), .A(n162), .ZN(
        O[11]) );
  INV_X1 U121 ( .A(\A_ns[9] ), .ZN(n735) );
  INV_X1 U122 ( .A(\A_s[9] ), .ZN(n737) );
  OAI221_X1 U123 ( .B1(n642), .B2(n738), .C1(n641), .C2(n740), .A(n161), .ZN(
        O[12]) );
  INV_X1 U124 ( .A(\A_ns[10] ), .ZN(n738) );
  INV_X1 U125 ( .A(\A_s[10] ), .ZN(n740) );
  OAI221_X1 U126 ( .B1(n642), .B2(n739), .C1(n641), .C2(n741), .A(n160), .ZN(
        O[13]) );
  INV_X1 U127 ( .A(\A_ns[11] ), .ZN(n739) );
  INV_X1 U128 ( .A(\A_s[11] ), .ZN(n741) );
  OAI221_X1 U129 ( .B1(n642), .B2(n742), .C1(n641), .C2(n744), .A(n159), .ZN(
        O[14]) );
  INV_X1 U130 ( .A(\A_ns[12] ), .ZN(n742) );
  INV_X1 U131 ( .A(\A_s[12] ), .ZN(n744) );
  OAI22_X1 U132 ( .A1(n108), .A2(n720), .B1(n109), .B2(n718), .ZN(O[1]) );
  OAI221_X1 U133 ( .B1(n718), .B2(n646), .C1(n720), .C2(n638), .A(n143), .ZN(
        O[2]) );
  AOI22_X1 U134 ( .A1(\A_ns[1] ), .A2(n632), .B1(\A_s[1] ), .B2(n625), .ZN(
        n143) );
  OAI221_X1 U135 ( .B1(n644), .B2(n719), .C1(n639), .C2(n721), .A(n132), .ZN(
        O[3]) );
  INV_X1 U136 ( .A(\A_ns[1] ), .ZN(n719) );
  INV_X1 U137 ( .A(\A_s[1] ), .ZN(n721) );
  OAI221_X1 U138 ( .B1(n645), .B2(n722), .C1(n638), .C2(n724), .A(n121), .ZN(
        O[4]) );
  INV_X1 U139 ( .A(\A_ns[2] ), .ZN(n722) );
  INV_X1 U140 ( .A(\A_s[2] ), .ZN(n724) );
  OAI221_X1 U141 ( .B1(n646), .B2(n723), .C1(n638), .C2(n725), .A(n116), .ZN(
        O[5]) );
  INV_X1 U142 ( .A(\A_ns[3] ), .ZN(n723) );
  INV_X1 U143 ( .A(\A_s[3] ), .ZN(n725) );
  OAI221_X1 U144 ( .B1(n645), .B2(n726), .C1(n638), .C2(n728), .A(n115), .ZN(
        O[6]) );
  INV_X1 U145 ( .A(\A_ns[4] ), .ZN(n726) );
  INV_X1 U146 ( .A(\A_s[4] ), .ZN(n728) );
  OAI221_X1 U147 ( .B1(n642), .B2(n746), .C1(n641), .C2(n748), .A(n157), .ZN(
        O[16]) );
  INV_X1 U148 ( .A(\A_ns[14] ), .ZN(n746) );
  INV_X1 U149 ( .A(\A_s[14] ), .ZN(n748) );
  AOI22_X1 U150 ( .A1(\A_ns[15] ), .A2(n631), .B1(\A_s[15] ), .B2(n624), .ZN(
        n157) );
  OAI221_X1 U151 ( .B1(n642), .B2(n747), .C1(n641), .C2(n749), .A(n156), .ZN(
        O[17]) );
  INV_X1 U152 ( .A(\A_ns[15] ), .ZN(n747) );
  INV_X1 U153 ( .A(\A_s[15] ), .ZN(n749) );
  AOI22_X1 U154 ( .A1(\A_ns[16] ), .A2(n631), .B1(\A_s[16] ), .B2(n624), .ZN(
        n156) );
  OAI221_X1 U155 ( .B1(n642), .B2(n750), .C1(n641), .C2(n752), .A(n155), .ZN(
        O[18]) );
  INV_X1 U156 ( .A(\A_ns[16] ), .ZN(n750) );
  INV_X1 U157 ( .A(\A_s[16] ), .ZN(n752) );
  AOI22_X1 U158 ( .A1(\A_ns[17] ), .A2(n631), .B1(\A_s[17] ), .B2(n624), .ZN(
        n155) );
  OAI221_X1 U159 ( .B1(n642), .B2(n751), .C1(n641), .C2(n753), .A(n154), .ZN(
        O[19]) );
  INV_X1 U160 ( .A(\A_ns[17] ), .ZN(n751) );
  INV_X1 U161 ( .A(\A_s[17] ), .ZN(n753) );
  AOI22_X1 U162 ( .A1(\A_ns[18] ), .A2(n631), .B1(\A_s[18] ), .B2(n624), .ZN(
        n154) );
  INV_X1 U163 ( .A(\A_ns[0] ), .ZN(n718) );
  INV_X1 U164 ( .A(\A_s[0] ), .ZN(n720) );
  AOI22_X1 U165 ( .A1(\A_ns[2] ), .A2(n633), .B1(\A_s[2] ), .B2(n626), .ZN(
        n132) );
  AOI22_X1 U166 ( .A1(\A_ns[3] ), .A2(n634), .B1(\A_s[3] ), .B2(n627), .ZN(
        n121) );
  AOI22_X1 U167 ( .A1(\A_ns[4] ), .A2(n634), .B1(\A_s[4] ), .B2(n627), .ZN(
        n116) );
  AOI22_X1 U168 ( .A1(\A_ns[5] ), .A2(n635), .B1(\A_s[5] ), .B2(n628), .ZN(
        n115) );
  AOI22_X1 U169 ( .A1(\A_ns[6] ), .A2(n635), .B1(\A_s[6] ), .B2(n628), .ZN(
        n114) );
  AOI22_X1 U170 ( .A1(\A_ns[7] ), .A2(n635), .B1(\A_s[7] ), .B2(n628), .ZN(
        n113) );
  AOI22_X1 U171 ( .A1(\A_ns[8] ), .A2(n635), .B1(\A_s[8] ), .B2(n628), .ZN(
        n112) );
  AOI22_X1 U172 ( .A1(\A_ns[9] ), .A2(n631), .B1(\A_s[9] ), .B2(n624), .ZN(
        n163) );
  AOI22_X1 U173 ( .A1(\A_ns[10] ), .A2(n631), .B1(\A_s[10] ), .B2(n624), .ZN(
        n162) );
  AOI22_X1 U174 ( .A1(\A_ns[11] ), .A2(n631), .B1(\A_s[11] ), .B2(n624), .ZN(
        n161) );
  AOI22_X1 U175 ( .A1(\A_ns[12] ), .A2(n631), .B1(\A_s[12] ), .B2(n624), .ZN(
        n160) );
  AOI22_X1 U176 ( .A1(\A_ns[13] ), .A2(n631), .B1(\A_s[13] ), .B2(n624), .ZN(
        n159) );
  AOI22_X1 U177 ( .A1(\A_ns[14] ), .A2(n631), .B1(\A_s[14] ), .B2(n624), .ZN(
        n158) );
  INV_X1 U178 ( .A(\A_ns[20] ), .ZN(n649) );
  INV_X1 U179 ( .A(\A_ns[21] ), .ZN(n650) );
  INV_X1 U180 ( .A(\A_ns[22] ), .ZN(n651) );
  INV_X1 U181 ( .A(\A_ns[23] ), .ZN(n652) );
  INV_X1 U182 ( .A(\A_ns[24] ), .ZN(n653) );
  INV_X1 U183 ( .A(\A_ns[25] ), .ZN(n654) );
  INV_X1 U184 ( .A(\A_ns[26] ), .ZN(n655) );
  INV_X1 U185 ( .A(\A_ns[27] ), .ZN(n656) );
  INV_X1 U186 ( .A(\A_ns[28] ), .ZN(n657) );
  INV_X1 U187 ( .A(\A_ns[29] ), .ZN(n658) );
  INV_X1 U188 ( .A(\A_ns[30] ), .ZN(n659) );
  INV_X1 U189 ( .A(\A_ns[31] ), .ZN(n660) );
  INV_X1 U190 ( .A(\A_ns[32] ), .ZN(n661) );
  INV_X1 U191 ( .A(\A_ns[33] ), .ZN(n662) );
  INV_X1 U192 ( .A(\A_ns[34] ), .ZN(n663) );
  INV_X1 U193 ( .A(\A_ns[35] ), .ZN(n664) );
  INV_X1 U194 ( .A(\A_ns[36] ), .ZN(n665) );
  INV_X1 U195 ( .A(\A_ns[37] ), .ZN(n666) );
  INV_X1 U196 ( .A(\A_ns[38] ), .ZN(n667) );
  INV_X1 U197 ( .A(n669), .ZN(A_nso[41]) );
  INV_X1 U198 ( .A(A_ns[39]), .ZN(n669) );
  INV_X1 U199 ( .A(\A_ns[40] ), .ZN(n670) );
  INV_X1 U200 ( .A(n672), .ZN(A_nso[43]) );
  INV_X1 U201 ( .A(A_ns[41]), .ZN(n672) );
  INV_X1 U202 ( .A(\A_ns[42] ), .ZN(n673) );
  INV_X1 U203 ( .A(\A_ns[43] ), .ZN(n674) );
  INV_X1 U204 ( .A(\A_ns[44] ), .ZN(n675) );
  INV_X1 U205 ( .A(\A_ns[45] ), .ZN(n676) );
  INV_X1 U206 ( .A(\A_ns[46] ), .ZN(n677) );
  INV_X1 U207 ( .A(\A_ns[47] ), .ZN(n678) );
  INV_X1 U208 ( .A(\A_ns[48] ), .ZN(n679) );
  INV_X1 U209 ( .A(\A_ns[49] ), .ZN(n680) );
  INV_X1 U210 ( .A(n682), .ZN(A_nso[52]) );
  INV_X1 U211 ( .A(A_ns[50]), .ZN(n682) );
  INV_X1 U212 ( .A(\A_ns[51] ), .ZN(n683) );
  INV_X1 U213 ( .A(\A_ns[19] ), .ZN(n684) );
  INV_X1 U214 ( .A(\A_s[19] ), .ZN(n685) );
  INV_X1 U215 ( .A(\A_s[20] ), .ZN(n686) );
  INV_X1 U216 ( .A(\A_s[21] ), .ZN(n687) );
  INV_X1 U219 ( .A(\A_s[22] ), .ZN(n688) );
  INV_X1 U220 ( .A(\A_s[23] ), .ZN(n689) );
  INV_X1 U221 ( .A(\A_s[24] ), .ZN(n690) );
  INV_X1 U222 ( .A(\A_s[25] ), .ZN(n691) );
  INV_X1 U223 ( .A(\A_s[26] ), .ZN(n692) );
  INV_X1 U224 ( .A(\A_s[27] ), .ZN(n693) );
  INV_X1 U225 ( .A(\A_s[28] ), .ZN(n694) );
  INV_X1 U226 ( .A(\A_s[29] ), .ZN(n695) );
  INV_X1 U227 ( .A(\A_s[30] ), .ZN(n696) );
  INV_X1 U228 ( .A(\A_s[31] ), .ZN(n697) );
  INV_X1 U229 ( .A(\A_s[32] ), .ZN(n698) );
  INV_X1 U230 ( .A(\A_s[33] ), .ZN(n699) );
  INV_X1 U231 ( .A(\A_s[34] ), .ZN(n700) );
  INV_X1 U232 ( .A(\A_s[35] ), .ZN(n701) );
  INV_X1 U233 ( .A(\A_s[36] ), .ZN(n702) );
  INV_X1 U234 ( .A(\A_s[37] ), .ZN(n703) );
  INV_X1 U235 ( .A(\A_s[38] ), .ZN(n704) );
  INV_X1 U236 ( .A(\A_s[39] ), .ZN(n705) );
  INV_X1 U237 ( .A(\A_s[40] ), .ZN(n706) );
  INV_X1 U238 ( .A(\A_s[41] ), .ZN(n707) );
  INV_X1 U239 ( .A(\A_s[42] ), .ZN(n708) );
  INV_X1 U240 ( .A(\A_s[43] ), .ZN(n709) );
  INV_X1 U241 ( .A(\A_s[44] ), .ZN(n710) );
  INV_X1 U242 ( .A(\A_s[45] ), .ZN(n711) );
  INV_X1 U243 ( .A(\A_s[46] ), .ZN(n712) );
  INV_X1 U244 ( .A(\A_s[47] ), .ZN(n713) );
  INV_X1 U245 ( .A(\A_s[48] ), .ZN(n714) );
  INV_X1 U246 ( .A(\A_s[49] ), .ZN(n715) );
  INV_X1 U247 ( .A(\A_s[50] ), .ZN(n716) );
  INV_X1 U248 ( .A(\A_s[51] ), .ZN(n717) );
endmodule


module BOOTHENC_NBIT56_i22 ( A_s, A_ns, B, O, A_so, A_nso );
  input [55:0] A_s;
  input [55:0] A_ns;
  input [55:0] B;
  output [55:0] O;
  output [55:0] A_so;
  output [55:0] A_nso;
  wire   \A_s[53] , \A_s[52] , \A_s[51] , \A_s[50] , \A_s[49] , \A_s[48] ,
         \A_s[47] , \A_s[46] , \A_s[45] , \A_s[44] , \A_s[43] , \A_s[42] ,
         \A_s[41] , \A_s[40] , \A_s[39] , \A_s[38] , \A_s[37] , \A_s[36] ,
         \A_s[35] , \A_s[34] , \A_s[33] , \A_s[32] , \A_s[31] , \A_s[30] ,
         \A_s[29] , \A_s[28] , \A_s[27] , \A_s[26] , \A_s[25] , \A_s[24] ,
         \A_s[23] , \A_s[22] , \A_s[21] , \A_s[20] , \A_s[19] , \A_s[18] ,
         \A_s[17] , \A_s[16] , \A_s[15] , \A_s[14] , \A_s[13] , \A_s[12] ,
         \A_s[11] , \A_s[10] , \A_s[9] , \A_s[8] , \A_s[7] , \A_s[6] ,
         \A_s[5] , \A_s[4] , \A_s[3] , \A_s[2] , \A_s[1] , \A_s[0] ,
         \A_ns[52] , \A_ns[51] , \A_ns[50] , \A_ns[49] , \A_ns[48] ,
         \A_ns[43] , \A_ns[42] , \A_ns[41] , \A_ns[40] , \A_ns[37] ,
         \A_ns[36] , \A_ns[35] , \A_ns[34] , \A_ns[33] , \A_ns[32] ,
         \A_ns[31] , \A_ns[30] , \A_ns[29] , \A_ns[28] , \A_ns[27] ,
         \A_ns[26] , \A_ns[25] , \A_ns[24] , \A_ns[23] , \A_ns[22] ,
         \A_ns[21] , \A_ns[20] , \A_ns[19] , \A_ns[18] , \A_ns[17] ,
         \A_ns[16] , \A_ns[15] , \A_ns[14] , \A_ns[13] , \A_ns[12] ,
         \A_ns[11] , \A_ns[10] , \A_ns[9] , \A_ns[8] , \A_ns[7] , \A_ns[6] ,
         \A_ns[5] , \A_ns[4] , \A_ns[3] , \A_ns[2] , \A_ns[1] , \A_ns[0] ,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n681, n683, n684, n685, n686, n687, n689,
         n691, n693, n695, n696, n697, n698, n699, n700, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781;
  assign A_nso[0] = 1'b0;
  assign A_nso[1] = 1'b0;
  assign A_so[0] = 1'b0;
  assign A_so[1] = 1'b0;
  assign O[0] = 1'b0;
  assign A_so[55] = \A_s[53] ;
  assign \A_s[53]  = A_s[53];
  assign A_so[54] = \A_s[52] ;
  assign \A_s[52]  = A_s[52];
  assign A_so[53] = \A_s[51] ;
  assign \A_s[51]  = A_s[51];
  assign A_so[52] = \A_s[50] ;
  assign \A_s[50]  = A_s[50];
  assign A_so[51] = \A_s[49] ;
  assign \A_s[49]  = A_s[49];
  assign A_so[50] = \A_s[48] ;
  assign \A_s[48]  = A_s[48];
  assign A_so[49] = \A_s[47] ;
  assign \A_s[47]  = A_s[47];
  assign A_so[48] = \A_s[46] ;
  assign \A_s[46]  = A_s[46];
  assign A_so[47] = \A_s[45] ;
  assign \A_s[45]  = A_s[45];
  assign A_so[46] = \A_s[44] ;
  assign \A_s[44]  = A_s[44];
  assign A_so[45] = \A_s[43] ;
  assign \A_s[43]  = A_s[43];
  assign A_so[44] = \A_s[42] ;
  assign \A_s[42]  = A_s[42];
  assign A_so[43] = \A_s[41] ;
  assign \A_s[41]  = A_s[41];
  assign A_so[42] = \A_s[40] ;
  assign \A_s[40]  = A_s[40];
  assign A_so[41] = \A_s[39] ;
  assign \A_s[39]  = A_s[39];
  assign A_so[40] = \A_s[38] ;
  assign \A_s[38]  = A_s[38];
  assign A_so[39] = \A_s[37] ;
  assign \A_s[37]  = A_s[37];
  assign A_so[38] = \A_s[36] ;
  assign \A_s[36]  = A_s[36];
  assign A_so[37] = \A_s[35] ;
  assign \A_s[35]  = A_s[35];
  assign A_so[36] = \A_s[34] ;
  assign \A_s[34]  = A_s[34];
  assign A_so[35] = \A_s[33] ;
  assign \A_s[33]  = A_s[33];
  assign A_so[34] = \A_s[32] ;
  assign \A_s[32]  = A_s[32];
  assign A_so[33] = \A_s[31] ;
  assign \A_s[31]  = A_s[31];
  assign A_so[32] = \A_s[30] ;
  assign \A_s[30]  = A_s[30];
  assign A_so[31] = \A_s[29] ;
  assign \A_s[29]  = A_s[29];
  assign A_so[30] = \A_s[28] ;
  assign \A_s[28]  = A_s[28];
  assign A_so[29] = \A_s[27] ;
  assign \A_s[27]  = A_s[27];
  assign A_so[28] = \A_s[26] ;
  assign \A_s[26]  = A_s[26];
  assign A_so[27] = \A_s[25] ;
  assign \A_s[25]  = A_s[25];
  assign A_so[26] = \A_s[24] ;
  assign \A_s[24]  = A_s[24];
  assign A_so[25] = \A_s[23] ;
  assign \A_s[23]  = A_s[23];
  assign A_so[24] = \A_s[22] ;
  assign \A_s[22]  = A_s[22];
  assign A_so[23] = \A_s[21] ;
  assign \A_s[21]  = A_s[21];
  assign A_so[22] = \A_s[20] ;
  assign \A_s[20]  = A_s[20];
  assign A_so[21] = \A_s[19] ;
  assign \A_s[19]  = A_s[19];
  assign A_so[20] = \A_s[18] ;
  assign \A_s[18]  = A_s[18];
  assign A_so[19] = \A_s[17] ;
  assign \A_s[17]  = A_s[17];
  assign A_so[18] = \A_s[16] ;
  assign \A_s[16]  = A_s[16];
  assign A_so[17] = \A_s[15] ;
  assign \A_s[15]  = A_s[15];
  assign A_so[16] = \A_s[14] ;
  assign \A_s[14]  = A_s[14];
  assign A_so[15] = \A_s[13] ;
  assign \A_s[13]  = A_s[13];
  assign A_so[14] = \A_s[12] ;
  assign \A_s[12]  = A_s[12];
  assign A_so[13] = \A_s[11] ;
  assign \A_s[11]  = A_s[11];
  assign A_so[12] = \A_s[10] ;
  assign \A_s[10]  = A_s[10];
  assign A_so[11] = \A_s[9] ;
  assign \A_s[9]  = A_s[9];
  assign A_so[10] = \A_s[8] ;
  assign \A_s[8]  = A_s[8];
  assign A_so[9] = \A_s[7] ;
  assign \A_s[7]  = A_s[7];
  assign A_so[8] = \A_s[6] ;
  assign \A_s[6]  = A_s[6];
  assign A_so[7] = \A_s[5] ;
  assign \A_s[5]  = A_s[5];
  assign A_so[6] = \A_s[4] ;
  assign \A_s[4]  = A_s[4];
  assign A_so[5] = \A_s[3] ;
  assign \A_s[3]  = A_s[3];
  assign A_so[4] = \A_s[2] ;
  assign \A_s[2]  = A_s[2];
  assign A_so[3] = \A_s[1] ;
  assign \A_s[1]  = A_s[1];
  assign A_so[2] = \A_s[0] ;
  assign \A_s[0]  = A_s[0];
  assign A_nso[54] = \A_ns[52] ;
  assign \A_ns[52]  = A_ns[52];
  assign A_nso[53] = \A_ns[51] ;
  assign \A_ns[51]  = A_ns[51];
  assign A_nso[52] = \A_ns[50] ;
  assign \A_ns[50]  = A_ns[50];
  assign A_nso[51] = \A_ns[49] ;
  assign \A_ns[49]  = A_ns[49];
  assign A_nso[50] = \A_ns[48] ;
  assign \A_ns[48]  = A_ns[48];
  assign A_nso[45] = \A_ns[43] ;
  assign \A_ns[43]  = A_ns[43];
  assign A_nso[44] = \A_ns[42] ;
  assign \A_ns[42]  = A_ns[42];
  assign A_nso[43] = \A_ns[41] ;
  assign \A_ns[41]  = A_ns[41];
  assign A_nso[42] = \A_ns[40] ;
  assign \A_ns[40]  = A_ns[40];
  assign A_nso[39] = \A_ns[37] ;
  assign \A_ns[37]  = A_ns[37];
  assign A_nso[38] = \A_ns[36] ;
  assign \A_ns[36]  = A_ns[36];
  assign A_nso[37] = \A_ns[35] ;
  assign \A_ns[35]  = A_ns[35];
  assign A_nso[36] = \A_ns[34] ;
  assign \A_ns[34]  = A_ns[34];
  assign A_nso[35] = \A_ns[33] ;
  assign \A_ns[33]  = A_ns[33];
  assign A_nso[34] = \A_ns[32] ;
  assign \A_ns[32]  = A_ns[32];
  assign A_nso[33] = \A_ns[31] ;
  assign \A_ns[31]  = A_ns[31];
  assign A_nso[32] = \A_ns[30] ;
  assign \A_ns[30]  = A_ns[30];
  assign A_nso[31] = \A_ns[29] ;
  assign \A_ns[29]  = A_ns[29];
  assign A_nso[30] = \A_ns[28] ;
  assign \A_ns[28]  = A_ns[28];
  assign A_nso[29] = \A_ns[27] ;
  assign \A_ns[27]  = A_ns[27];
  assign A_nso[28] = \A_ns[26] ;
  assign \A_ns[26]  = A_ns[26];
  assign A_nso[27] = \A_ns[25] ;
  assign \A_ns[25]  = A_ns[25];
  assign A_nso[26] = \A_ns[24] ;
  assign \A_ns[24]  = A_ns[24];
  assign A_nso[25] = \A_ns[23] ;
  assign \A_ns[23]  = A_ns[23];
  assign A_nso[24] = \A_ns[22] ;
  assign \A_ns[22]  = A_ns[22];
  assign A_nso[23] = \A_ns[21] ;
  assign \A_ns[21]  = A_ns[21];
  assign A_nso[22] = \A_ns[20] ;
  assign \A_ns[20]  = A_ns[20];
  assign A_nso[21] = \A_ns[19] ;
  assign \A_ns[19]  = A_ns[19];
  assign A_nso[20] = \A_ns[18] ;
  assign \A_ns[18]  = A_ns[18];
  assign A_nso[19] = \A_ns[17] ;
  assign \A_ns[17]  = A_ns[17];
  assign A_nso[18] = \A_ns[16] ;
  assign \A_ns[16]  = A_ns[16];
  assign A_nso[17] = \A_ns[15] ;
  assign \A_ns[15]  = A_ns[15];
  assign A_nso[16] = \A_ns[14] ;
  assign \A_ns[14]  = A_ns[14];
  assign A_nso[15] = \A_ns[13] ;
  assign \A_ns[13]  = A_ns[13];
  assign A_nso[14] = \A_ns[12] ;
  assign \A_ns[12]  = A_ns[12];
  assign A_nso[13] = \A_ns[11] ;
  assign \A_ns[11]  = A_ns[11];
  assign A_nso[12] = \A_ns[10] ;
  assign \A_ns[10]  = A_ns[10];
  assign A_nso[11] = \A_ns[9] ;
  assign \A_ns[9]  = A_ns[9];
  assign A_nso[10] = \A_ns[8] ;
  assign \A_ns[8]  = A_ns[8];
  assign A_nso[9] = \A_ns[7] ;
  assign \A_ns[7]  = A_ns[7];
  assign A_nso[8] = \A_ns[6] ;
  assign \A_ns[6]  = A_ns[6];
  assign A_nso[7] = \A_ns[5] ;
  assign \A_ns[5]  = A_ns[5];
  assign A_nso[6] = \A_ns[4] ;
  assign \A_ns[4]  = A_ns[4];
  assign A_nso[5] = \A_ns[3] ;
  assign \A_ns[3]  = A_ns[3];
  assign A_nso[4] = \A_ns[2] ;
  assign \A_ns[2]  = A_ns[2];
  assign A_nso[3] = \A_ns[1] ;
  assign \A_ns[1]  = A_ns[1];
  assign A_nso[2] = \A_ns[0] ;
  assign \A_ns[0]  = A_ns[0];

  XOR2_X1 U225 ( .A(B[21]), .B(B[22]), .Z(n170) );
  NAND3_X1 U226 ( .A1(B[22]), .A2(n781), .A3(B[21]), .ZN(n115) );
  OAI221_X1 U2 ( .B1(n658), .B2(n665), .C1(n655), .C2(n706), .A(n154), .ZN(
        O[25]) );
  OAI221_X1 U3 ( .B1(n658), .B2(n671), .C1(n654), .C2(n712), .A(n147), .ZN(
        O[31]) );
  OAI221_X1 U4 ( .B1(n659), .B2(n677), .C1(n654), .C2(n718), .A(n141), .ZN(
        O[37]) );
  OAI221_X1 U5 ( .B1(n659), .B2(n689), .C1(n653), .C2(n727), .A(n131), .ZN(
        O[46]) );
  OAI221_X1 U6 ( .B1(n660), .B2(n687), .C1(n653), .C2(n726), .A(n132), .ZN(
        O[45]) );
  OAI221_X1 U7 ( .B1(n660), .B2(n696), .C1(n652), .C2(n731), .A(n126), .ZN(
        O[50]) );
  AOI22_X1 U8 ( .A1(\A_ns[23] ), .A2(n646), .B1(\A_s[23] ), .B2(n639), .ZN(
        n155) );
  AOI22_X1 U9 ( .A1(A_ns[54]), .A2(n649), .B1(A_s[54]), .B2(n642), .ZN(n121)
         );
  BUF_X1 U10 ( .A(n643), .Z(n646) );
  BUF_X1 U11 ( .A(n636), .Z(n639) );
  BUF_X1 U12 ( .A(n643), .Z(n647) );
  BUF_X1 U13 ( .A(n636), .Z(n640) );
  BUF_X1 U14 ( .A(n644), .Z(n648) );
  BUF_X1 U15 ( .A(n637), .Z(n641) );
  BUF_X1 U16 ( .A(n644), .Z(n649) );
  BUF_X1 U17 ( .A(n637), .Z(n642) );
  BUF_X1 U18 ( .A(n643), .Z(n645) );
  BUF_X1 U19 ( .A(n636), .Z(n638) );
  OAI221_X1 U20 ( .B1(n661), .B2(n702), .C1(n652), .C2(n736), .A(n121), .ZN(
        O[55]) );
  AOI22_X1 U21 ( .A1(\A_ns[30] ), .A2(n646), .B1(\A_s[30] ), .B2(n639), .ZN(
        n147) );
  OAI221_X1 U22 ( .B1(n658), .B2(n703), .C1(n655), .C2(n704), .A(n156), .ZN(
        O[23]) );
  AOI22_X1 U23 ( .A1(\A_ns[22] ), .A2(n646), .B1(\A_s[22] ), .B2(n639), .ZN(
        n156) );
  AOI22_X1 U24 ( .A1(\A_ns[24] ), .A2(n646), .B1(\A_s[24] ), .B2(n639), .ZN(
        n154) );
  OAI221_X1 U25 ( .B1(n658), .B2(n666), .C1(n655), .C2(n707), .A(n153), .ZN(
        O[26]) );
  AOI22_X1 U26 ( .A1(\A_ns[25] ), .A2(n646), .B1(\A_s[25] ), .B2(n639), .ZN(
        n153) );
  OAI221_X1 U27 ( .B1(n658), .B2(n667), .C1(n654), .C2(n708), .A(n152), .ZN(
        O[27]) );
  AOI22_X1 U28 ( .A1(\A_ns[26] ), .A2(n646), .B1(\A_s[26] ), .B2(n639), .ZN(
        n152) );
  OAI221_X1 U29 ( .B1(n658), .B2(n668), .C1(n654), .C2(n709), .A(n151), .ZN(
        O[28]) );
  AOI22_X1 U30 ( .A1(\A_ns[27] ), .A2(n646), .B1(\A_s[27] ), .B2(n639), .ZN(
        n151) );
  OAI221_X1 U31 ( .B1(n658), .B2(n669), .C1(n654), .C2(n710), .A(n150), .ZN(
        O[29]) );
  AOI22_X1 U32 ( .A1(\A_ns[28] ), .A2(n646), .B1(\A_s[28] ), .B2(n639), .ZN(
        n150) );
  OAI221_X1 U33 ( .B1(n658), .B2(n670), .C1(n654), .C2(n711), .A(n148), .ZN(
        O[30]) );
  AOI22_X1 U34 ( .A1(\A_ns[29] ), .A2(n646), .B1(\A_s[29] ), .B2(n639), .ZN(
        n148) );
  BUF_X1 U35 ( .A(n779), .Z(n636) );
  BUF_X1 U36 ( .A(n780), .Z(n643) );
  AOI22_X1 U37 ( .A1(\A_ns[36] ), .A2(n647), .B1(\A_s[36] ), .B2(n640), .ZN(
        n141) );
  OAI221_X1 U38 ( .B1(n658), .B2(n674), .C1(n654), .C2(n715), .A(n144), .ZN(
        O[34]) );
  AOI22_X1 U39 ( .A1(\A_ns[33] ), .A2(n647), .B1(\A_s[33] ), .B2(n640), .ZN(
        n144) );
  OAI221_X1 U40 ( .B1(n659), .B2(n684), .C1(n653), .C2(n723), .A(n135), .ZN(
        O[42]) );
  AOI22_X1 U41 ( .A1(\A_ns[41] ), .A2(n647), .B1(\A_s[41] ), .B2(n640), .ZN(
        n135) );
  OAI221_X1 U42 ( .B1(n658), .B2(n672), .C1(n654), .C2(n713), .A(n146), .ZN(
        O[32]) );
  AOI22_X1 U43 ( .A1(\A_ns[31] ), .A2(n646), .B1(\A_s[31] ), .B2(n639), .ZN(
        n146) );
  OAI221_X1 U44 ( .B1(n659), .B2(n678), .C1(n654), .C2(n719), .A(n140), .ZN(
        O[38]) );
  AOI22_X1 U45 ( .A1(\A_ns[37] ), .A2(n647), .B1(\A_s[37] ), .B2(n640), .ZN(
        n140) );
  OAI221_X1 U46 ( .B1(n659), .B2(n681), .C1(n653), .C2(n721), .A(n137), .ZN(
        O[40]) );
  AOI22_X1 U47 ( .A1(A_nso[41]), .A2(n647), .B1(\A_s[39] ), .B2(n640), .ZN(
        n137) );
  OAI221_X1 U48 ( .B1(n659), .B2(n685), .C1(n653), .C2(n724), .A(n134), .ZN(
        O[43]) );
  AOI22_X1 U49 ( .A1(\A_ns[42] ), .A2(n647), .B1(\A_s[42] ), .B2(n640), .ZN(
        n134) );
  OAI221_X1 U50 ( .B1(n659), .B2(n675), .C1(n654), .C2(n716), .A(n143), .ZN(
        O[35]) );
  AOI22_X1 U51 ( .A1(\A_ns[34] ), .A2(n647), .B1(\A_s[34] ), .B2(n640), .ZN(
        n143) );
  OAI221_X1 U52 ( .B1(n659), .B2(n679), .C1(n653), .C2(n720), .A(n139), .ZN(
        O[39]) );
  AOI22_X1 U53 ( .A1(A_nso[40]), .A2(n647), .B1(\A_s[38] ), .B2(n640), .ZN(
        n139) );
  OAI221_X1 U54 ( .B1(n658), .B2(n673), .C1(n654), .C2(n714), .A(n145), .ZN(
        O[33]) );
  AOI22_X1 U55 ( .A1(\A_ns[32] ), .A2(n647), .B1(\A_s[32] ), .B2(n640), .ZN(
        n145) );
  OAI221_X1 U56 ( .B1(n659), .B2(n683), .C1(n653), .C2(n722), .A(n136), .ZN(
        O[41]) );
  AOI22_X1 U57 ( .A1(\A_ns[40] ), .A2(n647), .B1(\A_s[40] ), .B2(n640), .ZN(
        n136) );
  OAI221_X1 U58 ( .B1(n659), .B2(n676), .C1(n654), .C2(n717), .A(n142), .ZN(
        O[36]) );
  AOI22_X1 U59 ( .A1(\A_ns[35] ), .A2(n647), .B1(\A_s[35] ), .B2(n640), .ZN(
        n142) );
  OAI221_X1 U60 ( .B1(n660), .B2(n686), .C1(n653), .C2(n725), .A(n133), .ZN(
        O[44]) );
  AOI22_X1 U61 ( .A1(\A_ns[43] ), .A2(n648), .B1(\A_s[43] ), .B2(n641), .ZN(
        n133) );
  AOI22_X1 U62 ( .A1(A_nso[47]), .A2(n648), .B1(\A_s[45] ), .B2(n641), .ZN(
        n131) );
  OAI221_X1 U63 ( .B1(n660), .B2(n691), .C1(n653), .C2(n728), .A(n130), .ZN(
        O[47]) );
  AOI22_X1 U64 ( .A1(A_nso[48]), .A2(n648), .B1(\A_s[46] ), .B2(n641), .ZN(
        n130) );
  AOI22_X1 U65 ( .A1(A_nso[46]), .A2(n648), .B1(\A_s[44] ), .B2(n641), .ZN(
        n132) );
  OAI221_X1 U66 ( .B1(n660), .B2(n693), .C1(n653), .C2(n729), .A(n129), .ZN(
        O[48]) );
  AOI22_X1 U67 ( .A1(A_nso[49]), .A2(n648), .B1(\A_s[47] ), .B2(n641), .ZN(
        n129) );
  OAI221_X1 U68 ( .B1(n660), .B2(n695), .C1(n653), .C2(n730), .A(n128), .ZN(
        O[49]) );
  AOI22_X1 U69 ( .A1(\A_ns[48] ), .A2(n648), .B1(\A_s[48] ), .B2(n641), .ZN(
        n128) );
  AOI22_X1 U70 ( .A1(\A_ns[49] ), .A2(n648), .B1(\A_s[49] ), .B2(n641), .ZN(
        n126) );
  OAI221_X1 U71 ( .B1(n660), .B2(n697), .C1(n652), .C2(n732), .A(n125), .ZN(
        O[51]) );
  AOI22_X1 U72 ( .A1(\A_ns[50] ), .A2(n648), .B1(\A_s[50] ), .B2(n641), .ZN(
        n125) );
  OAI221_X1 U73 ( .B1(n660), .B2(n698), .C1(n652), .C2(n733), .A(n124), .ZN(
        O[52]) );
  AOI22_X1 U74 ( .A1(\A_ns[51] ), .A2(n648), .B1(\A_s[51] ), .B2(n641), .ZN(
        n124) );
  OAI221_X1 U75 ( .B1(n660), .B2(n700), .C1(n652), .C2(n735), .A(n122), .ZN(
        O[54]) );
  AOI22_X1 U76 ( .A1(A_nso[55]), .A2(n648), .B1(\A_s[53] ), .B2(n641), .ZN(
        n122) );
  OAI221_X1 U77 ( .B1(n660), .B2(n699), .C1(n652), .C2(n734), .A(n123), .ZN(
        O[53]) );
  AOI22_X1 U78 ( .A1(\A_ns[52] ), .A2(n648), .B1(\A_s[52] ), .B2(n641), .ZN(
        n123) );
  BUF_X1 U79 ( .A(n779), .Z(n637) );
  BUF_X1 U80 ( .A(n780), .Z(n644) );
  OAI221_X1 U81 ( .B1(n658), .B2(n664), .C1(n655), .C2(n705), .A(n155), .ZN(
        O[24]) );
  BUF_X1 U82 ( .A(n663), .Z(n658) );
  BUF_X1 U83 ( .A(n651), .Z(n655) );
  INV_X1 U84 ( .A(n112), .ZN(n779) );
  INV_X1 U85 ( .A(n113), .ZN(n780) );
  BUF_X1 U86 ( .A(n650), .Z(n654) );
  BUF_X1 U87 ( .A(n662), .Z(n659) );
  BUF_X1 U88 ( .A(n650), .Z(n653) );
  BUF_X1 U89 ( .A(n662), .Z(n660) );
  BUF_X1 U90 ( .A(n650), .Z(n652) );
  BUF_X1 U91 ( .A(n662), .Z(n661) );
  BUF_X1 U92 ( .A(n663), .Z(n657) );
  BUF_X1 U93 ( .A(n651), .Z(n656) );
  NAND2_X1 U94 ( .A1(n170), .A2(n781), .ZN(n112) );
  NAND2_X1 U95 ( .A1(n170), .A2(n112), .ZN(n113) );
  BUF_X1 U96 ( .A(n114), .Z(n663) );
  BUF_X1 U97 ( .A(n115), .Z(n651) );
  BUF_X1 U98 ( .A(n115), .Z(n650) );
  BUF_X1 U99 ( .A(n114), .Z(n662) );
  OAI221_X1 U100 ( .B1(n659), .B2(n777), .C1(n655), .C2(n778), .A(n157), .ZN(
        O[22]) );
  INV_X1 U101 ( .A(\A_ns[20] ), .ZN(n777) );
  INV_X1 U102 ( .A(\A_s[20] ), .ZN(n778) );
  AOI22_X1 U103 ( .A1(\A_ns[21] ), .A2(n646), .B1(\A_s[21] ), .B2(n639), .ZN(
        n157) );
  INV_X1 U104 ( .A(B[23]), .ZN(n781) );
  OR3_X1 U105 ( .A1(B[21]), .A2(B[22]), .A3(n781), .ZN(n114) );
  OAI221_X1 U106 ( .B1(n657), .B2(n774), .C1(n655), .C2(n776), .A(n158), .ZN(
        O[21]) );
  INV_X1 U107 ( .A(\A_ns[19] ), .ZN(n774) );
  OAI221_X1 U108 ( .B1(n657), .B2(n762), .C1(n655), .C2(n764), .A(n164), .ZN(
        O[15]) );
  INV_X1 U109 ( .A(\A_ns[13] ), .ZN(n762) );
  INV_X1 U110 ( .A(\A_s[13] ), .ZN(n764) );
  OAI221_X1 U111 ( .B1(n657), .B2(n765), .C1(n655), .C2(n767), .A(n163), .ZN(
        O[16]) );
  INV_X1 U112 ( .A(\A_ns[14] ), .ZN(n765) );
  OAI221_X1 U113 ( .B1(n657), .B2(n766), .C1(n655), .C2(n768), .A(n162), .ZN(
        O[17]) );
  INV_X1 U114 ( .A(\A_ns[15] ), .ZN(n766) );
  OAI221_X1 U115 ( .B1(n657), .B2(n769), .C1(n655), .C2(n771), .A(n161), .ZN(
        O[18]) );
  INV_X1 U116 ( .A(\A_ns[16] ), .ZN(n769) );
  OAI221_X1 U117 ( .B1(n657), .B2(n770), .C1(n655), .C2(n772), .A(n160), .ZN(
        O[19]) );
  INV_X1 U118 ( .A(\A_ns[17] ), .ZN(n770) );
  OAI221_X1 U119 ( .B1(n657), .B2(n773), .C1(n655), .C2(n775), .A(n159), .ZN(
        O[20]) );
  INV_X1 U120 ( .A(\A_ns[18] ), .ZN(n773) );
  OAI221_X1 U121 ( .B1(n661), .B2(n746), .C1(n652), .C2(n748), .A(n118), .ZN(
        O[7]) );
  INV_X1 U122 ( .A(\A_ns[5] ), .ZN(n746) );
  INV_X1 U123 ( .A(\A_s[5] ), .ZN(n748) );
  OAI221_X1 U124 ( .B1(n660), .B2(n749), .C1(n652), .C2(n751), .A(n117), .ZN(
        O[8]) );
  INV_X1 U125 ( .A(\A_ns[6] ), .ZN(n749) );
  INV_X1 U126 ( .A(\A_s[6] ), .ZN(n751) );
  OAI221_X1 U127 ( .B1(n657), .B2(n750), .C1(n654), .C2(n752), .A(n116), .ZN(
        O[9]) );
  INV_X1 U128 ( .A(\A_ns[7] ), .ZN(n750) );
  INV_X1 U129 ( .A(\A_s[7] ), .ZN(n752) );
  OAI221_X1 U130 ( .B1(n753), .B2(n661), .C1(n755), .C2(n652), .A(n169), .ZN(
        O[10]) );
  INV_X1 U131 ( .A(\A_s[8] ), .ZN(n755) );
  INV_X1 U132 ( .A(\A_ns[8] ), .ZN(n753) );
  OAI221_X1 U133 ( .B1(n657), .B2(n754), .C1(n652), .C2(n756), .A(n168), .ZN(
        O[11]) );
  INV_X1 U134 ( .A(\A_ns[9] ), .ZN(n754) );
  INV_X1 U135 ( .A(\A_s[9] ), .ZN(n756) );
  OAI221_X1 U136 ( .B1(n657), .B2(n757), .C1(n656), .C2(n759), .A(n167), .ZN(
        O[12]) );
  INV_X1 U137 ( .A(\A_ns[10] ), .ZN(n757) );
  INV_X1 U138 ( .A(\A_s[10] ), .ZN(n759) );
  OAI221_X1 U139 ( .B1(n657), .B2(n758), .C1(n656), .C2(n760), .A(n166), .ZN(
        O[13]) );
  INV_X1 U140 ( .A(\A_ns[11] ), .ZN(n758) );
  INV_X1 U141 ( .A(\A_s[11] ), .ZN(n760) );
  OAI221_X1 U142 ( .B1(n657), .B2(n761), .C1(n655), .C2(n763), .A(n165), .ZN(
        O[14]) );
  INV_X1 U143 ( .A(\A_ns[12] ), .ZN(n761) );
  INV_X1 U144 ( .A(\A_s[12] ), .ZN(n763) );
  OAI22_X1 U145 ( .A1(n112), .A2(n739), .B1(n113), .B2(n737), .ZN(O[1]) );
  OAI221_X1 U146 ( .B1(n737), .B2(n661), .C1(n739), .C2(n652), .A(n149), .ZN(
        O[2]) );
  AOI22_X1 U147 ( .A1(\A_ns[1] ), .A2(n646), .B1(\A_s[1] ), .B2(n639), .ZN(
        n149) );
  OAI221_X1 U148 ( .B1(n659), .B2(n738), .C1(n653), .C2(n740), .A(n138), .ZN(
        O[3]) );
  INV_X1 U149 ( .A(\A_ns[1] ), .ZN(n738) );
  INV_X1 U150 ( .A(\A_s[1] ), .ZN(n740) );
  OAI221_X1 U151 ( .B1(n660), .B2(n741), .C1(n653), .C2(n743), .A(n127), .ZN(
        O[4]) );
  INV_X1 U152 ( .A(\A_ns[2] ), .ZN(n741) );
  INV_X1 U153 ( .A(\A_s[2] ), .ZN(n743) );
  OAI221_X1 U154 ( .B1(n661), .B2(n742), .C1(n652), .C2(n744), .A(n120), .ZN(
        O[5]) );
  INV_X1 U155 ( .A(\A_ns[3] ), .ZN(n742) );
  INV_X1 U156 ( .A(\A_s[3] ), .ZN(n744) );
  OAI221_X1 U157 ( .B1(n661), .B2(n745), .C1(n652), .C2(n747), .A(n119), .ZN(
        O[6]) );
  INV_X1 U158 ( .A(\A_ns[4] ), .ZN(n745) );
  INV_X1 U159 ( .A(\A_s[4] ), .ZN(n747) );
  INV_X1 U160 ( .A(\A_ns[0] ), .ZN(n737) );
  INV_X1 U161 ( .A(\A_s[0] ), .ZN(n739) );
  AOI22_X1 U162 ( .A1(\A_ns[2] ), .A2(n647), .B1(\A_s[2] ), .B2(n640), .ZN(
        n138) );
  AOI22_X1 U163 ( .A1(\A_ns[3] ), .A2(n648), .B1(\A_s[3] ), .B2(n641), .ZN(
        n127) );
  AOI22_X1 U164 ( .A1(\A_ns[4] ), .A2(n649), .B1(\A_s[4] ), .B2(n642), .ZN(
        n120) );
  AOI22_X1 U165 ( .A1(\A_ns[5] ), .A2(n649), .B1(\A_s[5] ), .B2(n642), .ZN(
        n119) );
  AOI22_X1 U166 ( .A1(\A_ns[6] ), .A2(n649), .B1(\A_s[6] ), .B2(n642), .ZN(
        n118) );
  AOI22_X1 U167 ( .A1(\A_ns[7] ), .A2(n649), .B1(\A_s[7] ), .B2(n642), .ZN(
        n117) );
  AOI22_X1 U168 ( .A1(\A_ns[8] ), .A2(n649), .B1(\A_s[8] ), .B2(n642), .ZN(
        n116) );
  AOI22_X1 U169 ( .A1(\A_ns[9] ), .A2(n645), .B1(\A_s[9] ), .B2(n638), .ZN(
        n169) );
  AOI22_X1 U170 ( .A1(\A_ns[10] ), .A2(n645), .B1(\A_s[10] ), .B2(n638), .ZN(
        n168) );
  AOI22_X1 U171 ( .A1(\A_ns[11] ), .A2(n645), .B1(\A_s[11] ), .B2(n638), .ZN(
        n167) );
  AOI22_X1 U172 ( .A1(\A_ns[12] ), .A2(n645), .B1(\A_s[12] ), .B2(n638), .ZN(
        n166) );
  AOI22_X1 U173 ( .A1(\A_ns[13] ), .A2(n645), .B1(\A_s[13] ), .B2(n638), .ZN(
        n165) );
  AOI22_X1 U174 ( .A1(\A_ns[14] ), .A2(n645), .B1(\A_s[14] ), .B2(n638), .ZN(
        n164) );
  AOI22_X1 U175 ( .A1(\A_ns[15] ), .A2(n645), .B1(\A_s[15] ), .B2(n638), .ZN(
        n163) );
  AOI22_X1 U176 ( .A1(\A_ns[16] ), .A2(n645), .B1(\A_s[16] ), .B2(n638), .ZN(
        n162) );
  AOI22_X1 U177 ( .A1(\A_ns[17] ), .A2(n645), .B1(\A_s[17] ), .B2(n638), .ZN(
        n161) );
  AOI22_X1 U178 ( .A1(\A_ns[18] ), .A2(n645), .B1(\A_s[18] ), .B2(n638), .ZN(
        n160) );
  AOI22_X1 U179 ( .A1(\A_ns[19] ), .A2(n645), .B1(\A_s[19] ), .B2(n638), .ZN(
        n159) );
  AOI22_X1 U180 ( .A1(\A_ns[20] ), .A2(n645), .B1(\A_s[20] ), .B2(n638), .ZN(
        n158) );
  INV_X1 U181 ( .A(\A_s[14] ), .ZN(n767) );
  INV_X1 U182 ( .A(\A_s[15] ), .ZN(n768) );
  INV_X1 U183 ( .A(\A_s[16] ), .ZN(n771) );
  INV_X1 U184 ( .A(\A_s[17] ), .ZN(n772) );
  INV_X1 U185 ( .A(\A_s[18] ), .ZN(n775) );
  INV_X1 U186 ( .A(\A_s[19] ), .ZN(n776) );
  INV_X1 U187 ( .A(\A_ns[22] ), .ZN(n664) );
  INV_X1 U188 ( .A(\A_ns[23] ), .ZN(n665) );
  INV_X1 U189 ( .A(\A_ns[24] ), .ZN(n666) );
  INV_X1 U190 ( .A(\A_ns[25] ), .ZN(n667) );
  INV_X1 U191 ( .A(\A_ns[26] ), .ZN(n668) );
  INV_X1 U192 ( .A(\A_ns[27] ), .ZN(n669) );
  INV_X1 U193 ( .A(\A_ns[28] ), .ZN(n670) );
  INV_X1 U194 ( .A(\A_ns[29] ), .ZN(n671) );
  INV_X1 U195 ( .A(\A_ns[30] ), .ZN(n672) );
  INV_X1 U196 ( .A(\A_ns[31] ), .ZN(n673) );
  INV_X1 U197 ( .A(\A_ns[32] ), .ZN(n674) );
  INV_X1 U198 ( .A(\A_ns[33] ), .ZN(n675) );
  INV_X1 U199 ( .A(\A_ns[34] ), .ZN(n676) );
  INV_X1 U200 ( .A(\A_ns[35] ), .ZN(n677) );
  INV_X1 U201 ( .A(\A_ns[36] ), .ZN(n678) );
  INV_X1 U202 ( .A(\A_ns[37] ), .ZN(n679) );
  INV_X1 U203 ( .A(n681), .ZN(A_nso[40]) );
  INV_X1 U204 ( .A(A_ns[38]), .ZN(n681) );
  INV_X1 U205 ( .A(n683), .ZN(A_nso[41]) );
  INV_X1 U206 ( .A(A_ns[39]), .ZN(n683) );
  INV_X1 U207 ( .A(\A_ns[40] ), .ZN(n684) );
  INV_X1 U208 ( .A(\A_ns[41] ), .ZN(n685) );
  INV_X1 U209 ( .A(\A_ns[42] ), .ZN(n686) );
  INV_X1 U210 ( .A(\A_ns[43] ), .ZN(n687) );
  INV_X1 U211 ( .A(n689), .ZN(A_nso[46]) );
  INV_X1 U212 ( .A(A_ns[44]), .ZN(n689) );
  INV_X1 U213 ( .A(n691), .ZN(A_nso[47]) );
  INV_X1 U214 ( .A(A_ns[45]), .ZN(n691) );
  INV_X1 U215 ( .A(n693), .ZN(A_nso[48]) );
  INV_X1 U216 ( .A(A_ns[46]), .ZN(n693) );
  INV_X1 U217 ( .A(n695), .ZN(A_nso[49]) );
  INV_X1 U218 ( .A(A_ns[47]), .ZN(n695) );
  INV_X1 U219 ( .A(\A_ns[48] ), .ZN(n696) );
  INV_X1 U220 ( .A(\A_ns[49] ), .ZN(n697) );
  INV_X1 U221 ( .A(\A_ns[50] ), .ZN(n698) );
  INV_X1 U222 ( .A(\A_ns[51] ), .ZN(n699) );
  INV_X1 U223 ( .A(\A_ns[52] ), .ZN(n700) );
  INV_X1 U224 ( .A(n702), .ZN(A_nso[55]) );
  INV_X1 U227 ( .A(A_ns[53]), .ZN(n702) );
  INV_X1 U228 ( .A(\A_ns[21] ), .ZN(n703) );
  INV_X1 U229 ( .A(\A_s[21] ), .ZN(n704) );
  INV_X1 U230 ( .A(\A_s[22] ), .ZN(n705) );
  INV_X1 U231 ( .A(\A_s[23] ), .ZN(n706) );
  INV_X1 U232 ( .A(\A_s[24] ), .ZN(n707) );
  INV_X1 U233 ( .A(\A_s[25] ), .ZN(n708) );
  INV_X1 U234 ( .A(\A_s[26] ), .ZN(n709) );
  INV_X1 U235 ( .A(\A_s[27] ), .ZN(n710) );
  INV_X1 U236 ( .A(\A_s[28] ), .ZN(n711) );
  INV_X1 U237 ( .A(\A_s[29] ), .ZN(n712) );
  INV_X1 U238 ( .A(\A_s[30] ), .ZN(n713) );
  INV_X1 U239 ( .A(\A_s[31] ), .ZN(n714) );
  INV_X1 U240 ( .A(\A_s[32] ), .ZN(n715) );
  INV_X1 U241 ( .A(\A_s[33] ), .ZN(n716) );
  INV_X1 U242 ( .A(\A_s[34] ), .ZN(n717) );
  INV_X1 U243 ( .A(\A_s[35] ), .ZN(n718) );
  INV_X1 U244 ( .A(\A_s[36] ), .ZN(n719) );
  INV_X1 U245 ( .A(\A_s[37] ), .ZN(n720) );
  INV_X1 U246 ( .A(\A_s[38] ), .ZN(n721) );
  INV_X1 U247 ( .A(\A_s[39] ), .ZN(n722) );
  INV_X1 U248 ( .A(\A_s[40] ), .ZN(n723) );
  INV_X1 U249 ( .A(\A_s[41] ), .ZN(n724) );
  INV_X1 U250 ( .A(\A_s[42] ), .ZN(n725) );
  INV_X1 U251 ( .A(\A_s[43] ), .ZN(n726) );
  INV_X1 U252 ( .A(\A_s[44] ), .ZN(n727) );
  INV_X1 U253 ( .A(\A_s[45] ), .ZN(n728) );
  INV_X1 U254 ( .A(\A_s[46] ), .ZN(n729) );
  INV_X1 U255 ( .A(\A_s[47] ), .ZN(n730) );
  INV_X1 U256 ( .A(\A_s[48] ), .ZN(n731) );
  INV_X1 U257 ( .A(\A_s[49] ), .ZN(n732) );
  INV_X1 U258 ( .A(\A_s[50] ), .ZN(n733) );
  INV_X1 U259 ( .A(\A_s[51] ), .ZN(n734) );
  INV_X1 U260 ( .A(\A_s[52] ), .ZN(n735) );
  INV_X1 U261 ( .A(\A_s[53] ), .ZN(n736) );
endmodule


module BOOTHENC_NBIT58_i24 ( A_s, A_ns, B, O, A_so, A_nso );
  input [57:0] A_s;
  input [57:0] A_ns;
  input [57:0] B;
  output [57:0] O;
  output [57:0] A_so;
  output [57:0] A_nso;
  wire   \A_s[55] , \A_s[54] , \A_s[53] , \A_s[49] , \A_s[48] , \A_s[47] ,
         \A_s[46] , \A_s[45] , \A_s[44] , \A_s[43] , \A_s[42] , \A_s[41] ,
         \A_s[40] , \A_s[39] , \A_s[38] , \A_s[35] , \A_s[34] , \A_s[33] ,
         \A_s[32] , \A_s[31] , \A_s[30] , \A_s[29] , \A_s[28] , \A_s[27] ,
         \A_s[26] , \A_s[25] , \A_s[24] , \A_s[23] , \A_s[22] , \A_s[21] ,
         \A_s[20] , \A_s[19] , \A_s[18] , \A_s[17] , \A_s[16] , \A_s[15] ,
         \A_s[14] , \A_s[13] , \A_s[12] , \A_s[11] , \A_s[10] , \A_s[9] ,
         \A_s[8] , \A_s[7] , \A_s[6] , \A_s[5] , \A_s[4] , \A_s[3] , \A_s[2] ,
         \A_s[1] , \A_s[0] , \A_ns[55] , \A_ns[54] , \A_ns[53] , \A_ns[52] ,
         \A_ns[51] , \A_ns[50] , \A_ns[49] , \A_ns[48] , \A_ns[47] ,
         \A_ns[46] , \A_ns[45] , \A_ns[44] , \A_ns[43] , \A_ns[42] ,
         \A_ns[41] , \A_ns[40] , \A_ns[39] , \A_ns[37] , \A_ns[36] ,
         \A_ns[35] , \A_ns[34] , \A_ns[33] , \A_ns[32] , \A_ns[31] ,
         \A_ns[30] , \A_ns[29] , \A_ns[28] , \A_ns[27] , \A_ns[26] ,
         \A_ns[25] , \A_ns[24] , \A_ns[23] , \A_ns[22] , \A_ns[21] ,
         \A_ns[20] , \A_ns[19] , \A_ns[18] , \A_ns[17] , \A_ns[16] ,
         \A_ns[15] , \A_ns[14] , \A_ns[13] , \A_ns[12] , \A_ns[11] ,
         \A_ns[10] , \A_ns[9] , \A_ns[8] , \A_ns[7] , \A_ns[6] , \A_ns[5] ,
         \A_ns[4] , \A_ns[3] , \A_ns[2] , \A_ns[1] , \A_ns[0] , n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n754, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n770, n772, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826;
  assign A_nso[0] = 1'b0;
  assign A_nso[1] = 1'b0;
  assign A_so[0] = 1'b0;
  assign A_so[1] = 1'b0;
  assign O[0] = 1'b0;
  assign A_so[57] = \A_s[55] ;
  assign \A_s[55]  = A_s[55];
  assign A_so[56] = \A_s[54] ;
  assign \A_s[54]  = A_s[54];
  assign A_so[55] = \A_s[53] ;
  assign \A_s[53]  = A_s[53];
  assign A_so[51] = \A_s[49] ;
  assign \A_s[49]  = A_s[49];
  assign A_so[50] = \A_s[48] ;
  assign \A_s[48]  = A_s[48];
  assign A_so[49] = \A_s[47] ;
  assign \A_s[47]  = A_s[47];
  assign A_so[48] = \A_s[46] ;
  assign \A_s[46]  = A_s[46];
  assign A_so[47] = \A_s[45] ;
  assign \A_s[45]  = A_s[45];
  assign A_so[46] = \A_s[44] ;
  assign \A_s[44]  = A_s[44];
  assign A_so[45] = \A_s[43] ;
  assign \A_s[43]  = A_s[43];
  assign A_so[44] = \A_s[42] ;
  assign \A_s[42]  = A_s[42];
  assign A_so[43] = \A_s[41] ;
  assign \A_s[41]  = A_s[41];
  assign A_so[42] = \A_s[40] ;
  assign \A_s[40]  = A_s[40];
  assign A_so[41] = \A_s[39] ;
  assign \A_s[39]  = A_s[39];
  assign A_so[40] = \A_s[38] ;
  assign \A_s[38]  = A_s[38];
  assign A_so[37] = \A_s[35] ;
  assign \A_s[35]  = A_s[35];
  assign A_so[36] = \A_s[34] ;
  assign \A_s[34]  = A_s[34];
  assign A_so[35] = \A_s[33] ;
  assign \A_s[33]  = A_s[33];
  assign A_so[34] = \A_s[32] ;
  assign \A_s[32]  = A_s[32];
  assign A_so[33] = \A_s[31] ;
  assign \A_s[31]  = A_s[31];
  assign A_so[32] = \A_s[30] ;
  assign \A_s[30]  = A_s[30];
  assign A_so[31] = \A_s[29] ;
  assign \A_s[29]  = A_s[29];
  assign A_so[30] = \A_s[28] ;
  assign \A_s[28]  = A_s[28];
  assign A_so[29] = \A_s[27] ;
  assign \A_s[27]  = A_s[27];
  assign A_so[28] = \A_s[26] ;
  assign \A_s[26]  = A_s[26];
  assign A_so[27] = \A_s[25] ;
  assign \A_s[25]  = A_s[25];
  assign A_so[26] = \A_s[24] ;
  assign \A_s[24]  = A_s[24];
  assign A_so[25] = \A_s[23] ;
  assign \A_s[23]  = A_s[23];
  assign A_so[24] = \A_s[22] ;
  assign \A_s[22]  = A_s[22];
  assign A_so[23] = \A_s[21] ;
  assign \A_s[21]  = A_s[21];
  assign A_so[22] = \A_s[20] ;
  assign \A_s[20]  = A_s[20];
  assign A_so[21] = \A_s[19] ;
  assign \A_s[19]  = A_s[19];
  assign A_so[20] = \A_s[18] ;
  assign \A_s[18]  = A_s[18];
  assign A_so[19] = \A_s[17] ;
  assign \A_s[17]  = A_s[17];
  assign A_so[18] = \A_s[16] ;
  assign \A_s[16]  = A_s[16];
  assign A_so[17] = \A_s[15] ;
  assign \A_s[15]  = A_s[15];
  assign A_so[16] = \A_s[14] ;
  assign \A_s[14]  = A_s[14];
  assign A_so[15] = \A_s[13] ;
  assign \A_s[13]  = A_s[13];
  assign A_so[14] = \A_s[12] ;
  assign \A_s[12]  = A_s[12];
  assign A_so[13] = \A_s[11] ;
  assign \A_s[11]  = A_s[11];
  assign A_so[12] = \A_s[10] ;
  assign \A_s[10]  = A_s[10];
  assign A_so[11] = \A_s[9] ;
  assign \A_s[9]  = A_s[9];
  assign A_so[10] = \A_s[8] ;
  assign \A_s[8]  = A_s[8];
  assign A_so[9] = \A_s[7] ;
  assign \A_s[7]  = A_s[7];
  assign A_so[8] = \A_s[6] ;
  assign \A_s[6]  = A_s[6];
  assign A_so[7] = \A_s[5] ;
  assign \A_s[5]  = A_s[5];
  assign A_so[6] = \A_s[4] ;
  assign \A_s[4]  = A_s[4];
  assign A_so[5] = \A_s[3] ;
  assign \A_s[3]  = A_s[3];
  assign A_so[4] = \A_s[2] ;
  assign \A_s[2]  = A_s[2];
  assign A_so[3] = \A_s[1] ;
  assign \A_s[1]  = A_s[1];
  assign A_so[2] = \A_s[0] ;
  assign \A_s[0]  = A_s[0];
  assign A_nso[57] = \A_ns[55] ;
  assign \A_ns[55]  = A_ns[55];
  assign A_nso[56] = \A_ns[54] ;
  assign \A_ns[54]  = A_ns[54];
  assign A_nso[55] = \A_ns[53] ;
  assign \A_ns[53]  = A_ns[53];
  assign A_nso[54] = \A_ns[52] ;
  assign \A_ns[52]  = A_ns[52];
  assign A_nso[53] = \A_ns[51] ;
  assign \A_ns[51]  = A_ns[51];
  assign A_nso[52] = \A_ns[50] ;
  assign \A_ns[50]  = A_ns[50];
  assign A_nso[51] = \A_ns[49] ;
  assign \A_ns[49]  = A_ns[49];
  assign A_nso[50] = \A_ns[48] ;
  assign \A_ns[48]  = A_ns[48];
  assign A_nso[49] = \A_ns[47] ;
  assign \A_ns[47]  = A_ns[47];
  assign A_nso[48] = \A_ns[46] ;
  assign \A_ns[46]  = A_ns[46];
  assign A_nso[47] = \A_ns[45] ;
  assign \A_ns[45]  = A_ns[45];
  assign A_nso[46] = \A_ns[44] ;
  assign \A_ns[44]  = A_ns[44];
  assign A_nso[45] = \A_ns[43] ;
  assign \A_ns[43]  = A_ns[43];
  assign A_nso[44] = \A_ns[42] ;
  assign \A_ns[42]  = A_ns[42];
  assign A_nso[43] = \A_ns[41] ;
  assign \A_ns[41]  = A_ns[41];
  assign A_nso[42] = \A_ns[40] ;
  assign \A_ns[40]  = A_ns[40];
  assign A_nso[41] = \A_ns[39] ;
  assign \A_ns[39]  = A_ns[39];
  assign A_nso[39] = \A_ns[37] ;
  assign \A_ns[37]  = A_ns[37];
  assign A_nso[38] = \A_ns[36] ;
  assign \A_ns[36]  = A_ns[36];
  assign A_nso[37] = \A_ns[35] ;
  assign \A_ns[35]  = A_ns[35];
  assign A_nso[36] = \A_ns[34] ;
  assign \A_ns[34]  = A_ns[34];
  assign A_nso[35] = \A_ns[33] ;
  assign \A_ns[33]  = A_ns[33];
  assign A_nso[34] = \A_ns[32] ;
  assign \A_ns[32]  = A_ns[32];
  assign A_nso[33] = \A_ns[31] ;
  assign \A_ns[31]  = A_ns[31];
  assign A_nso[32] = \A_ns[30] ;
  assign \A_ns[30]  = A_ns[30];
  assign A_nso[31] = \A_ns[29] ;
  assign \A_ns[29]  = A_ns[29];
  assign A_nso[30] = \A_ns[28] ;
  assign \A_ns[28]  = A_ns[28];
  assign A_nso[29] = \A_ns[27] ;
  assign \A_ns[27]  = A_ns[27];
  assign A_nso[28] = \A_ns[26] ;
  assign \A_ns[26]  = A_ns[26];
  assign A_nso[27] = \A_ns[25] ;
  assign \A_ns[25]  = A_ns[25];
  assign A_nso[26] = \A_ns[24] ;
  assign \A_ns[24]  = A_ns[24];
  assign A_nso[25] = \A_ns[23] ;
  assign \A_ns[23]  = A_ns[23];
  assign A_nso[24] = \A_ns[22] ;
  assign \A_ns[22]  = A_ns[22];
  assign A_nso[23] = \A_ns[21] ;
  assign \A_ns[21]  = A_ns[21];
  assign A_nso[22] = \A_ns[20] ;
  assign \A_ns[20]  = A_ns[20];
  assign A_nso[21] = \A_ns[19] ;
  assign \A_ns[19]  = A_ns[19];
  assign A_nso[20] = \A_ns[18] ;
  assign \A_ns[18]  = A_ns[18];
  assign A_nso[19] = \A_ns[17] ;
  assign \A_ns[17]  = A_ns[17];
  assign A_nso[18] = \A_ns[16] ;
  assign \A_ns[16]  = A_ns[16];
  assign A_nso[17] = \A_ns[15] ;
  assign \A_ns[15]  = A_ns[15];
  assign A_nso[16] = \A_ns[14] ;
  assign \A_ns[14]  = A_ns[14];
  assign A_nso[15] = \A_ns[13] ;
  assign \A_ns[13]  = A_ns[13];
  assign A_nso[14] = \A_ns[12] ;
  assign \A_ns[12]  = A_ns[12];
  assign A_nso[13] = \A_ns[11] ;
  assign \A_ns[11]  = A_ns[11];
  assign A_nso[12] = \A_ns[10] ;
  assign \A_ns[10]  = A_ns[10];
  assign A_nso[11] = \A_ns[9] ;
  assign \A_ns[9]  = A_ns[9];
  assign A_nso[10] = \A_ns[8] ;
  assign \A_ns[8]  = A_ns[8];
  assign A_nso[9] = \A_ns[7] ;
  assign \A_ns[7]  = A_ns[7];
  assign A_nso[8] = \A_ns[6] ;
  assign \A_ns[6]  = A_ns[6];
  assign A_nso[7] = \A_ns[5] ;
  assign \A_ns[5]  = A_ns[5];
  assign A_nso[6] = \A_ns[4] ;
  assign \A_ns[4]  = A_ns[4];
  assign A_nso[5] = \A_ns[3] ;
  assign \A_ns[3]  = A_ns[3];
  assign A_nso[4] = \A_ns[2] ;
  assign \A_ns[2]  = A_ns[2];
  assign A_nso[3] = \A_ns[1] ;
  assign \A_ns[1]  = A_ns[1];
  assign A_nso[2] = \A_ns[0] ;
  assign \A_ns[0]  = A_ns[0];

  XOR2_X1 U233 ( .A(B[23]), .B(B[24]), .Z(n176) );
  NAND3_X1 U234 ( .A1(B[24]), .A2(n826), .A3(B[23]), .ZN(n117) );
  OAI221_X1 U2 ( .B1(n699), .B2(n737), .C1(n697), .C2(n776), .A(n124), .ZN(
        O[56]) );
  BUF_X1 U3 ( .A(n685), .Z(n688) );
  BUF_X1 U4 ( .A(n678), .Z(n681) );
  BUF_X1 U5 ( .A(n685), .Z(n689) );
  BUF_X1 U6 ( .A(n678), .Z(n682) );
  BUF_X1 U7 ( .A(n686), .Z(n690) );
  BUF_X1 U8 ( .A(n679), .Z(n683) );
  BUF_X1 U9 ( .A(n686), .Z(n691) );
  BUF_X1 U10 ( .A(n679), .Z(n684) );
  BUF_X1 U11 ( .A(n685), .Z(n687) );
  BUF_X1 U12 ( .A(n678), .Z(n680) );
  OAI221_X1 U13 ( .B1(n699), .B2(n738), .C1(n697), .C2(n777), .A(n123), .ZN(
        O[57]) );
  AOI22_X1 U14 ( .A1(A_ns[56]), .A2(n691), .B1(A_s[56]), .B2(n684), .ZN(n123)
         );
  AOI22_X1 U15 ( .A1(\A_ns[55] ), .A2(n691), .B1(\A_s[55] ), .B2(n684), .ZN(
        n124) );
  OAI221_X1 U16 ( .B1(n702), .B2(n739), .C1(n695), .C2(n740), .A(n158), .ZN(
        O[25]) );
  AOI22_X1 U17 ( .A1(\A_ns[24] ), .A2(n688), .B1(\A_s[24] ), .B2(n681), .ZN(
        n158) );
  OAI221_X1 U18 ( .B1(n702), .B2(n706), .C1(n695), .C2(n741), .A(n157), .ZN(
        O[26]) );
  AOI22_X1 U19 ( .A1(\A_ns[25] ), .A2(n688), .B1(\A_s[25] ), .B2(n681), .ZN(
        n157) );
  OAI221_X1 U20 ( .B1(n702), .B2(n707), .C1(n695), .C2(n742), .A(n156), .ZN(
        O[27]) );
  AOI22_X1 U21 ( .A1(\A_ns[26] ), .A2(n688), .B1(\A_s[26] ), .B2(n681), .ZN(
        n156) );
  BUF_X1 U22 ( .A(n824), .Z(n678) );
  BUF_X1 U23 ( .A(n825), .Z(n685) );
  OAI221_X1 U24 ( .B1(n702), .B2(n709), .C1(n695), .C2(n744), .A(n154), .ZN(
        O[29]) );
  AOI22_X1 U25 ( .A1(\A_ns[28] ), .A2(n688), .B1(\A_s[28] ), .B2(n681), .ZN(
        n154) );
  OAI221_X1 U26 ( .B1(n701), .B2(n711), .C1(n695), .C2(n746), .A(n151), .ZN(
        O[31]) );
  AOI22_X1 U27 ( .A1(\A_ns[30] ), .A2(n688), .B1(\A_s[30] ), .B2(n681), .ZN(
        n151) );
  OAI221_X1 U28 ( .B1(n701), .B2(n712), .C1(n695), .C2(n747), .A(n150), .ZN(
        O[32]) );
  AOI22_X1 U29 ( .A1(\A_ns[31] ), .A2(n688), .B1(\A_s[31] ), .B2(n681), .ZN(
        n150) );
  OAI221_X1 U30 ( .B1(n701), .B2(n713), .C1(n695), .C2(n748), .A(n149), .ZN(
        O[33]) );
  AOI22_X1 U31 ( .A1(\A_ns[32] ), .A2(n689), .B1(\A_s[32] ), .B2(n682), .ZN(
        n149) );
  OAI221_X1 U32 ( .B1(n701), .B2(n714), .C1(n695), .C2(n749), .A(n148), .ZN(
        O[34]) );
  AOI22_X1 U33 ( .A1(\A_ns[33] ), .A2(n689), .B1(\A_s[33] ), .B2(n682), .ZN(
        n148) );
  OAI221_X1 U34 ( .B1(n701), .B2(n715), .C1(n696), .C2(n750), .A(n147), .ZN(
        O[35]) );
  AOI22_X1 U35 ( .A1(\A_ns[34] ), .A2(n689), .B1(\A_s[34] ), .B2(n682), .ZN(
        n147) );
  OAI221_X1 U36 ( .B1(n701), .B2(n716), .C1(n696), .C2(n751), .A(n146), .ZN(
        O[36]) );
  AOI22_X1 U37 ( .A1(\A_ns[35] ), .A2(n689), .B1(\A_s[35] ), .B2(n682), .ZN(
        n146) );
  OAI221_X1 U38 ( .B1(n701), .B2(n717), .C1(n696), .C2(n752), .A(n145), .ZN(
        O[37]) );
  AOI22_X1 U39 ( .A1(\A_ns[36] ), .A2(n689), .B1(A_so[38]), .B2(n682), .ZN(
        n145) );
  OAI221_X1 U40 ( .B1(n701), .B2(n718), .C1(n696), .C2(n754), .A(n144), .ZN(
        O[38]) );
  AOI22_X1 U41 ( .A1(\A_ns[37] ), .A2(n689), .B1(A_so[39]), .B2(n682), .ZN(
        n144) );
  OAI221_X1 U42 ( .B1(n701), .B2(n719), .C1(n696), .C2(n756), .A(n143), .ZN(
        O[39]) );
  AOI22_X1 U43 ( .A1(A_nso[40]), .A2(n689), .B1(\A_s[38] ), .B2(n682), .ZN(
        n143) );
  OAI221_X1 U44 ( .B1(n700), .B2(n721), .C1(n696), .C2(n757), .A(n141), .ZN(
        O[40]) );
  AOI22_X1 U45 ( .A1(\A_ns[39] ), .A2(n689), .B1(\A_s[39] ), .B2(n682), .ZN(
        n141) );
  OAI221_X1 U46 ( .B1(n700), .B2(n722), .C1(n696), .C2(n758), .A(n140), .ZN(
        O[41]) );
  AOI22_X1 U47 ( .A1(\A_ns[40] ), .A2(n689), .B1(\A_s[40] ), .B2(n682), .ZN(
        n140) );
  OAI221_X1 U48 ( .B1(n702), .B2(n708), .C1(n695), .C2(n743), .A(n155), .ZN(
        O[28]) );
  AOI22_X1 U49 ( .A1(\A_ns[27] ), .A2(n688), .B1(\A_s[27] ), .B2(n681), .ZN(
        n155) );
  OAI221_X1 U50 ( .B1(n701), .B2(n710), .C1(n695), .C2(n745), .A(n152), .ZN(
        O[30]) );
  AOI22_X1 U51 ( .A1(\A_ns[29] ), .A2(n688), .B1(\A_s[29] ), .B2(n681), .ZN(
        n152) );
  OAI221_X1 U52 ( .B1(n700), .B2(n723), .C1(n696), .C2(n759), .A(n139), .ZN(
        O[42]) );
  AOI22_X1 U53 ( .A1(\A_ns[41] ), .A2(n689), .B1(\A_s[41] ), .B2(n682), .ZN(
        n139) );
  OAI221_X1 U54 ( .B1(n700), .B2(n724), .C1(n696), .C2(n760), .A(n138), .ZN(
        O[43]) );
  AOI22_X1 U55 ( .A1(\A_ns[42] ), .A2(n689), .B1(\A_s[42] ), .B2(n682), .ZN(
        n138) );
  OAI221_X1 U56 ( .B1(n700), .B2(n725), .C1(n696), .C2(n761), .A(n137), .ZN(
        O[44]) );
  AOI22_X1 U57 ( .A1(\A_ns[43] ), .A2(n690), .B1(\A_s[43] ), .B2(n683), .ZN(
        n137) );
  OAI221_X1 U58 ( .B1(n700), .B2(n726), .C1(n696), .C2(n762), .A(n136), .ZN(
        O[45]) );
  AOI22_X1 U59 ( .A1(\A_ns[44] ), .A2(n690), .B1(\A_s[44] ), .B2(n683), .ZN(
        n136) );
  OAI221_X1 U60 ( .B1(n700), .B2(n728), .C1(n697), .C2(n764), .A(n134), .ZN(
        O[47]) );
  AOI22_X1 U61 ( .A1(\A_ns[46] ), .A2(n690), .B1(\A_s[46] ), .B2(n683), .ZN(
        n134) );
  OAI221_X1 U62 ( .B1(n700), .B2(n729), .C1(n697), .C2(n765), .A(n133), .ZN(
        O[48]) );
  AOI22_X1 U63 ( .A1(\A_ns[47] ), .A2(n690), .B1(\A_s[47] ), .B2(n683), .ZN(
        n133) );
  OAI221_X1 U64 ( .B1(n700), .B2(n730), .C1(n697), .C2(n766), .A(n132), .ZN(
        O[49]) );
  AOI22_X1 U65 ( .A1(\A_ns[48] ), .A2(n690), .B1(\A_s[48] ), .B2(n683), .ZN(
        n132) );
  OAI221_X1 U66 ( .B1(n700), .B2(n731), .C1(n697), .C2(n767), .A(n130), .ZN(
        O[50]) );
  AOI22_X1 U67 ( .A1(\A_ns[49] ), .A2(n690), .B1(\A_s[49] ), .B2(n683), .ZN(
        n130) );
  OAI221_X1 U68 ( .B1(n699), .B2(n732), .C1(n697), .C2(n768), .A(n129), .ZN(
        O[51]) );
  AOI22_X1 U69 ( .A1(\A_ns[50] ), .A2(n690), .B1(A_so[52]), .B2(n683), .ZN(
        n129) );
  OAI221_X1 U70 ( .B1(n699), .B2(n733), .C1(n697), .C2(n770), .A(n128), .ZN(
        O[52]) );
  AOI22_X1 U71 ( .A1(\A_ns[51] ), .A2(n690), .B1(A_so[53]), .B2(n683), .ZN(
        n128) );
  OAI221_X1 U72 ( .B1(n699), .B2(n734), .C1(n697), .C2(n772), .A(n127), .ZN(
        O[53]) );
  AOI22_X1 U73 ( .A1(\A_ns[52] ), .A2(n690), .B1(A_so[54]), .B2(n683), .ZN(
        n127) );
  OAI221_X1 U74 ( .B1(n700), .B2(n727), .C1(n696), .C2(n763), .A(n135), .ZN(
        O[46]) );
  AOI22_X1 U75 ( .A1(\A_ns[45] ), .A2(n690), .B1(\A_s[45] ), .B2(n683), .ZN(
        n135) );
  OAI221_X1 U76 ( .B1(n699), .B2(n735), .C1(n697), .C2(n774), .A(n126), .ZN(
        O[54]) );
  AOI22_X1 U77 ( .A1(\A_ns[53] ), .A2(n690), .B1(\A_s[53] ), .B2(n683), .ZN(
        n126) );
  OAI221_X1 U78 ( .B1(n699), .B2(n736), .C1(n697), .C2(n775), .A(n125), .ZN(
        O[55]) );
  AOI22_X1 U79 ( .A1(\A_ns[54] ), .A2(n691), .B1(\A_s[54] ), .B2(n684), .ZN(
        n125) );
  BUF_X1 U80 ( .A(n824), .Z(n679) );
  BUF_X1 U81 ( .A(n825), .Z(n686) );
  INV_X1 U82 ( .A(n164), .ZN(n824) );
  INV_X1 U83 ( .A(n165), .ZN(n825) );
  BUF_X1 U84 ( .A(n704), .Z(n701) );
  BUF_X1 U85 ( .A(n704), .Z(n702) );
  BUF_X1 U86 ( .A(n692), .Z(n695) );
  BUF_X1 U87 ( .A(n692), .Z(n696) );
  BUF_X1 U88 ( .A(n705), .Z(n700) );
  BUF_X1 U89 ( .A(n705), .Z(n699) );
  BUF_X1 U90 ( .A(n693), .Z(n697) );
  BUF_X1 U91 ( .A(n692), .Z(n694) );
  BUF_X1 U92 ( .A(n704), .Z(n703) );
  BUF_X1 U93 ( .A(n693), .Z(n698) );
  NAND2_X1 U94 ( .A1(n176), .A2(n826), .ZN(n164) );
  NAND2_X1 U95 ( .A1(n176), .A2(n164), .ZN(n165) );
  BUF_X1 U96 ( .A(n117), .Z(n692) );
  BUF_X1 U97 ( .A(n116), .Z(n704) );
  BUF_X1 U98 ( .A(n116), .Z(n705) );
  BUF_X1 U99 ( .A(n117), .Z(n693) );
  OAI221_X1 U100 ( .B1(n702), .B2(n822), .C1(n695), .C2(n823), .A(n159), .ZN(
        O[24]) );
  INV_X1 U101 ( .A(\A_ns[22] ), .ZN(n822) );
  INV_X1 U102 ( .A(\A_s[22] ), .ZN(n823) );
  AOI22_X1 U103 ( .A1(\A_ns[23] ), .A2(n688), .B1(\A_s[23] ), .B2(n681), .ZN(
        n159) );
  INV_X1 U104 ( .A(B[25]), .ZN(n826) );
  OAI221_X1 U105 ( .B1(n702), .B2(n815), .C1(n694), .C2(n817), .A(n162), .ZN(
        O[21]) );
  INV_X1 U106 ( .A(\A_ns[19] ), .ZN(n815) );
  INV_X1 U107 ( .A(\A_s[19] ), .ZN(n817) );
  OAI221_X1 U108 ( .B1(n702), .B2(n818), .C1(n694), .C2(n820), .A(n161), .ZN(
        O[22]) );
  INV_X1 U109 ( .A(\A_ns[20] ), .ZN(n818) );
  OAI221_X1 U110 ( .B1(n702), .B2(n819), .C1(n695), .C2(n821), .A(n160), .ZN(
        O[23]) );
  INV_X1 U111 ( .A(\A_ns[21] ), .ZN(n819) );
  OR3_X1 U112 ( .A1(B[23]), .A2(B[24]), .A3(n826), .ZN(n116) );
  OAI221_X1 U113 ( .B1(n703), .B2(n803), .C1(n694), .C2(n805), .A(n170), .ZN(
        O[15]) );
  INV_X1 U114 ( .A(\A_ns[13] ), .ZN(n803) );
  INV_X1 U115 ( .A(\A_s[13] ), .ZN(n805) );
  OAI221_X1 U116 ( .B1(n703), .B2(n806), .C1(n694), .C2(n808), .A(n169), .ZN(
        O[16]) );
  INV_X1 U117 ( .A(\A_ns[14] ), .ZN(n806) );
  INV_X1 U118 ( .A(\A_s[14] ), .ZN(n808) );
  OAI221_X1 U119 ( .B1(n703), .B2(n807), .C1(n694), .C2(n809), .A(n168), .ZN(
        O[17]) );
  INV_X1 U120 ( .A(\A_ns[15] ), .ZN(n807) );
  INV_X1 U121 ( .A(\A_s[15] ), .ZN(n809) );
  OAI221_X1 U122 ( .B1(n702), .B2(n810), .C1(n694), .C2(n812), .A(n167), .ZN(
        O[18]) );
  INV_X1 U123 ( .A(\A_ns[16] ), .ZN(n810) );
  INV_X1 U124 ( .A(\A_s[16] ), .ZN(n812) );
  OAI221_X1 U125 ( .B1(n702), .B2(n811), .C1(n694), .C2(n813), .A(n166), .ZN(
        O[19]) );
  INV_X1 U126 ( .A(\A_ns[17] ), .ZN(n811) );
  INV_X1 U127 ( .A(\A_s[17] ), .ZN(n813) );
  OAI221_X1 U128 ( .B1(n702), .B2(n814), .C1(n694), .C2(n816), .A(n163), .ZN(
        O[20]) );
  INV_X1 U129 ( .A(\A_ns[18] ), .ZN(n814) );
  INV_X1 U130 ( .A(\A_s[18] ), .ZN(n816) );
  OAI221_X1 U131 ( .B1(n699), .B2(n787), .C1(n698), .C2(n789), .A(n120), .ZN(
        O[7]) );
  INV_X1 U132 ( .A(\A_ns[5] ), .ZN(n787) );
  INV_X1 U133 ( .A(\A_s[5] ), .ZN(n789) );
  OAI221_X1 U134 ( .B1(n699), .B2(n790), .C1(n698), .C2(n792), .A(n119), .ZN(
        O[8]) );
  INV_X1 U135 ( .A(\A_ns[6] ), .ZN(n790) );
  INV_X1 U136 ( .A(\A_s[6] ), .ZN(n792) );
  OAI221_X1 U137 ( .B1(n699), .B2(n791), .C1(n698), .C2(n793), .A(n118), .ZN(
        O[9]) );
  INV_X1 U138 ( .A(\A_ns[7] ), .ZN(n791) );
  INV_X1 U139 ( .A(\A_s[7] ), .ZN(n793) );
  OAI221_X1 U140 ( .B1(n794), .B2(n703), .C1(n796), .C2(n694), .A(n175), .ZN(
        O[10]) );
  INV_X1 U141 ( .A(\A_s[8] ), .ZN(n796) );
  INV_X1 U142 ( .A(\A_ns[8] ), .ZN(n794) );
  OAI221_X1 U143 ( .B1(n703), .B2(n795), .C1(n694), .C2(n797), .A(n174), .ZN(
        O[11]) );
  INV_X1 U144 ( .A(\A_ns[9] ), .ZN(n795) );
  INV_X1 U145 ( .A(\A_s[9] ), .ZN(n797) );
  OAI221_X1 U146 ( .B1(n703), .B2(n798), .C1(n694), .C2(n800), .A(n173), .ZN(
        O[12]) );
  INV_X1 U147 ( .A(\A_ns[10] ), .ZN(n798) );
  INV_X1 U148 ( .A(\A_s[10] ), .ZN(n800) );
  OAI221_X1 U149 ( .B1(n703), .B2(n799), .C1(n694), .C2(n801), .A(n172), .ZN(
        O[13]) );
  INV_X1 U150 ( .A(\A_ns[11] ), .ZN(n799) );
  INV_X1 U151 ( .A(\A_s[11] ), .ZN(n801) );
  OAI221_X1 U152 ( .B1(n703), .B2(n802), .C1(n694), .C2(n804), .A(n171), .ZN(
        O[14]) );
  INV_X1 U153 ( .A(\A_ns[12] ), .ZN(n802) );
  INV_X1 U154 ( .A(\A_s[12] ), .ZN(n804) );
  OAI22_X1 U155 ( .A1(n164), .A2(n780), .B1(n165), .B2(n778), .ZN(O[1]) );
  OAI221_X1 U156 ( .B1(n701), .B2(n778), .C1(n695), .C2(n780), .A(n153), .ZN(
        O[2]) );
  AOI22_X1 U157 ( .A1(\A_ns[1] ), .A2(n688), .B1(\A_s[1] ), .B2(n681), .ZN(
        n153) );
  OAI221_X1 U158 ( .B1(n701), .B2(n779), .C1(n696), .C2(n781), .A(n142), .ZN(
        O[3]) );
  INV_X1 U159 ( .A(\A_ns[1] ), .ZN(n779) );
  INV_X1 U160 ( .A(\A_s[1] ), .ZN(n781) );
  OAI221_X1 U161 ( .B1(n700), .B2(n782), .C1(n697), .C2(n784), .A(n131), .ZN(
        O[4]) );
  INV_X1 U162 ( .A(\A_ns[2] ), .ZN(n782) );
  INV_X1 U163 ( .A(\A_s[2] ), .ZN(n784) );
  OAI221_X1 U164 ( .B1(n699), .B2(n783), .C1(n697), .C2(n785), .A(n122), .ZN(
        O[5]) );
  INV_X1 U165 ( .A(\A_ns[3] ), .ZN(n783) );
  INV_X1 U166 ( .A(\A_s[3] ), .ZN(n785) );
  OAI221_X1 U167 ( .B1(n699), .B2(n786), .C1(n698), .C2(n788), .A(n121), .ZN(
        O[6]) );
  INV_X1 U168 ( .A(\A_ns[4] ), .ZN(n786) );
  INV_X1 U169 ( .A(\A_s[4] ), .ZN(n788) );
  INV_X1 U170 ( .A(\A_s[0] ), .ZN(n780) );
  INV_X1 U171 ( .A(\A_ns[0] ), .ZN(n778) );
  AOI22_X1 U172 ( .A1(\A_ns[2] ), .A2(n689), .B1(\A_s[2] ), .B2(n682), .ZN(
        n142) );
  AOI22_X1 U173 ( .A1(\A_ns[3] ), .A2(n690), .B1(\A_s[3] ), .B2(n683), .ZN(
        n131) );
  AOI22_X1 U174 ( .A1(\A_ns[4] ), .A2(n691), .B1(\A_s[4] ), .B2(n684), .ZN(
        n122) );
  AOI22_X1 U175 ( .A1(\A_ns[5] ), .A2(n691), .B1(\A_s[5] ), .B2(n684), .ZN(
        n121) );
  AOI22_X1 U176 ( .A1(\A_ns[6] ), .A2(n691), .B1(\A_s[6] ), .B2(n684), .ZN(
        n120) );
  AOI22_X1 U177 ( .A1(\A_ns[7] ), .A2(n691), .B1(\A_s[7] ), .B2(n684), .ZN(
        n119) );
  AOI22_X1 U178 ( .A1(\A_ns[8] ), .A2(n691), .B1(\A_s[8] ), .B2(n684), .ZN(
        n118) );
  AOI22_X1 U179 ( .A1(\A_ns[9] ), .A2(n687), .B1(\A_s[9] ), .B2(n680), .ZN(
        n175) );
  AOI22_X1 U180 ( .A1(\A_ns[10] ), .A2(n687), .B1(\A_s[10] ), .B2(n680), .ZN(
        n174) );
  AOI22_X1 U181 ( .A1(\A_ns[11] ), .A2(n687), .B1(\A_s[11] ), .B2(n680), .ZN(
        n173) );
  AOI22_X1 U182 ( .A1(\A_ns[12] ), .A2(n687), .B1(\A_s[12] ), .B2(n680), .ZN(
        n172) );
  AOI22_X1 U183 ( .A1(\A_ns[13] ), .A2(n687), .B1(\A_s[13] ), .B2(n680), .ZN(
        n171) );
  AOI22_X1 U184 ( .A1(\A_ns[14] ), .A2(n687), .B1(\A_s[14] ), .B2(n680), .ZN(
        n170) );
  AOI22_X1 U185 ( .A1(\A_ns[15] ), .A2(n687), .B1(\A_s[15] ), .B2(n680), .ZN(
        n169) );
  AOI22_X1 U186 ( .A1(\A_ns[16] ), .A2(n687), .B1(\A_s[16] ), .B2(n680), .ZN(
        n168) );
  AOI22_X1 U187 ( .A1(\A_ns[17] ), .A2(n687), .B1(\A_s[17] ), .B2(n680), .ZN(
        n167) );
  AOI22_X1 U188 ( .A1(\A_ns[18] ), .A2(n687), .B1(\A_s[18] ), .B2(n680), .ZN(
        n166) );
  AOI22_X1 U189 ( .A1(\A_ns[19] ), .A2(n687), .B1(\A_s[19] ), .B2(n680), .ZN(
        n163) );
  AOI22_X1 U190 ( .A1(\A_ns[20] ), .A2(n687), .B1(\A_s[20] ), .B2(n680), .ZN(
        n162) );
  AOI22_X1 U191 ( .A1(\A_ns[21] ), .A2(n688), .B1(\A_s[21] ), .B2(n681), .ZN(
        n161) );
  AOI22_X1 U192 ( .A1(\A_ns[22] ), .A2(n688), .B1(\A_s[22] ), .B2(n681), .ZN(
        n160) );
  INV_X1 U193 ( .A(\A_s[20] ), .ZN(n820) );
  INV_X1 U194 ( .A(\A_s[21] ), .ZN(n821) );
  INV_X1 U195 ( .A(\A_ns[24] ), .ZN(n706) );
  INV_X1 U196 ( .A(\A_ns[25] ), .ZN(n707) );
  INV_X1 U197 ( .A(\A_ns[26] ), .ZN(n708) );
  INV_X1 U198 ( .A(\A_ns[27] ), .ZN(n709) );
  INV_X1 U199 ( .A(\A_ns[28] ), .ZN(n710) );
  INV_X1 U200 ( .A(\A_ns[29] ), .ZN(n711) );
  INV_X1 U201 ( .A(\A_ns[30] ), .ZN(n712) );
  INV_X1 U202 ( .A(\A_ns[31] ), .ZN(n713) );
  INV_X1 U203 ( .A(\A_ns[32] ), .ZN(n714) );
  INV_X1 U204 ( .A(\A_ns[33] ), .ZN(n715) );
  INV_X1 U205 ( .A(\A_ns[34] ), .ZN(n716) );
  INV_X1 U206 ( .A(\A_ns[35] ), .ZN(n717) );
  INV_X1 U207 ( .A(\A_ns[36] ), .ZN(n718) );
  INV_X1 U208 ( .A(\A_ns[37] ), .ZN(n719) );
  INV_X1 U209 ( .A(n721), .ZN(A_nso[40]) );
  INV_X1 U210 ( .A(A_ns[38]), .ZN(n721) );
  INV_X1 U211 ( .A(\A_ns[39] ), .ZN(n722) );
  INV_X1 U212 ( .A(\A_ns[40] ), .ZN(n723) );
  INV_X1 U213 ( .A(\A_ns[41] ), .ZN(n724) );
  INV_X1 U214 ( .A(\A_ns[42] ), .ZN(n725) );
  INV_X1 U215 ( .A(\A_ns[43] ), .ZN(n726) );
  INV_X1 U216 ( .A(\A_ns[44] ), .ZN(n727) );
  INV_X1 U217 ( .A(\A_ns[45] ), .ZN(n728) );
  INV_X1 U218 ( .A(\A_ns[46] ), .ZN(n729) );
  INV_X1 U219 ( .A(\A_ns[47] ), .ZN(n730) );
  INV_X1 U220 ( .A(\A_ns[48] ), .ZN(n731) );
  INV_X1 U221 ( .A(\A_ns[49] ), .ZN(n732) );
  INV_X1 U222 ( .A(\A_ns[50] ), .ZN(n733) );
  INV_X1 U223 ( .A(\A_ns[51] ), .ZN(n734) );
  INV_X1 U224 ( .A(\A_ns[52] ), .ZN(n735) );
  INV_X1 U225 ( .A(\A_ns[53] ), .ZN(n736) );
  INV_X1 U226 ( .A(\A_ns[54] ), .ZN(n737) );
  INV_X1 U227 ( .A(\A_ns[55] ), .ZN(n738) );
  INV_X1 U228 ( .A(\A_ns[23] ), .ZN(n739) );
  INV_X1 U229 ( .A(\A_s[23] ), .ZN(n740) );
  INV_X1 U230 ( .A(\A_s[24] ), .ZN(n741) );
  INV_X1 U231 ( .A(\A_s[25] ), .ZN(n742) );
  INV_X1 U232 ( .A(\A_s[26] ), .ZN(n743) );
  INV_X1 U235 ( .A(\A_s[27] ), .ZN(n744) );
  INV_X1 U236 ( .A(\A_s[28] ), .ZN(n745) );
  INV_X1 U237 ( .A(\A_s[29] ), .ZN(n746) );
  INV_X1 U238 ( .A(\A_s[30] ), .ZN(n747) );
  INV_X1 U239 ( .A(\A_s[31] ), .ZN(n748) );
  INV_X1 U240 ( .A(\A_s[32] ), .ZN(n749) );
  INV_X1 U241 ( .A(\A_s[33] ), .ZN(n750) );
  INV_X1 U242 ( .A(\A_s[34] ), .ZN(n751) );
  INV_X1 U243 ( .A(\A_s[35] ), .ZN(n752) );
  INV_X1 U244 ( .A(n754), .ZN(A_so[38]) );
  INV_X1 U245 ( .A(A_s[36]), .ZN(n754) );
  INV_X1 U246 ( .A(n756), .ZN(A_so[39]) );
  INV_X1 U247 ( .A(A_s[37]), .ZN(n756) );
  INV_X1 U248 ( .A(\A_s[38] ), .ZN(n757) );
  INV_X1 U249 ( .A(\A_s[39] ), .ZN(n758) );
  INV_X1 U250 ( .A(\A_s[40] ), .ZN(n759) );
  INV_X1 U251 ( .A(\A_s[41] ), .ZN(n760) );
  INV_X1 U252 ( .A(\A_s[42] ), .ZN(n761) );
  INV_X1 U253 ( .A(\A_s[43] ), .ZN(n762) );
  INV_X1 U254 ( .A(\A_s[44] ), .ZN(n763) );
  INV_X1 U255 ( .A(\A_s[45] ), .ZN(n764) );
  INV_X1 U256 ( .A(\A_s[46] ), .ZN(n765) );
  INV_X1 U257 ( .A(\A_s[47] ), .ZN(n766) );
  INV_X1 U258 ( .A(\A_s[48] ), .ZN(n767) );
  INV_X1 U259 ( .A(\A_s[49] ), .ZN(n768) );
  INV_X1 U260 ( .A(n770), .ZN(A_so[52]) );
  INV_X1 U261 ( .A(A_s[50]), .ZN(n770) );
  INV_X1 U262 ( .A(n772), .ZN(A_so[53]) );
  INV_X1 U263 ( .A(A_s[51]), .ZN(n772) );
  INV_X1 U264 ( .A(n774), .ZN(A_so[54]) );
  INV_X1 U265 ( .A(A_s[52]), .ZN(n774) );
  INV_X1 U266 ( .A(\A_s[53] ), .ZN(n775) );
  INV_X1 U267 ( .A(\A_s[54] ), .ZN(n776) );
  INV_X1 U268 ( .A(\A_s[55] ), .ZN(n777) );
endmodule


module BOOTHENC_NBIT60_i26 ( A_s, A_ns, B, O, A_so, A_nso );
  input [59:0] A_s;
  input [59:0] A_ns;
  input [59:0] B;
  output [59:0] O;
  output [59:0] A_so;
  output [59:0] A_nso;
  wire   \A_s[57] , \A_s[56] , \A_s[55] , \A_s[54] , \A_s[53] , \A_s[52] ,
         \A_s[51] , \A_s[50] , \A_s[49] , \A_s[48] , \A_s[47] , \A_s[46] ,
         \A_s[45] , \A_s[44] , \A_s[43] , \A_s[42] , \A_s[41] , \A_s[40] ,
         \A_s[39] , \A_s[38] , \A_s[37] , \A_s[36] , \A_s[35] , \A_s[34] ,
         \A_s[33] , \A_s[32] , \A_s[31] , \A_s[30] , \A_s[29] , \A_s[28] ,
         \A_s[27] , \A_s[26] , \A_s[25] , \A_s[24] , \A_s[23] , \A_s[22] ,
         \A_s[21] , \A_s[20] , \A_s[19] , \A_s[18] , \A_s[17] , \A_s[16] ,
         \A_s[15] , \A_s[14] , \A_s[13] , \A_s[12] , \A_s[11] , \A_s[10] ,
         \A_s[9] , \A_s[8] , \A_s[7] , \A_s[6] , \A_s[5] , \A_s[4] , \A_s[3] ,
         \A_s[2] , \A_s[1] , \A_s[0] , \A_ns[57] , \A_ns[56] , \A_ns[55] ,
         \A_ns[54] , \A_ns[53] , \A_ns[52] , \A_ns[51] , \A_ns[50] ,
         \A_ns[49] , \A_ns[48] , \A_ns[47] , \A_ns[46] , \A_ns[45] ,
         \A_ns[44] , \A_ns[43] , \A_ns[42] , \A_ns[41] , \A_ns[40] ,
         \A_ns[39] , \A_ns[38] , \A_ns[37] , \A_ns[36] , \A_ns[35] ,
         \A_ns[34] , \A_ns[33] , \A_ns[32] , \A_ns[31] , \A_ns[30] ,
         \A_ns[29] , \A_ns[28] , \A_ns[27] , \A_ns[26] , \A_ns[25] ,
         \A_ns[24] , \A_ns[23] , \A_ns[22] , \A_ns[21] , \A_ns[20] ,
         \A_ns[19] , \A_ns[18] , \A_ns[17] , \A_ns[16] , \A_ns[15] ,
         \A_ns[14] , \A_ns[13] , \A_ns[12] , \A_ns[11] , \A_ns[10] , \A_ns[9] ,
         \A_ns[8] , \A_ns[7] , \A_ns[6] , \A_ns[5] , \A_ns[4] , \A_ns[3] ,
         \A_ns[2] , \A_ns[1] , \A_ns[0] , n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843;
  assign A_nso[0] = 1'b0;
  assign A_nso[1] = 1'b0;
  assign A_so[0] = 1'b0;
  assign A_so[1] = 1'b0;
  assign O[0] = 1'b0;
  assign A_so[59] = \A_s[57] ;
  assign \A_s[57]  = A_s[57];
  assign A_so[58] = \A_s[56] ;
  assign \A_s[56]  = A_s[56];
  assign A_so[57] = \A_s[55] ;
  assign \A_s[55]  = A_s[55];
  assign A_so[56] = \A_s[54] ;
  assign \A_s[54]  = A_s[54];
  assign A_so[55] = \A_s[53] ;
  assign \A_s[53]  = A_s[53];
  assign A_so[54] = \A_s[52] ;
  assign \A_s[52]  = A_s[52];
  assign A_so[53] = \A_s[51] ;
  assign \A_s[51]  = A_s[51];
  assign A_so[52] = \A_s[50] ;
  assign \A_s[50]  = A_s[50];
  assign A_so[51] = \A_s[49] ;
  assign \A_s[49]  = A_s[49];
  assign A_so[50] = \A_s[48] ;
  assign \A_s[48]  = A_s[48];
  assign A_so[49] = \A_s[47] ;
  assign \A_s[47]  = A_s[47];
  assign A_so[48] = \A_s[46] ;
  assign \A_s[46]  = A_s[46];
  assign A_so[47] = \A_s[45] ;
  assign \A_s[45]  = A_s[45];
  assign A_so[46] = \A_s[44] ;
  assign \A_s[44]  = A_s[44];
  assign A_so[45] = \A_s[43] ;
  assign \A_s[43]  = A_s[43];
  assign A_so[44] = \A_s[42] ;
  assign \A_s[42]  = A_s[42];
  assign A_so[43] = \A_s[41] ;
  assign \A_s[41]  = A_s[41];
  assign A_so[42] = \A_s[40] ;
  assign \A_s[40]  = A_s[40];
  assign A_so[41] = \A_s[39] ;
  assign \A_s[39]  = A_s[39];
  assign A_so[40] = \A_s[38] ;
  assign \A_s[38]  = A_s[38];
  assign A_so[39] = \A_s[37] ;
  assign \A_s[37]  = A_s[37];
  assign A_so[38] = \A_s[36] ;
  assign \A_s[36]  = A_s[36];
  assign A_so[37] = \A_s[35] ;
  assign \A_s[35]  = A_s[35];
  assign A_so[36] = \A_s[34] ;
  assign \A_s[34]  = A_s[34];
  assign A_so[35] = \A_s[33] ;
  assign \A_s[33]  = A_s[33];
  assign A_so[34] = \A_s[32] ;
  assign \A_s[32]  = A_s[32];
  assign A_so[33] = \A_s[31] ;
  assign \A_s[31]  = A_s[31];
  assign A_so[32] = \A_s[30] ;
  assign \A_s[30]  = A_s[30];
  assign A_so[31] = \A_s[29] ;
  assign \A_s[29]  = A_s[29];
  assign A_so[30] = \A_s[28] ;
  assign \A_s[28]  = A_s[28];
  assign A_so[29] = \A_s[27] ;
  assign \A_s[27]  = A_s[27];
  assign A_so[28] = \A_s[26] ;
  assign \A_s[26]  = A_s[26];
  assign A_so[27] = \A_s[25] ;
  assign \A_s[25]  = A_s[25];
  assign A_so[26] = \A_s[24] ;
  assign \A_s[24]  = A_s[24];
  assign A_so[25] = \A_s[23] ;
  assign \A_s[23]  = A_s[23];
  assign A_so[24] = \A_s[22] ;
  assign \A_s[22]  = A_s[22];
  assign A_so[23] = \A_s[21] ;
  assign \A_s[21]  = A_s[21];
  assign A_so[22] = \A_s[20] ;
  assign \A_s[20]  = A_s[20];
  assign A_so[21] = \A_s[19] ;
  assign \A_s[19]  = A_s[19];
  assign A_so[20] = \A_s[18] ;
  assign \A_s[18]  = A_s[18];
  assign A_so[19] = \A_s[17] ;
  assign \A_s[17]  = A_s[17];
  assign A_so[18] = \A_s[16] ;
  assign \A_s[16]  = A_s[16];
  assign A_so[17] = \A_s[15] ;
  assign \A_s[15]  = A_s[15];
  assign A_so[16] = \A_s[14] ;
  assign \A_s[14]  = A_s[14];
  assign A_so[15] = \A_s[13] ;
  assign \A_s[13]  = A_s[13];
  assign A_so[14] = \A_s[12] ;
  assign \A_s[12]  = A_s[12];
  assign A_so[13] = \A_s[11] ;
  assign \A_s[11]  = A_s[11];
  assign A_so[12] = \A_s[10] ;
  assign \A_s[10]  = A_s[10];
  assign A_so[11] = \A_s[9] ;
  assign \A_s[9]  = A_s[9];
  assign A_so[10] = \A_s[8] ;
  assign \A_s[8]  = A_s[8];
  assign A_so[9] = \A_s[7] ;
  assign \A_s[7]  = A_s[7];
  assign A_so[8] = \A_s[6] ;
  assign \A_s[6]  = A_s[6];
  assign A_so[7] = \A_s[5] ;
  assign \A_s[5]  = A_s[5];
  assign A_so[6] = \A_s[4] ;
  assign \A_s[4]  = A_s[4];
  assign A_so[5] = \A_s[3] ;
  assign \A_s[3]  = A_s[3];
  assign A_so[4] = \A_s[2] ;
  assign \A_s[2]  = A_s[2];
  assign A_so[3] = \A_s[1] ;
  assign \A_s[1]  = A_s[1];
  assign A_so[2] = \A_s[0] ;
  assign \A_s[0]  = A_s[0];
  assign A_nso[59] = \A_ns[57] ;
  assign \A_ns[57]  = A_ns[57];
  assign A_nso[58] = \A_ns[56] ;
  assign \A_ns[56]  = A_ns[56];
  assign A_nso[57] = \A_ns[55] ;
  assign \A_ns[55]  = A_ns[55];
  assign A_nso[56] = \A_ns[54] ;
  assign \A_ns[54]  = A_ns[54];
  assign A_nso[55] = \A_ns[53] ;
  assign \A_ns[53]  = A_ns[53];
  assign A_nso[54] = \A_ns[52] ;
  assign \A_ns[52]  = A_ns[52];
  assign A_nso[53] = \A_ns[51] ;
  assign \A_ns[51]  = A_ns[51];
  assign A_nso[52] = \A_ns[50] ;
  assign \A_ns[50]  = A_ns[50];
  assign A_nso[51] = \A_ns[49] ;
  assign \A_ns[49]  = A_ns[49];
  assign A_nso[50] = \A_ns[48] ;
  assign \A_ns[48]  = A_ns[48];
  assign A_nso[49] = \A_ns[47] ;
  assign \A_ns[47]  = A_ns[47];
  assign A_nso[48] = \A_ns[46] ;
  assign \A_ns[46]  = A_ns[46];
  assign A_nso[47] = \A_ns[45] ;
  assign \A_ns[45]  = A_ns[45];
  assign A_nso[46] = \A_ns[44] ;
  assign \A_ns[44]  = A_ns[44];
  assign A_nso[45] = \A_ns[43] ;
  assign \A_ns[43]  = A_ns[43];
  assign A_nso[44] = \A_ns[42] ;
  assign \A_ns[42]  = A_ns[42];
  assign A_nso[43] = \A_ns[41] ;
  assign \A_ns[41]  = A_ns[41];
  assign A_nso[42] = \A_ns[40] ;
  assign \A_ns[40]  = A_ns[40];
  assign A_nso[41] = \A_ns[39] ;
  assign \A_ns[39]  = A_ns[39];
  assign A_nso[40] = \A_ns[38] ;
  assign \A_ns[38]  = A_ns[38];
  assign A_nso[39] = \A_ns[37] ;
  assign \A_ns[37]  = A_ns[37];
  assign A_nso[38] = \A_ns[36] ;
  assign \A_ns[36]  = A_ns[36];
  assign A_nso[37] = \A_ns[35] ;
  assign \A_ns[35]  = A_ns[35];
  assign A_nso[36] = \A_ns[34] ;
  assign \A_ns[34]  = A_ns[34];
  assign A_nso[35] = \A_ns[33] ;
  assign \A_ns[33]  = A_ns[33];
  assign A_nso[34] = \A_ns[32] ;
  assign \A_ns[32]  = A_ns[32];
  assign A_nso[33] = \A_ns[31] ;
  assign \A_ns[31]  = A_ns[31];
  assign A_nso[32] = \A_ns[30] ;
  assign \A_ns[30]  = A_ns[30];
  assign A_nso[31] = \A_ns[29] ;
  assign \A_ns[29]  = A_ns[29];
  assign A_nso[30] = \A_ns[28] ;
  assign \A_ns[28]  = A_ns[28];
  assign A_nso[29] = \A_ns[27] ;
  assign \A_ns[27]  = A_ns[27];
  assign A_nso[28] = \A_ns[26] ;
  assign \A_ns[26]  = A_ns[26];
  assign A_nso[27] = \A_ns[25] ;
  assign \A_ns[25]  = A_ns[25];
  assign A_nso[26] = \A_ns[24] ;
  assign \A_ns[24]  = A_ns[24];
  assign A_nso[25] = \A_ns[23] ;
  assign \A_ns[23]  = A_ns[23];
  assign A_nso[24] = \A_ns[22] ;
  assign \A_ns[22]  = A_ns[22];
  assign A_nso[23] = \A_ns[21] ;
  assign \A_ns[21]  = A_ns[21];
  assign A_nso[22] = \A_ns[20] ;
  assign \A_ns[20]  = A_ns[20];
  assign A_nso[21] = \A_ns[19] ;
  assign \A_ns[19]  = A_ns[19];
  assign A_nso[20] = \A_ns[18] ;
  assign \A_ns[18]  = A_ns[18];
  assign A_nso[19] = \A_ns[17] ;
  assign \A_ns[17]  = A_ns[17];
  assign A_nso[18] = \A_ns[16] ;
  assign \A_ns[16]  = A_ns[16];
  assign A_nso[17] = \A_ns[15] ;
  assign \A_ns[15]  = A_ns[15];
  assign A_nso[16] = \A_ns[14] ;
  assign \A_ns[14]  = A_ns[14];
  assign A_nso[15] = \A_ns[13] ;
  assign \A_ns[13]  = A_ns[13];
  assign A_nso[14] = \A_ns[12] ;
  assign \A_ns[12]  = A_ns[12];
  assign A_nso[13] = \A_ns[11] ;
  assign \A_ns[11]  = A_ns[11];
  assign A_nso[12] = \A_ns[10] ;
  assign \A_ns[10]  = A_ns[10];
  assign A_nso[11] = \A_ns[9] ;
  assign \A_ns[9]  = A_ns[9];
  assign A_nso[10] = \A_ns[8] ;
  assign \A_ns[8]  = A_ns[8];
  assign A_nso[9] = \A_ns[7] ;
  assign \A_ns[7]  = A_ns[7];
  assign A_nso[8] = \A_ns[6] ;
  assign \A_ns[6]  = A_ns[6];
  assign A_nso[7] = \A_ns[5] ;
  assign \A_ns[5]  = A_ns[5];
  assign A_nso[6] = \A_ns[4] ;
  assign \A_ns[4]  = A_ns[4];
  assign A_nso[5] = \A_ns[3] ;
  assign \A_ns[3]  = A_ns[3];
  assign A_nso[4] = \A_ns[2] ;
  assign \A_ns[2]  = A_ns[2];
  assign A_nso[3] = \A_ns[1] ;
  assign \A_ns[1]  = A_ns[1];
  assign A_nso[2] = \A_ns[0] ;
  assign \A_ns[0]  = A_ns[0];

  XOR2_X1 U241 ( .A(B[25]), .B(B[26]), .Z(n182) );
  NAND3_X1 U242 ( .A1(B[26]), .A2(n843), .A3(B[25]), .ZN(n121) );
  OAI221_X1 U2 ( .B1(n722), .B2(n734), .C1(n715), .C2(n768), .A(n151), .ZN(
        O[37]) );
  OAI221_X1 U3 ( .B1(n721), .B2(n740), .C1(n715), .C2(n774), .A(n144), .ZN(
        O[43]) );
  OAI221_X1 U4 ( .B1(n723), .B2(n757), .C1(n714), .C2(n758), .A(n162), .ZN(
        O[27]) );
  OAI221_X1 U5 ( .B1(n723), .B2(n725), .C1(n714), .C2(n759), .A(n161), .ZN(
        O[28]) );
  OAI221_X1 U6 ( .B1(n723), .B2(n727), .C1(n714), .C2(n761), .A(n158), .ZN(
        O[30]) );
  OAI221_X1 U7 ( .B1(n721), .B2(n741), .C1(n715), .C2(n775), .A(n143), .ZN(
        O[44]) );
  OAI221_X1 U8 ( .B1(n721), .B2(n749), .C1(n716), .C2(n783), .A(n134), .ZN(
        O[52]) );
  AOI22_X1 U9 ( .A1(\A_ns[26] ), .A2(n707), .B1(\A_s[26] ), .B2(n700), .ZN(
        n162) );
  AOI22_X1 U10 ( .A1(A_ns[58]), .A2(n710), .B1(A_s[58]), .B2(n703), .ZN(n127)
         );
  BUF_X1 U11 ( .A(n704), .Z(n707) );
  BUF_X1 U12 ( .A(n697), .Z(n700) );
  BUF_X1 U13 ( .A(n704), .Z(n708) );
  BUF_X1 U14 ( .A(n697), .Z(n701) );
  BUF_X1 U15 ( .A(n705), .Z(n709) );
  BUF_X1 U16 ( .A(n698), .Z(n702) );
  BUF_X1 U17 ( .A(n705), .Z(n710) );
  BUF_X1 U18 ( .A(n698), .Z(n703) );
  BUF_X1 U19 ( .A(n704), .Z(n706) );
  BUF_X1 U20 ( .A(n697), .Z(n699) );
  OAI221_X1 U21 ( .B1(n720), .B2(n756), .C1(n717), .C2(n790), .A(n127), .ZN(
        O[59]) );
  OAI221_X1 U22 ( .B1(n723), .B2(n726), .C1(n714), .C2(n760), .A(n160), .ZN(
        O[29]) );
  AOI22_X1 U23 ( .A1(\A_ns[28] ), .A2(n707), .B1(\A_s[28] ), .B2(n700), .ZN(
        n160) );
  AOI22_X1 U24 ( .A1(\A_ns[27] ), .A2(n707), .B1(\A_s[27] ), .B2(n700), .ZN(
        n161) );
  AOI22_X1 U25 ( .A1(\A_ns[29] ), .A2(n707), .B1(\A_s[29] ), .B2(n700), .ZN(
        n158) );
  OAI221_X1 U26 ( .B1(n722), .B2(n730), .C1(n714), .C2(n764), .A(n155), .ZN(
        O[33]) );
  AOI22_X1 U27 ( .A1(\A_ns[32] ), .A2(n708), .B1(\A_s[32] ), .B2(n701), .ZN(
        n155) );
  OAI221_X1 U28 ( .B1(n722), .B2(n732), .C1(n715), .C2(n766), .A(n153), .ZN(
        O[35]) );
  AOI22_X1 U29 ( .A1(\A_ns[34] ), .A2(n708), .B1(\A_s[34] ), .B2(n701), .ZN(
        n153) );
  OAI221_X1 U30 ( .B1(n722), .B2(n728), .C1(n714), .C2(n762), .A(n157), .ZN(
        O[31]) );
  AOI22_X1 U31 ( .A1(\A_ns[30] ), .A2(n707), .B1(\A_s[30] ), .B2(n700), .ZN(
        n157) );
  AOI22_X1 U32 ( .A1(\A_ns[36] ), .A2(n708), .B1(\A_s[36] ), .B2(n701), .ZN(
        n151) );
  OAI221_X1 U33 ( .B1(n722), .B2(n733), .C1(n715), .C2(n767), .A(n152), .ZN(
        O[36]) );
  AOI22_X1 U34 ( .A1(\A_ns[35] ), .A2(n708), .B1(\A_s[35] ), .B2(n701), .ZN(
        n152) );
  OAI221_X1 U35 ( .B1(n722), .B2(n729), .C1(n714), .C2(n763), .A(n156), .ZN(
        O[32]) );
  AOI22_X1 U36 ( .A1(\A_ns[31] ), .A2(n707), .B1(\A_s[31] ), .B2(n700), .ZN(
        n156) );
  OAI221_X1 U37 ( .B1(n722), .B2(n731), .C1(n714), .C2(n765), .A(n154), .ZN(
        O[34]) );
  AOI22_X1 U38 ( .A1(\A_ns[33] ), .A2(n708), .B1(\A_s[33] ), .B2(n701), .ZN(
        n154) );
  OAI221_X1 U39 ( .B1(n722), .B2(n735), .C1(n715), .C2(n769), .A(n150), .ZN(
        O[38]) );
  AOI22_X1 U40 ( .A1(\A_ns[37] ), .A2(n708), .B1(\A_s[37] ), .B2(n701), .ZN(
        n150) );
  BUF_X1 U41 ( .A(n841), .Z(n697) );
  BUF_X1 U42 ( .A(n842), .Z(n704) );
  OAI221_X1 U43 ( .B1(n722), .B2(n736), .C1(n715), .C2(n770), .A(n149), .ZN(
        O[39]) );
  AOI22_X1 U44 ( .A1(\A_ns[38] ), .A2(n708), .B1(\A_s[38] ), .B2(n701), .ZN(
        n149) );
  AOI22_X1 U45 ( .A1(\A_ns[42] ), .A2(n708), .B1(\A_s[42] ), .B2(n701), .ZN(
        n144) );
  OAI221_X1 U46 ( .B1(n721), .B2(n746), .C1(n716), .C2(n780), .A(n138), .ZN(
        O[49]) );
  AOI22_X1 U47 ( .A1(\A_ns[48] ), .A2(n709), .B1(\A_s[48] ), .B2(n702), .ZN(
        n138) );
  OAI221_X1 U48 ( .B1(n722), .B2(n738), .C1(n715), .C2(n772), .A(n146), .ZN(
        O[41]) );
  AOI22_X1 U49 ( .A1(\A_ns[40] ), .A2(n708), .B1(\A_s[40] ), .B2(n701), .ZN(
        n146) );
  OAI221_X1 U50 ( .B1(n721), .B2(n739), .C1(n715), .C2(n773), .A(n145), .ZN(
        O[42]) );
  AOI22_X1 U51 ( .A1(\A_ns[41] ), .A2(n708), .B1(\A_s[41] ), .B2(n701), .ZN(
        n145) );
  OAI221_X1 U52 ( .B1(n721), .B2(n743), .C1(n715), .C2(n777), .A(n141), .ZN(
        O[46]) );
  AOI22_X1 U53 ( .A1(\A_ns[45] ), .A2(n709), .B1(\A_s[45] ), .B2(n702), .ZN(
        n141) );
  OAI221_X1 U54 ( .B1(n722), .B2(n737), .C1(n715), .C2(n771), .A(n147), .ZN(
        O[40]) );
  AOI22_X1 U55 ( .A1(\A_ns[39] ), .A2(n708), .B1(\A_s[39] ), .B2(n701), .ZN(
        n147) );
  OAI221_X1 U56 ( .B1(n721), .B2(n745), .C1(n716), .C2(n779), .A(n139), .ZN(
        O[48]) );
  AOI22_X1 U57 ( .A1(\A_ns[47] ), .A2(n709), .B1(\A_s[47] ), .B2(n702), .ZN(
        n139) );
  OAI221_X1 U58 ( .B1(n721), .B2(n747), .C1(n716), .C2(n781), .A(n136), .ZN(
        O[50]) );
  AOI22_X1 U59 ( .A1(\A_ns[49] ), .A2(n709), .B1(\A_s[49] ), .B2(n702), .ZN(
        n136) );
  AOI22_X1 U60 ( .A1(\A_ns[51] ), .A2(n709), .B1(\A_s[51] ), .B2(n702), .ZN(
        n134) );
  AOI22_X1 U61 ( .A1(\A_ns[43] ), .A2(n709), .B1(\A_s[43] ), .B2(n702), .ZN(
        n143) );
  OAI221_X1 U62 ( .B1(n721), .B2(n742), .C1(n715), .C2(n776), .A(n142), .ZN(
        O[45]) );
  AOI22_X1 U63 ( .A1(\A_ns[44] ), .A2(n709), .B1(\A_s[44] ), .B2(n702), .ZN(
        n142) );
  OAI221_X1 U64 ( .B1(n721), .B2(n744), .C1(n716), .C2(n778), .A(n140), .ZN(
        O[47]) );
  AOI22_X1 U65 ( .A1(\A_ns[46] ), .A2(n709), .B1(\A_s[46] ), .B2(n702), .ZN(
        n140) );
  OAI221_X1 U66 ( .B1(n721), .B2(n748), .C1(n716), .C2(n782), .A(n135), .ZN(
        O[51]) );
  AOI22_X1 U67 ( .A1(\A_ns[50] ), .A2(n709), .B1(\A_s[50] ), .B2(n702), .ZN(
        n135) );
  OAI221_X1 U68 ( .B1(n720), .B2(n750), .C1(n716), .C2(n784), .A(n133), .ZN(
        O[53]) );
  AOI22_X1 U69 ( .A1(\A_ns[52] ), .A2(n709), .B1(\A_s[52] ), .B2(n702), .ZN(
        n133) );
  OAI221_X1 U70 ( .B1(n720), .B2(n755), .C1(n716), .C2(n789), .A(n128), .ZN(
        O[58]) );
  AOI22_X1 U71 ( .A1(\A_ns[57] ), .A2(n710), .B1(\A_s[57] ), .B2(n703), .ZN(
        n128) );
  OAI221_X1 U72 ( .B1(n720), .B2(n751), .C1(n716), .C2(n785), .A(n132), .ZN(
        O[54]) );
  AOI22_X1 U73 ( .A1(\A_ns[53] ), .A2(n709), .B1(\A_s[53] ), .B2(n702), .ZN(
        n132) );
  OAI221_X1 U74 ( .B1(n720), .B2(n752), .C1(n716), .C2(n786), .A(n131), .ZN(
        O[55]) );
  AOI22_X1 U75 ( .A1(\A_ns[54] ), .A2(n710), .B1(\A_s[54] ), .B2(n703), .ZN(
        n131) );
  OAI221_X1 U76 ( .B1(n720), .B2(n754), .C1(n716), .C2(n788), .A(n129), .ZN(
        O[57]) );
  AOI22_X1 U77 ( .A1(\A_ns[56] ), .A2(n710), .B1(\A_s[56] ), .B2(n703), .ZN(
        n129) );
  OAI221_X1 U78 ( .B1(n720), .B2(n753), .C1(n716), .C2(n787), .A(n130), .ZN(
        O[56]) );
  AOI22_X1 U79 ( .A1(\A_ns[55] ), .A2(n710), .B1(\A_s[55] ), .B2(n703), .ZN(
        n130) );
  BUF_X1 U80 ( .A(n841), .Z(n698) );
  BUF_X1 U81 ( .A(n842), .Z(n705) );
  BUF_X1 U82 ( .A(n719), .Z(n723) );
  BUF_X1 U83 ( .A(n711), .Z(n714) );
  INV_X1 U84 ( .A(n170), .ZN(n841) );
  INV_X1 U85 ( .A(n171), .ZN(n842) );
  BUF_X1 U86 ( .A(n718), .Z(n722) );
  BUF_X1 U87 ( .A(n711), .Z(n715) );
  BUF_X1 U88 ( .A(n718), .Z(n721) );
  BUF_X1 U89 ( .A(n718), .Z(n720) );
  BUF_X1 U90 ( .A(n712), .Z(n716) );
  BUF_X1 U91 ( .A(n712), .Z(n717) );
  BUF_X1 U92 ( .A(n711), .Z(n713) );
  BUF_X1 U93 ( .A(n719), .Z(n724) );
  NAND2_X1 U94 ( .A1(n182), .A2(n843), .ZN(n170) );
  NAND2_X1 U95 ( .A1(n182), .A2(n170), .ZN(n171) );
  BUF_X1 U96 ( .A(n121), .Z(n711) );
  BUF_X1 U97 ( .A(n120), .Z(n719) );
  BUF_X1 U98 ( .A(n120), .Z(n718) );
  BUF_X1 U99 ( .A(n121), .Z(n712) );
  OAI221_X1 U100 ( .B1(n723), .B2(n839), .C1(n714), .C2(n840), .A(n163), .ZN(
        O[26]) );
  INV_X1 U101 ( .A(\A_ns[24] ), .ZN(n839) );
  INV_X1 U102 ( .A(\A_s[24] ), .ZN(n840) );
  AOI22_X1 U103 ( .A1(\A_ns[25] ), .A2(n707), .B1(\A_s[25] ), .B2(n700), .ZN(
        n163) );
  OAI221_X1 U104 ( .B1(n723), .B2(n828), .C1(n713), .C2(n830), .A(n168), .ZN(
        O[21]) );
  INV_X1 U105 ( .A(\A_ns[19] ), .ZN(n828) );
  INV_X1 U106 ( .A(\A_s[19] ), .ZN(n830) );
  OAI221_X1 U107 ( .B1(n723), .B2(n831), .C1(n713), .C2(n833), .A(n167), .ZN(
        O[22]) );
  INV_X1 U108 ( .A(\A_ns[20] ), .ZN(n831) );
  INV_X1 U109 ( .A(\A_s[20] ), .ZN(n833) );
  OAI221_X1 U110 ( .B1(n723), .B2(n832), .C1(n714), .C2(n834), .A(n166), .ZN(
        O[23]) );
  INV_X1 U111 ( .A(\A_ns[21] ), .ZN(n832) );
  INV_X1 U112 ( .A(\A_s[21] ), .ZN(n834) );
  OAI221_X1 U113 ( .B1(n723), .B2(n835), .C1(n714), .C2(n837), .A(n165), .ZN(
        O[24]) );
  INV_X1 U114 ( .A(\A_ns[22] ), .ZN(n835) );
  OAI221_X1 U115 ( .B1(n723), .B2(n836), .C1(n714), .C2(n838), .A(n164), .ZN(
        O[25]) );
  INV_X1 U116 ( .A(\A_ns[23] ), .ZN(n836) );
  INV_X1 U117 ( .A(B[27]), .ZN(n843) );
  OR3_X1 U118 ( .A1(B[25]), .A2(B[26]), .A3(n843), .ZN(n120) );
  OAI221_X1 U119 ( .B1(n724), .B2(n816), .C1(n713), .C2(n818), .A(n176), .ZN(
        O[15]) );
  INV_X1 U120 ( .A(\A_ns[13] ), .ZN(n816) );
  INV_X1 U121 ( .A(\A_s[13] ), .ZN(n818) );
  OAI221_X1 U122 ( .B1(n724), .B2(n819), .C1(n713), .C2(n821), .A(n175), .ZN(
        O[16]) );
  INV_X1 U123 ( .A(\A_ns[14] ), .ZN(n819) );
  INV_X1 U124 ( .A(\A_s[14] ), .ZN(n821) );
  OAI221_X1 U125 ( .B1(n724), .B2(n820), .C1(n713), .C2(n822), .A(n174), .ZN(
        O[17]) );
  INV_X1 U126 ( .A(\A_ns[15] ), .ZN(n820) );
  INV_X1 U127 ( .A(\A_s[15] ), .ZN(n822) );
  OAI221_X1 U128 ( .B1(n724), .B2(n823), .C1(n713), .C2(n825), .A(n173), .ZN(
        O[18]) );
  INV_X1 U129 ( .A(\A_ns[16] ), .ZN(n823) );
  INV_X1 U130 ( .A(\A_s[16] ), .ZN(n825) );
  OAI221_X1 U131 ( .B1(n724), .B2(n824), .C1(n713), .C2(n826), .A(n172), .ZN(
        O[19]) );
  INV_X1 U132 ( .A(\A_ns[17] ), .ZN(n824) );
  INV_X1 U133 ( .A(\A_s[17] ), .ZN(n826) );
  OAI221_X1 U134 ( .B1(n723), .B2(n827), .C1(n713), .C2(n829), .A(n169), .ZN(
        O[20]) );
  INV_X1 U135 ( .A(\A_ns[18] ), .ZN(n827) );
  INV_X1 U136 ( .A(\A_s[18] ), .ZN(n829) );
  OAI221_X1 U137 ( .B1(n720), .B2(n800), .C1(n717), .C2(n802), .A(n124), .ZN(
        O[7]) );
  INV_X1 U138 ( .A(\A_ns[5] ), .ZN(n800) );
  INV_X1 U139 ( .A(\A_s[5] ), .ZN(n802) );
  OAI221_X1 U140 ( .B1(n720), .B2(n803), .C1(n717), .C2(n805), .A(n123), .ZN(
        O[8]) );
  INV_X1 U141 ( .A(\A_ns[6] ), .ZN(n803) );
  INV_X1 U142 ( .A(\A_s[6] ), .ZN(n805) );
  OAI221_X1 U143 ( .B1(n720), .B2(n804), .C1(n717), .C2(n806), .A(n122), .ZN(
        O[9]) );
  INV_X1 U144 ( .A(\A_ns[7] ), .ZN(n804) );
  INV_X1 U145 ( .A(\A_s[7] ), .ZN(n806) );
  OAI221_X1 U146 ( .B1(n807), .B2(n724), .C1(n809), .C2(n713), .A(n181), .ZN(
        O[10]) );
  INV_X1 U147 ( .A(\A_s[8] ), .ZN(n809) );
  INV_X1 U148 ( .A(\A_ns[8] ), .ZN(n807) );
  OAI221_X1 U149 ( .B1(n724), .B2(n808), .C1(n713), .C2(n810), .A(n180), .ZN(
        O[11]) );
  INV_X1 U150 ( .A(\A_ns[9] ), .ZN(n808) );
  INV_X1 U151 ( .A(\A_s[9] ), .ZN(n810) );
  OAI221_X1 U152 ( .B1(n724), .B2(n811), .C1(n713), .C2(n813), .A(n179), .ZN(
        O[12]) );
  INV_X1 U153 ( .A(\A_ns[10] ), .ZN(n811) );
  INV_X1 U154 ( .A(\A_s[10] ), .ZN(n813) );
  OAI221_X1 U155 ( .B1(n724), .B2(n812), .C1(n713), .C2(n814), .A(n178), .ZN(
        O[13]) );
  INV_X1 U156 ( .A(\A_ns[11] ), .ZN(n812) );
  INV_X1 U157 ( .A(\A_s[11] ), .ZN(n814) );
  OAI221_X1 U158 ( .B1(n724), .B2(n815), .C1(n713), .C2(n817), .A(n177), .ZN(
        O[14]) );
  INV_X1 U159 ( .A(\A_ns[12] ), .ZN(n815) );
  INV_X1 U160 ( .A(\A_s[12] ), .ZN(n817) );
  OAI22_X1 U161 ( .A1(n170), .A2(n793), .B1(n171), .B2(n791), .ZN(O[1]) );
  OAI221_X1 U162 ( .B1(n723), .B2(n791), .C1(n714), .C2(n793), .A(n159), .ZN(
        O[2]) );
  AOI22_X1 U163 ( .A1(\A_ns[1] ), .A2(n707), .B1(\A_s[1] ), .B2(n700), .ZN(
        n159) );
  OAI221_X1 U164 ( .B1(n722), .B2(n792), .C1(n715), .C2(n794), .A(n148), .ZN(
        O[3]) );
  INV_X1 U165 ( .A(\A_ns[1] ), .ZN(n792) );
  INV_X1 U166 ( .A(\A_s[1] ), .ZN(n794) );
  OAI221_X1 U167 ( .B1(n721), .B2(n795), .C1(n716), .C2(n797), .A(n137), .ZN(
        O[4]) );
  INV_X1 U168 ( .A(\A_ns[2] ), .ZN(n795) );
  INV_X1 U169 ( .A(\A_s[2] ), .ZN(n797) );
  OAI221_X1 U170 ( .B1(n720), .B2(n796), .C1(n717), .C2(n798), .A(n126), .ZN(
        O[5]) );
  INV_X1 U171 ( .A(\A_ns[3] ), .ZN(n796) );
  INV_X1 U172 ( .A(\A_s[3] ), .ZN(n798) );
  OAI221_X1 U173 ( .B1(n720), .B2(n799), .C1(n717), .C2(n801), .A(n125), .ZN(
        O[6]) );
  INV_X1 U174 ( .A(\A_ns[4] ), .ZN(n799) );
  INV_X1 U175 ( .A(\A_s[4] ), .ZN(n801) );
  INV_X1 U176 ( .A(\A_s[0] ), .ZN(n793) );
  INV_X1 U177 ( .A(\A_ns[0] ), .ZN(n791) );
  AOI22_X1 U178 ( .A1(\A_ns[2] ), .A2(n708), .B1(\A_s[2] ), .B2(n701), .ZN(
        n148) );
  AOI22_X1 U179 ( .A1(\A_ns[3] ), .A2(n709), .B1(\A_s[3] ), .B2(n702), .ZN(
        n137) );
  AOI22_X1 U180 ( .A1(\A_ns[4] ), .A2(n710), .B1(\A_s[4] ), .B2(n703), .ZN(
        n126) );
  AOI22_X1 U181 ( .A1(\A_ns[5] ), .A2(n710), .B1(\A_s[5] ), .B2(n703), .ZN(
        n125) );
  AOI22_X1 U182 ( .A1(\A_ns[6] ), .A2(n710), .B1(\A_s[6] ), .B2(n703), .ZN(
        n124) );
  AOI22_X1 U183 ( .A1(\A_ns[7] ), .A2(n710), .B1(\A_s[7] ), .B2(n703), .ZN(
        n123) );
  AOI22_X1 U184 ( .A1(\A_ns[8] ), .A2(n710), .B1(\A_s[8] ), .B2(n703), .ZN(
        n122) );
  AOI22_X1 U185 ( .A1(\A_ns[9] ), .A2(n706), .B1(\A_s[9] ), .B2(n699), .ZN(
        n181) );
  AOI22_X1 U186 ( .A1(\A_ns[10] ), .A2(n706), .B1(\A_s[10] ), .B2(n699), .ZN(
        n180) );
  AOI22_X1 U187 ( .A1(\A_ns[11] ), .A2(n706), .B1(\A_s[11] ), .B2(n699), .ZN(
        n179) );
  AOI22_X1 U188 ( .A1(\A_ns[12] ), .A2(n706), .B1(\A_s[12] ), .B2(n699), .ZN(
        n178) );
  AOI22_X1 U189 ( .A1(\A_ns[13] ), .A2(n706), .B1(\A_s[13] ), .B2(n699), .ZN(
        n177) );
  AOI22_X1 U190 ( .A1(\A_ns[14] ), .A2(n706), .B1(\A_s[14] ), .B2(n699), .ZN(
        n176) );
  AOI22_X1 U191 ( .A1(\A_ns[15] ), .A2(n706), .B1(\A_s[15] ), .B2(n699), .ZN(
        n175) );
  AOI22_X1 U192 ( .A1(\A_ns[16] ), .A2(n706), .B1(\A_s[16] ), .B2(n699), .ZN(
        n174) );
  AOI22_X1 U193 ( .A1(\A_ns[17] ), .A2(n706), .B1(\A_s[17] ), .B2(n699), .ZN(
        n173) );
  AOI22_X1 U194 ( .A1(\A_ns[18] ), .A2(n706), .B1(\A_s[18] ), .B2(n699), .ZN(
        n172) );
  AOI22_X1 U195 ( .A1(\A_ns[19] ), .A2(n706), .B1(\A_s[19] ), .B2(n699), .ZN(
        n169) );
  AOI22_X1 U196 ( .A1(\A_ns[20] ), .A2(n706), .B1(\A_s[20] ), .B2(n699), .ZN(
        n168) );
  AOI22_X1 U197 ( .A1(\A_ns[21] ), .A2(n707), .B1(\A_s[21] ), .B2(n700), .ZN(
        n167) );
  AOI22_X1 U198 ( .A1(\A_ns[22] ), .A2(n707), .B1(\A_s[22] ), .B2(n700), .ZN(
        n166) );
  AOI22_X1 U199 ( .A1(\A_ns[23] ), .A2(n707), .B1(\A_s[23] ), .B2(n700), .ZN(
        n165) );
  AOI22_X1 U200 ( .A1(\A_ns[24] ), .A2(n707), .B1(\A_s[24] ), .B2(n700), .ZN(
        n164) );
  INV_X1 U201 ( .A(\A_s[22] ), .ZN(n837) );
  INV_X1 U202 ( .A(\A_s[23] ), .ZN(n838) );
  INV_X1 U203 ( .A(\A_ns[26] ), .ZN(n725) );
  INV_X1 U204 ( .A(\A_ns[27] ), .ZN(n726) );
  INV_X1 U205 ( .A(\A_ns[28] ), .ZN(n727) );
  INV_X1 U206 ( .A(\A_ns[29] ), .ZN(n728) );
  INV_X1 U207 ( .A(\A_ns[30] ), .ZN(n729) );
  INV_X1 U208 ( .A(\A_ns[31] ), .ZN(n730) );
  INV_X1 U209 ( .A(\A_ns[32] ), .ZN(n731) );
  INV_X1 U210 ( .A(\A_ns[33] ), .ZN(n732) );
  INV_X1 U211 ( .A(\A_ns[34] ), .ZN(n733) );
  INV_X1 U212 ( .A(\A_ns[35] ), .ZN(n734) );
  INV_X1 U213 ( .A(\A_ns[36] ), .ZN(n735) );
  INV_X1 U214 ( .A(\A_ns[37] ), .ZN(n736) );
  INV_X1 U215 ( .A(\A_ns[38] ), .ZN(n737) );
  INV_X1 U216 ( .A(\A_ns[39] ), .ZN(n738) );
  INV_X1 U217 ( .A(\A_ns[40] ), .ZN(n739) );
  INV_X1 U218 ( .A(\A_ns[41] ), .ZN(n740) );
  INV_X1 U219 ( .A(\A_ns[42] ), .ZN(n741) );
  INV_X1 U220 ( .A(\A_ns[43] ), .ZN(n742) );
  INV_X1 U221 ( .A(\A_ns[44] ), .ZN(n743) );
  INV_X1 U222 ( .A(\A_ns[45] ), .ZN(n744) );
  INV_X1 U223 ( .A(\A_ns[46] ), .ZN(n745) );
  INV_X1 U224 ( .A(\A_ns[47] ), .ZN(n746) );
  INV_X1 U225 ( .A(\A_ns[48] ), .ZN(n747) );
  INV_X1 U226 ( .A(\A_ns[49] ), .ZN(n748) );
  INV_X1 U227 ( .A(\A_ns[50] ), .ZN(n749) );
  INV_X1 U228 ( .A(\A_ns[51] ), .ZN(n750) );
  INV_X1 U229 ( .A(\A_ns[52] ), .ZN(n751) );
  INV_X1 U230 ( .A(\A_ns[53] ), .ZN(n752) );
  INV_X1 U231 ( .A(\A_ns[54] ), .ZN(n753) );
  INV_X1 U232 ( .A(\A_ns[55] ), .ZN(n754) );
  INV_X1 U233 ( .A(\A_ns[56] ), .ZN(n755) );
  INV_X1 U234 ( .A(\A_ns[57] ), .ZN(n756) );
  INV_X1 U235 ( .A(\A_ns[25] ), .ZN(n757) );
  INV_X1 U236 ( .A(\A_s[25] ), .ZN(n758) );
  INV_X1 U237 ( .A(\A_s[26] ), .ZN(n759) );
  INV_X1 U238 ( .A(\A_s[27] ), .ZN(n760) );
  INV_X1 U239 ( .A(\A_s[28] ), .ZN(n761) );
  INV_X1 U240 ( .A(\A_s[29] ), .ZN(n762) );
  INV_X1 U243 ( .A(\A_s[30] ), .ZN(n763) );
  INV_X1 U244 ( .A(\A_s[31] ), .ZN(n764) );
  INV_X1 U245 ( .A(\A_s[32] ), .ZN(n765) );
  INV_X1 U246 ( .A(\A_s[33] ), .ZN(n766) );
  INV_X1 U247 ( .A(\A_s[34] ), .ZN(n767) );
  INV_X1 U248 ( .A(\A_s[35] ), .ZN(n768) );
  INV_X1 U249 ( .A(\A_s[36] ), .ZN(n769) );
  INV_X1 U250 ( .A(\A_s[37] ), .ZN(n770) );
  INV_X1 U251 ( .A(\A_s[38] ), .ZN(n771) );
  INV_X1 U252 ( .A(\A_s[39] ), .ZN(n772) );
  INV_X1 U253 ( .A(\A_s[40] ), .ZN(n773) );
  INV_X1 U254 ( .A(\A_s[41] ), .ZN(n774) );
  INV_X1 U255 ( .A(\A_s[42] ), .ZN(n775) );
  INV_X1 U256 ( .A(\A_s[43] ), .ZN(n776) );
  INV_X1 U257 ( .A(\A_s[44] ), .ZN(n777) );
  INV_X1 U258 ( .A(\A_s[45] ), .ZN(n778) );
  INV_X1 U259 ( .A(\A_s[46] ), .ZN(n779) );
  INV_X1 U260 ( .A(\A_s[47] ), .ZN(n780) );
  INV_X1 U261 ( .A(\A_s[48] ), .ZN(n781) );
  INV_X1 U262 ( .A(\A_s[49] ), .ZN(n782) );
  INV_X1 U263 ( .A(\A_s[50] ), .ZN(n783) );
  INV_X1 U264 ( .A(\A_s[51] ), .ZN(n784) );
  INV_X1 U265 ( .A(\A_s[52] ), .ZN(n785) );
  INV_X1 U266 ( .A(\A_s[53] ), .ZN(n786) );
  INV_X1 U267 ( .A(\A_s[54] ), .ZN(n787) );
  INV_X1 U268 ( .A(\A_s[55] ), .ZN(n788) );
  INV_X1 U269 ( .A(\A_s[56] ), .ZN(n789) );
  INV_X1 U270 ( .A(\A_s[57] ), .ZN(n790) );
endmodule


module BOOTHENC_NBIT62_i28 ( A_s, A_ns, B, O, A_so, A_nso );
  input [61:0] A_s;
  input [61:0] A_ns;
  input [61:0] B;
  output [61:0] O;
  output [61:0] A_so;
  output [61:0] A_nso;
  wire   \A_s[59] , \A_s[58] , \A_s[57] , \A_s[56] , \A_s[55] , \A_s[54] ,
         \A_s[53] , \A_s[52] , \A_s[51] , \A_s[50] , \A_s[49] , \A_s[48] ,
         \A_s[47] , \A_s[46] , \A_s[45] , \A_s[44] , \A_s[43] , \A_s[42] ,
         \A_s[41] , \A_s[40] , \A_s[39] , \A_s[38] , \A_s[37] , \A_s[36] ,
         \A_s[35] , \A_s[34] , \A_s[33] , \A_s[32] , \A_s[31] , \A_s[30] ,
         \A_s[29] , \A_s[28] , \A_s[27] , \A_s[26] , \A_s[25] , \A_s[24] ,
         \A_s[23] , \A_s[22] , \A_s[21] , \A_s[20] , \A_s[19] , \A_s[18] ,
         \A_s[17] , \A_s[16] , \A_s[15] , \A_s[14] , \A_s[13] , \A_s[12] ,
         \A_s[11] , \A_s[10] , \A_s[9] , \A_s[8] , \A_s[7] , \A_s[6] ,
         \A_s[5] , \A_s[4] , \A_s[3] , \A_s[2] , \A_s[1] , \A_s[0] ,
         \A_ns[59] , \A_ns[58] , \A_ns[57] , \A_ns[56] , \A_ns[55] ,
         \A_ns[54] , \A_ns[53] , \A_ns[52] , \A_ns[51] , \A_ns[50] ,
         \A_ns[49] , \A_ns[48] , \A_ns[47] , \A_ns[46] , \A_ns[45] ,
         \A_ns[44] , \A_ns[43] , \A_ns[42] , \A_ns[41] , \A_ns[40] ,
         \A_ns[39] , \A_ns[38] , \A_ns[37] , \A_ns[36] , \A_ns[35] ,
         \A_ns[34] , \A_ns[33] , \A_ns[32] , \A_ns[31] , \A_ns[30] ,
         \A_ns[29] , \A_ns[28] , \A_ns[27] , \A_ns[26] , \A_ns[25] ,
         \A_ns[24] , \A_ns[23] , \A_ns[22] , \A_ns[21] , \A_ns[20] ,
         \A_ns[19] , \A_ns[18] , \A_ns[17] , \A_ns[16] , \A_ns[15] ,
         \A_ns[14] , \A_ns[13] , \A_ns[12] , \A_ns[11] , \A_ns[10] , \A_ns[9] ,
         \A_ns[8] , \A_ns[7] , \A_ns[6] , \A_ns[5] , \A_ns[4] , \A_ns[3] ,
         \A_ns[2] , \A_ns[1] , \A_ns[0] , n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869;
  assign A_nso[0] = 1'b0;
  assign A_nso[1] = 1'b0;
  assign A_so[0] = 1'b0;
  assign A_so[1] = 1'b0;
  assign O[0] = 1'b0;
  assign A_so[61] = \A_s[59] ;
  assign \A_s[59]  = A_s[59];
  assign A_so[60] = \A_s[58] ;
  assign \A_s[58]  = A_s[58];
  assign A_so[59] = \A_s[57] ;
  assign \A_s[57]  = A_s[57];
  assign A_so[58] = \A_s[56] ;
  assign \A_s[56]  = A_s[56];
  assign A_so[57] = \A_s[55] ;
  assign \A_s[55]  = A_s[55];
  assign A_so[56] = \A_s[54] ;
  assign \A_s[54]  = A_s[54];
  assign A_so[55] = \A_s[53] ;
  assign \A_s[53]  = A_s[53];
  assign A_so[54] = \A_s[52] ;
  assign \A_s[52]  = A_s[52];
  assign A_so[53] = \A_s[51] ;
  assign \A_s[51]  = A_s[51];
  assign A_so[52] = \A_s[50] ;
  assign \A_s[50]  = A_s[50];
  assign A_so[51] = \A_s[49] ;
  assign \A_s[49]  = A_s[49];
  assign A_so[50] = \A_s[48] ;
  assign \A_s[48]  = A_s[48];
  assign A_so[49] = \A_s[47] ;
  assign \A_s[47]  = A_s[47];
  assign A_so[48] = \A_s[46] ;
  assign \A_s[46]  = A_s[46];
  assign A_so[47] = \A_s[45] ;
  assign \A_s[45]  = A_s[45];
  assign A_so[46] = \A_s[44] ;
  assign \A_s[44]  = A_s[44];
  assign A_so[45] = \A_s[43] ;
  assign \A_s[43]  = A_s[43];
  assign A_so[44] = \A_s[42] ;
  assign \A_s[42]  = A_s[42];
  assign A_so[43] = \A_s[41] ;
  assign \A_s[41]  = A_s[41];
  assign A_so[42] = \A_s[40] ;
  assign \A_s[40]  = A_s[40];
  assign A_so[41] = \A_s[39] ;
  assign \A_s[39]  = A_s[39];
  assign A_so[40] = \A_s[38] ;
  assign \A_s[38]  = A_s[38];
  assign A_so[39] = \A_s[37] ;
  assign \A_s[37]  = A_s[37];
  assign A_so[38] = \A_s[36] ;
  assign \A_s[36]  = A_s[36];
  assign A_so[37] = \A_s[35] ;
  assign \A_s[35]  = A_s[35];
  assign A_so[36] = \A_s[34] ;
  assign \A_s[34]  = A_s[34];
  assign A_so[35] = \A_s[33] ;
  assign \A_s[33]  = A_s[33];
  assign A_so[34] = \A_s[32] ;
  assign \A_s[32]  = A_s[32];
  assign A_so[33] = \A_s[31] ;
  assign \A_s[31]  = A_s[31];
  assign A_so[32] = \A_s[30] ;
  assign \A_s[30]  = A_s[30];
  assign A_so[31] = \A_s[29] ;
  assign \A_s[29]  = A_s[29];
  assign A_so[30] = \A_s[28] ;
  assign \A_s[28]  = A_s[28];
  assign A_so[29] = \A_s[27] ;
  assign \A_s[27]  = A_s[27];
  assign A_so[28] = \A_s[26] ;
  assign \A_s[26]  = A_s[26];
  assign A_so[27] = \A_s[25] ;
  assign \A_s[25]  = A_s[25];
  assign A_so[26] = \A_s[24] ;
  assign \A_s[24]  = A_s[24];
  assign A_so[25] = \A_s[23] ;
  assign \A_s[23]  = A_s[23];
  assign A_so[24] = \A_s[22] ;
  assign \A_s[22]  = A_s[22];
  assign A_so[23] = \A_s[21] ;
  assign \A_s[21]  = A_s[21];
  assign A_so[22] = \A_s[20] ;
  assign \A_s[20]  = A_s[20];
  assign A_so[21] = \A_s[19] ;
  assign \A_s[19]  = A_s[19];
  assign A_so[20] = \A_s[18] ;
  assign \A_s[18]  = A_s[18];
  assign A_so[19] = \A_s[17] ;
  assign \A_s[17]  = A_s[17];
  assign A_so[18] = \A_s[16] ;
  assign \A_s[16]  = A_s[16];
  assign A_so[17] = \A_s[15] ;
  assign \A_s[15]  = A_s[15];
  assign A_so[16] = \A_s[14] ;
  assign \A_s[14]  = A_s[14];
  assign A_so[15] = \A_s[13] ;
  assign \A_s[13]  = A_s[13];
  assign A_so[14] = \A_s[12] ;
  assign \A_s[12]  = A_s[12];
  assign A_so[13] = \A_s[11] ;
  assign \A_s[11]  = A_s[11];
  assign A_so[12] = \A_s[10] ;
  assign \A_s[10]  = A_s[10];
  assign A_so[11] = \A_s[9] ;
  assign \A_s[9]  = A_s[9];
  assign A_so[10] = \A_s[8] ;
  assign \A_s[8]  = A_s[8];
  assign A_so[9] = \A_s[7] ;
  assign \A_s[7]  = A_s[7];
  assign A_so[8] = \A_s[6] ;
  assign \A_s[6]  = A_s[6];
  assign A_so[7] = \A_s[5] ;
  assign \A_s[5]  = A_s[5];
  assign A_so[6] = \A_s[4] ;
  assign \A_s[4]  = A_s[4];
  assign A_so[5] = \A_s[3] ;
  assign \A_s[3]  = A_s[3];
  assign A_so[4] = \A_s[2] ;
  assign \A_s[2]  = A_s[2];
  assign A_so[3] = \A_s[1] ;
  assign \A_s[1]  = A_s[1];
  assign A_so[2] = \A_s[0] ;
  assign \A_s[0]  = A_s[0];
  assign A_nso[61] = \A_ns[59] ;
  assign \A_ns[59]  = A_ns[59];
  assign A_nso[60] = \A_ns[58] ;
  assign \A_ns[58]  = A_ns[58];
  assign A_nso[59] = \A_ns[57] ;
  assign \A_ns[57]  = A_ns[57];
  assign A_nso[58] = \A_ns[56] ;
  assign \A_ns[56]  = A_ns[56];
  assign A_nso[57] = \A_ns[55] ;
  assign \A_ns[55]  = A_ns[55];
  assign A_nso[56] = \A_ns[54] ;
  assign \A_ns[54]  = A_ns[54];
  assign A_nso[55] = \A_ns[53] ;
  assign \A_ns[53]  = A_ns[53];
  assign A_nso[54] = \A_ns[52] ;
  assign \A_ns[52]  = A_ns[52];
  assign A_nso[53] = \A_ns[51] ;
  assign \A_ns[51]  = A_ns[51];
  assign A_nso[52] = \A_ns[50] ;
  assign \A_ns[50]  = A_ns[50];
  assign A_nso[51] = \A_ns[49] ;
  assign \A_ns[49]  = A_ns[49];
  assign A_nso[50] = \A_ns[48] ;
  assign \A_ns[48]  = A_ns[48];
  assign A_nso[49] = \A_ns[47] ;
  assign \A_ns[47]  = A_ns[47];
  assign A_nso[48] = \A_ns[46] ;
  assign \A_ns[46]  = A_ns[46];
  assign A_nso[47] = \A_ns[45] ;
  assign \A_ns[45]  = A_ns[45];
  assign A_nso[46] = \A_ns[44] ;
  assign \A_ns[44]  = A_ns[44];
  assign A_nso[45] = \A_ns[43] ;
  assign \A_ns[43]  = A_ns[43];
  assign A_nso[44] = \A_ns[42] ;
  assign \A_ns[42]  = A_ns[42];
  assign A_nso[43] = \A_ns[41] ;
  assign \A_ns[41]  = A_ns[41];
  assign A_nso[42] = \A_ns[40] ;
  assign \A_ns[40]  = A_ns[40];
  assign A_nso[41] = \A_ns[39] ;
  assign \A_ns[39]  = A_ns[39];
  assign A_nso[40] = \A_ns[38] ;
  assign \A_ns[38]  = A_ns[38];
  assign A_nso[39] = \A_ns[37] ;
  assign \A_ns[37]  = A_ns[37];
  assign A_nso[38] = \A_ns[36] ;
  assign \A_ns[36]  = A_ns[36];
  assign A_nso[37] = \A_ns[35] ;
  assign \A_ns[35]  = A_ns[35];
  assign A_nso[36] = \A_ns[34] ;
  assign \A_ns[34]  = A_ns[34];
  assign A_nso[35] = \A_ns[33] ;
  assign \A_ns[33]  = A_ns[33];
  assign A_nso[34] = \A_ns[32] ;
  assign \A_ns[32]  = A_ns[32];
  assign A_nso[33] = \A_ns[31] ;
  assign \A_ns[31]  = A_ns[31];
  assign A_nso[32] = \A_ns[30] ;
  assign \A_ns[30]  = A_ns[30];
  assign A_nso[31] = \A_ns[29] ;
  assign \A_ns[29]  = A_ns[29];
  assign A_nso[30] = \A_ns[28] ;
  assign \A_ns[28]  = A_ns[28];
  assign A_nso[29] = \A_ns[27] ;
  assign \A_ns[27]  = A_ns[27];
  assign A_nso[28] = \A_ns[26] ;
  assign \A_ns[26]  = A_ns[26];
  assign A_nso[27] = \A_ns[25] ;
  assign \A_ns[25]  = A_ns[25];
  assign A_nso[26] = \A_ns[24] ;
  assign \A_ns[24]  = A_ns[24];
  assign A_nso[25] = \A_ns[23] ;
  assign \A_ns[23]  = A_ns[23];
  assign A_nso[24] = \A_ns[22] ;
  assign \A_ns[22]  = A_ns[22];
  assign A_nso[23] = \A_ns[21] ;
  assign \A_ns[21]  = A_ns[21];
  assign A_nso[22] = \A_ns[20] ;
  assign \A_ns[20]  = A_ns[20];
  assign A_nso[21] = \A_ns[19] ;
  assign \A_ns[19]  = A_ns[19];
  assign A_nso[20] = \A_ns[18] ;
  assign \A_ns[18]  = A_ns[18];
  assign A_nso[19] = \A_ns[17] ;
  assign \A_ns[17]  = A_ns[17];
  assign A_nso[18] = \A_ns[16] ;
  assign \A_ns[16]  = A_ns[16];
  assign A_nso[17] = \A_ns[15] ;
  assign \A_ns[15]  = A_ns[15];
  assign A_nso[16] = \A_ns[14] ;
  assign \A_ns[14]  = A_ns[14];
  assign A_nso[15] = \A_ns[13] ;
  assign \A_ns[13]  = A_ns[13];
  assign A_nso[14] = \A_ns[12] ;
  assign \A_ns[12]  = A_ns[12];
  assign A_nso[13] = \A_ns[11] ;
  assign \A_ns[11]  = A_ns[11];
  assign A_nso[12] = \A_ns[10] ;
  assign \A_ns[10]  = A_ns[10];
  assign A_nso[11] = \A_ns[9] ;
  assign \A_ns[9]  = A_ns[9];
  assign A_nso[10] = \A_ns[8] ;
  assign \A_ns[8]  = A_ns[8];
  assign A_nso[9] = \A_ns[7] ;
  assign \A_ns[7]  = A_ns[7];
  assign A_nso[8] = \A_ns[6] ;
  assign \A_ns[6]  = A_ns[6];
  assign A_nso[7] = \A_ns[5] ;
  assign \A_ns[5]  = A_ns[5];
  assign A_nso[6] = \A_ns[4] ;
  assign \A_ns[4]  = A_ns[4];
  assign A_nso[5] = \A_ns[3] ;
  assign \A_ns[3]  = A_ns[3];
  assign A_nso[4] = \A_ns[2] ;
  assign \A_ns[2]  = A_ns[2];
  assign A_nso[3] = \A_ns[1] ;
  assign \A_ns[1]  = A_ns[1];
  assign A_nso[2] = \A_ns[0] ;
  assign \A_ns[0]  = A_ns[0];

  XOR2_X1 U249 ( .A(B[27]), .B(B[28]), .Z(n188) );
  NAND3_X1 U250 ( .A1(B[28]), .A2(n869), .A3(B[27]), .ZN(n125) );
  OAI221_X1 U2 ( .B1(n742), .B2(n776), .C1(n739), .C2(n810), .A(n133), .ZN(
        O[59]) );
  AOI22_X1 U3 ( .A1(\A_ns[27] ), .A2(n729), .B1(\A_s[27] ), .B2(n722), .ZN(
        n167) );
  AOI22_X1 U4 ( .A1(A_ns[60]), .A2(n732), .B1(A_s[60]), .B2(n725), .ZN(n130)
         );
  AOI22_X1 U5 ( .A1(\A_ns[56] ), .A2(n732), .B1(\A_s[56] ), .B2(n725), .ZN(
        n135) );
  BUF_X1 U6 ( .A(n726), .Z(n729) );
  BUF_X1 U7 ( .A(n719), .Z(n722) );
  BUF_X1 U8 ( .A(n726), .Z(n730) );
  BUF_X1 U9 ( .A(n719), .Z(n723) );
  BUF_X1 U10 ( .A(n727), .Z(n731) );
  BUF_X1 U11 ( .A(n720), .Z(n724) );
  BUF_X1 U12 ( .A(n727), .Z(n732) );
  BUF_X1 U13 ( .A(n720), .Z(n725) );
  BUF_X1 U14 ( .A(n726), .Z(n728) );
  BUF_X1 U15 ( .A(n719), .Z(n721) );
  OAI221_X1 U16 ( .B1(n742), .B2(n778), .C1(n739), .C2(n812), .A(n130), .ZN(
        O[61]) );
  OAI221_X1 U17 ( .B1(n742), .B2(n774), .C1(n738), .C2(n808), .A(n135), .ZN(
        O[57]) );
  OAI221_X1 U18 ( .B1(n742), .B2(n775), .C1(n738), .C2(n809), .A(n134), .ZN(
        O[58]) );
  AOI22_X1 U19 ( .A1(\A_ns[57] ), .A2(n732), .B1(\A_s[57] ), .B2(n725), .ZN(
        n134) );
  OAI221_X1 U20 ( .B1(n745), .B2(n779), .C1(n736), .C2(n780), .A(n166), .ZN(
        O[29]) );
  AOI22_X1 U21 ( .A1(\A_ns[28] ), .A2(n729), .B1(\A_s[28] ), .B2(n722), .ZN(
        n166) );
  OAI221_X1 U22 ( .B1(n744), .B2(n751), .C1(n736), .C2(n785), .A(n160), .ZN(
        O[34]) );
  AOI22_X1 U23 ( .A1(\A_ns[33] ), .A2(n730), .B1(\A_s[33] ), .B2(n723), .ZN(
        n160) );
  OAI221_X1 U24 ( .B1(n745), .B2(n749), .C1(n736), .C2(n783), .A(n162), .ZN(
        O[32]) );
  AOI22_X1 U25 ( .A1(\A_ns[31] ), .A2(n729), .B1(\A_s[31] ), .B2(n722), .ZN(
        n162) );
  OAI221_X1 U26 ( .B1(n745), .B2(n747), .C1(n736), .C2(n781), .A(n164), .ZN(
        O[30]) );
  AOI22_X1 U27 ( .A1(\A_ns[29] ), .A2(n729), .B1(\A_s[29] ), .B2(n722), .ZN(
        n164) );
  OAI221_X1 U28 ( .B1(n745), .B2(n748), .C1(n736), .C2(n782), .A(n163), .ZN(
        O[31]) );
  AOI22_X1 U29 ( .A1(\A_ns[30] ), .A2(n729), .B1(\A_s[30] ), .B2(n722), .ZN(
        n163) );
  OAI221_X1 U30 ( .B1(n744), .B2(n752), .C1(n737), .C2(n786), .A(n159), .ZN(
        O[35]) );
  AOI22_X1 U31 ( .A1(\A_ns[34] ), .A2(n730), .B1(\A_s[34] ), .B2(n723), .ZN(
        n159) );
  OAI221_X1 U32 ( .B1(n744), .B2(n750), .C1(n736), .C2(n784), .A(n161), .ZN(
        O[33]) );
  AOI22_X1 U33 ( .A1(\A_ns[32] ), .A2(n730), .B1(\A_s[32] ), .B2(n723), .ZN(
        n161) );
  BUF_X1 U34 ( .A(n867), .Z(n719) );
  BUF_X1 U35 ( .A(n868), .Z(n726) );
  OAI221_X1 U36 ( .B1(n744), .B2(n753), .C1(n737), .C2(n787), .A(n158), .ZN(
        O[36]) );
  AOI22_X1 U37 ( .A1(\A_ns[35] ), .A2(n730), .B1(\A_s[35] ), .B2(n723), .ZN(
        n158) );
  OAI221_X1 U38 ( .B1(n744), .B2(n755), .C1(n737), .C2(n789), .A(n156), .ZN(
        O[38]) );
  AOI22_X1 U39 ( .A1(\A_ns[37] ), .A2(n730), .B1(\A_s[37] ), .B2(n723), .ZN(
        n156) );
  OAI221_X1 U40 ( .B1(n743), .B2(n765), .C1(n738), .C2(n799), .A(n145), .ZN(
        O[48]) );
  AOI22_X1 U41 ( .A1(\A_ns[47] ), .A2(n731), .B1(\A_s[47] ), .B2(n724), .ZN(
        n145) );
  OAI221_X1 U42 ( .B1(n743), .B2(n764), .C1(n738), .C2(n798), .A(n146), .ZN(
        O[47]) );
  AOI22_X1 U43 ( .A1(\A_ns[46] ), .A2(n731), .B1(\A_s[46] ), .B2(n724), .ZN(
        n146) );
  OAI221_X1 U44 ( .B1(n744), .B2(n754), .C1(n737), .C2(n788), .A(n157), .ZN(
        O[37]) );
  AOI22_X1 U45 ( .A1(\A_ns[36] ), .A2(n730), .B1(\A_s[36] ), .B2(n723), .ZN(
        n157) );
  OAI221_X1 U46 ( .B1(n744), .B2(n759), .C1(n737), .C2(n793), .A(n151), .ZN(
        O[42]) );
  AOI22_X1 U47 ( .A1(\A_ns[41] ), .A2(n730), .B1(\A_s[41] ), .B2(n723), .ZN(
        n151) );
  OAI221_X1 U48 ( .B1(n744), .B2(n758), .C1(n737), .C2(n792), .A(n152), .ZN(
        O[41]) );
  AOI22_X1 U49 ( .A1(\A_ns[40] ), .A2(n730), .B1(\A_s[40] ), .B2(n723), .ZN(
        n152) );
  OAI221_X1 U50 ( .B1(n744), .B2(n757), .C1(n737), .C2(n791), .A(n153), .ZN(
        O[40]) );
  AOI22_X1 U51 ( .A1(\A_ns[39] ), .A2(n730), .B1(\A_s[39] ), .B2(n723), .ZN(
        n153) );
  OAI221_X1 U52 ( .B1(n744), .B2(n756), .C1(n737), .C2(n790), .A(n155), .ZN(
        O[39]) );
  AOI22_X1 U53 ( .A1(\A_ns[38] ), .A2(n730), .B1(\A_s[38] ), .B2(n723), .ZN(
        n155) );
  OAI221_X1 U54 ( .B1(n743), .B2(n761), .C1(n737), .C2(n795), .A(n149), .ZN(
        O[44]) );
  AOI22_X1 U55 ( .A1(\A_ns[43] ), .A2(n731), .B1(\A_s[43] ), .B2(n724), .ZN(
        n149) );
  OAI221_X1 U56 ( .B1(n744), .B2(n760), .C1(n737), .C2(n794), .A(n150), .ZN(
        O[43]) );
  AOI22_X1 U57 ( .A1(\A_ns[42] ), .A2(n730), .B1(\A_s[42] ), .B2(n723), .ZN(
        n150) );
  OAI221_X1 U58 ( .B1(n743), .B2(n762), .C1(n737), .C2(n796), .A(n148), .ZN(
        O[45]) );
  AOI22_X1 U59 ( .A1(\A_ns[44] ), .A2(n731), .B1(\A_s[44] ), .B2(n724), .ZN(
        n148) );
  OAI221_X1 U60 ( .B1(n743), .B2(n763), .C1(n737), .C2(n797), .A(n147), .ZN(
        O[46]) );
  AOI22_X1 U61 ( .A1(\A_ns[45] ), .A2(n731), .B1(\A_s[45] ), .B2(n724), .ZN(
        n147) );
  OAI221_X1 U62 ( .B1(n743), .B2(n766), .C1(n738), .C2(n800), .A(n144), .ZN(
        O[49]) );
  AOI22_X1 U63 ( .A1(\A_ns[48] ), .A2(n731), .B1(\A_s[48] ), .B2(n724), .ZN(
        n144) );
  OAI221_X1 U64 ( .B1(n743), .B2(n767), .C1(n738), .C2(n801), .A(n142), .ZN(
        O[50]) );
  AOI22_X1 U65 ( .A1(\A_ns[49] ), .A2(n731), .B1(\A_s[49] ), .B2(n724), .ZN(
        n142) );
  OAI221_X1 U66 ( .B1(n743), .B2(n768), .C1(n738), .C2(n802), .A(n141), .ZN(
        O[51]) );
  AOI22_X1 U67 ( .A1(\A_ns[50] ), .A2(n731), .B1(\A_s[50] ), .B2(n724), .ZN(
        n141) );
  OAI221_X1 U68 ( .B1(n743), .B2(n769), .C1(n738), .C2(n803), .A(n140), .ZN(
        O[52]) );
  AOI22_X1 U69 ( .A1(\A_ns[51] ), .A2(n731), .B1(\A_s[51] ), .B2(n724), .ZN(
        n140) );
  OAI221_X1 U70 ( .B1(n743), .B2(n770), .C1(n738), .C2(n804), .A(n139), .ZN(
        O[53]) );
  AOI22_X1 U71 ( .A1(\A_ns[52] ), .A2(n731), .B1(\A_s[52] ), .B2(n724), .ZN(
        n139) );
  OAI221_X1 U72 ( .B1(n743), .B2(n771), .C1(n738), .C2(n805), .A(n138), .ZN(
        O[54]) );
  AOI22_X1 U73 ( .A1(\A_ns[53] ), .A2(n731), .B1(\A_s[53] ), .B2(n724), .ZN(
        n138) );
  OAI221_X1 U74 ( .B1(n742), .B2(n772), .C1(n738), .C2(n806), .A(n137), .ZN(
        O[55]) );
  AOI22_X1 U75 ( .A1(\A_ns[54] ), .A2(n732), .B1(\A_s[54] ), .B2(n725), .ZN(
        n137) );
  AOI22_X1 U76 ( .A1(\A_ns[58] ), .A2(n732), .B1(\A_s[58] ), .B2(n725), .ZN(
        n133) );
  OAI221_X1 U77 ( .B1(n742), .B2(n773), .C1(n738), .C2(n807), .A(n136), .ZN(
        O[56]) );
  AOI22_X1 U78 ( .A1(\A_ns[55] ), .A2(n732), .B1(\A_s[55] ), .B2(n725), .ZN(
        n136) );
  OAI221_X1 U79 ( .B1(n742), .B2(n777), .C1(n739), .C2(n811), .A(n131), .ZN(
        O[60]) );
  AOI22_X1 U80 ( .A1(\A_ns[59] ), .A2(n732), .B1(\A_s[59] ), .B2(n725), .ZN(
        n131) );
  BUF_X1 U81 ( .A(n867), .Z(n720) );
  BUF_X1 U82 ( .A(n868), .Z(n727) );
  BUF_X1 U83 ( .A(n741), .Z(n745) );
  INV_X1 U84 ( .A(n176), .ZN(n867) );
  INV_X1 U85 ( .A(n177), .ZN(n868) );
  BUF_X1 U86 ( .A(n740), .Z(n744) );
  BUF_X1 U87 ( .A(n733), .Z(n736) );
  BUF_X1 U88 ( .A(n733), .Z(n737) );
  BUF_X1 U89 ( .A(n740), .Z(n743) );
  BUF_X1 U90 ( .A(n734), .Z(n738) );
  BUF_X1 U91 ( .A(n740), .Z(n742) );
  BUF_X1 U92 ( .A(n734), .Z(n739) );
  BUF_X1 U93 ( .A(n741), .Z(n746) );
  BUF_X1 U94 ( .A(n733), .Z(n735) );
  NAND2_X1 U95 ( .A1(n188), .A2(n869), .ZN(n176) );
  NAND2_X1 U96 ( .A1(n188), .A2(n176), .ZN(n177) );
  BUF_X1 U97 ( .A(n124), .Z(n741) );
  BUF_X1 U98 ( .A(n125), .Z(n733) );
  BUF_X1 U99 ( .A(n124), .Z(n740) );
  BUF_X1 U100 ( .A(n125), .Z(n734) );
  OAI221_X1 U101 ( .B1(n745), .B2(n865), .C1(n736), .C2(n866), .A(n167), .ZN(
        O[28]) );
  INV_X1 U102 ( .A(\A_ns[26] ), .ZN(n865) );
  INV_X1 U103 ( .A(\A_s[26] ), .ZN(n866) );
  OAI221_X1 U104 ( .B1(n745), .B2(n861), .C1(n736), .C2(n863), .A(n169), .ZN(
        O[26]) );
  INV_X1 U105 ( .A(\A_ns[24] ), .ZN(n861) );
  OAI221_X1 U106 ( .B1(n746), .B2(n850), .C1(n735), .C2(n852), .A(n174), .ZN(
        O[21]) );
  INV_X1 U107 ( .A(\A_ns[19] ), .ZN(n850) );
  INV_X1 U108 ( .A(\A_s[19] ), .ZN(n852) );
  OAI221_X1 U109 ( .B1(n745), .B2(n853), .C1(n735), .C2(n855), .A(n173), .ZN(
        O[22]) );
  INV_X1 U110 ( .A(\A_ns[20] ), .ZN(n853) );
  INV_X1 U111 ( .A(\A_s[20] ), .ZN(n855) );
  OAI221_X1 U112 ( .B1(n745), .B2(n854), .C1(n736), .C2(n856), .A(n172), .ZN(
        O[23]) );
  INV_X1 U113 ( .A(\A_ns[21] ), .ZN(n854) );
  INV_X1 U114 ( .A(\A_s[21] ), .ZN(n856) );
  OAI221_X1 U115 ( .B1(n745), .B2(n857), .C1(n736), .C2(n859), .A(n171), .ZN(
        O[24]) );
  INV_X1 U116 ( .A(\A_ns[22] ), .ZN(n857) );
  INV_X1 U117 ( .A(\A_s[22] ), .ZN(n859) );
  OAI221_X1 U118 ( .B1(n745), .B2(n858), .C1(n736), .C2(n860), .A(n170), .ZN(
        O[25]) );
  INV_X1 U119 ( .A(\A_ns[23] ), .ZN(n858) );
  INV_X1 U120 ( .A(\A_s[23] ), .ZN(n860) );
  OAI221_X1 U121 ( .B1(n745), .B2(n862), .C1(n736), .C2(n864), .A(n168), .ZN(
        O[27]) );
  INV_X1 U122 ( .A(\A_ns[25] ), .ZN(n862) );
  INV_X1 U123 ( .A(\A_s[25] ), .ZN(n864) );
  INV_X1 U124 ( .A(B[29]), .ZN(n869) );
  OR3_X1 U125 ( .A1(B[27]), .A2(B[28]), .A3(n869), .ZN(n124) );
  OAI221_X1 U126 ( .B1(n746), .B2(n838), .C1(n735), .C2(n840), .A(n182), .ZN(
        O[15]) );
  INV_X1 U127 ( .A(\A_ns[13] ), .ZN(n838) );
  INV_X1 U128 ( .A(\A_s[13] ), .ZN(n840) );
  OAI221_X1 U129 ( .B1(n746), .B2(n841), .C1(n735), .C2(n843), .A(n181), .ZN(
        O[16]) );
  INV_X1 U130 ( .A(\A_ns[14] ), .ZN(n841) );
  INV_X1 U131 ( .A(\A_s[14] ), .ZN(n843) );
  OAI221_X1 U132 ( .B1(n746), .B2(n842), .C1(n735), .C2(n844), .A(n180), .ZN(
        O[17]) );
  INV_X1 U133 ( .A(\A_ns[15] ), .ZN(n842) );
  INV_X1 U134 ( .A(\A_s[15] ), .ZN(n844) );
  OAI221_X1 U135 ( .B1(n746), .B2(n845), .C1(n735), .C2(n847), .A(n179), .ZN(
        O[18]) );
  INV_X1 U136 ( .A(\A_ns[16] ), .ZN(n845) );
  INV_X1 U137 ( .A(\A_s[16] ), .ZN(n847) );
  OAI221_X1 U138 ( .B1(n746), .B2(n846), .C1(n735), .C2(n848), .A(n178), .ZN(
        O[19]) );
  INV_X1 U139 ( .A(\A_ns[17] ), .ZN(n846) );
  INV_X1 U140 ( .A(\A_s[17] ), .ZN(n848) );
  OAI221_X1 U141 ( .B1(n746), .B2(n849), .C1(n735), .C2(n851), .A(n175), .ZN(
        O[20]) );
  INV_X1 U142 ( .A(\A_ns[18] ), .ZN(n849) );
  INV_X1 U143 ( .A(\A_s[18] ), .ZN(n851) );
  OAI221_X1 U144 ( .B1(n742), .B2(n822), .C1(n739), .C2(n824), .A(n128), .ZN(
        O[7]) );
  INV_X1 U145 ( .A(\A_ns[5] ), .ZN(n822) );
  INV_X1 U146 ( .A(\A_s[5] ), .ZN(n824) );
  OAI221_X1 U147 ( .B1(n742), .B2(n825), .C1(n739), .C2(n827), .A(n127), .ZN(
        O[8]) );
  INV_X1 U148 ( .A(\A_ns[6] ), .ZN(n825) );
  INV_X1 U149 ( .A(\A_s[6] ), .ZN(n827) );
  OAI221_X1 U150 ( .B1(n742), .B2(n826), .C1(n739), .C2(n828), .A(n126), .ZN(
        O[9]) );
  INV_X1 U151 ( .A(\A_ns[7] ), .ZN(n826) );
  INV_X1 U152 ( .A(\A_s[7] ), .ZN(n828) );
  OAI221_X1 U153 ( .B1(n829), .B2(n746), .C1(n831), .C2(n735), .A(n187), .ZN(
        O[10]) );
  INV_X1 U154 ( .A(\A_s[8] ), .ZN(n831) );
  INV_X1 U155 ( .A(\A_ns[8] ), .ZN(n829) );
  OAI221_X1 U156 ( .B1(n746), .B2(n830), .C1(n735), .C2(n832), .A(n186), .ZN(
        O[11]) );
  INV_X1 U157 ( .A(\A_ns[9] ), .ZN(n830) );
  INV_X1 U158 ( .A(\A_s[9] ), .ZN(n832) );
  OAI221_X1 U159 ( .B1(n746), .B2(n833), .C1(n735), .C2(n835), .A(n185), .ZN(
        O[12]) );
  INV_X1 U160 ( .A(\A_ns[10] ), .ZN(n833) );
  INV_X1 U161 ( .A(\A_s[10] ), .ZN(n835) );
  OAI221_X1 U162 ( .B1(n746), .B2(n834), .C1(n735), .C2(n836), .A(n184), .ZN(
        O[13]) );
  INV_X1 U163 ( .A(\A_ns[11] ), .ZN(n834) );
  INV_X1 U164 ( .A(\A_s[11] ), .ZN(n836) );
  OAI221_X1 U165 ( .B1(n746), .B2(n837), .C1(n735), .C2(n839), .A(n183), .ZN(
        O[14]) );
  INV_X1 U166 ( .A(\A_ns[12] ), .ZN(n837) );
  INV_X1 U167 ( .A(\A_s[12] ), .ZN(n839) );
  OAI22_X1 U168 ( .A1(n176), .A2(n815), .B1(n177), .B2(n813), .ZN(O[1]) );
  OAI221_X1 U169 ( .B1(n745), .B2(n813), .C1(n736), .C2(n815), .A(n165), .ZN(
        O[2]) );
  AOI22_X1 U170 ( .A1(\A_ns[1] ), .A2(n729), .B1(\A_s[1] ), .B2(n722), .ZN(
        n165) );
  OAI221_X1 U171 ( .B1(n744), .B2(n814), .C1(n737), .C2(n816), .A(n154), .ZN(
        O[3]) );
  INV_X1 U172 ( .A(\A_ns[1] ), .ZN(n814) );
  INV_X1 U173 ( .A(\A_s[1] ), .ZN(n816) );
  OAI221_X1 U174 ( .B1(n743), .B2(n817), .C1(n738), .C2(n819), .A(n143), .ZN(
        O[4]) );
  INV_X1 U175 ( .A(\A_ns[2] ), .ZN(n817) );
  INV_X1 U176 ( .A(\A_s[2] ), .ZN(n819) );
  OAI221_X1 U177 ( .B1(n742), .B2(n818), .C1(n739), .C2(n820), .A(n132), .ZN(
        O[5]) );
  INV_X1 U178 ( .A(\A_ns[3] ), .ZN(n818) );
  INV_X1 U179 ( .A(\A_s[3] ), .ZN(n820) );
  OAI221_X1 U180 ( .B1(n742), .B2(n821), .C1(n739), .C2(n823), .A(n129), .ZN(
        O[6]) );
  INV_X1 U181 ( .A(\A_ns[4] ), .ZN(n821) );
  INV_X1 U182 ( .A(\A_s[4] ), .ZN(n823) );
  INV_X1 U183 ( .A(\A_s[0] ), .ZN(n815) );
  INV_X1 U184 ( .A(\A_ns[0] ), .ZN(n813) );
  AOI22_X1 U185 ( .A1(\A_ns[2] ), .A2(n730), .B1(\A_s[2] ), .B2(n723), .ZN(
        n154) );
  AOI22_X1 U186 ( .A1(\A_ns[3] ), .A2(n731), .B1(\A_s[3] ), .B2(n724), .ZN(
        n143) );
  AOI22_X1 U187 ( .A1(\A_ns[4] ), .A2(n732), .B1(\A_s[4] ), .B2(n725), .ZN(
        n132) );
  AOI22_X1 U188 ( .A1(\A_ns[5] ), .A2(n732), .B1(\A_s[5] ), .B2(n725), .ZN(
        n129) );
  AOI22_X1 U189 ( .A1(\A_ns[6] ), .A2(n732), .B1(\A_s[6] ), .B2(n725), .ZN(
        n128) );
  AOI22_X1 U190 ( .A1(\A_ns[7] ), .A2(n732), .B1(\A_s[7] ), .B2(n725), .ZN(
        n127) );
  AOI22_X1 U191 ( .A1(\A_ns[8] ), .A2(n732), .B1(\A_s[8] ), .B2(n725), .ZN(
        n126) );
  AOI22_X1 U192 ( .A1(\A_ns[9] ), .A2(n728), .B1(\A_s[9] ), .B2(n721), .ZN(
        n187) );
  AOI22_X1 U193 ( .A1(\A_ns[10] ), .A2(n728), .B1(\A_s[10] ), .B2(n721), .ZN(
        n186) );
  AOI22_X1 U194 ( .A1(\A_ns[11] ), .A2(n728), .B1(\A_s[11] ), .B2(n721), .ZN(
        n185) );
  AOI22_X1 U195 ( .A1(\A_ns[12] ), .A2(n728), .B1(\A_s[12] ), .B2(n721), .ZN(
        n184) );
  AOI22_X1 U196 ( .A1(\A_ns[13] ), .A2(n728), .B1(\A_s[13] ), .B2(n721), .ZN(
        n183) );
  AOI22_X1 U197 ( .A1(\A_ns[14] ), .A2(n728), .B1(\A_s[14] ), .B2(n721), .ZN(
        n182) );
  AOI22_X1 U198 ( .A1(\A_ns[15] ), .A2(n728), .B1(\A_s[15] ), .B2(n721), .ZN(
        n181) );
  AOI22_X1 U199 ( .A1(\A_ns[16] ), .A2(n728), .B1(\A_s[16] ), .B2(n721), .ZN(
        n180) );
  AOI22_X1 U200 ( .A1(\A_ns[17] ), .A2(n728), .B1(\A_s[17] ), .B2(n721), .ZN(
        n179) );
  AOI22_X1 U201 ( .A1(\A_ns[18] ), .A2(n728), .B1(\A_s[18] ), .B2(n721), .ZN(
        n178) );
  AOI22_X1 U202 ( .A1(\A_ns[19] ), .A2(n728), .B1(\A_s[19] ), .B2(n721), .ZN(
        n175) );
  AOI22_X1 U203 ( .A1(\A_ns[20] ), .A2(n728), .B1(\A_s[20] ), .B2(n721), .ZN(
        n174) );
  AOI22_X1 U204 ( .A1(\A_ns[21] ), .A2(n729), .B1(\A_s[21] ), .B2(n722), .ZN(
        n173) );
  AOI22_X1 U205 ( .A1(\A_ns[22] ), .A2(n729), .B1(\A_s[22] ), .B2(n722), .ZN(
        n172) );
  AOI22_X1 U206 ( .A1(\A_ns[23] ), .A2(n729), .B1(\A_s[23] ), .B2(n722), .ZN(
        n171) );
  AOI22_X1 U207 ( .A1(\A_ns[24] ), .A2(n729), .B1(\A_s[24] ), .B2(n722), .ZN(
        n170) );
  AOI22_X1 U208 ( .A1(\A_ns[25] ), .A2(n729), .B1(\A_s[25] ), .B2(n722), .ZN(
        n169) );
  AOI22_X1 U209 ( .A1(\A_ns[26] ), .A2(n729), .B1(\A_s[26] ), .B2(n722), .ZN(
        n168) );
  INV_X1 U210 ( .A(\A_s[24] ), .ZN(n863) );
  INV_X1 U211 ( .A(\A_ns[28] ), .ZN(n747) );
  INV_X1 U212 ( .A(\A_ns[29] ), .ZN(n748) );
  INV_X1 U213 ( .A(\A_ns[30] ), .ZN(n749) );
  INV_X1 U214 ( .A(\A_ns[31] ), .ZN(n750) );
  INV_X1 U215 ( .A(\A_ns[32] ), .ZN(n751) );
  INV_X1 U216 ( .A(\A_ns[33] ), .ZN(n752) );
  INV_X1 U217 ( .A(\A_ns[34] ), .ZN(n753) );
  INV_X1 U218 ( .A(\A_ns[35] ), .ZN(n754) );
  INV_X1 U219 ( .A(\A_ns[36] ), .ZN(n755) );
  INV_X1 U220 ( .A(\A_ns[37] ), .ZN(n756) );
  INV_X1 U221 ( .A(\A_ns[38] ), .ZN(n757) );
  INV_X1 U222 ( .A(\A_ns[39] ), .ZN(n758) );
  INV_X1 U223 ( .A(\A_ns[40] ), .ZN(n759) );
  INV_X1 U224 ( .A(\A_ns[41] ), .ZN(n760) );
  INV_X1 U225 ( .A(\A_ns[42] ), .ZN(n761) );
  INV_X1 U226 ( .A(\A_ns[43] ), .ZN(n762) );
  INV_X1 U227 ( .A(\A_ns[44] ), .ZN(n763) );
  INV_X1 U228 ( .A(\A_ns[45] ), .ZN(n764) );
  INV_X1 U229 ( .A(\A_ns[46] ), .ZN(n765) );
  INV_X1 U230 ( .A(\A_ns[47] ), .ZN(n766) );
  INV_X1 U231 ( .A(\A_ns[48] ), .ZN(n767) );
  INV_X1 U232 ( .A(\A_ns[49] ), .ZN(n768) );
  INV_X1 U233 ( .A(\A_ns[50] ), .ZN(n769) );
  INV_X1 U234 ( .A(\A_ns[51] ), .ZN(n770) );
  INV_X1 U235 ( .A(\A_ns[52] ), .ZN(n771) );
  INV_X1 U236 ( .A(\A_ns[53] ), .ZN(n772) );
  INV_X1 U237 ( .A(\A_ns[54] ), .ZN(n773) );
  INV_X1 U238 ( .A(\A_ns[55] ), .ZN(n774) );
  INV_X1 U239 ( .A(\A_ns[56] ), .ZN(n775) );
  INV_X1 U240 ( .A(\A_ns[57] ), .ZN(n776) );
  INV_X1 U241 ( .A(\A_ns[58] ), .ZN(n777) );
  INV_X1 U242 ( .A(\A_ns[59] ), .ZN(n778) );
  INV_X1 U243 ( .A(\A_ns[27] ), .ZN(n779) );
  INV_X1 U244 ( .A(\A_s[27] ), .ZN(n780) );
  INV_X1 U245 ( .A(\A_s[28] ), .ZN(n781) );
  INV_X1 U246 ( .A(\A_s[29] ), .ZN(n782) );
  INV_X1 U247 ( .A(\A_s[30] ), .ZN(n783) );
  INV_X1 U248 ( .A(\A_s[31] ), .ZN(n784) );
  INV_X1 U251 ( .A(\A_s[32] ), .ZN(n785) );
  INV_X1 U252 ( .A(\A_s[33] ), .ZN(n786) );
  INV_X1 U253 ( .A(\A_s[34] ), .ZN(n787) );
  INV_X1 U254 ( .A(\A_s[35] ), .ZN(n788) );
  INV_X1 U255 ( .A(\A_s[36] ), .ZN(n789) );
  INV_X1 U256 ( .A(\A_s[37] ), .ZN(n790) );
  INV_X1 U257 ( .A(\A_s[38] ), .ZN(n791) );
  INV_X1 U258 ( .A(\A_s[39] ), .ZN(n792) );
  INV_X1 U259 ( .A(\A_s[40] ), .ZN(n793) );
  INV_X1 U260 ( .A(\A_s[41] ), .ZN(n794) );
  INV_X1 U261 ( .A(\A_s[42] ), .ZN(n795) );
  INV_X1 U262 ( .A(\A_s[43] ), .ZN(n796) );
  INV_X1 U263 ( .A(\A_s[44] ), .ZN(n797) );
  INV_X1 U264 ( .A(\A_s[45] ), .ZN(n798) );
  INV_X1 U265 ( .A(\A_s[46] ), .ZN(n799) );
  INV_X1 U266 ( .A(\A_s[47] ), .ZN(n800) );
  INV_X1 U267 ( .A(\A_s[48] ), .ZN(n801) );
  INV_X1 U268 ( .A(\A_s[49] ), .ZN(n802) );
  INV_X1 U269 ( .A(\A_s[50] ), .ZN(n803) );
  INV_X1 U270 ( .A(\A_s[51] ), .ZN(n804) );
  INV_X1 U271 ( .A(\A_s[52] ), .ZN(n805) );
  INV_X1 U272 ( .A(\A_s[53] ), .ZN(n806) );
  INV_X1 U273 ( .A(\A_s[54] ), .ZN(n807) );
  INV_X1 U274 ( .A(\A_s[55] ), .ZN(n808) );
  INV_X1 U275 ( .A(\A_s[56] ), .ZN(n809) );
  INV_X1 U276 ( .A(\A_s[57] ), .ZN(n810) );
  INV_X1 U277 ( .A(\A_s[58] ), .ZN(n811) );
  INV_X1 U278 ( .A(\A_s[59] ), .ZN(n812) );
endmodule


module BOOTHENC_NBIT64_i30 ( A_s, A_ns, B, O, A_so, A_nso );
  input [63:0] A_s;
  input [63:0] A_ns;
  input [63:0] B;
  output [63:0] O;
  output [63:0] A_so;
  output [63:0] A_nso;
  wire   \A_s[61] , \A_s[60] , \A_s[59] , \A_s[58] , \A_s[57] , \A_s[56] ,
         \A_s[55] , \A_s[54] , \A_s[53] , \A_s[52] , \A_s[51] , \A_s[50] ,
         \A_s[49] , \A_s[48] , \A_s[47] , \A_s[46] , \A_s[45] , \A_s[44] ,
         \A_s[43] , \A_s[42] , \A_s[41] , \A_s[40] , \A_s[39] , \A_s[38] ,
         \A_s[37] , \A_s[36] , \A_s[35] , \A_s[34] , \A_s[33] , \A_s[32] ,
         \A_s[31] , \A_s[30] , \A_s[29] , \A_s[28] , \A_s[27] , \A_s[26] ,
         \A_s[25] , \A_s[24] , \A_s[23] , \A_s[22] , \A_s[21] , \A_s[20] ,
         \A_s[19] , \A_s[18] , \A_s[17] , \A_s[16] , \A_s[15] , \A_s[14] ,
         \A_s[13] , \A_s[12] , \A_s[11] , \A_s[10] , \A_s[9] , \A_s[8] ,
         \A_s[7] , \A_s[6] , \A_s[5] , \A_s[4] , \A_s[3] , \A_s[2] , \A_s[1] ,
         \A_s[0] , \A_ns[61] , \A_ns[60] , \A_ns[59] , \A_ns[58] , \A_ns[57] ,
         \A_ns[56] , \A_ns[55] , \A_ns[54] , \A_ns[53] , \A_ns[52] ,
         \A_ns[51] , \A_ns[50] , \A_ns[49] , \A_ns[48] , \A_ns[47] ,
         \A_ns[46] , \A_ns[45] , \A_ns[44] , \A_ns[43] , \A_ns[42] ,
         \A_ns[41] , \A_ns[40] , \A_ns[39] , \A_ns[38] , \A_ns[37] ,
         \A_ns[36] , \A_ns[35] , \A_ns[34] , \A_ns[33] , \A_ns[32] ,
         \A_ns[31] , \A_ns[30] , \A_ns[29] , \A_ns[28] , \A_ns[27] ,
         \A_ns[26] , \A_ns[25] , \A_ns[24] , \A_ns[23] , \A_ns[22] ,
         \A_ns[21] , \A_ns[20] , \A_ns[19] , \A_ns[18] , \A_ns[17] ,
         \A_ns[16] , \A_ns[15] , \A_ns[14] , \A_ns[13] , \A_ns[12] ,
         \A_ns[11] , \A_ns[10] , \A_ns[9] , \A_ns[8] , \A_ns[7] , \A_ns[6] ,
         \A_ns[5] , \A_ns[4] , \A_ns[3] , \A_ns[2] , \A_ns[1] , \A_ns[0] ,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889;
  assign A_nso[0] = 1'b0;
  assign A_nso[1] = 1'b0;
  assign A_so[0] = 1'b0;
  assign A_so[1] = 1'b0;
  assign O[0] = 1'b0;
  assign A_so[63] = \A_s[61] ;
  assign \A_s[61]  = A_s[61];
  assign A_so[62] = \A_s[60] ;
  assign \A_s[60]  = A_s[60];
  assign A_so[61] = \A_s[59] ;
  assign \A_s[59]  = A_s[59];
  assign A_so[60] = \A_s[58] ;
  assign \A_s[58]  = A_s[58];
  assign A_so[59] = \A_s[57] ;
  assign \A_s[57]  = A_s[57];
  assign A_so[58] = \A_s[56] ;
  assign \A_s[56]  = A_s[56];
  assign A_so[57] = \A_s[55] ;
  assign \A_s[55]  = A_s[55];
  assign A_so[56] = \A_s[54] ;
  assign \A_s[54]  = A_s[54];
  assign A_so[55] = \A_s[53] ;
  assign \A_s[53]  = A_s[53];
  assign A_so[54] = \A_s[52] ;
  assign \A_s[52]  = A_s[52];
  assign A_so[53] = \A_s[51] ;
  assign \A_s[51]  = A_s[51];
  assign A_so[52] = \A_s[50] ;
  assign \A_s[50]  = A_s[50];
  assign A_so[51] = \A_s[49] ;
  assign \A_s[49]  = A_s[49];
  assign A_so[50] = \A_s[48] ;
  assign \A_s[48]  = A_s[48];
  assign A_so[49] = \A_s[47] ;
  assign \A_s[47]  = A_s[47];
  assign A_so[48] = \A_s[46] ;
  assign \A_s[46]  = A_s[46];
  assign A_so[47] = \A_s[45] ;
  assign \A_s[45]  = A_s[45];
  assign A_so[46] = \A_s[44] ;
  assign \A_s[44]  = A_s[44];
  assign A_so[45] = \A_s[43] ;
  assign \A_s[43]  = A_s[43];
  assign A_so[44] = \A_s[42] ;
  assign \A_s[42]  = A_s[42];
  assign A_so[43] = \A_s[41] ;
  assign \A_s[41]  = A_s[41];
  assign A_so[42] = \A_s[40] ;
  assign \A_s[40]  = A_s[40];
  assign A_so[41] = \A_s[39] ;
  assign \A_s[39]  = A_s[39];
  assign A_so[40] = \A_s[38] ;
  assign \A_s[38]  = A_s[38];
  assign A_so[39] = \A_s[37] ;
  assign \A_s[37]  = A_s[37];
  assign A_so[38] = \A_s[36] ;
  assign \A_s[36]  = A_s[36];
  assign A_so[37] = \A_s[35] ;
  assign \A_s[35]  = A_s[35];
  assign A_so[36] = \A_s[34] ;
  assign \A_s[34]  = A_s[34];
  assign A_so[35] = \A_s[33] ;
  assign \A_s[33]  = A_s[33];
  assign A_so[34] = \A_s[32] ;
  assign \A_s[32]  = A_s[32];
  assign A_so[33] = \A_s[31] ;
  assign \A_s[31]  = A_s[31];
  assign A_so[32] = \A_s[30] ;
  assign \A_s[30]  = A_s[30];
  assign A_so[31] = \A_s[29] ;
  assign \A_s[29]  = A_s[29];
  assign A_so[30] = \A_s[28] ;
  assign \A_s[28]  = A_s[28];
  assign A_so[29] = \A_s[27] ;
  assign \A_s[27]  = A_s[27];
  assign A_so[28] = \A_s[26] ;
  assign \A_s[26]  = A_s[26];
  assign A_so[27] = \A_s[25] ;
  assign \A_s[25]  = A_s[25];
  assign A_so[26] = \A_s[24] ;
  assign \A_s[24]  = A_s[24];
  assign A_so[25] = \A_s[23] ;
  assign \A_s[23]  = A_s[23];
  assign A_so[24] = \A_s[22] ;
  assign \A_s[22]  = A_s[22];
  assign A_so[23] = \A_s[21] ;
  assign \A_s[21]  = A_s[21];
  assign A_so[22] = \A_s[20] ;
  assign \A_s[20]  = A_s[20];
  assign A_so[21] = \A_s[19] ;
  assign \A_s[19]  = A_s[19];
  assign A_so[20] = \A_s[18] ;
  assign \A_s[18]  = A_s[18];
  assign A_so[19] = \A_s[17] ;
  assign \A_s[17]  = A_s[17];
  assign A_so[18] = \A_s[16] ;
  assign \A_s[16]  = A_s[16];
  assign A_so[17] = \A_s[15] ;
  assign \A_s[15]  = A_s[15];
  assign A_so[16] = \A_s[14] ;
  assign \A_s[14]  = A_s[14];
  assign A_so[15] = \A_s[13] ;
  assign \A_s[13]  = A_s[13];
  assign A_so[14] = \A_s[12] ;
  assign \A_s[12]  = A_s[12];
  assign A_so[13] = \A_s[11] ;
  assign \A_s[11]  = A_s[11];
  assign A_so[12] = \A_s[10] ;
  assign \A_s[10]  = A_s[10];
  assign A_so[11] = \A_s[9] ;
  assign \A_s[9]  = A_s[9];
  assign A_so[10] = \A_s[8] ;
  assign \A_s[8]  = A_s[8];
  assign A_so[9] = \A_s[7] ;
  assign \A_s[7]  = A_s[7];
  assign A_so[8] = \A_s[6] ;
  assign \A_s[6]  = A_s[6];
  assign A_so[7] = \A_s[5] ;
  assign \A_s[5]  = A_s[5];
  assign A_so[6] = \A_s[4] ;
  assign \A_s[4]  = A_s[4];
  assign A_so[5] = \A_s[3] ;
  assign \A_s[3]  = A_s[3];
  assign A_so[4] = \A_s[2] ;
  assign \A_s[2]  = A_s[2];
  assign A_so[3] = \A_s[1] ;
  assign \A_s[1]  = A_s[1];
  assign A_so[2] = \A_s[0] ;
  assign \A_s[0]  = A_s[0];
  assign A_nso[63] = \A_ns[61] ;
  assign \A_ns[61]  = A_ns[61];
  assign A_nso[62] = \A_ns[60] ;
  assign \A_ns[60]  = A_ns[60];
  assign A_nso[61] = \A_ns[59] ;
  assign \A_ns[59]  = A_ns[59];
  assign A_nso[60] = \A_ns[58] ;
  assign \A_ns[58]  = A_ns[58];
  assign A_nso[59] = \A_ns[57] ;
  assign \A_ns[57]  = A_ns[57];
  assign A_nso[58] = \A_ns[56] ;
  assign \A_ns[56]  = A_ns[56];
  assign A_nso[57] = \A_ns[55] ;
  assign \A_ns[55]  = A_ns[55];
  assign A_nso[56] = \A_ns[54] ;
  assign \A_ns[54]  = A_ns[54];
  assign A_nso[55] = \A_ns[53] ;
  assign \A_ns[53]  = A_ns[53];
  assign A_nso[54] = \A_ns[52] ;
  assign \A_ns[52]  = A_ns[52];
  assign A_nso[53] = \A_ns[51] ;
  assign \A_ns[51]  = A_ns[51];
  assign A_nso[52] = \A_ns[50] ;
  assign \A_ns[50]  = A_ns[50];
  assign A_nso[51] = \A_ns[49] ;
  assign \A_ns[49]  = A_ns[49];
  assign A_nso[50] = \A_ns[48] ;
  assign \A_ns[48]  = A_ns[48];
  assign A_nso[49] = \A_ns[47] ;
  assign \A_ns[47]  = A_ns[47];
  assign A_nso[48] = \A_ns[46] ;
  assign \A_ns[46]  = A_ns[46];
  assign A_nso[47] = \A_ns[45] ;
  assign \A_ns[45]  = A_ns[45];
  assign A_nso[46] = \A_ns[44] ;
  assign \A_ns[44]  = A_ns[44];
  assign A_nso[45] = \A_ns[43] ;
  assign \A_ns[43]  = A_ns[43];
  assign A_nso[44] = \A_ns[42] ;
  assign \A_ns[42]  = A_ns[42];
  assign A_nso[43] = \A_ns[41] ;
  assign \A_ns[41]  = A_ns[41];
  assign A_nso[42] = \A_ns[40] ;
  assign \A_ns[40]  = A_ns[40];
  assign A_nso[41] = \A_ns[39] ;
  assign \A_ns[39]  = A_ns[39];
  assign A_nso[40] = \A_ns[38] ;
  assign \A_ns[38]  = A_ns[38];
  assign A_nso[39] = \A_ns[37] ;
  assign \A_ns[37]  = A_ns[37];
  assign A_nso[38] = \A_ns[36] ;
  assign \A_ns[36]  = A_ns[36];
  assign A_nso[37] = \A_ns[35] ;
  assign \A_ns[35]  = A_ns[35];
  assign A_nso[36] = \A_ns[34] ;
  assign \A_ns[34]  = A_ns[34];
  assign A_nso[35] = \A_ns[33] ;
  assign \A_ns[33]  = A_ns[33];
  assign A_nso[34] = \A_ns[32] ;
  assign \A_ns[32]  = A_ns[32];
  assign A_nso[33] = \A_ns[31] ;
  assign \A_ns[31]  = A_ns[31];
  assign A_nso[32] = \A_ns[30] ;
  assign \A_ns[30]  = A_ns[30];
  assign A_nso[31] = \A_ns[29] ;
  assign \A_ns[29]  = A_ns[29];
  assign A_nso[30] = \A_ns[28] ;
  assign \A_ns[28]  = A_ns[28];
  assign A_nso[29] = \A_ns[27] ;
  assign \A_ns[27]  = A_ns[27];
  assign A_nso[28] = \A_ns[26] ;
  assign \A_ns[26]  = A_ns[26];
  assign A_nso[27] = \A_ns[25] ;
  assign \A_ns[25]  = A_ns[25];
  assign A_nso[26] = \A_ns[24] ;
  assign \A_ns[24]  = A_ns[24];
  assign A_nso[25] = \A_ns[23] ;
  assign \A_ns[23]  = A_ns[23];
  assign A_nso[24] = \A_ns[22] ;
  assign \A_ns[22]  = A_ns[22];
  assign A_nso[23] = \A_ns[21] ;
  assign \A_ns[21]  = A_ns[21];
  assign A_nso[22] = \A_ns[20] ;
  assign \A_ns[20]  = A_ns[20];
  assign A_nso[21] = \A_ns[19] ;
  assign \A_ns[19]  = A_ns[19];
  assign A_nso[20] = \A_ns[18] ;
  assign \A_ns[18]  = A_ns[18];
  assign A_nso[19] = \A_ns[17] ;
  assign \A_ns[17]  = A_ns[17];
  assign A_nso[18] = \A_ns[16] ;
  assign \A_ns[16]  = A_ns[16];
  assign A_nso[17] = \A_ns[15] ;
  assign \A_ns[15]  = A_ns[15];
  assign A_nso[16] = \A_ns[14] ;
  assign \A_ns[14]  = A_ns[14];
  assign A_nso[15] = \A_ns[13] ;
  assign \A_ns[13]  = A_ns[13];
  assign A_nso[14] = \A_ns[12] ;
  assign \A_ns[12]  = A_ns[12];
  assign A_nso[13] = \A_ns[11] ;
  assign \A_ns[11]  = A_ns[11];
  assign A_nso[12] = \A_ns[10] ;
  assign \A_ns[10]  = A_ns[10];
  assign A_nso[11] = \A_ns[9] ;
  assign \A_ns[9]  = A_ns[9];
  assign A_nso[10] = \A_ns[8] ;
  assign \A_ns[8]  = A_ns[8];
  assign A_nso[9] = \A_ns[7] ;
  assign \A_ns[7]  = A_ns[7];
  assign A_nso[8] = \A_ns[6] ;
  assign \A_ns[6]  = A_ns[6];
  assign A_nso[7] = \A_ns[5] ;
  assign \A_ns[5]  = A_ns[5];
  assign A_nso[6] = \A_ns[4] ;
  assign \A_ns[4]  = A_ns[4];
  assign A_nso[5] = \A_ns[3] ;
  assign \A_ns[3]  = A_ns[3];
  assign A_nso[4] = \A_ns[2] ;
  assign \A_ns[2]  = A_ns[2];
  assign A_nso[3] = \A_ns[1] ;
  assign \A_ns[1]  = A_ns[1];
  assign A_nso[2] = \A_ns[0] ;
  assign \A_ns[0]  = A_ns[0];

  XOR2_X1 U257 ( .A(B[29]), .B(B[30]), .Z(n194) );
  NAND3_X1 U258 ( .A1(B[30]), .A2(n889), .A3(B[29]), .ZN(n129) );
  OAI221_X1 U2 ( .B1(n757), .B2(n788), .C1(n755), .C2(n822), .A(n141), .ZN(
        O[57]) );
  AOI22_X1 U3 ( .A1(A_ns[62]), .A2(n748), .B1(A_s[62]), .B2(n742), .ZN(n134)
         );
  BUF_X1 U4 ( .A(n888), .Z(n745) );
  BUF_X1 U5 ( .A(n888), .Z(n746) );
  BUF_X1 U6 ( .A(n887), .Z(n739) );
  BUF_X1 U7 ( .A(n887), .Z(n740) );
  BUF_X1 U8 ( .A(n888), .Z(n747) );
  BUF_X1 U9 ( .A(n887), .Z(n741) );
  BUF_X1 U10 ( .A(n887), .Z(n742) );
  BUF_X1 U11 ( .A(n888), .Z(n748) );
  BUF_X1 U12 ( .A(n888), .Z(n744) );
  BUF_X1 U13 ( .A(n887), .Z(n738) );
  OAI221_X1 U14 ( .B1(n757), .B2(n794), .C1(n756), .C2(n828), .A(n134), .ZN(
        O[63]) );
  OAI221_X1 U15 ( .B1(n760), .B2(n795), .C1(n753), .C2(n796), .A(n169), .ZN(
        O[31]) );
  AOI22_X1 U16 ( .A1(\A_ns[30] ), .A2(n745), .B1(\A_s[30] ), .B2(n739), .ZN(
        n169) );
  OAI221_X1 U17 ( .B1(n760), .B2(n763), .C1(n753), .C2(n797), .A(n168), .ZN(
        O[32]) );
  AOI22_X1 U18 ( .A1(\A_ns[31] ), .A2(n745), .B1(\A_s[31] ), .B2(n739), .ZN(
        n168) );
  OAI221_X1 U19 ( .B1(n760), .B2(n765), .C1(n753), .C2(n799), .A(n166), .ZN(
        O[34]) );
  AOI22_X1 U20 ( .A1(\A_ns[33] ), .A2(n746), .B1(\A_s[33] ), .B2(n740), .ZN(
        n166) );
  OAI221_X1 U21 ( .B1(n759), .B2(n767), .C1(n754), .C2(n801), .A(n164), .ZN(
        O[36]) );
  AOI22_X1 U22 ( .A1(\A_ns[35] ), .A2(n746), .B1(\A_s[35] ), .B2(n740), .ZN(
        n164) );
  OAI221_X1 U23 ( .B1(n759), .B2(n769), .C1(n754), .C2(n803), .A(n162), .ZN(
        O[38]) );
  AOI22_X1 U24 ( .A1(\A_ns[37] ), .A2(n746), .B1(\A_s[37] ), .B2(n740), .ZN(
        n162) );
  OAI221_X1 U25 ( .B1(n760), .B2(n764), .C1(n753), .C2(n798), .A(n167), .ZN(
        O[33]) );
  AOI22_X1 U26 ( .A1(\A_ns[32] ), .A2(n746), .B1(\A_s[32] ), .B2(n740), .ZN(
        n167) );
  OAI221_X1 U27 ( .B1(n759), .B2(n768), .C1(n754), .C2(n802), .A(n163), .ZN(
        O[37]) );
  AOI22_X1 U28 ( .A1(\A_ns[36] ), .A2(n746), .B1(\A_s[36] ), .B2(n740), .ZN(
        n163) );
  OAI221_X1 U29 ( .B1(n759), .B2(n770), .C1(n754), .C2(n804), .A(n161), .ZN(
        O[39]) );
  AOI22_X1 U30 ( .A1(\A_ns[38] ), .A2(n746), .B1(\A_s[38] ), .B2(n740), .ZN(
        n161) );
  OAI221_X1 U31 ( .B1(n759), .B2(n773), .C1(n754), .C2(n807), .A(n157), .ZN(
        O[42]) );
  AOI22_X1 U32 ( .A1(\A_ns[41] ), .A2(n746), .B1(\A_s[41] ), .B2(n740), .ZN(
        n157) );
  OAI221_X1 U33 ( .B1(n759), .B2(n766), .C1(n754), .C2(n800), .A(n165), .ZN(
        O[35]) );
  AOI22_X1 U34 ( .A1(\A_ns[34] ), .A2(n746), .B1(\A_s[34] ), .B2(n740), .ZN(
        n165) );
  OAI221_X1 U35 ( .B1(n759), .B2(n772), .C1(n754), .C2(n806), .A(n158), .ZN(
        O[41]) );
  AOI22_X1 U36 ( .A1(\A_ns[40] ), .A2(n746), .B1(\A_s[40] ), .B2(n740), .ZN(
        n158) );
  OAI221_X1 U37 ( .B1(n759), .B2(n774), .C1(n754), .C2(n808), .A(n156), .ZN(
        O[43]) );
  AOI22_X1 U38 ( .A1(\A_ns[42] ), .A2(n746), .B1(\A_s[42] ), .B2(n740), .ZN(
        n156) );
  OAI221_X1 U39 ( .B1(n759), .B2(n771), .C1(n754), .C2(n805), .A(n159), .ZN(
        O[40]) );
  AOI22_X1 U40 ( .A1(\A_ns[39] ), .A2(n746), .B1(\A_s[39] ), .B2(n740), .ZN(
        n159) );
  BUF_X1 U41 ( .A(n750), .Z(n753) );
  OAI221_X1 U42 ( .B1(n759), .B2(n775), .C1(n754), .C2(n809), .A(n155), .ZN(
        O[44]) );
  AOI22_X1 U43 ( .A1(\A_ns[43] ), .A2(n747), .B1(\A_s[43] ), .B2(n741), .ZN(
        n155) );
  OAI221_X1 U44 ( .B1(n759), .B2(n776), .C1(n754), .C2(n810), .A(n154), .ZN(
        O[45]) );
  AOI22_X1 U45 ( .A1(\A_ns[44] ), .A2(n747), .B1(\A_s[44] ), .B2(n741), .ZN(
        n154) );
  INV_X1 U46 ( .A(n183), .ZN(n888) );
  INV_X1 U47 ( .A(n182), .ZN(n887) );
  AOI22_X1 U48 ( .A1(\A_ns[56] ), .A2(n748), .B1(\A_s[56] ), .B2(n742), .ZN(
        n141) );
  OAI221_X1 U49 ( .B1(n757), .B2(n792), .C1(n756), .C2(n826), .A(n136), .ZN(
        O[61]) );
  AOI22_X1 U50 ( .A1(\A_ns[60] ), .A2(n748), .B1(\A_s[60] ), .B2(n742), .ZN(
        n136) );
  OAI221_X1 U51 ( .B1(n757), .B2(n790), .C1(n756), .C2(n824), .A(n139), .ZN(
        O[59]) );
  AOI22_X1 U52 ( .A1(\A_ns[58] ), .A2(n748), .B1(\A_s[58] ), .B2(n742), .ZN(
        n139) );
  OAI221_X1 U53 ( .B1(n758), .B2(n779), .C1(n755), .C2(n813), .A(n151), .ZN(
        O[48]) );
  AOI22_X1 U54 ( .A1(\A_ns[47] ), .A2(n747), .B1(\A_s[47] ), .B2(n741), .ZN(
        n151) );
  OAI221_X1 U55 ( .B1(n758), .B2(n780), .C1(n755), .C2(n814), .A(n150), .ZN(
        O[49]) );
  AOI22_X1 U56 ( .A1(\A_ns[48] ), .A2(n747), .B1(\A_s[48] ), .B2(n741), .ZN(
        n150) );
  OAI221_X1 U57 ( .B1(n758), .B2(n777), .C1(n754), .C2(n811), .A(n153), .ZN(
        O[46]) );
  AOI22_X1 U58 ( .A1(\A_ns[45] ), .A2(n747), .B1(\A_s[45] ), .B2(n741), .ZN(
        n153) );
  BUF_X1 U59 ( .A(n750), .Z(n754) );
  OAI221_X1 U60 ( .B1(n758), .B2(n778), .C1(n755), .C2(n812), .A(n152), .ZN(
        O[47]) );
  AOI22_X1 U61 ( .A1(\A_ns[46] ), .A2(n747), .B1(\A_s[46] ), .B2(n741), .ZN(
        n152) );
  OAI221_X1 U62 ( .B1(n758), .B2(n781), .C1(n755), .C2(n815), .A(n148), .ZN(
        O[50]) );
  AOI22_X1 U63 ( .A1(\A_ns[49] ), .A2(n747), .B1(\A_s[49] ), .B2(n741), .ZN(
        n148) );
  OAI221_X1 U64 ( .B1(n758), .B2(n782), .C1(n755), .C2(n816), .A(n147), .ZN(
        O[51]) );
  AOI22_X1 U65 ( .A1(\A_ns[50] ), .A2(n747), .B1(\A_s[50] ), .B2(n741), .ZN(
        n147) );
  OAI221_X1 U66 ( .B1(n758), .B2(n783), .C1(n755), .C2(n817), .A(n146), .ZN(
        O[52]) );
  AOI22_X1 U67 ( .A1(\A_ns[51] ), .A2(n747), .B1(\A_s[51] ), .B2(n741), .ZN(
        n146) );
  OAI221_X1 U68 ( .B1(n758), .B2(n784), .C1(n755), .C2(n818), .A(n145), .ZN(
        O[53]) );
  AOI22_X1 U69 ( .A1(\A_ns[52] ), .A2(n747), .B1(\A_s[52] ), .B2(n741), .ZN(
        n145) );
  OAI221_X1 U70 ( .B1(n758), .B2(n785), .C1(n755), .C2(n819), .A(n144), .ZN(
        O[54]) );
  AOI22_X1 U71 ( .A1(\A_ns[53] ), .A2(n747), .B1(\A_s[53] ), .B2(n741), .ZN(
        n144) );
  OAI221_X1 U72 ( .B1(n758), .B2(n786), .C1(n755), .C2(n820), .A(n143), .ZN(
        O[55]) );
  AOI22_X1 U73 ( .A1(\A_ns[54] ), .A2(n748), .B1(\A_s[54] ), .B2(n742), .ZN(
        n143) );
  OAI221_X1 U74 ( .B1(n758), .B2(n787), .C1(n755), .C2(n821), .A(n142), .ZN(
        O[56]) );
  AOI22_X1 U75 ( .A1(\A_ns[55] ), .A2(n748), .B1(\A_s[55] ), .B2(n742), .ZN(
        n142) );
  OAI221_X1 U76 ( .B1(n757), .B2(n789), .C1(n755), .C2(n823), .A(n140), .ZN(
        O[58]) );
  AOI22_X1 U77 ( .A1(\A_ns[57] ), .A2(n748), .B1(\A_s[57] ), .B2(n742), .ZN(
        n140) );
  OAI221_X1 U78 ( .B1(n757), .B2(n791), .C1(n756), .C2(n825), .A(n137), .ZN(
        O[60]) );
  AOI22_X1 U79 ( .A1(\A_ns[59] ), .A2(n748), .B1(\A_s[59] ), .B2(n742), .ZN(
        n137) );
  OAI221_X1 U80 ( .B1(n757), .B2(n793), .C1(n756), .C2(n827), .A(n135), .ZN(
        O[62]) );
  AOI22_X1 U81 ( .A1(\A_ns[61] ), .A2(n748), .B1(\A_s[61] ), .B2(n742), .ZN(
        n135) );
  BUF_X1 U82 ( .A(n751), .Z(n755) );
  BUF_X1 U83 ( .A(n751), .Z(n756) );
  BUF_X1 U84 ( .A(n750), .Z(n752) );
  BUF_X1 U85 ( .A(n128), .Z(n760) );
  NAND2_X1 U86 ( .A1(n194), .A2(n889), .ZN(n182) );
  NAND2_X1 U87 ( .A1(n194), .A2(n182), .ZN(n183) );
  BUF_X1 U88 ( .A(n129), .Z(n750) );
  BUF_X1 U89 ( .A(n128), .Z(n759) );
  BUF_X1 U90 ( .A(n128), .Z(n758) );
  BUF_X1 U91 ( .A(n129), .Z(n751) );
  BUF_X1 U92 ( .A(n128), .Z(n757) );
  BUF_X1 U93 ( .A(n128), .Z(n761) );
  OAI221_X1 U94 ( .B1(n760), .B2(n881), .C1(n753), .C2(n883), .A(n173), .ZN(
        O[28]) );
  INV_X1 U95 ( .A(\A_ns[26] ), .ZN(n881) );
  INV_X1 U96 ( .A(\A_s[26] ), .ZN(n883) );
  OAI221_X1 U97 ( .B1(n760), .B2(n885), .C1(n753), .C2(n886), .A(n170), .ZN(
        O[30]) );
  INV_X1 U98 ( .A(\A_ns[28] ), .ZN(n885) );
  INV_X1 U99 ( .A(\A_s[28] ), .ZN(n886) );
  AOI22_X1 U100 ( .A1(\A_ns[29] ), .A2(n745), .B1(\A_s[29] ), .B2(n739), .ZN(
        n170) );
  OAI221_X1 U101 ( .B1(n761), .B2(n866), .C1(n752), .C2(n868), .A(n180), .ZN(
        O[21]) );
  INV_X1 U102 ( .A(\A_ns[19] ), .ZN(n866) );
  INV_X1 U103 ( .A(\A_s[19] ), .ZN(n868) );
  OAI221_X1 U104 ( .B1(n761), .B2(n869), .C1(n752), .C2(n871), .A(n179), .ZN(
        O[22]) );
  INV_X1 U105 ( .A(\A_ns[20] ), .ZN(n869) );
  INV_X1 U106 ( .A(\A_s[20] ), .ZN(n871) );
  OAI221_X1 U107 ( .B1(n761), .B2(n870), .C1(n753), .C2(n872), .A(n178), .ZN(
        O[23]) );
  INV_X1 U108 ( .A(\A_ns[21] ), .ZN(n870) );
  INV_X1 U109 ( .A(\A_s[21] ), .ZN(n872) );
  OAI221_X1 U110 ( .B1(n760), .B2(n873), .C1(n753), .C2(n875), .A(n177), .ZN(
        O[24]) );
  INV_X1 U111 ( .A(\A_ns[22] ), .ZN(n873) );
  INV_X1 U112 ( .A(\A_s[22] ), .ZN(n875) );
  OAI221_X1 U113 ( .B1(n760), .B2(n874), .C1(n753), .C2(n876), .A(n176), .ZN(
        O[25]) );
  INV_X1 U114 ( .A(\A_ns[23] ), .ZN(n874) );
  INV_X1 U115 ( .A(\A_s[23] ), .ZN(n876) );
  OAI221_X1 U116 ( .B1(n760), .B2(n877), .C1(n753), .C2(n879), .A(n175), .ZN(
        O[26]) );
  INV_X1 U117 ( .A(\A_ns[24] ), .ZN(n877) );
  INV_X1 U118 ( .A(\A_s[24] ), .ZN(n879) );
  OAI221_X1 U119 ( .B1(n760), .B2(n878), .C1(n753), .C2(n880), .A(n174), .ZN(
        O[27]) );
  INV_X1 U120 ( .A(\A_ns[25] ), .ZN(n878) );
  INV_X1 U121 ( .A(\A_s[25] ), .ZN(n880) );
  OR3_X1 U122 ( .A1(B[29]), .A2(B[30]), .A3(n889), .ZN(n128) );
  INV_X1 U123 ( .A(B[31]), .ZN(n889) );
  OAI221_X1 U124 ( .B1(n761), .B2(n854), .C1(n752), .C2(n856), .A(n188), .ZN(
        O[15]) );
  INV_X1 U125 ( .A(\A_ns[13] ), .ZN(n854) );
  INV_X1 U126 ( .A(\A_s[13] ), .ZN(n856) );
  OAI221_X1 U127 ( .B1(n761), .B2(n857), .C1(n752), .C2(n859), .A(n187), .ZN(
        O[16]) );
  INV_X1 U128 ( .A(\A_ns[14] ), .ZN(n857) );
  INV_X1 U129 ( .A(\A_s[14] ), .ZN(n859) );
  OAI221_X1 U130 ( .B1(n761), .B2(n858), .C1(n752), .C2(n860), .A(n186), .ZN(
        O[17]) );
  INV_X1 U131 ( .A(\A_ns[15] ), .ZN(n858) );
  INV_X1 U132 ( .A(\A_s[15] ), .ZN(n860) );
  OAI221_X1 U133 ( .B1(n761), .B2(n861), .C1(n752), .C2(n863), .A(n185), .ZN(
        O[18]) );
  INV_X1 U134 ( .A(\A_ns[16] ), .ZN(n861) );
  INV_X1 U135 ( .A(\A_s[16] ), .ZN(n863) );
  OAI221_X1 U136 ( .B1(n761), .B2(n862), .C1(n752), .C2(n864), .A(n184), .ZN(
        O[19]) );
  INV_X1 U137 ( .A(\A_ns[17] ), .ZN(n862) );
  INV_X1 U138 ( .A(\A_s[17] ), .ZN(n864) );
  OAI221_X1 U139 ( .B1(n761), .B2(n865), .C1(n752), .C2(n867), .A(n181), .ZN(
        O[20]) );
  INV_X1 U140 ( .A(\A_ns[18] ), .ZN(n865) );
  INV_X1 U141 ( .A(\A_s[18] ), .ZN(n867) );
  OAI221_X1 U142 ( .B1(n757), .B2(n838), .C1(n756), .C2(n840), .A(n132), .ZN(
        O[7]) );
  INV_X1 U143 ( .A(\A_ns[5] ), .ZN(n838) );
  INV_X1 U144 ( .A(\A_s[5] ), .ZN(n840) );
  OAI221_X1 U145 ( .B1(n757), .B2(n841), .C1(n756), .C2(n843), .A(n131), .ZN(
        O[8]) );
  INV_X1 U146 ( .A(\A_ns[6] ), .ZN(n841) );
  INV_X1 U147 ( .A(\A_s[6] ), .ZN(n843) );
  OAI221_X1 U148 ( .B1(n757), .B2(n842), .C1(n756), .C2(n844), .A(n130), .ZN(
        O[9]) );
  INV_X1 U149 ( .A(\A_ns[7] ), .ZN(n842) );
  INV_X1 U150 ( .A(\A_s[7] ), .ZN(n844) );
  OAI221_X1 U151 ( .B1(n845), .B2(n762), .C1(n847), .C2(n752), .A(n193), .ZN(
        O[10]) );
  INV_X1 U152 ( .A(\A_s[8] ), .ZN(n847) );
  INV_X1 U153 ( .A(\A_ns[8] ), .ZN(n845) );
  OAI221_X1 U154 ( .B1(n762), .B2(n846), .C1(n752), .C2(n848), .A(n192), .ZN(
        O[11]) );
  INV_X1 U155 ( .A(\A_ns[9] ), .ZN(n846) );
  INV_X1 U156 ( .A(\A_s[9] ), .ZN(n848) );
  OAI221_X1 U157 ( .B1(n761), .B2(n849), .C1(n752), .C2(n851), .A(n191), .ZN(
        O[12]) );
  INV_X1 U158 ( .A(\A_ns[10] ), .ZN(n849) );
  INV_X1 U159 ( .A(\A_s[10] ), .ZN(n851) );
  OAI221_X1 U160 ( .B1(n761), .B2(n850), .C1(n752), .C2(n852), .A(n190), .ZN(
        O[13]) );
  INV_X1 U161 ( .A(\A_ns[11] ), .ZN(n850) );
  INV_X1 U162 ( .A(\A_s[11] ), .ZN(n852) );
  OAI221_X1 U163 ( .B1(n761), .B2(n853), .C1(n752), .C2(n855), .A(n189), .ZN(
        O[14]) );
  INV_X1 U164 ( .A(\A_ns[12] ), .ZN(n853) );
  INV_X1 U165 ( .A(\A_s[12] ), .ZN(n855) );
  OAI22_X1 U166 ( .A1(n182), .A2(n831), .B1(n183), .B2(n829), .ZN(O[1]) );
  OAI221_X1 U167 ( .B1(n760), .B2(n829), .C1(n753), .C2(n831), .A(n171), .ZN(
        O[2]) );
  AOI22_X1 U168 ( .A1(\A_ns[1] ), .A2(n745), .B1(\A_s[1] ), .B2(n739), .ZN(
        n171) );
  OAI221_X1 U169 ( .B1(n759), .B2(n830), .C1(n754), .C2(n832), .A(n160), .ZN(
        O[3]) );
  INV_X1 U170 ( .A(\A_ns[1] ), .ZN(n830) );
  INV_X1 U171 ( .A(\A_s[1] ), .ZN(n832) );
  OAI221_X1 U172 ( .B1(n758), .B2(n833), .C1(n755), .C2(n835), .A(n149), .ZN(
        O[4]) );
  INV_X1 U173 ( .A(\A_ns[2] ), .ZN(n833) );
  INV_X1 U174 ( .A(\A_s[2] ), .ZN(n835) );
  OAI221_X1 U175 ( .B1(n757), .B2(n834), .C1(n756), .C2(n836), .A(n138), .ZN(
        O[5]) );
  INV_X1 U176 ( .A(\A_ns[3] ), .ZN(n834) );
  INV_X1 U177 ( .A(\A_s[3] ), .ZN(n836) );
  OAI221_X1 U178 ( .B1(n757), .B2(n837), .C1(n756), .C2(n839), .A(n133), .ZN(
        O[6]) );
  INV_X1 U179 ( .A(\A_ns[4] ), .ZN(n837) );
  INV_X1 U180 ( .A(\A_s[4] ), .ZN(n839) );
  OAI221_X1 U181 ( .B1(n760), .B2(n882), .C1(n753), .C2(n884), .A(n172), .ZN(
        O[29]) );
  INV_X1 U182 ( .A(\A_ns[27] ), .ZN(n882) );
  INV_X1 U183 ( .A(\A_s[27] ), .ZN(n884) );
  AOI22_X1 U184 ( .A1(\A_ns[28] ), .A2(n745), .B1(\A_s[28] ), .B2(n739), .ZN(
        n172) );
  INV_X1 U185 ( .A(\A_s[0] ), .ZN(n831) );
  INV_X1 U186 ( .A(\A_ns[0] ), .ZN(n829) );
  AOI22_X1 U187 ( .A1(\A_ns[2] ), .A2(n746), .B1(\A_s[2] ), .B2(n740), .ZN(
        n160) );
  AOI22_X1 U188 ( .A1(\A_ns[3] ), .A2(n747), .B1(\A_s[3] ), .B2(n741), .ZN(
        n149) );
  AOI22_X1 U189 ( .A1(\A_ns[4] ), .A2(n748), .B1(\A_s[4] ), .B2(n742), .ZN(
        n138) );
  AOI22_X1 U190 ( .A1(\A_ns[5] ), .A2(n748), .B1(\A_s[5] ), .B2(n742), .ZN(
        n133) );
  AOI22_X1 U191 ( .A1(\A_ns[6] ), .A2(n748), .B1(\A_s[6] ), .B2(n742), .ZN(
        n132) );
  AOI22_X1 U192 ( .A1(\A_ns[7] ), .A2(n749), .B1(\A_s[7] ), .B2(n743), .ZN(
        n131) );
  AOI22_X1 U193 ( .A1(\A_ns[8] ), .A2(n749), .B1(\A_s[8] ), .B2(n743), .ZN(
        n130) );
  AOI22_X1 U194 ( .A1(\A_ns[9] ), .A2(n744), .B1(\A_s[9] ), .B2(n738), .ZN(
        n193) );
  AOI22_X1 U195 ( .A1(\A_ns[10] ), .A2(n744), .B1(\A_s[10] ), .B2(n738), .ZN(
        n192) );
  AOI22_X1 U196 ( .A1(\A_ns[11] ), .A2(n744), .B1(\A_s[11] ), .B2(n738), .ZN(
        n191) );
  AOI22_X1 U197 ( .A1(\A_ns[12] ), .A2(n744), .B1(\A_s[12] ), .B2(n738), .ZN(
        n190) );
  AOI22_X1 U198 ( .A1(\A_ns[13] ), .A2(n744), .B1(\A_s[13] ), .B2(n738), .ZN(
        n189) );
  AOI22_X1 U199 ( .A1(\A_ns[14] ), .A2(n744), .B1(\A_s[14] ), .B2(n738), .ZN(
        n188) );
  AOI22_X1 U200 ( .A1(\A_ns[15] ), .A2(n744), .B1(\A_s[15] ), .B2(n738), .ZN(
        n187) );
  AOI22_X1 U201 ( .A1(\A_ns[16] ), .A2(n744), .B1(\A_s[16] ), .B2(n738), .ZN(
        n186) );
  AOI22_X1 U202 ( .A1(\A_ns[17] ), .A2(n744), .B1(\A_s[17] ), .B2(n738), .ZN(
        n185) );
  AOI22_X1 U203 ( .A1(\A_ns[18] ), .A2(n744), .B1(\A_s[18] ), .B2(n738), .ZN(
        n184) );
  AOI22_X1 U204 ( .A1(\A_ns[19] ), .A2(n744), .B1(\A_s[19] ), .B2(n738), .ZN(
        n181) );
  AOI22_X1 U205 ( .A1(\A_ns[20] ), .A2(n744), .B1(\A_s[20] ), .B2(n738), .ZN(
        n180) );
  AOI22_X1 U206 ( .A1(\A_ns[21] ), .A2(n745), .B1(\A_s[21] ), .B2(n739), .ZN(
        n179) );
  AOI22_X1 U207 ( .A1(\A_ns[22] ), .A2(n745), .B1(\A_s[22] ), .B2(n739), .ZN(
        n178) );
  AOI22_X1 U208 ( .A1(\A_ns[23] ), .A2(n745), .B1(\A_s[23] ), .B2(n739), .ZN(
        n177) );
  AOI22_X1 U209 ( .A1(\A_ns[24] ), .A2(n745), .B1(\A_s[24] ), .B2(n739), .ZN(
        n176) );
  AOI22_X1 U210 ( .A1(\A_ns[25] ), .A2(n745), .B1(\A_s[25] ), .B2(n739), .ZN(
        n175) );
  AOI22_X1 U211 ( .A1(\A_ns[26] ), .A2(n745), .B1(\A_s[26] ), .B2(n739), .ZN(
        n174) );
  AOI22_X1 U212 ( .A1(\A_ns[27] ), .A2(n745), .B1(\A_s[27] ), .B2(n739), .ZN(
        n173) );
  CLKBUF_X1 U213 ( .A(n887), .Z(n743) );
  CLKBUF_X1 U214 ( .A(n888), .Z(n749) );
  CLKBUF_X1 U215 ( .A(n128), .Z(n762) );
  INV_X1 U216 ( .A(\A_ns[30] ), .ZN(n763) );
  INV_X1 U217 ( .A(\A_ns[31] ), .ZN(n764) );
  INV_X1 U218 ( .A(\A_ns[32] ), .ZN(n765) );
  INV_X1 U219 ( .A(\A_ns[33] ), .ZN(n766) );
  INV_X1 U220 ( .A(\A_ns[34] ), .ZN(n767) );
  INV_X1 U221 ( .A(\A_ns[35] ), .ZN(n768) );
  INV_X1 U222 ( .A(\A_ns[36] ), .ZN(n769) );
  INV_X1 U223 ( .A(\A_ns[37] ), .ZN(n770) );
  INV_X1 U224 ( .A(\A_ns[38] ), .ZN(n771) );
  INV_X1 U225 ( .A(\A_ns[39] ), .ZN(n772) );
  INV_X1 U226 ( .A(\A_ns[40] ), .ZN(n773) );
  INV_X1 U227 ( .A(\A_ns[41] ), .ZN(n774) );
  INV_X1 U228 ( .A(\A_ns[42] ), .ZN(n775) );
  INV_X1 U229 ( .A(\A_ns[43] ), .ZN(n776) );
  INV_X1 U230 ( .A(\A_ns[44] ), .ZN(n777) );
  INV_X1 U231 ( .A(\A_ns[45] ), .ZN(n778) );
  INV_X1 U232 ( .A(\A_ns[46] ), .ZN(n779) );
  INV_X1 U233 ( .A(\A_ns[47] ), .ZN(n780) );
  INV_X1 U234 ( .A(\A_ns[48] ), .ZN(n781) );
  INV_X1 U235 ( .A(\A_ns[49] ), .ZN(n782) );
  INV_X1 U236 ( .A(\A_ns[50] ), .ZN(n783) );
  INV_X1 U237 ( .A(\A_ns[51] ), .ZN(n784) );
  INV_X1 U238 ( .A(\A_ns[52] ), .ZN(n785) );
  INV_X1 U239 ( .A(\A_ns[53] ), .ZN(n786) );
  INV_X1 U240 ( .A(\A_ns[54] ), .ZN(n787) );
  INV_X1 U241 ( .A(\A_ns[55] ), .ZN(n788) );
  INV_X1 U242 ( .A(\A_ns[56] ), .ZN(n789) );
  INV_X1 U243 ( .A(\A_ns[57] ), .ZN(n790) );
  INV_X1 U244 ( .A(\A_ns[58] ), .ZN(n791) );
  INV_X1 U245 ( .A(\A_ns[59] ), .ZN(n792) );
  INV_X1 U246 ( .A(\A_ns[60] ), .ZN(n793) );
  INV_X1 U247 ( .A(\A_ns[61] ), .ZN(n794) );
  INV_X1 U248 ( .A(\A_ns[29] ), .ZN(n795) );
  INV_X1 U249 ( .A(\A_s[29] ), .ZN(n796) );
  INV_X1 U250 ( .A(\A_s[30] ), .ZN(n797) );
  INV_X1 U251 ( .A(\A_s[31] ), .ZN(n798) );
  INV_X1 U252 ( .A(\A_s[32] ), .ZN(n799) );
  INV_X1 U253 ( .A(\A_s[33] ), .ZN(n800) );
  INV_X1 U254 ( .A(\A_s[34] ), .ZN(n801) );
  INV_X1 U255 ( .A(\A_s[35] ), .ZN(n802) );
  INV_X1 U256 ( .A(\A_s[36] ), .ZN(n803) );
  INV_X1 U259 ( .A(\A_s[37] ), .ZN(n804) );
  INV_X1 U260 ( .A(\A_s[38] ), .ZN(n805) );
  INV_X1 U261 ( .A(\A_s[39] ), .ZN(n806) );
  INV_X1 U262 ( .A(\A_s[40] ), .ZN(n807) );
  INV_X1 U263 ( .A(\A_s[41] ), .ZN(n808) );
  INV_X1 U264 ( .A(\A_s[42] ), .ZN(n809) );
  INV_X1 U265 ( .A(\A_s[43] ), .ZN(n810) );
  INV_X1 U266 ( .A(\A_s[44] ), .ZN(n811) );
  INV_X1 U267 ( .A(\A_s[45] ), .ZN(n812) );
  INV_X1 U268 ( .A(\A_s[46] ), .ZN(n813) );
  INV_X1 U269 ( .A(\A_s[47] ), .ZN(n814) );
  INV_X1 U270 ( .A(\A_s[48] ), .ZN(n815) );
  INV_X1 U271 ( .A(\A_s[49] ), .ZN(n816) );
  INV_X1 U272 ( .A(\A_s[50] ), .ZN(n817) );
  INV_X1 U273 ( .A(\A_s[51] ), .ZN(n818) );
  INV_X1 U274 ( .A(\A_s[52] ), .ZN(n819) );
  INV_X1 U275 ( .A(\A_s[53] ), .ZN(n820) );
  INV_X1 U276 ( .A(\A_s[54] ), .ZN(n821) );
  INV_X1 U277 ( .A(\A_s[55] ), .ZN(n822) );
  INV_X1 U278 ( .A(\A_s[56] ), .ZN(n823) );
  INV_X1 U279 ( .A(\A_s[57] ), .ZN(n824) );
  INV_X1 U280 ( .A(\A_s[58] ), .ZN(n825) );
  INV_X1 U281 ( .A(\A_s[59] ), .ZN(n826) );
  INV_X1 U282 ( .A(\A_s[60] ), .ZN(n827) );
  INV_X1 U283 ( .A(\A_s[61] ), .ZN(n828) );
endmodule


module RCA_NBIT36_DW01_add_0 ( A, B, CI, SUM, CO );
  input [35:0] A;
  input [35:0] B;
  output [35:0] SUM;
  input CI;
  output CO;
  wire   n1, n267, n268, n269, n270, n272, n273, n274, n278, n284, n286, n287,
         n288, n290, n291, n293, n294, n295, n296, n297, n299, n300, n302,
         n303, n304, n305, n306, n308, n309, n312, n314, n315, n316, n317,
         n318, n320, n321, n323, n324, n326, n327, n329, n330, n331, n332,
         n333, n334, n336, n337, n338, n339, n341, n342, n349, n350, net176420,
         net182748, net182821, net183238, net183235, net185506, net185591,
         net187523, net187529, net188161, net193306, net188172, net187659,
         net187351, net187324, net182759, n348, n347, n281, net187162,
         net184546, net182643, net176417, net176416, net176400, n346, n345,
         n344, n343, n283, n279, n277, n275, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n271, n276, n280, n282, n285, n289, n292, n298,
         n301, n307, n310, n311, n313, n319, n322, n325, n328, n335, n340,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402;
  wire   [35:1] carry;

  FA_X1 U1_35 ( .A(A[35]), .B(B[35]), .CI(n349), .S(SUM[35]) );
  FA_X1 U1_32 ( .A(A[32]), .B(B[32]), .CI(n383), .CO(carry[33]), .S(SUM[32])
         );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U133 ( .A(n268), .B(n267), .Z(SUM[34]) );
  XOR2_X1 U134 ( .A(carry[33]), .B(n287), .Z(SUM[33]) );
  XOR2_X1 U135 ( .A(A[33]), .B(B[33]), .Z(n287) );
  XOR2_X1 U136 ( .A(carry[31]), .B(n270), .Z(SUM[31]) );
  XOR2_X1 U137 ( .A(A[31]), .B(B[31]), .Z(n270) );
  XOR2_X1 U138 ( .A(net187523), .B(n288), .Z(SUM[2]) );
  XOR2_X1 U144 ( .A(n302), .B(n304), .Z(SUM[22]) );
  XOR2_X1 U145 ( .A(B[22]), .B(A[22]), .Z(n304) );
  XOR2_X1 U149 ( .A(B[18]), .B(A[18]), .Z(n316) );
  XOR2_X1 U153 ( .A(B[13]), .B(A[13]), .Z(n331) );
  XOR2_X1 U156 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  XOR2_X1 U139 ( .A(carry[2]), .B(n252), .Z(n288) );
  XOR2_X1 U132 ( .A(B[3]), .B(net187351), .Z(n286) );
  XOR2_X1 U131 ( .A(A[4]), .B(B[4]), .Z(n284) );
  OR2_X1 U1 ( .A1(n273), .A2(n402), .ZN(n292) );
  NAND2_X1 U2 ( .A1(n292), .A2(n307), .ZN(n226) );
  AOI21_X1 U3 ( .B1(n232), .B2(A[8]), .A(B[8]), .ZN(n227) );
  OR2_X1 U4 ( .A1(n299), .A2(n395), .ZN(n228) );
  NAND2_X1 U5 ( .A1(n228), .A2(n300), .ZN(n296) );
  AND2_X1 U6 ( .A1(n234), .A2(net183235), .ZN(n229) );
  NOR2_X1 U7 ( .A1(n229), .A2(n227), .ZN(n363) );
  BUF_X1 U8 ( .A(n281), .Z(n230) );
  AND2_X1 U9 ( .A1(n386), .A2(n358), .ZN(n352) );
  OAI21_X1 U10 ( .B1(n357), .B2(A[17]), .A(B[17]), .ZN(n318) );
  OR2_X1 U11 ( .A1(n317), .A2(n398), .ZN(n365) );
  XNOR2_X1 U12 ( .A(A[23]), .B(B[23]), .ZN(n231) );
  NAND2_X1 U13 ( .A1(n343), .A2(n247), .ZN(n232) );
  CLKBUF_X1 U14 ( .A(n307), .Z(n233) );
  BUF_X1 U15 ( .A(net187529), .Z(net182748) );
  AND2_X1 U16 ( .A1(n343), .A2(n247), .ZN(n234) );
  OAI21_X1 U17 ( .B1(A[10]), .B2(n226), .A(n391), .ZN(n235) );
  OAI21_X1 U18 ( .B1(A[10]), .B2(n226), .A(n391), .ZN(n335) );
  INV_X1 U19 ( .A(n316), .ZN(n374) );
  AND2_X1 U20 ( .A1(n256), .A2(n388), .ZN(n236) );
  AND2_X2 U21 ( .A1(n335), .A2(n401), .ZN(n372) );
  AND2_X1 U22 ( .A1(n391), .A2(n238), .ZN(n237) );
  NAND2_X1 U23 ( .A1(n233), .A2(n239), .ZN(n238) );
  AND2_X1 U24 ( .A1(n292), .A2(n240), .ZN(n239) );
  INV_X1 U25 ( .A(A[10]), .ZN(n240) );
  NOR2_X1 U26 ( .A1(n294), .A2(n370), .ZN(n290) );
  OR2_X1 U27 ( .A1(n327), .A2(n362), .ZN(n323) );
  AND3_X1 U28 ( .A1(net176420), .A2(n368), .A3(A[9]), .ZN(n241) );
  INV_X1 U29 ( .A(n241), .ZN(n364) );
  AOI21_X1 U30 ( .B1(n277), .B2(n244), .A(n242), .ZN(n243) );
  INV_X1 U31 ( .A(B[7]), .ZN(n242) );
  INV_X1 U32 ( .A(n243), .ZN(n343) );
  XNOR2_X1 U33 ( .A(n275), .B(n246), .ZN(SUM[8]) );
  XNOR2_X1 U34 ( .A(B[8]), .B(A[8]), .ZN(n246) );
  NAND2_X1 U35 ( .A1(n343), .A2(n247), .ZN(n275) );
  AOI21_X1 U36 ( .B1(n232), .B2(A[8]), .A(B[8]), .ZN(n342) );
  OR2_X1 U37 ( .A1(net183238), .A2(n244), .ZN(n247) );
  INV_X1 U38 ( .A(A[7]), .ZN(n244) );
  XNOR2_X1 U39 ( .A(B[7]), .B(n244), .ZN(n278) );
  OAI21_X1 U40 ( .B1(A[6]), .B2(net182748), .A(n245), .ZN(n277) );
  INV_X1 U41 ( .A(n344), .ZN(n245) );
  OAI21_X1 U42 ( .B1(A[6]), .B2(net182748), .A(n245), .ZN(net183238) );
  AOI21_X1 U43 ( .B1(n279), .B2(A[6]), .A(B[6]), .ZN(n344) );
  NAND2_X1 U44 ( .A1(n345), .A2(net187162), .ZN(n279) );
  OR2_X1 U45 ( .A1(n281), .A2(net176400), .ZN(net187162) );
  INV_X1 U46 ( .A(A[5]), .ZN(net176400) );
  OR2_X1 U47 ( .A1(net176400), .A2(n281), .ZN(net193306) );
  OAI21_X1 U48 ( .B1(net176417), .B2(A[5]), .A(B[5]), .ZN(n345) );
  INV_X1 U49 ( .A(net184546), .ZN(net176417) );
  OAI21_X1 U50 ( .B1(A[5]), .B2(net176417), .A(B[5]), .ZN(net188161) );
  OAI22_X1 U51 ( .A1(n248), .A2(net182643), .B1(n346), .B2(B[4]), .ZN(
        net184546) );
  AND2_X1 U52 ( .A1(net176416), .A2(n248), .ZN(n346) );
  BUF_X1 U53 ( .A(A[4]), .Z(n248) );
  AND2_X1 U54 ( .A1(net176416), .A2(n248), .ZN(n249) );
  OAI22_X1 U55 ( .A1(n248), .A2(net182643), .B1(n249), .B2(net188172), .ZN(
        n281) );
  INV_X1 U56 ( .A(n283), .ZN(net176416) );
  BUF_X1 U57 ( .A(net176416), .Z(net182643) );
  OAI22_X1 U58 ( .A1(net187659), .A2(net182759), .B1(n347), .B2(B[3]), .ZN(
        n283) );
  BUF_X1 U59 ( .A(net187324), .Z(net182759) );
  AND2_X1 U60 ( .A1(n255), .A2(n387), .ZN(n250) );
  XNOR2_X1 U61 ( .A(n230), .B(net185591), .ZN(SUM[5]) );
  CLKBUF_X1 U62 ( .A(B[4]), .Z(net188172) );
  OAI22_X1 U63 ( .A1(net187659), .A2(net182759), .B1(B[3]), .B2(n347), .ZN(
        net182821) );
  INV_X1 U64 ( .A(net182759), .ZN(net185506) );
  BUF_X1 U65 ( .A(A[3]), .Z(net187659) );
  CLKBUF_X1 U66 ( .A(net187659), .Z(net187351) );
  AND2_X1 U67 ( .A1(net187324), .A2(A[3]), .ZN(n347) );
  NOR2_X1 U68 ( .A1(n348), .A2(n251), .ZN(net187324) );
  NOR2_X1 U69 ( .A1(A[2]), .A2(B[2]), .ZN(n251) );
  AOI21_X1 U70 ( .B1(A[2]), .B2(B[2]), .A(carry[2]), .ZN(n348) );
  CLKBUF_X1 U71 ( .A(A[2]), .Z(net187523) );
  CLKBUF_X1 U72 ( .A(B[2]), .Z(n252) );
  NAND2_X1 U73 ( .A1(n253), .A2(n254), .ZN(n255) );
  NAND2_X1 U74 ( .A1(n255), .A2(n387), .ZN(n305) );
  INV_X1 U75 ( .A(A[20]), .ZN(n253) );
  INV_X1 U76 ( .A(n353), .ZN(n254) );
  XNOR2_X1 U77 ( .A(n351), .B(n231), .ZN(SUM[23]) );
  OR2_X1 U78 ( .A1(A[18]), .A2(n354), .ZN(n256) );
  NAND2_X1 U79 ( .A1(n256), .A2(n388), .ZN(n301) );
  OAI21_X1 U80 ( .B1(n352), .B2(A[23]), .A(B[23]), .ZN(n257) );
  BUF_X1 U81 ( .A(n352), .Z(n351) );
  XOR2_X1 U82 ( .A(A[30]), .B(B[30]), .Z(n258) );
  XOR2_X1 U83 ( .A(carry[30]), .B(n258), .Z(SUM[30]) );
  NAND2_X1 U84 ( .A1(carry[30]), .A2(A[30]), .ZN(n259) );
  NAND2_X1 U85 ( .A1(carry[30]), .A2(B[30]), .ZN(n260) );
  NAND2_X1 U86 ( .A1(A[30]), .A2(B[30]), .ZN(n261) );
  NAND3_X1 U87 ( .A1(n259), .A2(n260), .A3(n261), .ZN(carry[31]) );
  OR2_X1 U88 ( .A1(n390), .A2(n356), .ZN(n340) );
  OAI21_X1 U89 ( .B1(n299), .B2(n395), .A(n257), .ZN(n262) );
  XNOR2_X1 U90 ( .A(n298), .B(n376), .ZN(SUM[14]) );
  XOR2_X1 U91 ( .A(A[28]), .B(B[28]), .Z(n263) );
  XOR2_X1 U92 ( .A(n350), .B(n263), .Z(SUM[28]) );
  NAND2_X1 U93 ( .A1(A[28]), .A2(B[28]), .ZN(n264) );
  NAND2_X1 U94 ( .A1(A[28]), .A2(n350), .ZN(n265) );
  NAND2_X1 U95 ( .A1(B[28]), .A2(n350), .ZN(n266) );
  NAND3_X1 U96 ( .A1(n264), .A2(n265), .A3(n266), .ZN(carry[29]) );
  XOR2_X1 U97 ( .A(A[29]), .B(B[29]), .Z(n271) );
  XOR2_X1 U98 ( .A(n271), .B(carry[29]), .Z(SUM[29]) );
  NAND2_X1 U99 ( .A1(A[29]), .A2(B[29]), .ZN(n276) );
  NAND2_X1 U100 ( .A1(A[29]), .A2(carry[29]), .ZN(n280) );
  NAND2_X1 U101 ( .A1(B[29]), .A2(carry[29]), .ZN(n282) );
  NAND3_X1 U102 ( .A1(n276), .A2(n280), .A3(n282), .ZN(carry[30]) );
  AOI21_X1 U103 ( .B1(n340), .B2(A[13]), .A(B[13]), .ZN(n285) );
  CLKBUF_X1 U104 ( .A(n262), .Z(n289) );
  NOR2_X1 U105 ( .A1(n285), .A2(n369), .ZN(n298) );
  OAI21_X1 U106 ( .B1(n363), .B2(A[9]), .A(B[9]), .ZN(n307) );
  NAND2_X1 U107 ( .A1(n292), .A2(n307), .ZN(n310) );
  NAND2_X1 U108 ( .A1(net188161), .A2(net193306), .ZN(net187529) );
  XNOR2_X1 U109 ( .A(n301), .B(n382), .ZN(SUM[19]) );
  NAND2_X1 U110 ( .A1(n291), .A2(n311), .ZN(n361) );
  NAND2_X1 U111 ( .A1(n290), .A2(A[26]), .ZN(n311) );
  XNOR2_X1 U112 ( .A(n290), .B(n313), .ZN(SUM[26]) );
  XNOR2_X1 U113 ( .A(A[26]), .B(B[26]), .ZN(n313) );
  NAND2_X1 U114 ( .A1(n361), .A2(A[27]), .ZN(n355) );
  AOI21_X1 U115 ( .B1(n237), .B2(A[11]), .A(B[11]), .ZN(n319) );
  OAI21_X1 U116 ( .B1(A[19]), .B2(n236), .A(B[19]), .ZN(n322) );
  NOR2_X1 U117 ( .A1(n390), .A2(n356), .ZN(n329) );
  NOR2_X1 U118 ( .A1(n319), .A2(n372), .ZN(n325) );
  NOR2_X1 U119 ( .A1(n336), .A2(n372), .ZN(n332) );
  OAI21_X1 U120 ( .B1(A[24]), .B2(n289), .A(n385), .ZN(n328) );
  XOR2_X1 U121 ( .A(B[5]), .B(A[5]), .Z(net185591) );
  NAND2_X1 U122 ( .A1(n322), .A2(n359), .ZN(n353) );
  NAND2_X1 U123 ( .A1(n365), .A2(n318), .ZN(n354) );
  NAND2_X1 U124 ( .A1(n355), .A2(n272), .ZN(n350) );
  AND2_X1 U125 ( .A1(n325), .A2(A[12]), .ZN(n356) );
  AND2_X1 U126 ( .A1(n389), .A2(n366), .ZN(n357) );
  OR2_X1 U127 ( .A1(A[22]), .A2(n302), .ZN(n358) );
  NAND2_X1 U128 ( .A1(n386), .A2(n358), .ZN(n299) );
  OR2_X1 U129 ( .A1(n301), .A2(n397), .ZN(n359) );
  NAND2_X1 U130 ( .A1(n312), .A2(n359), .ZN(n308) );
  XNOR2_X1 U140 ( .A(n328), .B(n295), .ZN(SUM[25]) );
  NOR2_X1 U141 ( .A1(n362), .A2(n327), .ZN(n360) );
  NOR2_X1 U142 ( .A1(A[14]), .A2(n326), .ZN(n362) );
  NAND2_X1 U143 ( .A1(n364), .A2(n341), .ZN(n338) );
  NAND2_X1 U146 ( .A1(n365), .A2(n318), .ZN(n314) );
  OR2_X1 U147 ( .A1(A[16]), .A2(n320), .ZN(n366) );
  NAND2_X1 U148 ( .A1(n389), .A2(n366), .ZN(n317) );
  XOR2_X1 U150 ( .A(n305), .B(n377), .Z(SUM[21]) );
  XNOR2_X1 U151 ( .A(n320), .B(n367), .ZN(SUM[16]) );
  XNOR2_X1 U152 ( .A(B[16]), .B(A[16]), .ZN(n367) );
  NAND2_X1 U154 ( .A1(net183235), .A2(n234), .ZN(n368) );
  NAND2_X1 U155 ( .A1(net176420), .A2(n368), .ZN(n273) );
  INV_X1 U157 ( .A(A[8]), .ZN(net183235) );
  AND2_X1 U158 ( .A1(n329), .A2(n400), .ZN(n369) );
  NOR2_X1 U159 ( .A1(n330), .A2(n369), .ZN(n326) );
  AND2_X1 U160 ( .A1(n394), .A2(n328), .ZN(n370) );
  XNOR2_X1 U161 ( .A(n262), .B(n371), .ZN(SUM[24]) );
  XNOR2_X1 U162 ( .A(B[24]), .B(A[24]), .ZN(n371) );
  XNOR2_X1 U163 ( .A(n323), .B(n373), .ZN(SUM[15]) );
  XOR2_X1 U164 ( .A(A[15]), .B(B[15]), .Z(n373) );
  XNOR2_X1 U165 ( .A(n354), .B(n374), .ZN(SUM[18]) );
  XNOR2_X1 U166 ( .A(n317), .B(n375), .ZN(SUM[17]) );
  XOR2_X1 U167 ( .A(A[17]), .B(B[17]), .Z(n375) );
  XNOR2_X1 U168 ( .A(n329), .B(n331), .ZN(SUM[13]) );
  XNOR2_X1 U169 ( .A(A[14]), .B(B[14]), .ZN(n376) );
  XNOR2_X1 U170 ( .A(A[21]), .B(B[21]), .ZN(n377) );
  XNOR2_X1 U171 ( .A(B[25]), .B(n394), .ZN(n295) );
  XNOR2_X1 U172 ( .A(B[11]), .B(n401), .ZN(n337) );
  XNOR2_X1 U173 ( .A(B[9]), .B(n402), .ZN(n274) );
  INV_X1 U174 ( .A(B[34]), .ZN(n392) );
  INV_X1 U175 ( .A(n297), .ZN(n385) );
  XNOR2_X1 U176 ( .A(n361), .B(n378), .ZN(SUM[27]) );
  XNOR2_X1 U177 ( .A(B[27]), .B(A[27]), .ZN(n378) );
  XNOR2_X1 U178 ( .A(n310), .B(n379), .ZN(SUM[10]) );
  XNOR2_X1 U179 ( .A(B[10]), .B(A[10]), .ZN(n379) );
  XNOR2_X1 U180 ( .A(net187529), .B(n380), .ZN(SUM[6]) );
  XNOR2_X1 U181 ( .A(B[6]), .B(A[6]), .ZN(n380) );
  INV_X1 U182 ( .A(A[13]), .ZN(n400) );
  INV_X1 U183 ( .A(A[15]), .ZN(n399) );
  INV_X1 U184 ( .A(A[21]), .ZN(n396) );
  OAI21_X1 U185 ( .B1(n250), .B2(A[21]), .A(B[21]), .ZN(n306) );
  INV_X1 U186 ( .A(A[23]), .ZN(n395) );
  OAI21_X1 U187 ( .B1(n352), .B2(A[23]), .A(B[23]), .ZN(n300) );
  INV_X1 U188 ( .A(A[19]), .ZN(n397) );
  OAI21_X1 U189 ( .B1(n236), .B2(A[19]), .A(B[19]), .ZN(n312) );
  INV_X1 U190 ( .A(A[17]), .ZN(n398) );
  OAI22_X1 U191 ( .A1(n392), .A2(n393), .B1(n267), .B2(n268), .ZN(n349) );
  XNOR2_X1 U192 ( .A(n353), .B(n381), .ZN(SUM[20]) );
  XNOR2_X1 U193 ( .A(B[20]), .B(A[20]), .ZN(n381) );
  XNOR2_X1 U194 ( .A(A[12]), .B(B[12]), .ZN(n334) );
  AOI22_X1 U195 ( .A1(B[33]), .A2(A[33]), .B1(n287), .B2(carry[33]), .ZN(n267)
         );
  INV_X1 U196 ( .A(n303), .ZN(n386) );
  XOR2_X1 U197 ( .A(A[19]), .B(B[19]), .Z(n382) );
  AOI22_X1 U198 ( .A1(B[31]), .A2(A[31]), .B1(carry[31]), .B2(n270), .ZN(n269)
         );
  OAI21_X1 U199 ( .B1(n361), .B2(A[27]), .A(B[27]), .ZN(n272) );
  INV_X1 U200 ( .A(n269), .ZN(n383) );
  AOI21_X1 U201 ( .B1(n384), .B2(A[25]), .A(B[25]), .ZN(n294) );
  INV_X1 U202 ( .A(n293), .ZN(n384) );
  INV_X1 U203 ( .A(A[9]), .ZN(n402) );
  OAI21_X1 U204 ( .B1(A[26]), .B2(n290), .A(B[26]), .ZN(n291) );
  INV_X1 U205 ( .A(A[11]), .ZN(n401) );
  XNOR2_X1 U206 ( .A(A[34]), .B(B[34]), .ZN(n268) );
  INV_X1 U207 ( .A(A[25]), .ZN(n394) );
  INV_X1 U208 ( .A(A[34]), .ZN(n393) );
  AND2_X1 U209 ( .A1(A[0]), .A2(B[0]), .ZN(n1) );
  XNOR2_X1 U210 ( .A(net185506), .B(n286), .ZN(SUM[3]) );
  XNOR2_X1 U211 ( .A(n235), .B(n337), .ZN(SUM[11]) );
  XNOR2_X1 U212 ( .A(n325), .B(n334), .ZN(SUM[12]) );
  OAI21_X1 U213 ( .B1(n305), .B2(n396), .A(n306), .ZN(n302) );
  INV_X1 U214 ( .A(n309), .ZN(n387) );
  INV_X1 U215 ( .A(n321), .ZN(n389) );
  XNOR2_X1 U216 ( .A(n284), .B(net182821), .ZN(SUM[4]) );
  OAI21_X1 U217 ( .B1(n360), .B2(A[15]), .A(B[15]), .ZN(n324) );
  AOI21_X1 U218 ( .B1(n320), .B2(A[16]), .A(B[16]), .ZN(n321) );
  AOI21_X1 U219 ( .B1(n237), .B2(A[11]), .A(B[11]), .ZN(n336) );
  OAI21_X1 U220 ( .B1(n399), .B2(n323), .A(n324), .ZN(n320) );
  AOI21_X1 U221 ( .B1(n308), .B2(A[20]), .A(B[20]), .ZN(n309) );
  AOI21_X1 U222 ( .B1(n314), .B2(A[18]), .A(B[18]), .ZN(n315) );
  AOI21_X1 U223 ( .B1(n340), .B2(A[13]), .A(B[13]), .ZN(n330) );
  OAI21_X1 U224 ( .B1(n363), .B2(A[9]), .A(B[9]), .ZN(n341) );
  OAI21_X1 U225 ( .B1(A[24]), .B2(n289), .A(n385), .ZN(n293) );
  AOI21_X1 U226 ( .B1(n296), .B2(A[24]), .A(B[24]), .ZN(n297) );
  AOI21_X1 U227 ( .B1(n302), .B2(A[22]), .A(B[22]), .ZN(n303) );
  INV_X1 U228 ( .A(n315), .ZN(n388) );
  INV_X1 U229 ( .A(n333), .ZN(n390) );
  OAI21_X1 U230 ( .B1(n332), .B2(A[12]), .A(B[12]), .ZN(n333) );
  INV_X1 U231 ( .A(n342), .ZN(net176420) );
  XNOR2_X1 U232 ( .A(n273), .B(n274), .ZN(SUM[9]) );
  AOI21_X1 U233 ( .B1(n326), .B2(A[14]), .A(B[14]), .ZN(n327) );
  INV_X1 U234 ( .A(n339), .ZN(n391) );
  AOI21_X1 U235 ( .B1(n338), .B2(A[10]), .A(B[10]), .ZN(n339) );
  XNOR2_X1 U236 ( .A(net183238), .B(n278), .ZN(SUM[7]) );
endmodule


module RCA_NBIT36 ( A, B, Ci, S, Co );
  input [35:0] A;
  input [35:0] B;
  output [35:0] S;
  input Ci;
  output Co;

  assign Co = 1'b0;

  RCA_NBIT36_DW01_add_0 add_95 ( .A(A), .B(B), .CI(1'b0), .SUM(S) );
endmodule


module RCA_NBIT38_DW01_add_0 ( A, B, CI, SUM, CO );
  input [37:0] A;
  input [37:0] B;
  output [37:0] SUM;
  input CI;
  output CO;
  wire   n1, net63979, n237, n238, n240, n243, n245, n246, n248, n249, n251,
         n253, n254, n255, n256, n257, n258, n259, n260, n262, n263, n264,
         n265, n266, n267, n268, n269, n272, n277, n279, n280, n281, n283,
         n284, n285, n286, n290, n292, n293, n294, n295, n296, n299, n300,
         n301, n302, n303, n305, n306, n307, n309, n310, net176441, net176451,
         net184369, net184368, net184367, net185867, net191042, net191664,
         n244, n242, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n239, n241, n247, n250, n252, n261, n270, n271, n273,
         n274, n275, n276, n278, n282, n287, n288, n289, n291, n297, n298,
         n304, n308, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392;
  wire   [37:1] carry;

  FA_X1 U1_35 ( .A(A[35]), .B(B[35]), .CI(n372), .CO(carry[36]), .S(SUM[35])
         );
  FA_X1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FA_X1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U104 ( .A(n352), .B(n254), .Z(SUM[6]) );
  XOR2_X1 U106 ( .A(B[5]), .B(n334), .Z(n256) );
  XOR2_X1 U107 ( .A(A[4]), .B(n257), .Z(SUM[4]) );
  XOR2_X1 U108 ( .A(carry[4]), .B(B[4]), .Z(n257) );
  XOR2_X1 U110 ( .A(carry[36]), .B(n260), .Z(SUM[36]) );
  XOR2_X1 U111 ( .A(A[36]), .B(B[36]), .Z(n260) );
  XOR2_X1 U112 ( .A(carry[34]), .B(n238), .Z(SUM[34]) );
  XOR2_X1 U116 ( .A(n331), .B(n264), .Z(SUM[27]) );
  XOR2_X1 U117 ( .A(B[27]), .B(A[27]), .Z(n264) );
  XOR2_X1 U136 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U1 ( .A(n302), .Z(n368) );
  AND2_X2 U2 ( .A1(A[14]), .A2(B[14]), .ZN(net191664) );
  CLKBUF_X1 U3 ( .A(A[13]), .Z(n204) );
  CLKBUF_X1 U4 ( .A(n255), .Z(n333) );
  CLKBUF_X1 U5 ( .A(n262), .Z(n331) );
  INV_X1 U6 ( .A(B[24]), .ZN(n361) );
  INV_X1 U7 ( .A(B[12]), .ZN(n271) );
  INV_X1 U8 ( .A(B[34]), .ZN(n304) );
  NAND2_X1 U9 ( .A1(n291), .A2(net176441), .ZN(n288) );
  CLKBUF_X1 U10 ( .A(n249), .Z(n205) );
  BUF_X1 U11 ( .A(n280), .Z(n344) );
  OAI21_X1 U12 ( .B1(n212), .B2(n213), .A(n214), .ZN(n206) );
  MUX2_X1 U13 ( .A(n288), .B(n274), .S(net176451), .Z(n252) );
  INV_X1 U14 ( .A(n208), .ZN(n207) );
  NOR2_X1 U15 ( .A1(n209), .A2(n306), .ZN(n208) );
  NOR2_X1 U16 ( .A1(n249), .A2(A[8]), .ZN(n209) );
  BUF_X1 U17 ( .A(n240), .Z(n234) );
  XOR2_X1 U18 ( .A(A[7]), .B(B[7]), .Z(n369) );
  XNOR2_X1 U19 ( .A(A[6]), .B(n214), .ZN(n254) );
  INV_X1 U20 ( .A(B[26]), .ZN(n318) );
  AND2_X1 U21 ( .A1(n216), .A2(n210), .ZN(n243) );
  NAND2_X1 U22 ( .A1(n230), .A2(n387), .ZN(n210) );
  INV_X1 U23 ( .A(B[14]), .ZN(net176441) );
  INV_X1 U24 ( .A(B[18]), .ZN(n366) );
  INV_X1 U25 ( .A(B[29]), .ZN(n323) );
  INV_X1 U26 ( .A(B[9]), .ZN(n315) );
  INV_X1 U27 ( .A(B[11]), .ZN(n365) );
  INV_X1 U28 ( .A(B[17]), .ZN(n367) );
  NAND2_X1 U29 ( .A1(n213), .A2(n211), .ZN(n359) );
  INV_X1 U30 ( .A(n253), .ZN(n211) );
  OAI21_X1 U31 ( .B1(n212), .B2(n213), .A(n214), .ZN(n381) );
  INV_X1 U32 ( .A(n253), .ZN(n212) );
  INV_X1 U33 ( .A(A[6]), .ZN(n213) );
  INV_X1 U34 ( .A(B[6]), .ZN(n214) );
  OR2_X1 U35 ( .A1(A[13]), .A2(B[13]), .ZN(n287) );
  OAI21_X1 U36 ( .B1(n330), .B2(n387), .A(n215), .ZN(n216) );
  INV_X1 U37 ( .A(B[20]), .ZN(n215) );
  XOR2_X2 U38 ( .A(n258), .B(n259), .Z(SUM[37]) );
  XNOR2_X1 U39 ( .A(n218), .B(n227), .ZN(SUM[23]) );
  CLKBUF_X1 U40 ( .A(A[23]), .Z(n227) );
  XNOR2_X1 U41 ( .A(n222), .B(B[23]), .ZN(n218) );
  NAND3_X1 U42 ( .A1(n219), .A2(n220), .A3(n221), .ZN(n222) );
  OR2_X1 U43 ( .A1(B[23]), .A2(A[23]), .ZN(net191042) );
  NAND2_X1 U44 ( .A1(A[23]), .A2(B[23]), .ZN(net184369) );
  NAND2_X1 U45 ( .A1(n217), .A2(A[22]), .ZN(n219) );
  AND3_X1 U46 ( .A1(n219), .A2(n220), .A3(n221), .ZN(net184368) );
  INV_X1 U47 ( .A(n242), .ZN(n217) );
  XNOR2_X1 U48 ( .A(n217), .B(n223), .ZN(SUM[22]) );
  NAND2_X1 U49 ( .A1(n217), .A2(B[22]), .ZN(n220) );
  AOI22_X1 U50 ( .A1(n224), .A2(n226), .B1(n244), .B2(B[21]), .ZN(n242) );
  OR2_X1 U51 ( .A1(n243), .A2(A[21]), .ZN(n244) );
  CLKBUF_X1 U52 ( .A(A[21]), .Z(n226) );
  CLKBUF_X1 U53 ( .A(n243), .Z(n224) );
  XNOR2_X1 U54 ( .A(n224), .B(n225), .ZN(SUM[21]) );
  NAND2_X1 U55 ( .A1(A[22]), .A2(B[22]), .ZN(n221) );
  XNOR2_X1 U56 ( .A(A[22]), .B(B[22]), .ZN(n223) );
  XNOR2_X1 U57 ( .A(A[21]), .B(B[21]), .ZN(n225) );
  AND2_X1 U58 ( .A1(net191042), .A2(net184367), .ZN(n228) );
  INV_X1 U59 ( .A(n384), .ZN(n229) );
  CLKBUF_X1 U60 ( .A(n377), .Z(n339) );
  AOI22_X1 U61 ( .A1(n344), .A2(n340), .B1(n281), .B2(B[19]), .ZN(n230) );
  CLKBUF_X1 U62 ( .A(A[15]), .Z(n231) );
  NAND3_X1 U63 ( .A1(n325), .A2(n326), .A3(n327), .ZN(n232) );
  NAND2_X1 U64 ( .A1(net191042), .A2(net184367), .ZN(net185867) );
  XNOR2_X1 U65 ( .A(A[20]), .B(n215), .ZN(n279) );
  XNOR2_X1 U66 ( .A(n233), .B(n368), .ZN(SUM[10]) );
  XNOR2_X1 U67 ( .A(A[10]), .B(B[10]), .ZN(n233) );
  BUF_X1 U68 ( .A(A[11]), .Z(n332) );
  INV_X1 U69 ( .A(n240), .ZN(n278) );
  XNOR2_X1 U70 ( .A(A[12]), .B(B[12]), .ZN(n276) );
  NAND2_X1 U71 ( .A1(A[12]), .A2(B[12]), .ZN(n282) );
  INV_X1 U72 ( .A(A[12]), .ZN(n270) );
  NAND2_X1 U73 ( .A1(A[13]), .A2(B[13]), .ZN(n247) );
  INV_X1 U74 ( .A(n204), .ZN(n273) );
  NAND2_X1 U75 ( .A1(n287), .A2(n297), .ZN(n250) );
  NAND2_X1 U76 ( .A1(n250), .A2(n247), .ZN(n241) );
  NAND2_X1 U77 ( .A1(n289), .A2(n247), .ZN(net63979) );
  NAND2_X1 U78 ( .A1(net191664), .A2(net63979), .ZN(n261) );
  NAND2_X1 U79 ( .A1(n239), .A2(n236), .ZN(n235) );
  XNOR2_X1 U80 ( .A(n235), .B(B[13]), .ZN(n275) );
  XNOR2_X1 U81 ( .A(n275), .B(n273), .ZN(SUM[13]) );
  INV_X1 U82 ( .A(A[14]), .ZN(net176451) );
  NAND2_X1 U83 ( .A1(n287), .A2(n297), .ZN(n289) );
  NAND2_X1 U84 ( .A1(n278), .A2(n282), .ZN(n239) );
  XNOR2_X1 U85 ( .A(n241), .B(B[14]), .ZN(n274) );
  AND2_X1 U86 ( .A1(n289), .A2(n247), .ZN(n291) );
  XNOR2_X1 U87 ( .A(n276), .B(n234), .ZN(SUM[12]) );
  NAND2_X1 U88 ( .A1(n252), .A2(n261), .ZN(SUM[14]) );
  NAND2_X1 U89 ( .A1(n270), .A2(n271), .ZN(n236) );
  AND2_X1 U90 ( .A1(n239), .A2(n236), .ZN(n297) );
  OAI21_X1 U91 ( .B1(A[27]), .B2(n331), .A(n374), .ZN(n298) );
  XNOR2_X1 U92 ( .A(A[34]), .B(n304), .ZN(n238) );
  BUF_X1 U93 ( .A(n299), .Z(n360) );
  NOR2_X1 U94 ( .A1(net191664), .A2(net63979), .ZN(n296) );
  NAND2_X1 U95 ( .A1(n293), .A2(n292), .ZN(n308) );
  NOR2_X1 U96 ( .A1(net63979), .A2(net191664), .ZN(n314) );
  XNOR2_X1 U97 ( .A(A[30]), .B(B[30]), .ZN(n319) );
  INV_X1 U98 ( .A(n245), .ZN(n311) );
  CLKBUF_X1 U99 ( .A(n378), .Z(n338) );
  CLKBUF_X1 U100 ( .A(n320), .Z(n312) );
  OR2_X1 U101 ( .A1(n312), .A2(n338), .ZN(n313) );
  XNOR2_X1 U102 ( .A(A[9]), .B(n315), .ZN(n248) );
  OR2_X1 U103 ( .A1(n280), .A2(n340), .ZN(n316) );
  CLKBUF_X1 U105 ( .A(n308), .Z(n357) );
  OR2_X1 U109 ( .A1(n378), .A2(n320), .ZN(n317) );
  XNOR2_X1 U113 ( .A(A[26]), .B(n318), .ZN(n267) );
  XNOR2_X1 U114 ( .A(n319), .B(n232), .ZN(SUM[30]) );
  AND2_X1 U115 ( .A1(n308), .A2(A[16]), .ZN(n320) );
  CLKBUF_X1 U118 ( .A(n253), .Z(n352) );
  NAND3_X1 U119 ( .A1(n348), .A2(n347), .A3(n346), .ZN(n321) );
  OR2_X1 U120 ( .A1(net185867), .A2(n386), .ZN(n322) );
  NAND2_X1 U121 ( .A1(n272), .A2(n322), .ZN(n268) );
  XNOR2_X1 U122 ( .A(A[29]), .B(n323), .ZN(n324) );
  XOR2_X1 U123 ( .A(carry[29]), .B(n324), .Z(SUM[29]) );
  NAND2_X1 U124 ( .A1(carry[29]), .A2(A[29]), .ZN(n325) );
  NAND2_X1 U125 ( .A1(carry[29]), .A2(B[29]), .ZN(n326) );
  NAND2_X1 U126 ( .A1(A[29]), .A2(B[29]), .ZN(n327) );
  NAND3_X1 U127 ( .A1(n326), .A2(n325), .A3(n327), .ZN(carry[30]) );
  XNOR2_X1 U128 ( .A(n337), .B(n328), .ZN(SUM[25]) );
  XNOR2_X1 U129 ( .A(B[25]), .B(A[25]), .ZN(n328) );
  NOR2_X1 U130 ( .A1(n314), .A2(n343), .ZN(n329) );
  AOI22_X1 U131 ( .A1(n344), .A2(n340), .B1(n281), .B2(B[19]), .ZN(n330) );
  AOI22_X1 U132 ( .A1(n344), .A2(n340), .B1(n316), .B2(B[19]), .ZN(n277) );
  CLKBUF_X1 U133 ( .A(A[5]), .Z(n334) );
  XNOR2_X1 U134 ( .A(n373), .B(n335), .ZN(SUM[28]) );
  XNOR2_X1 U135 ( .A(B[28]), .B(A[28]), .ZN(n335) );
  CLKBUF_X1 U137 ( .A(n268), .Z(n337) );
  XNOR2_X1 U138 ( .A(n336), .B(n321), .ZN(SUM[31]) );
  XNOR2_X1 U139 ( .A(A[31]), .B(B[31]), .ZN(n336) );
  BUF_X1 U140 ( .A(A[19]), .Z(n340) );
  AOI21_X1 U141 ( .B1(n357), .B2(A[16]), .A(n338), .ZN(n341) );
  OAI21_X1 U142 ( .B1(A[17]), .B2(n313), .A(n339), .ZN(n342) );
  AND2_X1 U143 ( .A1(net176441), .A2(net176451), .ZN(n343) );
  NOR2_X1 U144 ( .A1(n296), .A2(n343), .ZN(n294) );
  OR2_X1 U145 ( .A1(n265), .A2(n384), .ZN(n345) );
  NAND2_X1 U146 ( .A1(n266), .A2(n345), .ZN(n262) );
  NAND2_X1 U147 ( .A1(A[30]), .A2(B[30]), .ZN(n346) );
  NAND2_X1 U148 ( .A1(A[30]), .A2(carry[30]), .ZN(n347) );
  NAND2_X1 U149 ( .A1(B[30]), .A2(carry[30]), .ZN(n348) );
  NAND3_X1 U150 ( .A1(n348), .A2(n347), .A3(n346), .ZN(carry[31]) );
  NAND2_X1 U151 ( .A1(A[31]), .A2(B[31]), .ZN(n349) );
  NAND2_X1 U152 ( .A1(A[31]), .A2(carry[31]), .ZN(n350) );
  NAND2_X1 U153 ( .A1(B[31]), .A2(carry[31]), .ZN(n351) );
  NAND3_X1 U154 ( .A1(n349), .A2(n350), .A3(n351), .ZN(carry[32]) );
  XNOR2_X1 U155 ( .A(n357), .B(n353), .ZN(SUM[16]) );
  XNOR2_X1 U156 ( .A(A[16]), .B(B[16]), .ZN(n353) );
  AND2_X1 U157 ( .A1(n375), .A2(n356), .ZN(n354) );
  XNOR2_X1 U158 ( .A(n355), .B(n205), .ZN(SUM[8]) );
  XNOR2_X1 U159 ( .A(A[8]), .B(B[8]), .ZN(n355) );
  NAND2_X1 U160 ( .A1(net184368), .A2(net184369), .ZN(net184367) );
  OR2_X1 U161 ( .A1(A[25]), .A2(n268), .ZN(n356) );
  NAND2_X1 U162 ( .A1(n375), .A2(n356), .ZN(n265) );
  AND2_X1 U163 ( .A1(n381), .A2(n359), .ZN(n358) );
  NAND2_X1 U164 ( .A1(n206), .A2(n359), .ZN(n251) );
  XNOR2_X1 U165 ( .A(n361), .B(A[24]), .ZN(n371) );
  INV_X1 U166 ( .A(n386), .ZN(n362) );
  XNOR2_X1 U167 ( .A(n344), .B(n363), .ZN(SUM[19]) );
  XNOR2_X1 U168 ( .A(B[19]), .B(A[19]), .ZN(n363) );
  CLKBUF_X1 U169 ( .A(A[10]), .Z(n364) );
  XNOR2_X1 U170 ( .A(A[11]), .B(n365), .ZN(n301) );
  XNOR2_X1 U171 ( .A(n366), .B(A[18]), .ZN(n285) );
  XNOR2_X1 U172 ( .A(A[17]), .B(n367), .ZN(n370) );
  XNOR2_X1 U173 ( .A(n369), .B(n251), .ZN(SUM[7]) );
  XNOR2_X1 U174 ( .A(n370), .B(n341), .ZN(SUM[17]) );
  XNOR2_X1 U175 ( .A(net185867), .B(n371), .ZN(SUM[24]) );
  XNOR2_X1 U176 ( .A(n342), .B(n285), .ZN(SUM[18]) );
  XNOR2_X1 U177 ( .A(n277), .B(n279), .ZN(SUM[20]) );
  AOI22_X1 U178 ( .A1(B[34]), .A2(A[34]), .B1(n238), .B2(carry[34]), .ZN(n237)
         );
  XNOR2_X1 U179 ( .A(n267), .B(n265), .ZN(SUM[26]) );
  INV_X1 U180 ( .A(n298), .ZN(n373) );
  INV_X1 U181 ( .A(n269), .ZN(n375) );
  AOI21_X1 U182 ( .B1(n268), .B2(A[25]), .A(B[25]), .ZN(n269) );
  OAI21_X1 U183 ( .B1(n376), .B2(A[18]), .A(B[18]), .ZN(n284) );
  INV_X1 U184 ( .A(n283), .ZN(n376) );
  XNOR2_X1 U185 ( .A(n295), .B(B[15]), .ZN(SUM[15]) );
  OAI21_X1 U186 ( .B1(n229), .B2(n354), .A(B[26]), .ZN(n266) );
  INV_X1 U187 ( .A(A[24]), .ZN(n386) );
  OAI21_X1 U188 ( .B1(n228), .B2(n362), .A(B[24]), .ZN(n272) );
  OAI21_X1 U189 ( .B1(A[27]), .B2(n331), .A(n374), .ZN(n245) );
  INV_X1 U190 ( .A(n263), .ZN(n374) );
  AOI21_X1 U191 ( .B1(n262), .B2(A[27]), .A(B[27]), .ZN(n263) );
  OAI21_X1 U192 ( .B1(n311), .B2(A[28]), .A(B[28]), .ZN(n246) );
  INV_X1 U193 ( .A(n237), .ZN(n372) );
  INV_X1 U194 ( .A(A[26]), .ZN(n384) );
  INV_X1 U195 ( .A(A[20]), .ZN(n387) );
  OAI21_X1 U196 ( .B1(A[17]), .B2(n313), .A(n377), .ZN(n283) );
  AOI21_X1 U197 ( .B1(n317), .B2(A[17]), .A(B[17]), .ZN(n286) );
  INV_X1 U198 ( .A(A[28]), .ZN(n385) );
  XNOR2_X1 U199 ( .A(B[37]), .B(A[37]), .ZN(n258) );
  AOI22_X1 U200 ( .A1(carry[36]), .A2(n260), .B1(A[36]), .B2(B[36]), .ZN(n259)
         );
  OAI21_X1 U201 ( .B1(B[4]), .B2(A[4]), .A(n383), .ZN(n255) );
  INV_X1 U202 ( .A(n310), .ZN(n383) );
  AOI21_X1 U203 ( .B1(A[4]), .B2(B[4]), .A(carry[4]), .ZN(n310) );
  OAI21_X1 U204 ( .B1(n333), .B2(n392), .A(n309), .ZN(n253) );
  INV_X1 U205 ( .A(A[5]), .ZN(n392) );
  OAI21_X1 U206 ( .B1(A[5]), .B2(n382), .A(B[5]), .ZN(n309) );
  INV_X1 U207 ( .A(n255), .ZN(n382) );
  OAI21_X1 U208 ( .B1(n298), .B2(n385), .A(n246), .ZN(carry[29]) );
  XNOR2_X1 U209 ( .A(n333), .B(n256), .ZN(SUM[5]) );
  AND2_X1 U210 ( .A1(A[0]), .A2(B[0]), .ZN(n1) );
  OAI21_X1 U211 ( .B1(n342), .B2(n388), .A(n284), .ZN(n280) );
  OAI21_X1 U212 ( .B1(A[9]), .B2(n208), .A(B[9]), .ZN(n305) );
  INV_X1 U213 ( .A(A[9]), .ZN(n390) );
  INV_X1 U214 ( .A(n290), .ZN(n378) );
  OAI21_X1 U215 ( .B1(n231), .B2(n294), .A(n292), .ZN(n295) );
  NAND2_X1 U216 ( .A1(A[15]), .A2(n294), .ZN(n292) );
  OAI21_X1 U217 ( .B1(A[15]), .B2(n329), .A(B[15]), .ZN(n293) );
  OAI21_X1 U218 ( .B1(n308), .B2(A[16]), .A(B[16]), .ZN(n290) );
  OAI21_X1 U219 ( .B1(n358), .B2(A[7]), .A(B[7]), .ZN(n307) );
  INV_X1 U220 ( .A(A[7]), .ZN(n391) );
  INV_X1 U221 ( .A(n286), .ZN(n377) );
  OR2_X1 U222 ( .A1(n280), .A2(n340), .ZN(n281) );
  AOI21_X1 U223 ( .B1(n302), .B2(A[10]), .A(B[10]), .ZN(n303) );
  AOI21_X1 U224 ( .B1(A[8]), .B2(n249), .A(B[8]), .ZN(n306) );
  OAI21_X1 U225 ( .B1(n379), .B2(n332), .A(B[11]), .ZN(n300) );
  INV_X1 U226 ( .A(n332), .ZN(n389) );
  INV_X1 U227 ( .A(A[18]), .ZN(n388) );
  XNOR2_X1 U228 ( .A(n360), .B(n301), .ZN(SUM[11]) );
  OAI21_X1 U229 ( .B1(n360), .B2(n389), .A(n300), .ZN(n240) );
  INV_X1 U230 ( .A(n299), .ZN(n379) );
  XNOR2_X1 U231 ( .A(n248), .B(n207), .ZN(SUM[9]) );
  OAI21_X1 U232 ( .B1(n207), .B2(n390), .A(n305), .ZN(n302) );
  OAI21_X1 U233 ( .B1(n251), .B2(n391), .A(n307), .ZN(n249) );
  OAI21_X1 U234 ( .B1(n364), .B2(n368), .A(n380), .ZN(n299) );
  INV_X1 U235 ( .A(n303), .ZN(n380) );
endmodule


module RCA_NBIT38 ( A, B, Ci, S, Co );
  input [37:0] A;
  input [37:0] B;
  output [37:0] S;
  input Ci;
  output Co;

  assign Co = 1'b0;

  RCA_NBIT38_DW01_add_0 add_95 ( .A(A), .B(B), .CI(1'b0), .SUM(S) );
endmodule


module RCA_NBIT40_DW01_add_0 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, net88456, n238, n211, n212, n215, n216, n218, n219, n220, n222,
         n224, n225, n227, n228, n230, n239, n240, n242, n243, n245, n246,
         n255, n257, n260, n261, n263, n264, n265, n266, n267, n268, net176492,
         net176493, net176501, net183387, net184530, net184527, net184854,
         net187179, net183098, net183017, n214, net193275, n252, n248, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n213, n217, n221, n223, n226,
         n229, n231, n232, n233, n234, n235, n236, n237, n241, n244, n247,
         n249, n250, n251, n253, n254, n256, n258, n259, n262, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325;
  wire   [39:1] carry;
  assign net88456 = A[10];

  FA_X1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FA_X1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FA_X1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FA_X1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FA_X1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FA_X1 U1_32 ( .A(B[32]), .B(n268), .CI(A[32]), .CO(carry[33]), .S(SUM[32])
         );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U75 ( .A(n316), .B(n224), .Z(SUM[7]) );
  XOR2_X1 U76 ( .A(B[7]), .B(n291), .Z(n224) );
  XOR2_X1 U77 ( .A(A[6]), .B(n225), .Z(SUM[6]) );
  XOR2_X1 U78 ( .A(carry[6]), .B(B[6]), .Z(n225) );
  XOR2_X1 U81 ( .A(n187), .B(n211), .Z(SUM[31]) );
  XOR2_X1 U83 ( .A(carry[30]), .B(n227), .Z(SUM[30]) );
  XOR2_X1 U110 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  NAND2_X1 U1 ( .A1(n232), .A2(n231), .ZN(n182) );
  XNOR2_X1 U2 ( .A(n296), .B(n183), .ZN(SUM[8]) );
  XOR2_X1 U3 ( .A(A[8]), .B(n193), .Z(n183) );
  BUF_X1 U4 ( .A(A[26]), .Z(n287) );
  XNOR2_X1 U5 ( .A(n184), .B(n185), .ZN(SUM[24]) );
  AND2_X1 U6 ( .A1(n208), .A2(n209), .ZN(n184) );
  XOR2_X1 U7 ( .A(B[24]), .B(A[24]), .Z(n185) );
  NAND2_X1 U8 ( .A1(n188), .A2(n210), .ZN(net184854) );
  INV_X1 U9 ( .A(net183387), .ZN(n210) );
  NAND2_X1 U10 ( .A1(n244), .A2(n237), .ZN(n207) );
  NAND2_X1 U11 ( .A1(n229), .A2(n241), .ZN(n206) );
  XNOR2_X1 U12 ( .A(n233), .B(n203), .ZN(SUM[22]) );
  INV_X1 U13 ( .A(B[20]), .ZN(net183017) );
  INV_X1 U14 ( .A(n203), .ZN(n241) );
  INV_X1 U15 ( .A(B[22]), .ZN(n229) );
  NAND2_X1 U16 ( .A1(n203), .A2(B[22]), .ZN(n244) );
  INV_X1 U17 ( .A(B[9]), .ZN(n292) );
  INV_X1 U18 ( .A(B[23]), .ZN(n232) );
  INV_X1 U19 ( .A(B[8]), .ZN(n193) );
  INV_X1 U20 ( .A(B[30]), .ZN(n288) );
  AND2_X1 U21 ( .A1(n206), .A2(n207), .ZN(n186) );
  CLKBUF_X1 U22 ( .A(n212), .Z(n187) );
  AND2_X1 U23 ( .A1(n209), .A2(n208), .ZN(n188) );
  OR2_X1 U24 ( .A1(n299), .A2(n311), .ZN(net193275) );
  OR2_X2 U25 ( .A1(n299), .A2(n311), .ZN(n297) );
  XOR2_X1 U26 ( .A(A[34]), .B(B[34]), .Z(n189) );
  XOR2_X1 U27 ( .A(carry[34]), .B(n189), .Z(SUM[34]) );
  NAND2_X1 U28 ( .A1(carry[34]), .A2(A[34]), .ZN(n190) );
  NAND2_X1 U29 ( .A1(carry[34]), .A2(B[34]), .ZN(n191) );
  NAND2_X1 U30 ( .A1(A[34]), .A2(B[34]), .ZN(n192) );
  NAND3_X1 U31 ( .A1(n190), .A2(n191), .A3(n192), .ZN(carry[35]) );
  XNOR2_X1 U32 ( .A(A[39]), .B(n196), .ZN(SUM[39]) );
  CLKBUF_X1 U33 ( .A(n222), .Z(n296) );
  NAND2_X1 U34 ( .A1(n289), .A2(n313), .ZN(n194) );
  INV_X1 U35 ( .A(B[39]), .ZN(n271) );
  OR2_X2 U36 ( .A1(n201), .A2(n195), .ZN(n277) );
  NOR2_X1 U37 ( .A1(n194), .A2(n322), .ZN(n195) );
  XOR2_X1 U38 ( .A(carry[39]), .B(n271), .Z(n196) );
  NAND2_X1 U39 ( .A1(B[20]), .A2(A[20]), .ZN(n226) );
  BUF_X1 U40 ( .A(n248), .Z(n262) );
  NAND2_X1 U41 ( .A1(n204), .A2(n205), .ZN(n203) );
  OAI21_X1 U42 ( .B1(B[21]), .B2(n221), .A(A[21]), .ZN(n205) );
  BUF_X1 U43 ( .A(n220), .Z(n285) );
  BUF_X1 U44 ( .A(A[13]), .Z(n259) );
  BUF_X1 U45 ( .A(net176493), .Z(net184527) );
  BUF_X1 U46 ( .A(A[12]), .Z(n280) );
  OAI21_X1 U47 ( .B1(n198), .B2(n197), .A(n199), .ZN(net176492) );
  INV_X1 U48 ( .A(A[14]), .ZN(n197) );
  INV_X1 U49 ( .A(n248), .ZN(n198) );
  INV_X1 U50 ( .A(B[14]), .ZN(n199) );
  AOI21_X1 U51 ( .B1(n257), .B2(n322), .A(n200), .ZN(n201) );
  INV_X1 U52 ( .A(B[11]), .ZN(n200) );
  XOR2_X1 U53 ( .A(n235), .B(n214), .Z(SUM[20]) );
  AND2_X1 U54 ( .A1(net176501), .A2(net184854), .ZN(n202) );
  OAI21_X1 U55 ( .B1(n213), .B2(n217), .A(net184530), .ZN(n235) );
  NAND2_X1 U56 ( .A1(n235), .A2(n214), .ZN(n223) );
  NOR2_X1 U57 ( .A1(net193275), .A2(B[19]), .ZN(n213) );
  INV_X1 U58 ( .A(A[23]), .ZN(n231) );
  NAND2_X1 U59 ( .A1(n223), .A2(n226), .ZN(n221) );
  NAND2_X1 U60 ( .A1(n223), .A2(n226), .ZN(n250) );
  NAND2_X1 U61 ( .A1(B[23]), .A2(n249), .ZN(n208) );
  XNOR2_X1 U62 ( .A(n249), .B(B[23]), .ZN(net183098) );
  NAND2_X1 U63 ( .A1(n247), .A2(n186), .ZN(n209) );
  NAND2_X1 U64 ( .A1(n253), .A2(n208), .ZN(n251) );
  XNOR2_X1 U65 ( .A(n250), .B(B[21]), .ZN(n234) );
  NAND2_X1 U66 ( .A1(B[21]), .A2(n221), .ZN(n204) );
  AOI21_X1 U67 ( .B1(n251), .B2(net183387), .A(B[24]), .ZN(n230) );
  XNOR2_X1 U68 ( .A(B[19]), .B(A[19]), .ZN(n236) );
  INV_X1 U69 ( .A(A[19]), .ZN(n217) );
  XNOR2_X1 U70 ( .A(B[22]), .B(A[22]), .ZN(n233) );
  INV_X1 U71 ( .A(A[22]), .ZN(n237) );
  NAND2_X1 U72 ( .A1(n232), .A2(n231), .ZN(n247) );
  XNOR2_X1 U73 ( .A(n234), .B(A[21]), .ZN(SUM[21]) );
  BUF_X1 U74 ( .A(A[23]), .Z(n249) );
  XNOR2_X1 U79 ( .A(n297), .B(n236), .ZN(SUM[19]) );
  NAND2_X1 U80 ( .A1(n182), .A2(n186), .ZN(n253) );
  OR2_X1 U82 ( .A1(n276), .A2(n255), .ZN(n254) );
  BUF_X1 U84 ( .A(A[18]), .Z(n274) );
  XNOR2_X1 U85 ( .A(n269), .B(n262), .ZN(SUM[14]) );
  OAI21_X1 U86 ( .B1(n262), .B2(n270), .A(net176492), .ZN(n245) );
  XNOR2_X1 U87 ( .A(A[14]), .B(B[14]), .ZN(n269) );
  OAI21_X1 U88 ( .B1(n254), .B2(n256), .A(n252), .ZN(n248) );
  OAI21_X1 U89 ( .B1(n259), .B2(net187179), .A(B[13]), .ZN(n252) );
  INV_X1 U90 ( .A(n259), .ZN(n256) );
  CLKBUF_X1 U91 ( .A(A[14]), .Z(n270) );
  XNOR2_X1 U92 ( .A(n258), .B(net187179), .ZN(SUM[13]) );
  XNOR2_X1 U93 ( .A(A[13]), .B(B[13]), .ZN(n258) );
  OAI21_X1 U94 ( .B1(n279), .B2(A[25]), .A(B[25]), .ZN(n272) );
  NAND2_X1 U95 ( .A1(n272), .A2(n275), .ZN(n273) );
  OR2_X1 U96 ( .A1(n215), .A2(n320), .ZN(n275) );
  NAND2_X1 U97 ( .A1(n216), .A2(n275), .ZN(n238) );
  XNOR2_X1 U98 ( .A(net183098), .B(n186), .ZN(SUM[23]) );
  XNOR2_X1 U99 ( .A(A[20]), .B(net183017), .ZN(n214) );
  NOR2_X1 U100 ( .A1(n255), .A2(n276), .ZN(net187179) );
  NOR2_X1 U101 ( .A1(n277), .A2(n280), .ZN(n276) );
  INV_X1 U102 ( .A(n321), .ZN(n278) );
  AND2_X1 U103 ( .A1(net176501), .A2(net184854), .ZN(n279) );
  CLKBUF_X1 U104 ( .A(n260), .Z(n281) );
  XNOR2_X1 U105 ( .A(n282), .B(n238), .ZN(SUM[26]) );
  XNOR2_X1 U106 ( .A(A[26]), .B(B[26]), .ZN(n282) );
  CLKBUF_X1 U107 ( .A(n303), .Z(n283) );
  CLKBUF_X1 U108 ( .A(n312), .Z(n284) );
  AND2_X1 U109 ( .A1(n312), .A2(n303), .ZN(n286) );
  XNOR2_X1 U111 ( .A(A[30]), .B(n288), .ZN(n227) );
  NAND2_X1 U112 ( .A1(net184854), .A2(net176501), .ZN(n215) );
  OR2_X1 U113 ( .A1(B[10]), .A2(n260), .ZN(n289) );
  NAND2_X1 U114 ( .A1(n313), .A2(n289), .ZN(n257) );
  CLKBUF_X1 U115 ( .A(A[8]), .Z(n290) );
  INV_X1 U116 ( .A(n324), .ZN(n291) );
  XNOR2_X1 U117 ( .A(n279), .B(n228), .ZN(SUM[25]) );
  NAND2_X1 U118 ( .A1(n297), .A2(B[19]), .ZN(net184530) );
  XNOR2_X1 U119 ( .A(A[9]), .B(n292), .ZN(n307) );
  NAND2_X1 U120 ( .A1(n273), .A2(n287), .ZN(n293) );
  NAND2_X1 U121 ( .A1(n273), .A2(B[26]), .ZN(n294) );
  NAND2_X1 U122 ( .A1(n287), .A2(B[26]), .ZN(n295) );
  NAND3_X1 U123 ( .A1(n294), .A2(n293), .A3(n295), .ZN(carry[27]) );
  XNOR2_X1 U124 ( .A(A[11]), .B(n200), .ZN(n306) );
  BUF_X1 U125 ( .A(A[31]), .Z(n298) );
  CLKBUF_X1 U126 ( .A(A[24]), .Z(net183387) );
  XNOR2_X1 U127 ( .A(A[31]), .B(B[31]), .ZN(n212) );
  XNOR2_X1 U128 ( .A(A[25]), .B(B[25]), .ZN(n228) );
  AND2_X1 U129 ( .A1(n218), .A2(n274), .ZN(n299) );
  OR2_X1 U130 ( .A1(n318), .A2(n245), .ZN(n300) );
  NAND2_X1 U131 ( .A1(n246), .A2(n300), .ZN(n242) );
  AND2_X1 U132 ( .A1(n312), .A2(n303), .ZN(n301) );
  XNOR2_X1 U133 ( .A(n301), .B(n302), .ZN(SUM[17]) );
  XNOR2_X1 U134 ( .A(A[17]), .B(B[17]), .ZN(n302) );
  OR2_X1 U135 ( .A1(A[16]), .A2(n242), .ZN(n303) );
  NAND2_X1 U136 ( .A1(n283), .A2(n284), .ZN(n239) );
  XNOR2_X1 U137 ( .A(B[16]), .B(A[16]), .ZN(n304) );
  XNOR2_X1 U138 ( .A(n242), .B(n304), .ZN(SUM[16]) );
  XNOR2_X1 U139 ( .A(n218), .B(n305), .ZN(SUM[18]) );
  XNOR2_X1 U140 ( .A(A[18]), .B(B[18]), .ZN(n305) );
  INV_X1 U141 ( .A(A[25]), .ZN(n320) );
  INV_X1 U142 ( .A(n230), .ZN(net176501) );
  XNOR2_X1 U143 ( .A(n306), .B(n257), .ZN(SUM[11]) );
  XNOR2_X1 U144 ( .A(n307), .B(n285), .ZN(SUM[9]) );
  INV_X1 U145 ( .A(A[17]), .ZN(n321) );
  INV_X1 U146 ( .A(n261), .ZN(n313) );
  INV_X1 U147 ( .A(A[15]), .ZN(n318) );
  OAI21_X1 U148 ( .B1(net176493), .B2(A[15]), .A(B[15]), .ZN(n246) );
  XNOR2_X1 U149 ( .A(n281), .B(n308), .ZN(SUM[10]) );
  XNOR2_X1 U150 ( .A(net88456), .B(B[10]), .ZN(n308) );
  XNOR2_X1 U151 ( .A(n309), .B(n277), .ZN(SUM[12]) );
  XNOR2_X1 U152 ( .A(A[12]), .B(B[12]), .ZN(n309) );
  INV_X1 U153 ( .A(n243), .ZN(n312) );
  XNOR2_X1 U154 ( .A(net184527), .B(n310), .ZN(SUM[15]) );
  XNOR2_X1 U155 ( .A(A[15]), .B(B[15]), .ZN(n310) );
  OAI21_X1 U156 ( .B1(n202), .B2(A[25]), .A(B[25]), .ZN(n216) );
  OAI21_X1 U157 ( .B1(n314), .B2(A[9]), .A(B[9]), .ZN(n263) );
  INV_X1 U158 ( .A(B[31]), .ZN(n325) );
  AOI22_X1 U159 ( .A1(B[30]), .A2(A[30]), .B1(n227), .B2(carry[30]), .ZN(n211)
         );
  OAI22_X1 U160 ( .A1(n325), .A2(n319), .B1(n211), .B2(n212), .ZN(n268) );
  INV_X1 U161 ( .A(n265), .ZN(n316) );
  INV_X1 U162 ( .A(n298), .ZN(n319) );
  AOI21_X1 U163 ( .B1(A[6]), .B2(B[6]), .A(n317), .ZN(n265) );
  INV_X1 U164 ( .A(n267), .ZN(n317) );
  OAI21_X1 U165 ( .B1(A[6]), .B2(B[6]), .A(carry[6]), .ZN(n267) );
  AOI21_X1 U166 ( .B1(n324), .B2(n265), .A(n266), .ZN(n222) );
  INV_X1 U167 ( .A(A[7]), .ZN(n324) );
  AOI21_X1 U168 ( .B1(n316), .B2(A[7]), .A(B[7]), .ZN(n266) );
  AND2_X1 U169 ( .A1(A[0]), .A2(B[0]), .ZN(n1) );
  INV_X1 U170 ( .A(n264), .ZN(n315) );
  AOI21_X1 U171 ( .B1(n286), .B2(n278), .A(B[17]), .ZN(n240) );
  AOI21_X1 U172 ( .B1(n277), .B2(n280), .A(B[12]), .ZN(n255) );
  AOI21_X1 U173 ( .B1(n321), .B2(n239), .A(n240), .ZN(n218) );
  AOI21_X1 U174 ( .B1(n242), .B2(A[16]), .A(B[16]), .ZN(n243) );
  INV_X1 U175 ( .A(n245), .ZN(net176493) );
  OAI21_X1 U176 ( .B1(n290), .B2(n296), .A(n315), .ZN(n220) );
  AOI21_X1 U177 ( .B1(A[8]), .B2(n222), .A(B[8]), .ZN(n264) );
  OAI21_X1 U178 ( .B1(n218), .B2(n274), .A(B[18]), .ZN(n219) );
  AOI21_X1 U179 ( .B1(n260), .B2(B[10]), .A(net88456), .ZN(n261) );
  OAI21_X1 U180 ( .B1(n285), .B2(n323), .A(n263), .ZN(n260) );
  INV_X1 U181 ( .A(n220), .ZN(n314) );
  INV_X1 U182 ( .A(A[11]), .ZN(n322) );
  INV_X1 U183 ( .A(n219), .ZN(n311) );
  INV_X1 U184 ( .A(A[9]), .ZN(n323) );
endmodule


module RCA_NBIT40 ( A, B, Ci, S, Co );
  input [39:0] A;
  input [39:0] B;
  output [39:0] S;
  input Ci;
  output Co;

  assign Co = 1'b0;

  RCA_NBIT40_DW01_add_0 add_95 ( .A(A), .B(B), .CI(1'b0), .SUM(S) );
endmodule


module RCA_NBIT42_DW01_add_0 ( A, B, CI, SUM, CO );
  input [41:0] A;
  input [41:0] B;
  output [41:0] SUM;
  input CI;
  output CO;
  wire   \carry[32] , \carry[31] , \carry[30] , \carry[29] , \carry[28] ,
         \carry[26] , \carry[24] , \carry[23] , \carry[22] , n223, n224, n225,
         n226, n227, n228, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n253, n256, n257, n258, n259, n261, n262, n263,
         n266, n268, n269, n271, n272, n277, n279, n280, n281, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, net183027, net184427, net186686, net187832, n278, n274, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n229, n252, n254, n255, n260, n264, n265, n267, n270, n273,
         n275, n276, n282, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350;
  wire   [41:1] carry;

  FA_X1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FA_X1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FA_X1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FA_X1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(n275), .CO(\carry[22] ), .S(SUM[21])
         );
  FA_X1 U1_22 ( .A(B[22]), .B(A[22]), .CI(\carry[22] ), .CO(\carry[23] ), .S(
        SUM[22]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(n326), .CO(\carry[26] ), .S(SUM[25])
         );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(n325), .CO(\carry[28] ), .S(SUM[27])
         );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(\carry[28] ), .CO(\carry[29] ), .S(
        SUM[28]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(\carry[29] ), .CO(\carry[30] ), .S(
        SUM[29]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(\carry[30] ), .CO(\carry[31] ), .S(
        SUM[30]) );
  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(\carry[31] ), .CO(\carry[32] ), .S(
        SUM[31]) );
  XNOR2_X2 U6 ( .A(n244), .B(n245), .ZN(SUM[41]) );
  XOR2_X1 U89 ( .A(n232), .B(n233), .Z(SUM[9]) );
  XOR2_X1 U90 ( .A(B[9]), .B(n305), .Z(n233) );
  XOR2_X1 U91 ( .A(n234), .B(n235), .Z(SUM[8]) );
  XOR2_X1 U92 ( .A(n345), .B(B[8]), .Z(n235) );
  XOR2_X1 U93 ( .A(n236), .B(n237), .Z(SUM[7]) );
  XOR2_X1 U94 ( .A(B[7]), .B(A[7]), .Z(n237) );
  XOR2_X1 U95 ( .A(n238), .B(n239), .Z(SUM[6]) );
  XOR2_X1 U96 ( .A(n346), .B(B[6]), .Z(n239) );
  XOR2_X1 U97 ( .A(n240), .B(n241), .Z(SUM[5]) );
  XOR2_X1 U98 ( .A(B[5]), .B(A[5]), .Z(n241) );
  XOR2_X1 U99 ( .A(n242), .B(n243), .Z(SUM[4]) );
  XOR2_X1 U100 ( .A(n347), .B(B[4]), .Z(n243) );
  XOR2_X1 U101 ( .A(B[41]), .B(A[41]), .Z(n245) );
  XOR2_X1 U102 ( .A(n247), .B(n248), .Z(SUM[40]) );
  XOR2_X1 U103 ( .A(B[40]), .B(A[40]), .Z(n248) );
  XOR2_X1 U108 ( .A(n338), .B(n253), .Z(SUM[2]) );
  XOR2_X1 U109 ( .A(n348), .B(B[2]), .Z(n253) );
  XOR2_X1 U110 ( .A(n226), .B(\carry[26] ), .Z(SUM[26]) );
  XOR2_X1 U112 ( .A(n228), .B(n213), .Z(SUM[24]) );
  XOR2_X1 U116 ( .A(n339), .B(n257), .Z(SUM[1]) );
  XOR2_X1 U117 ( .A(B[1]), .B(A[1]), .Z(n257) );
  XOR2_X1 U134 ( .A(n315), .B(n285), .Z(SUM[10]) );
  XOR2_X1 U135 ( .A(n344), .B(B[10]), .Z(n285) );
  XOR2_X1 U136 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  NAND3_X1 U1 ( .A1(n220), .A2(n221), .A3(n222), .ZN(n188) );
  BUF_X1 U2 ( .A(n204), .Z(net186686) );
  BUF_X1 U3 ( .A(n230), .Z(n189) );
  BUF_X1 U4 ( .A(n283), .Z(n315) );
  AND2_X1 U5 ( .A1(n330), .A2(n218), .ZN(n190) );
  AND2_X1 U7 ( .A1(n330), .A2(n218), .ZN(net187832) );
  CLKBUF_X1 U8 ( .A(\carry[23] ), .Z(n299) );
  CLKBUF_X1 U9 ( .A(n268), .Z(n273) );
  BUF_X1 U10 ( .A(n327), .Z(n191) );
  INV_X1 U11 ( .A(B[33]), .ZN(n193) );
  AOI21_X1 U12 ( .B1(n350), .B2(n340), .A(n249), .ZN(n247) );
  OAI21_X1 U13 ( .B1(A[7]), .B2(n236), .A(n334), .ZN(n234) );
  INV_X1 U14 ( .A(B[24]), .ZN(n260) );
  AND2_X1 U15 ( .A1(n197), .A2(n196), .ZN(n192) );
  BUF_X1 U16 ( .A(A[11]), .Z(n298) );
  CLKBUF_X1 U17 ( .A(A[9]), .Z(n305) );
  XNOR2_X1 U18 ( .A(A[33]), .B(n193), .ZN(n219) );
  CLKBUF_X1 U19 ( .A(n218), .Z(n194) );
  OR2_X1 U20 ( .A1(n269), .A2(n301), .ZN(n195) );
  XNOR2_X1 U21 ( .A(B[20]), .B(A[20]), .ZN(n300) );
  CLKBUF_X1 U22 ( .A(A[20]), .Z(n311) );
  NAND2_X1 U23 ( .A1(n191), .A2(n264), .ZN(n196) );
  NAND2_X1 U24 ( .A1(n259), .A2(B[18]), .ZN(n197) );
  NAND2_X1 U25 ( .A1(n197), .A2(n196), .ZN(n198) );
  BUF_X1 U26 ( .A(n327), .Z(n307) );
  INV_X1 U27 ( .A(B[32]), .ZN(n308) );
  CLKBUF_X1 U28 ( .A(A[17]), .Z(n282) );
  NOR2_X1 U29 ( .A1(n200), .A2(n201), .ZN(n199) );
  NOR2_X1 U30 ( .A1(net184427), .A2(B[13]), .ZN(n200) );
  NOR2_X1 U31 ( .A1(n274), .A2(B[13]), .ZN(n201) );
  BUF_X1 U32 ( .A(A[13]), .Z(net184427) );
  INV_X1 U33 ( .A(B[26]), .ZN(n313) );
  XNOR2_X1 U34 ( .A(n188), .B(n202), .ZN(SUM[34]) );
  XNOR2_X1 U35 ( .A(A[34]), .B(B[34]), .ZN(n202) );
  INV_X1 U36 ( .A(B[16]), .ZN(n316) );
  INV_X1 U37 ( .A(B[12]), .ZN(n208) );
  INV_X1 U38 ( .A(B[19]), .ZN(n312) );
  OAI21_X1 U39 ( .B1(n270), .B2(A[14]), .A(B[14]), .ZN(n272) );
  OAI21_X1 U40 ( .B1(n190), .B2(n209), .A(B[12]), .ZN(n203) );
  OAI21_X1 U41 ( .B1(n210), .B2(n211), .A(n203), .ZN(n204) );
  INV_X1 U42 ( .A(n340), .ZN(n205) );
  XNOR2_X1 U43 ( .A(n207), .B(n204), .ZN(SUM[13]) );
  XNOR2_X1 U44 ( .A(A[13]), .B(B[13]), .ZN(n207) );
  OAI21_X1 U45 ( .B1(n210), .B2(n211), .A(n278), .ZN(n274) );
  OAI21_X1 U46 ( .B1(net187832), .B2(n209), .A(B[12]), .ZN(n278) );
  INV_X1 U47 ( .A(n206), .ZN(n209) );
  INV_X1 U48 ( .A(A[12]), .ZN(n206) );
  CLKBUF_X1 U49 ( .A(n206), .Z(n211) );
  INV_X1 U50 ( .A(n190), .ZN(n210) );
  XNOR2_X1 U51 ( .A(A[12]), .B(n208), .ZN(n279) );
  OR2_X1 U52 ( .A1(n234), .A2(n345), .ZN(n212) );
  NAND2_X1 U53 ( .A1(n212), .A2(n287), .ZN(n232) );
  NAND3_X1 U54 ( .A1(n302), .A2(n304), .A3(n303), .ZN(n213) );
  XNOR2_X1 U55 ( .A(n297), .B(A[23]), .ZN(SUM[23]) );
  NAND2_X1 U56 ( .A1(n188), .A2(A[34]), .ZN(n214) );
  NAND2_X1 U57 ( .A1(carry[34]), .A2(B[34]), .ZN(n215) );
  NAND2_X1 U58 ( .A1(A[34]), .A2(B[34]), .ZN(n216) );
  NAND3_X1 U59 ( .A1(n214), .A2(n215), .A3(n216), .ZN(carry[35]) );
  XNOR2_X1 U60 ( .A(A[32]), .B(B[32]), .ZN(n252) );
  CLKBUF_X1 U61 ( .A(A[26]), .Z(n217) );
  XNOR2_X1 U62 ( .A(n205), .B(n323), .ZN(SUM[39]) );
  OR2_X1 U63 ( .A1(n276), .A2(n298), .ZN(n218) );
  NAND2_X1 U64 ( .A1(n194), .A2(n330), .ZN(n277) );
  XOR2_X1 U65 ( .A(n324), .B(n219), .Z(SUM[33]) );
  NAND2_X1 U66 ( .A1(n324), .A2(A[33]), .ZN(n220) );
  NAND2_X1 U67 ( .A1(n324), .A2(B[33]), .ZN(n221) );
  NAND2_X1 U68 ( .A1(A[33]), .A2(B[33]), .ZN(n222) );
  NAND3_X1 U69 ( .A1(n220), .A2(n221), .A3(n222), .ZN(carry[34]) );
  XNOR2_X1 U70 ( .A(n307), .B(n229), .ZN(SUM[18]) );
  XNOR2_X1 U71 ( .A(A[18]), .B(B[18]), .ZN(n229) );
  XNOR2_X1 U72 ( .A(\carry[32] ), .B(n252), .ZN(SUM[32]) );
  CLKBUF_X1 U73 ( .A(A[19]), .Z(n254) );
  NAND2_X1 U74 ( .A1(n231), .A2(n255), .ZN(n275) );
  NAND2_X1 U75 ( .A1(n230), .A2(n311), .ZN(n255) );
  XNOR2_X1 U76 ( .A(A[24]), .B(n260), .ZN(n228) );
  CLKBUF_X1 U77 ( .A(A[18]), .Z(n264) );
  OAI21_X1 U78 ( .B1(n331), .B2(A[10]), .A(B[10]), .ZN(n265) );
  OAI21_X1 U79 ( .B1(net183027), .B2(net186686), .A(n199), .ZN(n267) );
  INV_X1 U80 ( .A(n271), .ZN(n270) );
  CLKBUF_X1 U81 ( .A(n262), .Z(n317) );
  OAI21_X1 U82 ( .B1(n315), .B2(n344), .A(n265), .ZN(n276) );
  XNOR2_X1 U83 ( .A(\carry[23] ), .B(B[23]), .ZN(n297) );
  XNOR2_X1 U84 ( .A(n189), .B(n300), .ZN(SUM[20]) );
  NOR2_X1 U85 ( .A1(n269), .A2(n301), .ZN(n309) );
  NOR2_X1 U86 ( .A1(n268), .A2(A[15]), .ZN(n301) );
  NAND2_X1 U87 ( .A1(A[23]), .A2(n299), .ZN(n302) );
  NAND2_X1 U88 ( .A1(A[23]), .A2(B[23]), .ZN(n303) );
  NAND2_X1 U104 ( .A1(n299), .A2(B[23]), .ZN(n304) );
  NAND3_X1 U105 ( .A1(n302), .A2(n303), .A3(n304), .ZN(\carry[24] ) );
  AOI21_X1 U106 ( .B1(n192), .B2(n341), .A(n256), .ZN(n230) );
  XNOR2_X1 U107 ( .A(n306), .B(n273), .ZN(SUM[15]) );
  XNOR2_X1 U111 ( .A(A[15]), .B(B[15]), .ZN(n306) );
  CLKBUF_X1 U113 ( .A(net184427), .Z(net183027) );
  XNOR2_X1 U114 ( .A(A[32]), .B(n308), .ZN(n224) );
  XNOR2_X1 U115 ( .A(n192), .B(n258), .ZN(SUM[19]) );
  CLKBUF_X1 U118 ( .A(A[32]), .Z(n310) );
  XNOR2_X1 U119 ( .A(A[19]), .B(n312), .ZN(n258) );
  XNOR2_X1 U120 ( .A(n195), .B(n320), .ZN(SUM[16]) );
  XNOR2_X1 U121 ( .A(A[26]), .B(n313), .ZN(n226) );
  OR2_X1 U122 ( .A1(n267), .A2(n343), .ZN(n314) );
  NAND2_X1 U123 ( .A1(n272), .A2(n314), .ZN(n268) );
  XNOR2_X1 U124 ( .A(A[16]), .B(n316), .ZN(n320) );
  XNOR2_X1 U125 ( .A(n277), .B(n279), .ZN(SUM[12]) );
  CLKBUF_X1 U126 ( .A(A[24]), .Z(n318) );
  XNOR2_X1 U127 ( .A(n317), .B(n319), .ZN(SUM[17]) );
  XNOR2_X1 U128 ( .A(A[17]), .B(B[17]), .ZN(n319) );
  INV_X1 U129 ( .A(n254), .ZN(n341) );
  INV_X1 U130 ( .A(n267), .ZN(n329) );
  INV_X1 U131 ( .A(A[10]), .ZN(n344) );
  XNOR2_X1 U132 ( .A(n321), .B(n329), .ZN(SUM[14]) );
  XNOR2_X1 U133 ( .A(A[14]), .B(B[14]), .ZN(n321) );
  INV_X1 U137 ( .A(A[14]), .ZN(n343) );
  INV_X1 U138 ( .A(A[16]), .ZN(n342) );
  XNOR2_X1 U139 ( .A(n322), .B(n276), .ZN(SUM[11]) );
  XNOR2_X1 U140 ( .A(A[11]), .B(B[11]), .ZN(n322) );
  AOI22_X1 U141 ( .A1(B[32]), .A2(n310), .B1(n224), .B2(\carry[32] ), .ZN(n223) );
  AOI22_X1 U142 ( .A1(B[26]), .A2(n217), .B1(\carry[26] ), .B2(n226), .ZN(n225) );
  AOI22_X1 U143 ( .A1(B[24]), .A2(n318), .B1(n228), .B2(\carry[24] ), .ZN(n227) );
  INV_X1 U144 ( .A(n227), .ZN(n326) );
  INV_X1 U145 ( .A(A[8]), .ZN(n345) );
  XNOR2_X1 U146 ( .A(carry[39]), .B(B[39]), .ZN(n323) );
  INV_X1 U147 ( .A(B[39]), .ZN(n350) );
  INV_X1 U148 ( .A(A[39]), .ZN(n340) );
  AOI21_X1 U149 ( .B1(A[39]), .B2(B[39]), .A(carry[39]), .ZN(n249) );
  INV_X1 U150 ( .A(n223), .ZN(n324) );
  INV_X1 U151 ( .A(n225), .ZN(n325) );
  AND2_X1 U152 ( .A1(A[40]), .A2(n247), .ZN(n246) );
  INV_X1 U153 ( .A(A[6]), .ZN(n346) );
  INV_X1 U154 ( .A(n294), .ZN(n338) );
  INV_X1 U155 ( .A(n286), .ZN(n332) );
  OAI22_X1 U156 ( .A1(n246), .A2(B[40]), .B1(n247), .B2(A[40]), .ZN(n244) );
  OAI21_X1 U157 ( .B1(A[8]), .B2(n333), .A(B[8]), .ZN(n287) );
  INV_X1 U158 ( .A(n234), .ZN(n333) );
  XNOR2_X1 U159 ( .A(A[3]), .B(B[3]), .ZN(n250) );
  INV_X1 U160 ( .A(A[2]), .ZN(n348) );
  INV_X1 U161 ( .A(A[4]), .ZN(n347) );
  OAI22_X1 U162 ( .A1(A[3]), .A2(n251), .B1(B[3]), .B2(n292), .ZN(n242) );
  AND2_X1 U163 ( .A1(n251), .A2(A[3]), .ZN(n292) );
  OAI21_X1 U164 ( .B1(n338), .B2(n348), .A(n293), .ZN(n251) );
  OAI21_X1 U165 ( .B1(n294), .B2(A[2]), .A(B[2]), .ZN(n293) );
  OAI21_X1 U166 ( .B1(A[5]), .B2(n240), .A(n336), .ZN(n238) );
  INV_X1 U167 ( .A(n290), .ZN(n336) );
  AOI21_X1 U168 ( .B1(n240), .B2(A[5]), .A(B[5]), .ZN(n290) );
  INV_X1 U169 ( .A(n288), .ZN(n334) );
  AOI21_X1 U170 ( .B1(n236), .B2(A[7]), .A(B[7]), .ZN(n288) );
  OAI21_X1 U171 ( .B1(n238), .B2(n346), .A(n289), .ZN(n236) );
  OAI21_X1 U172 ( .B1(n335), .B2(A[6]), .A(B[6]), .ZN(n289) );
  INV_X1 U173 ( .A(n238), .ZN(n335) );
  OAI21_X1 U174 ( .B1(n242), .B2(n347), .A(n291), .ZN(n240) );
  OAI21_X1 U175 ( .B1(n337), .B2(A[4]), .A(B[4]), .ZN(n291) );
  INV_X1 U176 ( .A(n242), .ZN(n337) );
  AOI21_X1 U177 ( .B1(n349), .B2(n295), .A(n296), .ZN(n294) );
  INV_X1 U178 ( .A(A[1]), .ZN(n349) );
  AOI21_X1 U179 ( .B1(n339), .B2(A[1]), .A(B[1]), .ZN(n296) );
  INV_X1 U180 ( .A(n295), .ZN(n339) );
  XNOR2_X1 U181 ( .A(n250), .B(n251), .ZN(SUM[3]) );
  NAND2_X1 U182 ( .A1(B[0]), .A2(A[0]), .ZN(n295) );
  OAI21_X1 U183 ( .B1(n309), .B2(A[16]), .A(B[16]), .ZN(n266) );
  INV_X1 U184 ( .A(n263), .ZN(n328) );
  OAI21_X1 U185 ( .B1(n305), .B2(n232), .A(n332), .ZN(n283) );
  AOI21_X1 U186 ( .B1(n232), .B2(A[9]), .A(B[9]), .ZN(n286) );
  OR2_X1 U187 ( .A1(n327), .A2(A[18]), .ZN(n259) );
  INV_X1 U188 ( .A(n283), .ZN(n331) );
  INV_X1 U189 ( .A(n281), .ZN(n330) );
  INV_X1 U190 ( .A(n261), .ZN(n327) );
  AOI21_X1 U191 ( .B1(n280), .B2(n298), .A(B[11]), .ZN(n281) );
  OAI21_X1 U192 ( .B1(n195), .B2(n342), .A(n266), .ZN(n262) );
  OAI21_X1 U193 ( .B1(n315), .B2(n344), .A(n284), .ZN(n280) );
  OAI21_X1 U194 ( .B1(n331), .B2(A[10]), .A(B[10]), .ZN(n284) );
  AOI21_X1 U195 ( .B1(n198), .B2(A[19]), .A(B[19]), .ZN(n256) );
  OAI21_X1 U196 ( .B1(net183027), .B2(net186686), .A(n199), .ZN(n271) );
  OAI21_X1 U197 ( .B1(n230), .B2(A[20]), .A(B[20]), .ZN(n231) );
  OAI21_X1 U198 ( .B1(n282), .B2(n317), .A(n328), .ZN(n261) );
  AOI21_X1 U199 ( .B1(n262), .B2(A[17]), .A(B[17]), .ZN(n263) );
  AOI21_X1 U200 ( .B1(n268), .B2(A[15]), .A(B[15]), .ZN(n269) );
endmodule


module RCA_NBIT42 ( A, B, Ci, S, Co );
  input [41:0] A;
  input [41:0] B;
  output [41:0] S;
  input Ci;
  output Co;

  assign Co = 1'b0;

  RCA_NBIT42_DW01_add_0 add_95 ( .A(A), .B(B), .CI(1'b0), .SUM(S) );
endmodule


module RCA_NBIT44_DW01_add_0 ( A, B, CI, SUM, CO );
  input [43:0] A;
  input [43:0] B;
  output [43:0] SUM;
  input CI;
  output CO;
  wire   \carry[43] , n1, \carry[9] , \carry[8] , \carry[7] , \carry[6] ,
         \carry[5] , \carry[4] , \carry[3] , \carry[2] , \carry[10] , n305,
         n306, n310, n311, n312, n313, n316, n317, n318, n319, n321, n322,
         n323, n324, n325, n327, n328, n329, n330, n331, n333, n334, n335,
         n336, n337, n339, n340, n341, n342, n343, n345, n346, n347, n348,
         n349, n351, n352, n353, n354, n355, n356, n357, n358, n361, n362,
         n363, n364, n366, n367, n368, n369, n370, n372, n373, n374, n375,
         n376, n378, n379, n380, n381, n382, net176555, net186695, n389, n302,
         n390, n387, n386, n384, n303, \carry[14] , \carry[13] , n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n304, n307, n308, n309, n314,
         n315, n320, n326, n332, n338, n344, n350, n359, n360, n365, n371,
         n377, n383, n385, n388, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477;

  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(\carry[2] ), .S(SUM[1]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(\carry[5] ), .CO(\carry[6] ), .S(SUM[5]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(\carry[6] ), .CO(\carry[7] ), .S(SUM[6]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(\carry[7] ), .CO(\carry[8] ), .S(SUM[7]) );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(\carry[8] ), .CO(\carry[9] ), .S(SUM[8]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(\carry[9] ), .CO(\carry[10] ), .S(
        SUM[9]) );
  XOR2_X1 U163 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  XOR2_X1 U161 ( .A(\carry[10] ), .B(n389), .Z(SUM[10]) );
  XOR2_X1 U162 ( .A(A[10]), .B(B[10]), .Z(n389) );
  XOR2_X1 U160 ( .A(n303), .B(n302), .Z(SUM[11]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(n390), .CO(\carry[13] ), .S(SUM[12])
         );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(\carry[13] ), .CO(\carry[14] ), .S(
        SUM[13]) );
  CLKBUF_X1 U1 ( .A(n354), .Z(n411) );
  BUF_X1 U2 ( .A(n364), .Z(n263) );
  NAND2_X1 U3 ( .A1(n274), .A2(n275), .ZN(n261) );
  BUF_X1 U4 ( .A(n330), .Z(n403) );
  CLKBUF_X1 U5 ( .A(A[31]), .Z(n262) );
  CLKBUF_X1 U6 ( .A(n439), .Z(n292) );
  OR2_X1 U7 ( .A1(n330), .A2(n383), .ZN(n331) );
  INV_X1 U8 ( .A(B[15]), .ZN(n298) );
  INV_X1 U9 ( .A(B[19]), .ZN(n393) );
  INV_X1 U10 ( .A(B[23]), .ZN(n442) );
  INV_X1 U11 ( .A(B[16]), .ZN(n408) );
  INV_X1 U12 ( .A(B[34]), .ZN(n417) );
  CLKBUF_X1 U13 ( .A(n305), .Z(n264) );
  NOR2_X1 U14 ( .A1(n328), .A2(n407), .ZN(n265) );
  OR2_X1 U15 ( .A1(n433), .A2(n477), .ZN(n437) );
  CLKBUF_X1 U16 ( .A(n372), .Z(n320) );
  BUF_X1 U17 ( .A(A[18]), .Z(n436) );
  OAI22_X1 U18 ( .A1(n304), .A2(n299), .B1(B[15]), .B2(n384), .ZN(n266) );
  CLKBUF_X1 U19 ( .A(A[29]), .Z(n267) );
  CLKBUF_X1 U20 ( .A(n383), .Z(n326) );
  AOI21_X1 U21 ( .B1(n385), .B2(n474), .A(n271), .ZN(n268) );
  OAI21_X1 U22 ( .B1(A[35]), .B2(n324), .A(B[35]), .ZN(n269) );
  CLKBUF_X1 U23 ( .A(n339), .Z(n429) );
  OR2_X1 U24 ( .A1(n426), .A2(n349), .ZN(n270) );
  AOI21_X1 U25 ( .B1(n460), .B2(A[25]), .A(B[25]), .ZN(n271) );
  BUF_X1 U26 ( .A(A[16]), .Z(n402) );
  NOR2_X1 U27 ( .A1(n287), .A2(n414), .ZN(n272) );
  NOR2_X1 U28 ( .A1(n272), .A2(n263), .ZN(n273) );
  BUF_X1 U29 ( .A(n363), .Z(n414) );
  NAND2_X1 U30 ( .A1(n264), .A2(A[41]), .ZN(n274) );
  NAND2_X1 U31 ( .A1(n306), .A2(B[41]), .ZN(n275) );
  NAND2_X1 U32 ( .A1(n274), .A2(n275), .ZN(n276) );
  INV_X1 U33 ( .A(B[28]), .ZN(n398) );
  INV_X1 U34 ( .A(B[30]), .ZN(n418) );
  BUF_X1 U35 ( .A(n336), .Z(n405) );
  INV_X1 U36 ( .A(B[36]), .ZN(n344) );
  INV_X1 U37 ( .A(B[37]), .ZN(n314) );
  INV_X1 U38 ( .A(B[21]), .ZN(n430) );
  INV_X1 U39 ( .A(B[25]), .ZN(n415) );
  INV_X1 U40 ( .A(B[17]), .ZN(n443) );
  AND2_X1 U41 ( .A1(n432), .A2(n463), .ZN(n413) );
  NOR2_X1 U42 ( .A1(n359), .A2(n338), .ZN(n404) );
  XNOR2_X1 U43 ( .A(n446), .B(n281), .ZN(SUM[20]) );
  XNOR2_X1 U44 ( .A(n288), .B(n335), .ZN(SUM[32]) );
  AOI21_X1 U45 ( .B1(n277), .B2(n278), .A(n387), .ZN(n296) );
  INV_X1 U46 ( .A(B[14]), .ZN(n277) );
  INV_X1 U47 ( .A(A[14]), .ZN(n278) );
  NOR2_X1 U48 ( .A1(n316), .A2(n434), .ZN(n312) );
  OAI21_X1 U49 ( .B1(n397), .B2(n279), .A(n417), .ZN(n280) );
  INV_X1 U50 ( .A(A[34]), .ZN(n279) );
  INV_X1 U51 ( .A(n280), .ZN(n328) );
  CLKBUF_X1 U52 ( .A(A[23]), .Z(n290) );
  NAND2_X1 U53 ( .A1(n440), .A2(n373), .ZN(n281) );
  INV_X1 U54 ( .A(n469), .ZN(n282) );
  XNOR2_X1 U55 ( .A(n265), .B(n449), .ZN(SUM[35]) );
  INV_X1 U56 ( .A(n286), .ZN(n283) );
  AOI21_X1 U57 ( .B1(n350), .B2(n282), .A(B[36]), .ZN(n284) );
  AND2_X1 U58 ( .A1(n285), .A2(n269), .ZN(n410) );
  AND2_X1 U59 ( .A1(n394), .A2(n469), .ZN(n285) );
  OAI21_X1 U60 ( .B1(n287), .B2(n414), .A(n462), .ZN(n286) );
  CLKBUF_X1 U61 ( .A(A[22]), .Z(n287) );
  AOI22_X1 U62 ( .A1(n405), .A2(n262), .B1(n337), .B2(B[31]), .ZN(n288) );
  OR2_X1 U63 ( .A1(n360), .A2(n454), .ZN(n289) );
  OR2_X1 U64 ( .A1(n365), .A2(n454), .ZN(n293) );
  XNOR2_X1 U65 ( .A(n261), .B(n291), .ZN(SUM[42]) );
  XNOR2_X1 U66 ( .A(A[42]), .B(B[42]), .ZN(n291) );
  CLKBUF_X1 U67 ( .A(A[15]), .Z(n304) );
  XNOR2_X1 U68 ( .A(n300), .B(n386), .ZN(SUM[15]) );
  XNOR2_X1 U69 ( .A(A[15]), .B(n298), .ZN(n386) );
  INV_X1 U70 ( .A(n299), .ZN(n300) );
  BUF_X1 U71 ( .A(n296), .Z(n299) );
  OAI22_X1 U72 ( .A1(n304), .A2(n299), .B1(n384), .B2(B[15]), .ZN(n382) );
  AND2_X1 U73 ( .A1(A[15]), .A2(n296), .ZN(n384) );
  AOI21_X1 U74 ( .B1(A[14]), .B2(B[14]), .A(\carry[14] ), .ZN(n387) );
  CLKBUF_X1 U75 ( .A(A[14]), .Z(n301) );
  XNOR2_X1 U76 ( .A(n301), .B(n297), .ZN(SUM[14]) );
  XNOR2_X1 U77 ( .A(\carry[14] ), .B(B[14]), .ZN(n297) );
  OAI22_X1 U78 ( .A1(n294), .A2(n295), .B1(n302), .B2(n303), .ZN(n390) );
  INV_X1 U79 ( .A(A[11]), .ZN(n295) );
  INV_X1 U80 ( .A(B[11]), .ZN(n294) );
  XNOR2_X1 U81 ( .A(A[11]), .B(B[11]), .ZN(n303) );
  XNOR2_X1 U82 ( .A(n305), .B(n307), .ZN(SUM[41]) );
  XNOR2_X1 U83 ( .A(B[41]), .B(A[41]), .ZN(n307) );
  XNOR2_X1 U84 ( .A(n332), .B(n308), .ZN(SUM[37]) );
  XOR2_X1 U85 ( .A(n314), .B(A[37]), .Z(n308) );
  AND2_X1 U86 ( .A1(n268), .A2(A[26]), .ZN(n309) );
  CLKBUF_X1 U87 ( .A(A[24]), .Z(n315) );
  XOR2_X1 U88 ( .A(B[38]), .B(A[38]), .Z(n317) );
  NOR2_X1 U89 ( .A1(n284), .A2(n410), .ZN(n332) );
  AOI22_X1 U90 ( .A1(B[10]), .A2(A[10]), .B1(n389), .B2(\carry[10] ), .ZN(n302) );
  AOI21_X1 U91 ( .B1(n375), .B2(n436), .A(B[18]), .ZN(n338) );
  CLKBUF_X1 U92 ( .A(n286), .Z(n401) );
  BUF_X1 U93 ( .A(n411), .Z(n385) );
  XNOR2_X1 U94 ( .A(A[36]), .B(n344), .ZN(n323) );
  NAND2_X1 U95 ( .A1(n325), .A2(n394), .ZN(n350) );
  AND2_X1 U96 ( .A1(n394), .A2(n269), .ZN(n321) );
  NOR2_X1 U97 ( .A1(n436), .A2(n399), .ZN(n359) );
  BUF_X1 U98 ( .A(A[30]), .Z(n377) );
  AND2_X1 U99 ( .A1(n406), .A2(A[39]), .ZN(n360) );
  NOR2_X1 U100 ( .A1(n360), .A2(n454), .ZN(n400) );
  BUF_X1 U101 ( .A(n312), .Z(n406) );
  AND2_X1 U102 ( .A1(n406), .A2(A[39]), .ZN(n365) );
  CLKBUF_X1 U103 ( .A(n330), .Z(n371) );
  BUF_X1 U104 ( .A(A[33]), .Z(n383) );
  BUF_X1 U105 ( .A(n342), .Z(n409) );
  OAI21_X1 U106 ( .B1(n465), .B2(n391), .A(B[17]), .ZN(n388) );
  INV_X1 U107 ( .A(n477), .ZN(n391) );
  OAI21_X1 U108 ( .B1(n273), .B2(A[23]), .A(B[23]), .ZN(n392) );
  XNOR2_X1 U109 ( .A(A[19]), .B(n393), .ZN(n374) );
  NAND2_X1 U110 ( .A1(n324), .A2(A[35]), .ZN(n394) );
  BUF_X1 U111 ( .A(n288), .Z(n428) );
  OR2_X1 U112 ( .A1(n459), .A2(n427), .ZN(n395) );
  OR2_X1 U113 ( .A1(n459), .A2(n427), .ZN(n423) );
  OR2_X1 U114 ( .A1(n399), .A2(n436), .ZN(n396) );
  XOR2_X1 U115 ( .A(B[32]), .B(A[32]), .Z(n335) );
  AOI22_X1 U116 ( .A1(n371), .A2(n383), .B1(n331), .B2(B[33]), .ZN(n397) );
  XNOR2_X1 U117 ( .A(n398), .B(A[28]), .ZN(n347) );
  CLKBUF_X1 U118 ( .A(net176555), .Z(net186695) );
  NAND2_X1 U119 ( .A1(n388), .A2(n437), .ZN(n399) );
  AOI22_X1 U120 ( .A1(n371), .A2(n326), .B1(n331), .B2(B[33]), .ZN(n327) );
  XNOR2_X1 U121 ( .A(n453), .B(A[43]), .ZN(SUM[43]) );
  AND2_X1 U122 ( .A1(n279), .A2(n327), .ZN(n407) );
  NOR2_X1 U123 ( .A1(n407), .A2(n328), .ZN(n324) );
  XNOR2_X1 U124 ( .A(n408), .B(A[16]), .ZN(n441) );
  XNOR2_X1 U125 ( .A(n406), .B(n447), .ZN(SUM[39]) );
  NOR2_X1 U126 ( .A1(n410), .A2(n322), .ZN(n318) );
  AOI21_X1 U127 ( .B1(n385), .B2(n474), .A(n271), .ZN(n412) );
  XNOR2_X1 U128 ( .A(A[25]), .B(n415), .ZN(n356) );
  OR2_X1 U129 ( .A1(n455), .A2(n424), .ZN(n416) );
  XNOR2_X1 U130 ( .A(A[34]), .B(n417), .ZN(n329) );
  XNOR2_X1 U131 ( .A(A[30]), .B(n418), .ZN(n341) );
  NAND2_X1 U132 ( .A1(n276), .A2(A[42]), .ZN(n419) );
  NAND2_X1 U133 ( .A1(n261), .A2(B[42]), .ZN(n420) );
  NAND2_X1 U134 ( .A1(A[42]), .A2(B[42]), .ZN(n421) );
  NAND3_X1 U135 ( .A1(n420), .A2(n419), .A3(n421), .ZN(\carry[43] ) );
  NOR2_X1 U136 ( .A1(n455), .A2(n424), .ZN(n422) );
  AND2_X1 U137 ( .A1(n332), .A2(A[37]), .ZN(n424) );
  INV_X1 U138 ( .A(n289), .ZN(n425) );
  AND2_X1 U139 ( .A1(n348), .A2(n473), .ZN(n426) );
  NOR2_X1 U140 ( .A1(n349), .A2(n426), .ZN(n346) );
  AND2_X1 U141 ( .A1(n412), .A2(A[26]), .ZN(n427) );
  NOR2_X1 U142 ( .A1(n309), .A2(n459), .ZN(n348) );
  AOI22_X1 U143 ( .A1(n405), .A2(n262), .B1(n337), .B2(B[31]), .ZN(n333) );
  XNOR2_X1 U144 ( .A(A[21]), .B(n430), .ZN(n368) );
  NAND2_X1 U145 ( .A1(n361), .A2(n292), .ZN(n431) );
  NAND2_X1 U146 ( .A1(n464), .A2(n396), .ZN(n372) );
  OR2_X1 U147 ( .A1(n281), .A2(A[20]), .ZN(n432) );
  NAND2_X1 U148 ( .A1(n463), .A2(n432), .ZN(n366) );
  OAI22_X1 U149 ( .A1(n402), .A2(net186695), .B1(n381), .B2(B[16]), .ZN(n433)
         );
  XNOR2_X1 U150 ( .A(n405), .B(n451), .ZN(SUM[31]) );
  AND2_X1 U151 ( .A1(n422), .A2(n468), .ZN(n434) );
  XNOR2_X1 U152 ( .A(n414), .B(n435), .ZN(SUM[22]) );
  XNOR2_X1 U153 ( .A(A[22]), .B(B[22]), .ZN(n435) );
  XNOR2_X1 U154 ( .A(n452), .B(n409), .ZN(SUM[29]) );
  NAND2_X1 U155 ( .A1(n379), .A2(n437), .ZN(n375) );
  OR2_X1 U156 ( .A1(n476), .A2(n366), .ZN(n438) );
  NAND2_X1 U157 ( .A1(n367), .A2(n438), .ZN(n363) );
  OR2_X1 U158 ( .A1(n286), .A2(n475), .ZN(n439) );
  NAND2_X1 U159 ( .A1(n439), .A2(n392), .ZN(n357) );
  OR2_X1 U164 ( .A1(n372), .A2(n466), .ZN(n440) );
  NAND2_X1 U165 ( .A1(n440), .A2(n373), .ZN(n369) );
  XNOR2_X1 U166 ( .A(n266), .B(n441), .ZN(SUM[16]) );
  XNOR2_X1 U167 ( .A(A[23]), .B(n442), .ZN(n362) );
  XNOR2_X1 U168 ( .A(A[17]), .B(n443), .ZN(n380) );
  XNOR2_X1 U169 ( .A(n431), .B(n444), .ZN(SUM[24]) );
  XNOR2_X1 U170 ( .A(A[24]), .B(B[24]), .ZN(n444) );
  XNOR2_X1 U171 ( .A(n399), .B(n445), .ZN(SUM[18]) );
  XNOR2_X1 U172 ( .A(A[18]), .B(B[18]), .ZN(n445) );
  XNOR2_X1 U173 ( .A(A[20]), .B(B[20]), .ZN(n446) );
  INV_X1 U174 ( .A(A[32]), .ZN(n470) );
  INV_X1 U175 ( .A(A[25]), .ZN(n474) );
  AOI21_X1 U176 ( .B1(n416), .B2(A[38]), .A(B[38]), .ZN(n316) );
  XNOR2_X1 U177 ( .A(B[39]), .B(A[39]), .ZN(n447) );
  XNOR2_X1 U178 ( .A(n403), .B(n448), .ZN(SUM[33]) );
  XNOR2_X1 U179 ( .A(A[33]), .B(B[33]), .ZN(n448) );
  XNOR2_X1 U180 ( .A(B[35]), .B(A[35]), .ZN(n449) );
  XNOR2_X1 U181 ( .A(n450), .B(n423), .ZN(SUM[27]) );
  XNOR2_X1 U182 ( .A(A[27]), .B(B[27]), .ZN(n450) );
  AOI21_X1 U183 ( .B1(n350), .B2(n282), .A(B[36]), .ZN(n322) );
  XNOR2_X1 U184 ( .A(B[31]), .B(A[31]), .ZN(n451) );
  XNOR2_X1 U185 ( .A(B[40]), .B(n467), .ZN(n311) );
  AOI21_X1 U186 ( .B1(n293), .B2(A[40]), .A(B[40]), .ZN(n310) );
  OAI21_X1 U187 ( .B1(n290), .B2(n283), .A(B[23]), .ZN(n361) );
  OAI21_X1 U188 ( .B1(n413), .B2(A[21]), .A(B[21]), .ZN(n367) );
  INV_X1 U189 ( .A(A[17]), .ZN(n477) );
  OAI21_X1 U190 ( .B1(n465), .B2(n391), .A(B[17]), .ZN(n379) );
  OAI21_X1 U191 ( .B1(n270), .B2(n472), .A(n345), .ZN(n342) );
  INV_X1 U192 ( .A(A[28]), .ZN(n472) );
  AOI21_X1 U193 ( .B1(n428), .B2(n470), .A(n334), .ZN(n330) );
  AOI21_X1 U194 ( .B1(n456), .B2(A[32]), .A(B[32]), .ZN(n334) );
  INV_X1 U195 ( .A(n313), .ZN(n454) );
  OAI21_X1 U196 ( .B1(n312), .B2(A[39]), .A(B[39]), .ZN(n313) );
  INV_X1 U197 ( .A(n364), .ZN(n462) );
  INV_X1 U198 ( .A(n319), .ZN(n455) );
  XNOR2_X1 U199 ( .A(A[29]), .B(B[29]), .ZN(n452) );
  OAI21_X1 U200 ( .B1(n267), .B2(n409), .A(n458), .ZN(n339) );
  INV_X1 U201 ( .A(n343), .ZN(n458) );
  AOI21_X1 U202 ( .B1(n342), .B2(A[29]), .A(B[29]), .ZN(n343) );
  XNOR2_X1 U203 ( .A(n270), .B(n347), .ZN(SUM[28]) );
  INV_X1 U204 ( .A(n354), .ZN(n460) );
  XNOR2_X1 U205 ( .A(n356), .B(n411), .ZN(SUM[25]) );
  OAI21_X1 U206 ( .B1(n265), .B2(A[35]), .A(B[35]), .ZN(n325) );
  XNOR2_X1 U207 ( .A(A[26]), .B(B[26]), .ZN(n353) );
  OAI21_X1 U208 ( .B1(n457), .B2(A[30]), .A(B[30]), .ZN(n340) );
  INV_X1 U209 ( .A(A[40]), .ZN(n467) );
  INV_X1 U210 ( .A(A[38]), .ZN(n468) );
  INV_X1 U211 ( .A(A[36]), .ZN(n469) );
  INV_X1 U212 ( .A(n377), .ZN(n471) );
  OR2_X1 U213 ( .A1(n336), .A2(A[31]), .ZN(n337) );
  XNOR2_X1 U214 ( .A(\carry[43] ), .B(B[43]), .ZN(n453) );
  AND2_X1 U215 ( .A1(A[0]), .A2(B[0]), .ZN(n1) );
  AOI21_X1 U216 ( .B1(n395), .B2(A[27]), .A(B[27]), .ZN(n349) );
  INV_X1 U217 ( .A(A[27]), .ZN(n473) );
  OR2_X1 U218 ( .A1(n305), .A2(A[41]), .ZN(n306) );
  AOI21_X1 U219 ( .B1(n467), .B2(n425), .A(n310), .ZN(n305) );
  XNOR2_X1 U220 ( .A(n400), .B(n311), .ZN(SUM[40]) );
  XNOR2_X1 U221 ( .A(n422), .B(n317), .ZN(SUM[38]) );
  XNOR2_X1 U222 ( .A(n321), .B(n323), .ZN(SUM[36]) );
  OAI21_X1 U223 ( .B1(n318), .B2(A[37]), .A(B[37]), .ZN(n319) );
  XNOR2_X1 U224 ( .A(n327), .B(n329), .ZN(SUM[34]) );
  INV_X1 U225 ( .A(n333), .ZN(n456) );
  XNOR2_X1 U226 ( .A(n429), .B(n341), .ZN(SUM[30]) );
  OAI21_X1 U227 ( .B1(n429), .B2(n471), .A(n340), .ZN(n336) );
  INV_X1 U228 ( .A(n339), .ZN(n457) );
  OAI21_X1 U229 ( .B1(n346), .B2(A[28]), .A(B[28]), .ZN(n345) );
  XNOR2_X1 U230 ( .A(n268), .B(n353), .ZN(SUM[26]) );
  OAI21_X1 U231 ( .B1(n351), .B2(A[26]), .A(B[26]), .ZN(n352) );
  AOI21_X1 U232 ( .B1(n369), .B2(A[20]), .A(B[20]), .ZN(n370) );
  AOI21_X1 U233 ( .B1(n375), .B2(n436), .A(B[18]), .ZN(n376) );
  AOI21_X1 U234 ( .B1(n363), .B2(A[22]), .A(B[22]), .ZN(n364) );
  XNOR2_X1 U235 ( .A(n368), .B(n366), .ZN(SUM[21]) );
  XNOR2_X1 U236 ( .A(n320), .B(n374), .ZN(SUM[19]) );
  INV_X1 U237 ( .A(n378), .ZN(n465) );
  INV_X1 U238 ( .A(n382), .ZN(net176555) );
  OAI22_X1 U239 ( .A1(n402), .A2(net186695), .B1(n381), .B2(B[16]), .ZN(n378)
         );
  INV_X1 U240 ( .A(n358), .ZN(n461) );
  INV_X1 U241 ( .A(n352), .ZN(n459) );
  INV_X1 U242 ( .A(n376), .ZN(n464) );
  INV_X1 U243 ( .A(n370), .ZN(n463) );
  AOI21_X1 U244 ( .B1(n411), .B2(n474), .A(n355), .ZN(n351) );
  AOI21_X1 U245 ( .B1(n460), .B2(A[25]), .A(B[25]), .ZN(n355) );
  AND2_X1 U246 ( .A1(net176555), .A2(n402), .ZN(n381) );
  INV_X1 U247 ( .A(A[23]), .ZN(n475) );
  OAI21_X1 U248 ( .B1(n404), .B2(A[19]), .A(B[19]), .ZN(n373) );
  XNOR2_X1 U249 ( .A(n362), .B(n401), .ZN(SUM[23]) );
  XNOR2_X1 U250 ( .A(n433), .B(n380), .ZN(SUM[17]) );
  OAI21_X1 U251 ( .B1(n431), .B2(n315), .A(n461), .ZN(n354) );
  AOI21_X1 U252 ( .B1(n357), .B2(A[24]), .A(B[24]), .ZN(n358) );
  INV_X1 U253 ( .A(A[19]), .ZN(n466) );
  INV_X1 U254 ( .A(A[21]), .ZN(n476) );
endmodule


module RCA_NBIT44 ( A, B, Ci, S, Co );
  input [43:0] A;
  input [43:0] B;
  output [43:0] S;
  input Ci;
  output Co;

  assign Co = 1'b0;

  RCA_NBIT44_DW01_add_0 add_95 ( .A(A), .B(B), .CI(1'b0), .SUM(S) );
endmodule


module RCA_NBIT46_DW01_add_0 ( A, B, CI, SUM, CO );
  input [45:0] A;
  input [45:0] B;
  output [45:0] SUM;
  input CI;
  output CO;
  wire   n1, n193, n194, n195, n202, n203, n205, n206, n207, n208, n209, n212,
         n213, n215, n217, n223, n229, n232, n233, n235, n236, n239, n245,
         n256, n259, n260, n261, n265, n266, n267, n268, n269, n271, n272,
         n274, n275, n276, n277, n278, net176583, net176584, net176585,
         net176604, net176614, net180672, net182635, net182663, net182738,
         net182805, net182801, net182839, net182959, net183097, net183284,
         net183394, net183573, net183647, net183674, net183836, net184160,
         net184862, net184972, net184977, net185361, net185811, net186087,
         net187757, n242, n238, net191673, net194375, net194454, net197603,
         net197636, net201007, net201277, n230, n224, n221, n220, n218, n214,
         net186622, net183136, net182694, net182693, n190, n188, n187, n200,
         n197, n184, n183, \carry[42] , net185256, net183182, net182883,
         net176602, n251, n248, net184940, net184399, net183088, net176581,
         n257, n255, n254, n250, n325, n326, n327, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481;
  wire   [45:1] carry;

  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U169 ( .A(A[18]), .B(B[18]), .Z(n261) );
  XOR2_X1 U175 ( .A(n455), .B(B[13]), .Z(n276) );
  XOR2_X1 U176 ( .A(A[12]), .B(n278), .Z(SUM[12]) );
  XOR2_X1 U177 ( .A(carry[12]), .B(B[12]), .Z(n278) );
  XOR2_X1 U178 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  NAND2_X1 U1 ( .A1(n326), .A2(n254), .ZN(n325) );
  OR2_X1 U2 ( .A1(net176581), .A2(n360), .ZN(n326) );
  NAND2_X1 U3 ( .A1(n326), .A2(n254), .ZN(n250) );
  AND2_X1 U4 ( .A1(n194), .A2(net194454), .ZN(n327) );
  XOR2_X1 U5 ( .A(n401), .B(n217), .Z(SUM[32]) );
  BUF_X1 U6 ( .A(n205), .Z(n412) );
  BUF_X1 U7 ( .A(n448), .Z(n329) );
  BUF_X1 U8 ( .A(A[29]), .Z(net187757) );
  CLKBUF_X1 U9 ( .A(A[34]), .Z(n330) );
  OR2_X1 U10 ( .A1(net185256), .A2(net176602), .ZN(n365) );
  AOI21_X1 U11 ( .B1(n341), .B2(n350), .A(n351), .ZN(n390) );
  INV_X1 U12 ( .A(B[15]), .ZN(n406) );
  INV_X1 U13 ( .A(B[44]), .ZN(n385) );
  NAND2_X1 U14 ( .A1(n248), .A2(n342), .ZN(n331) );
  CLKBUF_X1 U15 ( .A(A[33]), .Z(n396) );
  OR2_X1 U16 ( .A1(n468), .A2(n465), .ZN(n332) );
  OR2_X1 U17 ( .A1(n468), .A2(n465), .ZN(net183573) );
  BUF_X1 U18 ( .A(A[21]), .Z(net183182) );
  OAI21_X1 U19 ( .B1(n470), .B2(n433), .A(B[18]), .ZN(n333) );
  OR2_X1 U20 ( .A1(net176604), .A2(net184972), .ZN(net183394) );
  OAI21_X1 U21 ( .B1(n256), .B2(n358), .A(B[19]), .ZN(n334) );
  INV_X1 U22 ( .A(n344), .ZN(n335) );
  NOR2_X1 U23 ( .A1(net191673), .A2(net176614), .ZN(n336) );
  BUF_X1 U24 ( .A(A[24]), .Z(n419) );
  BUF_X1 U25 ( .A(A[25]), .Z(n418) );
  NAND2_X1 U26 ( .A1(n260), .A2(n424), .ZN(n337) );
  NAND2_X1 U27 ( .A1(n215), .A2(n338), .ZN(n416) );
  NAND2_X1 U28 ( .A1(n396), .A2(n395), .ZN(n338) );
  NAND2_X1 U29 ( .A1(n340), .A2(B[28]), .ZN(n339) );
  NAND2_X1 U30 ( .A1(n229), .A2(net176584), .ZN(n340) );
  AND2_X1 U31 ( .A1(n230), .A2(net182839), .ZN(n341) );
  INV_X1 U32 ( .A(B[26]), .ZN(n409) );
  NAND2_X1 U33 ( .A1(n365), .A2(n364), .ZN(n342) );
  NAND2_X1 U34 ( .A1(n343), .A2(B[40]), .ZN(n374) );
  INV_X1 U35 ( .A(A[40]), .ZN(n344) );
  NAND2_X1 U36 ( .A1(n345), .A2(n344), .ZN(n343) );
  NOR2_X1 U37 ( .A1(n368), .A2(n369), .ZN(n345) );
  AOI22_X1 U38 ( .A1(n443), .A2(n450), .B1(n268), .B2(B[15]), .ZN(n346) );
  BUF_X1 U39 ( .A(n473), .Z(n450) );
  INV_X1 U40 ( .A(B[40]), .ZN(net194375) );
  INV_X1 U41 ( .A(B[38]), .ZN(n347) );
  XNOR2_X1 U42 ( .A(A[38]), .B(n347), .ZN(n349) );
  CLKBUF_X1 U43 ( .A(n208), .Z(n413) );
  BUF_X1 U44 ( .A(A[41]), .Z(n371) );
  AND2_X1 U45 ( .A1(n266), .A2(n451), .ZN(n348) );
  INV_X1 U46 ( .A(B[34]), .ZN(n432) );
  XNOR2_X1 U47 ( .A(net182959), .B(n349), .ZN(SUM[38]) );
  INV_X1 U48 ( .A(B[36]), .ZN(n425) );
  INV_X1 U49 ( .A(B[20]), .ZN(n359) );
  INV_X1 U50 ( .A(B[16]), .ZN(n415) );
  BUF_X1 U51 ( .A(n474), .Z(n458) );
  INV_X1 U52 ( .A(B[24]), .ZN(n408) );
  INV_X1 U53 ( .A(B[30]), .ZN(net185811) );
  INV_X1 U54 ( .A(A[29]), .ZN(n350) );
  INV_X1 U55 ( .A(B[29]), .ZN(n351) );
  AND2_X1 U56 ( .A1(n208), .A2(A[35]), .ZN(n445) );
  AOI21_X1 U57 ( .B1(n346), .B2(n481), .A(n415), .ZN(n352) );
  INV_X1 U58 ( .A(n352), .ZN(n437) );
  AOI21_X1 U59 ( .B1(n348), .B2(n353), .A(n354), .ZN(n471) );
  INV_X1 U60 ( .A(A[17]), .ZN(n353) );
  INV_X1 U61 ( .A(B[17]), .ZN(n354) );
  AOI22_X1 U62 ( .A1(n271), .A2(B[14]), .B1(n458), .B2(A[14]), .ZN(n269) );
  XNOR2_X1 U63 ( .A(n355), .B(n356), .ZN(SUM[45]) );
  NAND2_X1 U64 ( .A1(n379), .A2(n378), .ZN(n355) );
  XNOR2_X1 U65 ( .A(B[45]), .B(A[45]), .ZN(n356) );
  XNOR2_X1 U66 ( .A(net182883), .B(n325), .ZN(SUM[21]) );
  AND2_X1 U67 ( .A1(n325), .A2(net183182), .ZN(net185256) );
  OAI21_X1 U68 ( .B1(n250), .B2(net183182), .A(B[21]), .ZN(n251) );
  OAI21_X1 U69 ( .B1(net184940), .B2(net183088), .A(B[20]), .ZN(n254) );
  INV_X1 U70 ( .A(net176581), .ZN(net183088) );
  INV_X1 U71 ( .A(A[20]), .ZN(net176581) );
  NAND2_X1 U72 ( .A1(n334), .A2(net184399), .ZN(net184940) );
  AND2_X1 U73 ( .A1(n257), .A2(net184399), .ZN(n360) );
  XNOR2_X1 U74 ( .A(n360), .B(n255), .ZN(SUM[20]) );
  XNOR2_X1 U75 ( .A(A[20]), .B(n359), .ZN(n255) );
  OAI21_X1 U76 ( .B1(n256), .B2(n358), .A(B[19]), .ZN(n257) );
  CLKBUF_X1 U77 ( .A(A[19]), .Z(n358) );
  NAND2_X1 U78 ( .A1(n337), .A2(n358), .ZN(net184399) );
  XNOR2_X1 U79 ( .A(n337), .B(n357), .ZN(SUM[19]) );
  XNOR2_X1 U80 ( .A(A[19]), .B(B[19]), .ZN(n357) );
  AND2_X1 U81 ( .A1(n331), .A2(net180672), .ZN(net184972) );
  OAI21_X1 U82 ( .B1(n331), .B2(net180672), .A(B[23]), .ZN(n245) );
  XNOR2_X1 U83 ( .A(n331), .B(net183097), .ZN(SUM[23]) );
  OAI21_X1 U84 ( .B1(n363), .B2(n364), .A(B[22]), .ZN(n248) );
  INV_X1 U85 ( .A(n361), .ZN(n364) );
  INV_X1 U86 ( .A(A[22]), .ZN(n361) );
  OR2_X1 U87 ( .A1(net176602), .A2(net185256), .ZN(n363) );
  INV_X1 U88 ( .A(n251), .ZN(net176602) );
  XNOR2_X1 U89 ( .A(A[22]), .B(B[22]), .ZN(n362) );
  XNOR2_X1 U90 ( .A(A[21]), .B(B[21]), .ZN(net182883) );
  XNOR2_X1 U91 ( .A(n365), .B(n362), .ZN(SUM[22]) );
  OAI21_X1 U92 ( .B1(n327), .B2(n367), .A(n183), .ZN(\carry[42] ) );
  NAND2_X1 U93 ( .A1(\carry[42] ), .A2(B[42]), .ZN(net182694) );
  NAND2_X1 U94 ( .A1(\carry[42] ), .A2(net186622), .ZN(net182693) );
  XNOR2_X1 U95 ( .A(\carry[42] ), .B(net183136), .ZN(SUM[42]) );
  OAI21_X1 U96 ( .B1(n184), .B2(n371), .A(B[41]), .ZN(n183) );
  INV_X1 U97 ( .A(n371), .ZN(n367) );
  NAND2_X1 U98 ( .A1(n374), .A2(n376), .ZN(n184) );
  OR2_X1 U99 ( .A1(n373), .A2(n344), .ZN(n376) );
  OR2_X1 U100 ( .A1(n373), .A2(n344), .ZN(net194454) );
  INV_X1 U101 ( .A(n197), .ZN(n368) );
  OR2_X1 U102 ( .A1(n369), .A2(n368), .ZN(n377) );
  NOR2_X1 U103 ( .A1(n369), .A2(n368), .ZN(n373) );
  NOR2_X1 U104 ( .A1(n369), .A2(n368), .ZN(n193) );
  OAI21_X1 U105 ( .B1(n370), .B2(n375), .A(B[39]), .ZN(n197) );
  BUF_X1 U106 ( .A(A[39]), .Z(n375) );
  AND2_X1 U107 ( .A1(n375), .A2(net197603), .ZN(n369) );
  NAND2_X1 U108 ( .A1(n200), .A2(net182805), .ZN(n370) );
  OAI21_X1 U109 ( .B1(net183573), .B2(n372), .A(B[38]), .ZN(n200) );
  INV_X1 U110 ( .A(n366), .ZN(n372) );
  OAI21_X1 U111 ( .B1(n372), .B2(n332), .A(B[38]), .ZN(net197636) );
  INV_X1 U112 ( .A(A[38]), .ZN(n366) );
  OR2_X1 U113 ( .A1(net182959), .A2(n366), .ZN(net182805) );
  XNOR2_X1 U114 ( .A(B[41]), .B(A[41]), .ZN(net182738) );
  XNOR2_X1 U115 ( .A(net194375), .B(A[40]), .ZN(n195) );
  OAI21_X1 U116 ( .B1(n377), .B2(n335), .A(B[40]), .ZN(n194) );
  NAND2_X1 U117 ( .A1(A[44]), .A2(n384), .ZN(n378) );
  NAND2_X1 U118 ( .A1(n187), .A2(B[44]), .ZN(n379) );
  OR2_X1 U119 ( .A1(n381), .A2(A[44]), .ZN(n187) );
  INV_X1 U120 ( .A(n188), .ZN(n381) );
  CLKBUF_X1 U121 ( .A(n381), .Z(n384) );
  AOI21_X1 U122 ( .B1(n387), .B2(B[43]), .A(n380), .ZN(n188) );
  INV_X1 U123 ( .A(n190), .ZN(n380) );
  AOI21_X1 U124 ( .B1(n387), .B2(B[43]), .A(n380), .ZN(net185361) );
  OAI21_X1 U125 ( .B1(A[43]), .B2(B[43]), .A(n386), .ZN(n190) );
  NAND3_X1 U126 ( .A1(net182694), .A2(net182693), .A3(n382), .ZN(n386) );
  BUF_X1 U127 ( .A(n383), .Z(n387) );
  BUF_X1 U128 ( .A(A[43]), .Z(n383) );
  XNOR2_X1 U129 ( .A(net183674), .B(n383), .ZN(SUM[43]) );
  XNOR2_X1 U130 ( .A(n385), .B(A[44]), .ZN(net183647) );
  NAND3_X1 U131 ( .A1(net182693), .A2(net182694), .A3(n382), .ZN(carry[43]) );
  BUF_X1 U132 ( .A(A[42]), .Z(net186622) );
  NAND2_X1 U133 ( .A1(net186622), .A2(B[42]), .ZN(n382) );
  XNOR2_X1 U134 ( .A(A[42]), .B(B[42]), .ZN(net183136) );
  OR2_X1 U135 ( .A1(n469), .A2(n445), .ZN(n388) );
  OR2_X1 U136 ( .A1(n469), .A2(n445), .ZN(n441) );
  XNOR2_X1 U137 ( .A(n397), .B(n395), .ZN(SUM[33]) );
  BUF_X1 U138 ( .A(n214), .Z(n395) );
  AND2_X1 U139 ( .A1(n214), .A2(n396), .ZN(net191673) );
  XNOR2_X1 U140 ( .A(A[33]), .B(B[33]), .ZN(n397) );
  NAND2_X1 U141 ( .A1(n218), .A2(n392), .ZN(n214) );
  OAI21_X1 U142 ( .B1(n214), .B2(A[33]), .A(B[33]), .ZN(n215) );
  OR2_X1 U143 ( .A1(n217), .A2(n389), .ZN(n392) );
  INV_X1 U144 ( .A(A[32]), .ZN(n389) );
  OAI21_X1 U145 ( .B1(n394), .B2(A[32]), .A(B[32]), .ZN(n218) );
  OR2_X1 U146 ( .A1(n391), .A2(net182635), .ZN(n394) );
  INV_X1 U147 ( .A(n221), .ZN(n391) );
  NOR2_X1 U148 ( .A1(net182635), .A2(n391), .ZN(n217) );
  OAI21_X1 U149 ( .B1(n220), .B2(A[31]), .A(B[31]), .ZN(n221) );
  NAND2_X1 U150 ( .A1(n224), .A2(net184977), .ZN(n220) );
  OAI21_X1 U151 ( .B1(n393), .B2(A[30]), .A(B[30]), .ZN(n224) );
  OR2_X1 U152 ( .A1(net182801), .A2(n390), .ZN(n393) );
  OR2_X1 U153 ( .A1(n390), .A2(net182801), .ZN(net201277) );
  NOR2_X1 U154 ( .A1(net201007), .A2(n390), .ZN(n223) );
  OAI21_X1 U155 ( .B1(n399), .B2(A[28]), .A(B[28]), .ZN(n230) );
  NAND2_X1 U156 ( .A1(net184160), .A2(n400), .ZN(n399) );
  OAI21_X1 U157 ( .B1(n398), .B2(n232), .A(B[27]), .ZN(n400) );
  BUF_X1 U158 ( .A(A[27]), .Z(n398) );
  NAND2_X1 U159 ( .A1(net183836), .A2(n398), .ZN(net184160) );
  OAI21_X1 U160 ( .B1(n232), .B2(n398), .A(B[27]), .ZN(n233) );
  XNOR2_X1 U161 ( .A(A[32]), .B(B[32]), .ZN(n401) );
  BUF_X1 U162 ( .A(A[15]), .Z(n443) );
  AND2_X1 U163 ( .A1(n448), .A2(net187757), .ZN(net201007) );
  OR2_X1 U164 ( .A1(n477), .A2(n235), .ZN(n402) );
  AND2_X1 U165 ( .A1(n239), .A2(net184862), .ZN(n403) );
  NAND2_X1 U166 ( .A1(net197636), .A2(net182805), .ZN(net197603) );
  OAI21_X1 U167 ( .B1(n238), .B2(n418), .A(B[25]), .ZN(n404) );
  NAND2_X1 U168 ( .A1(n194), .A2(net194454), .ZN(net186087) );
  AND2_X1 U170 ( .A1(n239), .A2(net184862), .ZN(n235) );
  AND2_X1 U171 ( .A1(n233), .A2(net184160), .ZN(n229) );
  OR2_X1 U172 ( .A1(n473), .A2(A[15]), .ZN(n405) );
  OR2_X1 U173 ( .A1(n473), .A2(A[15]), .ZN(n268) );
  XNOR2_X1 U174 ( .A(A[15]), .B(n406), .ZN(n414) );
  NAND2_X1 U179 ( .A1(n404), .A2(net184862), .ZN(n407) );
  NOR2_X1 U180 ( .A1(net176614), .A2(net191673), .ZN(n442) );
  XNOR2_X1 U181 ( .A(A[24]), .B(n408), .ZN(net182663) );
  XNOR2_X1 U182 ( .A(A[26]), .B(n409), .ZN(n427) );
  NAND2_X1 U183 ( .A1(n411), .A2(net184977), .ZN(n410) );
  OAI21_X1 U184 ( .B1(net201277), .B2(A[30]), .A(B[30]), .ZN(n411) );
  NOR2_X1 U185 ( .A1(n469), .A2(n445), .ZN(n205) );
  XNOR2_X1 U186 ( .A(n439), .B(n414), .ZN(SUM[15]) );
  XNOR2_X1 U187 ( .A(n415), .B(A[16]), .ZN(n267) );
  XNOR2_X1 U188 ( .A(n417), .B(n420), .ZN(SUM[25]) );
  XNOR2_X1 U189 ( .A(A[25]), .B(B[25]), .ZN(n417) );
  NAND2_X1 U190 ( .A1(n421), .A2(net183284), .ZN(n420) );
  NAND2_X1 U191 ( .A1(n420), .A2(n418), .ZN(net184862) );
  OAI21_X1 U192 ( .B1(net183394), .B2(n422), .A(B[24]), .ZN(n421) );
  BUF_X1 U193 ( .A(n419), .Z(n422) );
  OAI21_X1 U194 ( .B1(net183394), .B2(n422), .A(B[24]), .ZN(n242) );
  INV_X1 U195 ( .A(n419), .ZN(net176583) );
  OAI21_X1 U196 ( .B1(n238), .B2(n418), .A(B[25]), .ZN(n239) );
  NAND2_X1 U197 ( .A1(n242), .A2(net183284), .ZN(n238) );
  BUF_X1 U198 ( .A(A[17]), .Z(n435) );
  INV_X1 U199 ( .A(n229), .ZN(n423) );
  OR2_X1 U200 ( .A1(n480), .A2(n259), .ZN(n424) );
  NAND2_X1 U201 ( .A1(n333), .A2(n424), .ZN(n256) );
  XNOR2_X1 U202 ( .A(A[36]), .B(n425), .ZN(n207) );
  AOI21_X1 U203 ( .B1(n428), .B2(n435), .A(n471), .ZN(n426) );
  XNOR2_X1 U204 ( .A(n466), .B(n423), .ZN(SUM[28]) );
  XNOR2_X1 U205 ( .A(n403), .B(n427), .ZN(SUM[26]) );
  CLKBUF_X1 U206 ( .A(n438), .Z(n428) );
  OAI21_X1 U207 ( .B1(n388), .B2(n431), .A(B[36]), .ZN(n429) );
  INV_X1 U208 ( .A(n452), .ZN(n430) );
  XNOR2_X1 U209 ( .A(A[23]), .B(B[23]), .ZN(net183097) );
  INV_X1 U210 ( .A(n478), .ZN(n431) );
  XNOR2_X1 U211 ( .A(A[34]), .B(n432), .ZN(n213) );
  INV_X1 U212 ( .A(n480), .ZN(n433) );
  OAI21_X1 U213 ( .B1(n412), .B2(n478), .A(n429), .ZN(n434) );
  XNOR2_X1 U214 ( .A(A[30]), .B(net185811), .ZN(n449) );
  INV_X1 U215 ( .A(n481), .ZN(n436) );
  NAND2_X1 U216 ( .A1(n437), .A2(n451), .ZN(n438) );
  INV_X1 U217 ( .A(n450), .ZN(n439) );
  CLKBUF_X1 U218 ( .A(A[23]), .Z(net180672) );
  CLKBUF_X1 U219 ( .A(A[13]), .Z(n455) );
  INV_X1 U220 ( .A(n477), .ZN(n440) );
  OR2_X1 U221 ( .A1(n223), .A2(net176585), .ZN(net184977) );
  NOR2_X1 U222 ( .A1(net176604), .A2(net184972), .ZN(n456) );
  OAI21_X1 U223 ( .B1(n407), .B2(n440), .A(B[26]), .ZN(n444) );
  OR2_X1 U224 ( .A1(n442), .A2(n479), .ZN(n446) );
  NAND2_X1 U225 ( .A1(n446), .A2(n212), .ZN(n208) );
  AOI22_X1 U226 ( .A1(n443), .A2(n450), .B1(n268), .B2(B[15]), .ZN(n447) );
  XNOR2_X1 U227 ( .A(carry[43]), .B(B[43]), .ZN(net183674) );
  NAND2_X1 U228 ( .A1(n339), .A2(net182839), .ZN(n448) );
  XNOR2_X1 U229 ( .A(n449), .B(n223), .ZN(SUM[30]) );
  XNOR2_X1 U230 ( .A(net197603), .B(n460), .ZN(SUM[39]) );
  NAND2_X1 U231 ( .A1(n402), .A2(n444), .ZN(net183836) );
  XNOR2_X1 U232 ( .A(net185361), .B(net183647), .ZN(SUM[44]) );
  OR2_X1 U233 ( .A1(net176583), .A2(n456), .ZN(net183284) );
  AOI21_X1 U234 ( .B1(n428), .B2(n435), .A(n471), .ZN(n259) );
  OR2_X1 U235 ( .A1(n481), .A2(n265), .ZN(n451) );
  AOI22_X1 U236 ( .A1(n443), .A2(n450), .B1(n405), .B2(B[15]), .ZN(n265) );
  CLKBUF_X1 U237 ( .A(n475), .Z(n452) );
  XNOR2_X1 U238 ( .A(n453), .B(net183836), .ZN(SUM[27]) );
  XNOR2_X1 U239 ( .A(A[27]), .B(B[27]), .ZN(n453) );
  XNOR2_X1 U240 ( .A(n438), .B(n454), .ZN(SUM[17]) );
  XNOR2_X1 U241 ( .A(A[17]), .B(B[17]), .ZN(n454) );
  NOR2_X1 U242 ( .A1(n468), .A2(n465), .ZN(net182959) );
  XNOR2_X1 U243 ( .A(n193), .B(n195), .ZN(SUM[40]) );
  OR2_X1 U244 ( .A1(net176584), .A2(n229), .ZN(net182839) );
  OR2_X1 U245 ( .A1(n235), .A2(n477), .ZN(n457) );
  NAND2_X1 U246 ( .A1(n457), .A2(n236), .ZN(n232) );
  AND2_X1 U247 ( .A1(n448), .A2(net187757), .ZN(net182801) );
  INV_X1 U248 ( .A(n458), .ZN(n459) );
  XNOR2_X1 U249 ( .A(A[39]), .B(B[39]), .ZN(n460) );
  XNOR2_X1 U250 ( .A(net186087), .B(net182738), .ZN(SUM[41]) );
  XNOR2_X1 U251 ( .A(n329), .B(n461), .ZN(SUM[29]) );
  XNOR2_X1 U252 ( .A(A[29]), .B(B[29]), .ZN(n461) );
  XNOR2_X1 U253 ( .A(n462), .B(n410), .ZN(SUM[31]) );
  XNOR2_X1 U254 ( .A(A[31]), .B(B[31]), .ZN(n462) );
  XNOR2_X1 U255 ( .A(n463), .B(n413), .ZN(SUM[35]) );
  XNOR2_X1 U256 ( .A(A[35]), .B(B[35]), .ZN(n463) );
  XNOR2_X1 U257 ( .A(n434), .B(n464), .ZN(SUM[37]) );
  XNOR2_X1 U258 ( .A(B[37]), .B(A[37]), .ZN(n464) );
  XNOR2_X1 U259 ( .A(n456), .B(net182663), .ZN(SUM[24]) );
  AND2_X1 U260 ( .A1(A[31]), .A2(n410), .ZN(net182635) );
  AND2_X1 U261 ( .A1(n434), .A2(A[37]), .ZN(n465) );
  INV_X1 U262 ( .A(A[34]), .ZN(n479) );
  INV_X1 U263 ( .A(A[18]), .ZN(n480) );
  XNOR2_X1 U264 ( .A(A[28]), .B(B[28]), .ZN(n466) );
  XOR2_X1 U265 ( .A(n459), .B(n467), .Z(SUM[14]) );
  XNOR2_X1 U266 ( .A(A[14]), .B(B[14]), .ZN(n467) );
  INV_X1 U267 ( .A(n277), .ZN(n476) );
  OAI21_X1 U268 ( .B1(A[12]), .B2(B[12]), .A(carry[12]), .ZN(n277) );
  AND2_X1 U269 ( .A1(A[0]), .A2(B[0]), .ZN(n1) );
  XNOR2_X1 U270 ( .A(n205), .B(n207), .ZN(SUM[36]) );
  INV_X1 U271 ( .A(A[26]), .ZN(n477) );
  INV_X1 U272 ( .A(A[30]), .ZN(net176585) );
  XNOR2_X1 U273 ( .A(n259), .B(n261), .ZN(SUM[18]) );
  OAI21_X1 U274 ( .B1(n208), .B2(A[35]), .A(B[35]), .ZN(n209) );
  AOI22_X1 U275 ( .A1(n452), .A2(n455), .B1(n274), .B2(B[13]), .ZN(n272) );
  OR2_X1 U276 ( .A1(n474), .A2(A[14]), .ZN(n271) );
  XNOR2_X1 U277 ( .A(n213), .B(n336), .ZN(SUM[34]) );
  INV_X1 U278 ( .A(n426), .ZN(n470) );
  OAI21_X1 U279 ( .B1(n202), .B2(A[37]), .A(B[37]), .ZN(n203) );
  XNOR2_X1 U280 ( .A(n265), .B(n267), .ZN(SUM[16]) );
  INV_X1 U281 ( .A(n269), .ZN(n473) );
  AOI21_X1 U282 ( .B1(A[12]), .B2(B[12]), .A(n476), .ZN(n275) );
  OAI21_X1 U283 ( .B1(n407), .B2(n440), .A(B[26]), .ZN(n236) );
  OR2_X1 U284 ( .A1(n475), .A2(A[13]), .ZN(n274) );
  INV_X1 U285 ( .A(n203), .ZN(n468) );
  INV_X1 U286 ( .A(A[16]), .ZN(n481) );
  OAI21_X1 U287 ( .B1(n472), .B2(n436), .A(B[16]), .ZN(n266) );
  OAI21_X1 U288 ( .B1(n412), .B2(n478), .A(n206), .ZN(n202) );
  INV_X1 U289 ( .A(A[36]), .ZN(n478) );
  OAI21_X1 U290 ( .B1(n441), .B2(n431), .A(B[36]), .ZN(n206) );
  INV_X1 U291 ( .A(A[28]), .ZN(net176584) );
  XNOR2_X1 U292 ( .A(n430), .B(n276), .ZN(SUM[13]) );
  INV_X1 U293 ( .A(n275), .ZN(n475) );
  INV_X1 U294 ( .A(n209), .ZN(n469) );
  INV_X1 U295 ( .A(n245), .ZN(net176604) );
  INV_X1 U296 ( .A(n272), .ZN(n474) );
  INV_X1 U297 ( .A(n447), .ZN(n472) );
  OAI21_X1 U298 ( .B1(n470), .B2(n433), .A(B[18]), .ZN(n260) );
  OAI21_X1 U299 ( .B1(n330), .B2(n416), .A(B[34]), .ZN(n212) );
  INV_X1 U300 ( .A(n215), .ZN(net176614) );
endmodule


module RCA_NBIT46 ( A, B, Ci, S, Co );
  input [45:0] A;
  input [45:0] B;
  output [45:0] S;
  input Ci;
  output Co;

  assign Co = 1'b0;

  RCA_NBIT46_DW01_add_0 add_95 ( .A(A), .B(B), .CI(1'b0), .SUM(S) );
endmodule


module RCA_NBIT48_DW01_add_0 ( A, B, CI, SUM, CO );
  input [47:0] A;
  input [47:0] B;
  output [47:0] SUM;
  input CI;
  output CO;
  wire   n1, n348, n352, n358, n359, n365, n392, n409, n413, n414, n415, n416,
         net176633, net176634, net176648, net176649, net180698, net180758,
         net182679, net182928, net182927, net182926, net184167, net184414,
         net184470, net185338, net185572, net185671, net185696, net185904,
         net186038, net186732, net186735, net187284, net187879, net184860,
         net190457, net190619, n410, n407, n403, net190341, net187564,
         net191693, net185916, net184075, net176630, n377, n373, net185965,
         net192749, net191647, net186708, net186707, net186706, net185440,
         n386, n382, net197568, net199347, net186737, net185472, net185000,
         net176627, n404, n401, n397, net183444, net183443, net183442,
         \carry[47] , net182215, net188944, net184640, net182753, net180728,
         n344, n343, n342, n341, n337, net183918, net182925, net182923,
         net176666, net176664, n338, n335, n334, n331, n329, n328, n326, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n327, n330, n332, n333, n336,
         n339, n340, n345, n346, n347, n349, n350, n351, n353, n354, n355,
         n356, n357, n360, n361, n362, n363, n364, n366, n367, n368, n369,
         n370, n371, n372, n374, n375, n376, n378, n379, n380, n381, n383,
         n384, n385, n387, n388, n389, n390, n391, n393, n394, n395, n396,
         n398, n399, n400, n402, n405, n406, n408, n411, n412, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462;
  wire   [47:1] carry;

  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U174 ( .A(n429), .B(n414), .Z(SUM[15]) );
  XOR2_X1 U175 ( .A(A[14]), .B(n416), .Z(SUM[14]) );
  XOR2_X1 U176 ( .A(carry[14]), .B(B[14]), .Z(n416) );
  XOR2_X1 U177 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U1 ( .A(net184470), .Z(net197568) );
  BUF_X1 U2 ( .A(n409), .Z(net185671) );
  CLKBUF_X1 U3 ( .A(A[28]), .Z(net184414) );
  OAI21_X1 U4 ( .B1(n380), .B2(n381), .A(B[36]), .ZN(n275) );
  AND2_X1 U5 ( .A1(n357), .A2(n356), .ZN(n276) );
  AND2_X1 U6 ( .A1(n357), .A2(n356), .ZN(n380) );
  AOI21_X1 U7 ( .B1(n319), .B2(n318), .A(B[43]), .ZN(n277) );
  AOI21_X1 U8 ( .B1(net176630), .B2(net184075), .A(n377), .ZN(n373) );
  NAND2_X1 U9 ( .A1(n364), .A2(B[33]), .ZN(n374) );
  NAND2_X1 U10 ( .A1(n327), .A2(n330), .ZN(n320) );
  INV_X1 U11 ( .A(B[20]), .ZN(n330) );
  INV_X1 U12 ( .A(B[25]), .ZN(n412) );
  INV_X1 U13 ( .A(B[29]), .ZN(n437) );
  BUF_X1 U14 ( .A(n343), .Z(net184640) );
  NAND2_X1 U15 ( .A1(n443), .A2(n432), .ZN(n435) );
  INV_X1 U16 ( .A(B[35]), .ZN(n368) );
  INV_X1 U17 ( .A(B[23]), .ZN(net186706) );
  AND2_X1 U18 ( .A1(n376), .A2(n367), .ZN(n278) );
  INV_X1 U19 ( .A(B[26]), .ZN(n399) );
  NOR2_X1 U20 ( .A1(n277), .A2(n316), .ZN(n279) );
  NAND2_X1 U21 ( .A1(n324), .A2(n325), .ZN(n280) );
  XNOR2_X1 U22 ( .A(n281), .B(net184075), .ZN(SUM[27]) );
  XOR2_X1 U23 ( .A(A[27]), .B(B[27]), .Z(n281) );
  CLKBUF_X1 U24 ( .A(A[17]), .Z(n282) );
  BUF_X1 U25 ( .A(n431), .Z(n285) );
  CLKBUF_X1 U26 ( .A(A[21]), .Z(n347) );
  CLKBUF_X1 U27 ( .A(n462), .Z(n283) );
  BUF_X1 U28 ( .A(A[40]), .Z(net183918) );
  AND2_X1 U29 ( .A1(n320), .A2(n321), .ZN(n349) );
  NAND2_X1 U30 ( .A1(net176648), .A2(n323), .ZN(net187879) );
  CLKBUF_X1 U31 ( .A(A[19]), .Z(net186737) );
  AOI21_X1 U32 ( .B1(n290), .B2(n384), .A(B[39]), .ZN(n284) );
  BUF_X1 U33 ( .A(n403), .Z(n396) );
  CLKBUF_X1 U34 ( .A(n382), .Z(n419) );
  AOI21_X1 U35 ( .B1(n291), .B2(n292), .A(n293), .ZN(n286) );
  NOR2_X1 U36 ( .A1(n341), .A2(n385), .ZN(n287) );
  OR2_X1 U37 ( .A1(n343), .A2(A[38]), .ZN(n344) );
  NAND2_X1 U38 ( .A1(net184640), .A2(n387), .ZN(n288) );
  NAND2_X1 U39 ( .A1(n344), .A2(B[38]), .ZN(n289) );
  NAND2_X1 U40 ( .A1(n288), .A2(n289), .ZN(n290) );
  INV_X1 U41 ( .A(B[46]), .ZN(n312) );
  INV_X1 U42 ( .A(B[45]), .ZN(n305) );
  CLKBUF_X1 U43 ( .A(A[38]), .Z(n387) );
  MUX2_X1 U44 ( .A(n309), .B(n313), .S(n302), .Z(SUM[46]) );
  BUF_X1 U45 ( .A(A[27]), .Z(net185916) );
  NOR2_X1 U46 ( .A1(n329), .A2(n316), .ZN(n326) );
  AOI21_X1 U47 ( .B1(n291), .B2(n292), .A(n293), .ZN(net176666) );
  INV_X1 U48 ( .A(n331), .ZN(n291) );
  INV_X1 U49 ( .A(A[42]), .ZN(n292) );
  INV_X1 U50 ( .A(B[42]), .ZN(n293) );
  AOI21_X1 U51 ( .B1(n317), .B2(A[41]), .A(B[41]), .ZN(n335) );
  OAI21_X1 U52 ( .B1(net176627), .B2(n398), .A(n401), .ZN(n397) );
  AOI21_X1 U53 ( .B1(n294), .B2(n295), .A(n415), .ZN(n460) );
  INV_X1 U54 ( .A(B[14]), .ZN(n294) );
  INV_X1 U55 ( .A(A[14]), .ZN(n295) );
  XNOR2_X1 U56 ( .A(n336), .B(n397), .ZN(SUM[20]) );
  XNOR2_X1 U57 ( .A(net188944), .B(n342), .ZN(SUM[39]) );
  AND2_X1 U58 ( .A1(n304), .A2(n303), .ZN(n296) );
  NAND2_X1 U59 ( .A1(n305), .A2(n298), .ZN(n303) );
  NOR2_X1 U60 ( .A1(n359), .A2(n389), .ZN(n297) );
  AND2_X1 U61 ( .A1(n301), .A2(n300), .ZN(n298) );
  OAI21_X1 U62 ( .B1(B[44]), .B2(A[44]), .A(n326), .ZN(n301) );
  XNOR2_X1 U63 ( .A(n279), .B(n308), .ZN(SUM[44]) );
  XNOR2_X1 U64 ( .A(A[46]), .B(B[46]), .ZN(n309) );
  NAND2_X1 U65 ( .A1(n296), .A2(n311), .ZN(net183442) );
  NAND2_X1 U66 ( .A1(n311), .A2(B[46]), .ZN(net183444) );
  INV_X1 U67 ( .A(A[45]), .ZN(n307) );
  NAND2_X1 U68 ( .A1(n310), .A2(n307), .ZN(n304) );
  XNOR2_X1 U69 ( .A(n306), .B(n307), .ZN(SUM[45]) );
  CLKBUF_X1 U70 ( .A(A[46]), .Z(n311) );
  NAND2_X1 U71 ( .A1(n301), .A2(n300), .ZN(n299) );
  XNOR2_X1 U72 ( .A(n299), .B(n305), .ZN(n306) );
  NAND2_X1 U73 ( .A1(n299), .A2(B[45]), .ZN(n310) );
  XNOR2_X1 U74 ( .A(A[46]), .B(n312), .ZN(n313) );
  NAND2_X1 U75 ( .A1(n303), .A2(n304), .ZN(n302) );
  XNOR2_X1 U76 ( .A(B[44]), .B(A[44]), .ZN(n308) );
  NAND2_X1 U77 ( .A1(B[44]), .A2(A[44]), .ZN(n300) );
  NAND2_X1 U78 ( .A1(B[46]), .A2(n296), .ZN(net183443) );
  AND2_X1 U79 ( .A1(n315), .A2(n328), .ZN(n316) );
  NOR2_X1 U80 ( .A1(net182923), .A2(n286), .ZN(n328) );
  OR2_X1 U81 ( .A1(n286), .A2(net182923), .ZN(n319) );
  OR2_X1 U82 ( .A1(net176666), .A2(net182923), .ZN(net191693) );
  INV_X1 U83 ( .A(A[43]), .ZN(n315) );
  INV_X1 U84 ( .A(n315), .ZN(n318) );
  AOI21_X1 U85 ( .B1(n319), .B2(n318), .A(B[43]), .ZN(n329) );
  AND2_X1 U86 ( .A1(n331), .A2(A[42]), .ZN(net182923) );
  AOI21_X1 U87 ( .B1(n314), .B2(n334), .A(n335), .ZN(n331) );
  INV_X1 U88 ( .A(A[41]), .ZN(n314) );
  OR2_X1 U89 ( .A1(net176664), .A2(net182925), .ZN(n317) );
  INV_X1 U90 ( .A(n338), .ZN(net176664) );
  OR2_X1 U91 ( .A1(net176664), .A2(net182925), .ZN(net185965) );
  OAI21_X1 U92 ( .B1(n337), .B2(net183918), .A(B[40]), .ZN(n338) );
  AND2_X1 U93 ( .A1(n287), .A2(net183918), .ZN(net182925) );
  INV_X1 U94 ( .A(net185965), .ZN(n334) );
  XNOR2_X1 U95 ( .A(A[42]), .B(B[42]), .ZN(net185338) );
  XNOR2_X1 U96 ( .A(A[43]), .B(B[43]), .ZN(net185696) );
  XNOR2_X1 U97 ( .A(A[41]), .B(B[41]), .ZN(net180698) );
  XNOR2_X1 U98 ( .A(net182215), .B(n287), .ZN(SUM[40]) );
  NAND2_X1 U99 ( .A1(n345), .A2(n332), .ZN(n323) );
  INV_X1 U100 ( .A(n397), .ZN(n339) );
  XNOR2_X1 U101 ( .A(A[20]), .B(B[20]), .ZN(n336) );
  NAND2_X1 U102 ( .A1(A[20]), .A2(B[20]), .ZN(n340) );
  INV_X1 U103 ( .A(A[20]), .ZN(n327) );
  XNOR2_X1 U104 ( .A(n322), .B(B[22]), .ZN(n333) );
  XNOR2_X1 U105 ( .A(n333), .B(n351), .ZN(SUM[22]) );
  XNOR2_X1 U106 ( .A(A[21]), .B(B[21]), .ZN(n346) );
  OAI21_X1 U107 ( .B1(n350), .B2(B[21]), .A(n347), .ZN(n325) );
  NAND2_X1 U108 ( .A1(n324), .A2(n325), .ZN(n322) );
  INV_X1 U109 ( .A(n280), .ZN(n345) );
  AOI21_X1 U110 ( .B1(n280), .B2(A[22]), .A(B[22]), .ZN(n392) );
  XNOR2_X1 U111 ( .A(n346), .B(n349), .ZN(SUM[21]) );
  AND2_X1 U112 ( .A1(n320), .A2(n321), .ZN(n350) );
  INV_X1 U113 ( .A(A[22]), .ZN(n332) );
  INV_X1 U114 ( .A(n332), .ZN(n351) );
  NAND2_X1 U115 ( .A1(B[21]), .A2(n349), .ZN(n324) );
  NAND2_X1 U116 ( .A1(n339), .A2(n340), .ZN(n321) );
  OAI21_X1 U117 ( .B1(A[32]), .B2(n379), .A(B[32]), .ZN(n354) );
  BUF_X1 U118 ( .A(net199347), .Z(n379) );
  NAND2_X1 U119 ( .A1(n354), .A2(n353), .ZN(net187284) );
  INV_X1 U120 ( .A(net182926), .ZN(n353) );
  AND2_X1 U121 ( .A1(n354), .A2(n353), .ZN(n358) );
  INV_X1 U122 ( .A(A[34]), .ZN(n366) );
  OAI21_X1 U123 ( .B1(n380), .B2(n381), .A(B[36]), .ZN(n363) );
  NAND2_X1 U124 ( .A1(n275), .A2(n362), .ZN(n361) );
  NAND2_X1 U125 ( .A1(n352), .A2(net176634), .ZN(n356) );
  NAND2_X1 U126 ( .A1(n361), .A2(A[37]), .ZN(n372) );
  OAI21_X1 U127 ( .B1(n278), .B2(net176634), .A(n368), .ZN(n357) );
  OAI211_X1 U128 ( .C1(n358), .C2(n355), .A(n366), .B(n374), .ZN(n375) );
  NAND2_X1 U129 ( .A1(n375), .A2(B[34]), .ZN(n376) );
  NAND2_X1 U130 ( .A1(n276), .A2(n381), .ZN(n362) );
  NAND2_X1 U131 ( .A1(n372), .A2(n369), .ZN(n371) );
  INV_X1 U132 ( .A(net184470), .ZN(n367) );
  INV_X1 U133 ( .A(A[37]), .ZN(n360) );
  NAND2_X1 U134 ( .A1(net186038), .A2(n360), .ZN(n370) );
  AND2_X1 U135 ( .A1(n375), .A2(B[34]), .ZN(net185904) );
  INV_X1 U136 ( .A(B[37]), .ZN(n369) );
  XNOR2_X1 U137 ( .A(A[37]), .B(n369), .ZN(n348) );
  NOR2_X1 U138 ( .A1(n364), .A2(B[33]), .ZN(n355) );
  XNOR2_X1 U139 ( .A(A[36]), .B(B[36]), .ZN(n378) );
  INV_X1 U140 ( .A(net176633), .ZN(n364) );
  AND2_X1 U141 ( .A1(n363), .A2(n362), .ZN(net186038) );
  AND2_X1 U142 ( .A1(n371), .A2(n370), .ZN(n343) );
  CLKBUF_X1 U143 ( .A(A[36]), .Z(n381) );
  XNOR2_X1 U144 ( .A(n276), .B(n378), .ZN(SUM[36]) );
  NOR2_X1 U145 ( .A1(n385), .A2(n284), .ZN(n337) );
  AND2_X1 U146 ( .A1(n383), .A2(net188944), .ZN(n385) );
  INV_X1 U147 ( .A(A[39]), .ZN(n383) );
  INV_X1 U148 ( .A(n383), .ZN(n384) );
  AOI21_X1 U149 ( .B1(n290), .B2(n384), .A(B[39]), .ZN(n341) );
  AOI22_X1 U150 ( .A1(net184640), .A2(n387), .B1(n344), .B2(B[38]), .ZN(
        net188944) );
  XNOR2_X1 U151 ( .A(net184640), .B(net182753), .ZN(SUM[38]) );
  XNOR2_X1 U152 ( .A(A[39]), .B(net180728), .ZN(n342) );
  INV_X1 U153 ( .A(B[39]), .ZN(net180728) );
  XNOR2_X1 U154 ( .A(A[38]), .B(B[38]), .ZN(net182753) );
  XNOR2_X1 U155 ( .A(A[40]), .B(B[40]), .ZN(net182215) );
  XNOR2_X1 U156 ( .A(n388), .B(A[47]), .ZN(SUM[47]) );
  XNOR2_X1 U157 ( .A(\carry[47] ), .B(B[47]), .ZN(n388) );
  NAND3_X1 U158 ( .A1(net183442), .A2(net183443), .A3(net183444), .ZN(
        \carry[47] ) );
  AND2_X1 U159 ( .A1(n358), .A2(net176633), .ZN(n389) );
  CLKBUF_X1 U160 ( .A(A[23]), .Z(net185440) );
  OAI21_X1 U161 ( .B1(net185000), .B2(A[19]), .A(B[19]), .ZN(n401) );
  INV_X1 U162 ( .A(net185472), .ZN(net185000) );
  OAI21_X1 U163 ( .B1(n394), .B2(n396), .A(n390), .ZN(net185472) );
  INV_X1 U164 ( .A(n404), .ZN(n390) );
  OAI21_X1 U165 ( .B1(n394), .B2(n396), .A(n390), .ZN(n398) );
  AOI21_X1 U166 ( .B1(A[18]), .B2(n403), .A(B[18]), .ZN(n404) );
  XNOR2_X1 U167 ( .A(n395), .B(n396), .ZN(SUM[18]) );
  CLKBUF_X1 U168 ( .A(A[18]), .Z(n394) );
  INV_X1 U169 ( .A(net186737), .ZN(net176627) );
  INV_X1 U170 ( .A(n398), .ZN(n391) );
  XNOR2_X1 U171 ( .A(n393), .B(n391), .ZN(SUM[19]) );
  XNOR2_X1 U172 ( .A(A[19]), .B(B[19]), .ZN(n393) );
  XNOR2_X1 U173 ( .A(A[18]), .B(B[18]), .ZN(n395) );
  AOI21_X1 U178 ( .B1(n461), .B2(net182928), .A(n365), .ZN(net199347) );
  XNOR2_X1 U179 ( .A(A[26]), .B(n399), .ZN(n422) );
  XNOR2_X1 U180 ( .A(n411), .B(n419), .ZN(SUM[25]) );
  OR2_X1 U181 ( .A1(n382), .A2(B[25]), .ZN(n420) );
  OR2_X1 U182 ( .A1(n382), .A2(A[25]), .ZN(n421) );
  AND2_X1 U183 ( .A1(n421), .A2(n420), .ZN(n402) );
  NAND2_X1 U184 ( .A1(n402), .A2(n405), .ZN(n400) );
  NAND2_X1 U185 ( .A1(n425), .A2(n399), .ZN(n406) );
  OAI21_X1 U186 ( .B1(n399), .B2(n425), .A(n418), .ZN(n408) );
  INV_X1 U187 ( .A(n424), .ZN(n418) );
  NAND2_X1 U188 ( .A1(n406), .A2(n408), .ZN(net184075) );
  XNOR2_X1 U189 ( .A(A[25]), .B(B[25]), .ZN(n411) );
  INV_X1 U190 ( .A(A[25]), .ZN(n417) );
  AOI21_X1 U191 ( .B1(net185916), .B2(n423), .A(B[27]), .ZN(n377) );
  XNOR2_X1 U192 ( .A(n422), .B(n400), .ZN(SUM[26]) );
  AND2_X1 U193 ( .A1(n406), .A2(n408), .ZN(n423) );
  CLKBUF_X1 U194 ( .A(A[26]), .Z(n424) );
  NAND2_X1 U195 ( .A1(n417), .A2(n412), .ZN(n405) );
  NAND2_X1 U196 ( .A1(n402), .A2(n405), .ZN(n425) );
  AND2_X1 U197 ( .A1(n441), .A2(n440), .ZN(n426) );
  NAND2_X1 U198 ( .A1(net190457), .A2(n282), .ZN(n448) );
  NAND2_X1 U199 ( .A1(n444), .A2(n435), .ZN(n427) );
  INV_X1 U200 ( .A(net182928), .ZN(n428) );
  INV_X1 U201 ( .A(n453), .ZN(n429) );
  XNOR2_X1 U202 ( .A(n427), .B(n445), .ZN(SUM[30]) );
  OAI21_X1 U203 ( .B1(net187564), .B2(net182927), .A(n386), .ZN(n382) );
  OAI21_X1 U204 ( .B1(net190341), .B2(n430), .A(B[24]), .ZN(n386) );
  OAI22_X1 U205 ( .A1(net186735), .A2(net186707), .B1(net191647), .B2(
        net186706), .ZN(n430) );
  OAI22_X1 U206 ( .A1(net186735), .A2(net186707), .B1(net186708), .B2(
        net186706), .ZN(net192749) );
  OAI22_X1 U207 ( .A1(net186735), .A2(net186707), .B1(net186708), .B2(
        net186706), .ZN(net190619) );
  NOR2_X1 U208 ( .A1(net176649), .A2(net185440), .ZN(net191647) );
  INV_X1 U209 ( .A(net185440), .ZN(net186707) );
  NOR2_X1 U210 ( .A1(net176649), .A2(net185440), .ZN(net186708) );
  NAND2_X1 U211 ( .A1(n438), .A2(n437), .ZN(n436) );
  NAND2_X1 U212 ( .A1(n436), .A2(n435), .ZN(n434) );
  NAND2_X1 U213 ( .A1(n435), .A2(n444), .ZN(n442) );
  NAND2_X1 U214 ( .A1(n442), .A2(n433), .ZN(n441) );
  OAI21_X1 U215 ( .B1(n433), .B2(n434), .A(n439), .ZN(n440) );
  NAND2_X1 U216 ( .A1(net185572), .A2(net184167), .ZN(n431) );
  INV_X1 U217 ( .A(A[30]), .ZN(n439) );
  NAND2_X1 U218 ( .A1(n431), .A2(A[29]), .ZN(n438) );
  XNOR2_X1 U219 ( .A(A[29]), .B(B[29]), .ZN(net180758) );
  INV_X1 U220 ( .A(A[29]), .ZN(n432) );
  AND2_X1 U221 ( .A1(net185572), .A2(net184167), .ZN(n443) );
  NAND2_X1 U222 ( .A1(n438), .A2(n437), .ZN(n444) );
  INV_X1 U223 ( .A(B[30]), .ZN(n433) );
  XNOR2_X1 U224 ( .A(A[30]), .B(n433), .ZN(n445) );
  XNOR2_X1 U225 ( .A(n331), .B(net185338), .ZN(SUM[42]) );
  NAND2_X1 U226 ( .A1(n373), .A2(net184414), .ZN(net184167) );
  OAI21_X1 U227 ( .B1(net184414), .B2(n373), .A(B[28]), .ZN(net185572) );
  XNOR2_X1 U228 ( .A(n373), .B(net182679), .ZN(SUM[28]) );
  INV_X1 U229 ( .A(net185916), .ZN(net176630) );
  BUF_X1 U230 ( .A(A[24]), .Z(net190341) );
  INV_X1 U231 ( .A(net190341), .ZN(net187564) );
  OR2_X1 U232 ( .A1(net197568), .A2(net185904), .ZN(n446) );
  XNOR2_X1 U233 ( .A(A[28]), .B(B[28]), .ZN(net182679) );
  NAND2_X1 U234 ( .A1(n407), .A2(n448), .ZN(n403) );
  INV_X1 U235 ( .A(n410), .ZN(n447) );
  AND2_X1 U236 ( .A1(n447), .A2(n449), .ZN(net190457) );
  AND2_X1 U237 ( .A1(n447), .A2(n449), .ZN(n450) );
  AOI21_X1 U238 ( .B1(n409), .B2(A[16]), .A(B[16]), .ZN(n410) );
  OAI21_X1 U239 ( .B1(n450), .B2(A[17]), .A(B[17]), .ZN(n407) );
  XNOR2_X1 U240 ( .A(A[17]), .B(B[17]), .ZN(net184860) );
  OR2_X1 U241 ( .A1(n409), .A2(A[16]), .ZN(n449) );
  XNOR2_X1 U242 ( .A(A[16]), .B(B[16]), .ZN(net186732) );
  NOR2_X1 U243 ( .A1(n389), .A2(n359), .ZN(n451) );
  XNOR2_X1 U244 ( .A(net184860), .B(net190457), .ZN(SUM[17]) );
  CLKBUF_X1 U245 ( .A(net187879), .Z(net186735) );
  XNOR2_X1 U246 ( .A(net186732), .B(net185671), .ZN(SUM[16]) );
  XNOR2_X1 U247 ( .A(n452), .B(n297), .ZN(SUM[34]) );
  XNOR2_X1 U248 ( .A(A[34]), .B(B[34]), .ZN(n452) );
  INV_X1 U249 ( .A(n460), .ZN(n453) );
  XNOR2_X1 U250 ( .A(net185696), .B(net191693), .ZN(SUM[43]) );
  AND2_X1 U251 ( .A1(A[34]), .A2(n451), .ZN(net184470) );
  NOR2_X1 U252 ( .A1(net185904), .A2(net197568), .ZN(n352) );
  XNOR2_X1 U253 ( .A(net186038), .B(n348), .ZN(SUM[37]) );
  XNOR2_X1 U254 ( .A(A[24]), .B(B[24]), .ZN(n455) );
  XNOR2_X1 U255 ( .A(A[32]), .B(B[32]), .ZN(n454) );
  XNOR2_X1 U256 ( .A(n379), .B(n454), .ZN(SUM[32]) );
  XNOR2_X1 U257 ( .A(n428), .B(n457), .ZN(SUM[31]) );
  XNOR2_X1 U258 ( .A(n456), .B(n446), .ZN(SUM[35]) );
  XNOR2_X1 U259 ( .A(n455), .B(net192749), .ZN(SUM[24]) );
  AND2_X1 U260 ( .A1(net199347), .A2(A[32]), .ZN(net182926) );
  INV_X1 U261 ( .A(net190619), .ZN(net182927) );
  INV_X1 U262 ( .A(n426), .ZN(net182928) );
  INV_X1 U263 ( .A(A[15]), .ZN(n462) );
  XNOR2_X1 U264 ( .A(A[35]), .B(B[35]), .ZN(n456) );
  XNOR2_X1 U265 ( .A(A[31]), .B(B[31]), .ZN(n457) );
  XNOR2_X1 U266 ( .A(A[33]), .B(B[33]), .ZN(n459) );
  INV_X1 U267 ( .A(net187879), .ZN(net176649) );
  XNOR2_X1 U268 ( .A(n458), .B(net176649), .ZN(SUM[23]) );
  XNOR2_X1 U269 ( .A(A[23]), .B(B[23]), .ZN(n458) );
  OAI21_X1 U270 ( .B1(n462), .B2(n453), .A(n413), .ZN(n409) );
  OAI21_X1 U271 ( .B1(A[15]), .B2(n460), .A(B[15]), .ZN(n413) );
  AOI21_X1 U272 ( .B1(A[14]), .B2(B[14]), .A(carry[14]), .ZN(n415) );
  XNOR2_X1 U273 ( .A(B[15]), .B(n283), .ZN(n414) );
  AND2_X1 U274 ( .A1(A[0]), .A2(B[0]), .ZN(n1) );
  XNOR2_X1 U275 ( .A(n285), .B(net180758), .ZN(SUM[29]) );
  XNOR2_X1 U276 ( .A(n459), .B(net187284), .ZN(SUM[33]) );
  XNOR2_X1 U277 ( .A(net180698), .B(net185965), .ZN(SUM[41]) );
  INV_X1 U278 ( .A(A[31]), .ZN(n461) );
  AOI21_X1 U279 ( .B1(n426), .B2(A[31]), .A(B[31]), .ZN(n365) );
  AOI21_X1 U280 ( .B1(A[33]), .B2(net187284), .A(B[33]), .ZN(n359) );
  INV_X1 U281 ( .A(A[33]), .ZN(net176633) );
  INV_X1 U282 ( .A(A[35]), .ZN(net176634) );
  INV_X1 U283 ( .A(n392), .ZN(net176648) );
endmodule


module RCA_NBIT48 ( A, B, Ci, S, Co );
  input [47:0] A;
  input [47:0] B;
  output [47:0] S;
  input Ci;
  output Co;

  assign Co = 1'b0;

  RCA_NBIT48_DW01_add_0 add_95 ( .A(A), .B(B), .CI(1'b0), .SUM(S) );
endmodule


module RCA_NBIT50_DW01_add_0 ( A, B, CI, SUM, CO );
  input [49:0] A;
  input [49:0] B;
  output [49:0] SUM;
  input CI;
  output CO;
  wire   n1, \carry[44] , \carry[16] , \carry[43] , \carry[42] , net76696,
         n304, n306, n307, n308, n309, n310, n311, n331, n334, n338, n360,
         n364, n367, n378, n381, n382, n384, n386, n387, n388, n389, n390,
         n391, net176691, net176705, net176708, net180780, net182414,
         net182425, net182464, net182465, net182656, net182664, net182676,
         net182726, net183202, net183664, net184159, net184620, net185094,
         net185161, net185264, net185453, net185452, net185898, net185908,
         net187723, net180768, net184622, net190661, net190992, net183946,
         net182434, net176675, net176674, n355, n351, net197646, n352, n349,
         n346, n345, n343, net183591, n312, n379, n376, n375, n373, n372, n370,
         n369, n366, net193269, net187480, net184093, net183901, net182455,
         n361, n318, n315, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n305, n313,
         n314, n316, n317, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n332, n333, n335, n336, n337, n339, n340,
         n341, n342, n344, n347, n348, n350, n353, n354, n356, n357, n358,
         n359, n362, n363, n365, n368, n371, n374, n377, n380, n383, n385,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425;
  wire   [49:1] carry;

  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(\carry[16] ), .S(
        SUM[15]) );
  FA_X1 U1_44 ( .A(A[44]), .B(B[44]), .CI(\carry[44] ), .CO(net76696), .S(
        SUM[44]) );
  FA_X1 U1_41 ( .A(B[41]), .B(A[41]), .CI(n419), .CO(\carry[42] ), .S(SUM[41])
         );
  FA_X1 U1_43 ( .A(A[43]), .B(B[43]), .CI(\carry[43] ), .CO(\carry[44] ), .S(
        SUM[43]) );
  FA_X1 U1_42 ( .A(A[42]), .B(B[42]), .CI(\carry[42] ), .CO(\carry[43] ), .S(
        SUM[42]) );
  XOR2_X1 U101 ( .A(B[49]), .B(A[49]), .Z(n308) );
  XOR2_X1 U102 ( .A(net176708), .B(n310), .Z(SUM[48]) );
  XOR2_X1 U155 ( .A(n413), .B(n389), .Z(SUM[17]) );
  XOR2_X1 U156 ( .A(B[17]), .B(n399), .Z(n389) );
  XOR2_X1 U157 ( .A(n402), .B(n391), .Z(SUM[16]) );
  XOR2_X1 U158 ( .A(\carry[16] ), .B(B[16]), .Z(n391) );
  XOR2_X1 U159 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  CLKBUF_X1 U1 ( .A(A[24]), .Z(net180780) );
  BUF_X1 U2 ( .A(n351), .Z(n357) );
  AND2_X1 U3 ( .A1(n341), .A2(n342), .ZN(n265) );
  NAND2_X1 U4 ( .A1(n345), .A2(n268), .ZN(n266) );
  AND2_X1 U5 ( .A1(n348), .A2(n342), .ZN(n267) );
  CLKBUF_X1 U6 ( .A(A[28]), .Z(n300) );
  BUF_X1 U7 ( .A(A[31]), .Z(n268) );
  AOI21_X1 U8 ( .B1(net176675), .B2(n356), .A(n349), .ZN(n269) );
  AOI21_X1 U9 ( .B1(net176675), .B2(n356), .A(n349), .ZN(n345) );
  CLKBUF_X1 U10 ( .A(A[26]), .Z(n270) );
  AOI21_X1 U11 ( .B1(n406), .B2(n408), .A(B[36]), .ZN(n271) );
  CLKBUF_X1 U12 ( .A(n323), .Z(n272) );
  CLKBUF_X1 U13 ( .A(A[29]), .Z(n358) );
  AND2_X1 U14 ( .A1(n398), .A2(A[18]), .ZN(n273) );
  OAI22_X1 U15 ( .A1(n395), .A2(n413), .B1(B[17]), .B2(n388), .ZN(n274) );
  BUF_X1 U16 ( .A(A[25]), .Z(n332) );
  CLKBUF_X1 U17 ( .A(A[21]), .Z(n275) );
  CLKBUF_X1 U18 ( .A(A[23]), .Z(n322) );
  CLKBUF_X1 U19 ( .A(A[45]), .Z(net197646) );
  INV_X1 U20 ( .A(B[48]), .ZN(n401) );
  NAND2_X1 U21 ( .A1(n265), .A2(net187723), .ZN(net184159) );
  INV_X1 U22 ( .A(B[46]), .ZN(n278) );
  NAND2_X1 U23 ( .A1(n278), .A2(n280), .ZN(n276) );
  AND2_X1 U24 ( .A1(n276), .A2(n277), .ZN(n279) );
  NAND2_X1 U25 ( .A1(A[46]), .A2(n292), .ZN(n280) );
  OR2_X1 U26 ( .A1(n315), .A2(A[46]), .ZN(n277) );
  INV_X1 U27 ( .A(n298), .ZN(n281) );
  INV_X1 U28 ( .A(net187480), .ZN(n282) );
  NAND2_X1 U29 ( .A1(n284), .A2(n285), .ZN(n283) );
  OR2_X1 U30 ( .A1(n281), .A2(n282), .ZN(n284) );
  NAND2_X1 U31 ( .A1(net193269), .A2(B[27]), .ZN(n285) );
  XNOR2_X1 U32 ( .A(B[31]), .B(A[31]), .ZN(net182414) );
  NAND2_X1 U33 ( .A1(n298), .A2(net187480), .ZN(n286) );
  NAND2_X1 U34 ( .A1(n299), .A2(B[27]), .ZN(n287) );
  NAND2_X1 U35 ( .A1(n286), .A2(n287), .ZN(n288) );
  XNOR2_X1 U36 ( .A(n291), .B(n315), .ZN(SUM[46]) );
  XNOR2_X1 U37 ( .A(A[46]), .B(B[46]), .ZN(n291) );
  AOI21_X1 U38 ( .B1(n289), .B2(n290), .A(n318), .ZN(n315) );
  INV_X1 U39 ( .A(A[45]), .ZN(n290) );
  AOI21_X1 U40 ( .B1(n289), .B2(n290), .A(n318), .ZN(n292) );
  INV_X1 U41 ( .A(B[45]), .ZN(n289) );
  AOI21_X1 U42 ( .B1(A[45]), .B2(B[45]), .A(net76696), .ZN(n318) );
  XNOR2_X1 U43 ( .A(net76696), .B(B[45]), .ZN(net182425) );
  NAND2_X1 U44 ( .A1(n365), .A2(n368), .ZN(n293) );
  NAND2_X1 U45 ( .A1(n335), .A2(n333), .ZN(n294) );
  NOR2_X1 U46 ( .A1(n271), .A2(n409), .ZN(n295) );
  BUF_X1 U47 ( .A(n393), .Z(net184620) );
  XNOR2_X1 U48 ( .A(net182455), .B(n283), .ZN(SUM[28]) );
  XNOR2_X1 U49 ( .A(A[28]), .B(B[28]), .ZN(net182455) );
  CLKBUF_X1 U50 ( .A(A[27]), .Z(n298) );
  AOI22_X1 U51 ( .A1(net187480), .A2(n298), .B1(net193269), .B2(B[27]), .ZN(
        net184622) );
  INV_X1 U52 ( .A(A[28]), .ZN(net176674) );
  AOI21_X1 U53 ( .B1(n288), .B2(n300), .A(B[28]), .ZN(n355) );
  AND2_X1 U54 ( .A1(n296), .A2(n297), .ZN(net187480) );
  XNOR2_X1 U55 ( .A(net183901), .B(net187480), .ZN(SUM[27]) );
  INV_X1 U56 ( .A(n361), .ZN(n296) );
  AND2_X1 U57 ( .A1(n296), .A2(n297), .ZN(net184093) );
  AOI21_X1 U58 ( .B1(n360), .B2(A[26]), .A(B[26]), .ZN(n361) );
  OR2_X1 U59 ( .A1(net184093), .A2(A[27]), .ZN(net193269) );
  OR2_X1 U60 ( .A1(net184093), .A2(A[27]), .ZN(n299) );
  XNOR2_X1 U61 ( .A(A[27]), .B(B[27]), .ZN(net183901) );
  OR2_X1 U62 ( .A1(n360), .A2(n270), .ZN(n297) );
  BUF_X1 U63 ( .A(n360), .Z(net190992) );
  XNOR2_X1 U64 ( .A(A[26]), .B(B[26]), .ZN(net180768) );
  OAI21_X1 U65 ( .B1(n272), .B2(n320), .A(n370), .ZN(n366) );
  OR2_X1 U66 ( .A1(net180780), .A2(n366), .ZN(net183664) );
  XNOR2_X1 U67 ( .A(n366), .B(net182664), .ZN(SUM[24]) );
  AOI21_X1 U68 ( .B1(n366), .B2(net180780), .A(B[24]), .ZN(n367) );
  OAI21_X1 U69 ( .B1(n321), .B2(n322), .A(B[23]), .ZN(n370) );
  INV_X1 U70 ( .A(n322), .ZN(n320) );
  INV_X1 U71 ( .A(n369), .ZN(n321) );
  OAI21_X1 U72 ( .B1(n317), .B2(n316), .A(n305), .ZN(n369) );
  INV_X1 U73 ( .A(n373), .ZN(n305) );
  OAI21_X1 U74 ( .B1(n317), .B2(n316), .A(n305), .ZN(n323) );
  AOI21_X1 U75 ( .B1(n372), .B2(A[22]), .A(B[22]), .ZN(n373) );
  CLKBUF_X1 U76 ( .A(A[22]), .Z(n316) );
  CLKBUF_X1 U77 ( .A(n372), .Z(n317) );
  XNOR2_X1 U78 ( .A(n317), .B(net182726), .ZN(SUM[22]) );
  INV_X1 U79 ( .A(n323), .ZN(n313) );
  XNOR2_X1 U80 ( .A(n313), .B(n314), .ZN(SUM[23]) );
  XNOR2_X1 U81 ( .A(A[23]), .B(B[23]), .ZN(n314) );
  OAI21_X1 U82 ( .B1(net185264), .B2(n301), .A(n376), .ZN(n372) );
  OAI21_X1 U83 ( .B1(n303), .B2(n275), .A(B[21]), .ZN(n376) );
  INV_X1 U84 ( .A(A[21]), .ZN(n301) );
  INV_X1 U85 ( .A(n375), .ZN(n303) );
  OAI21_X1 U86 ( .B1(net185094), .B2(n319), .A(n302), .ZN(n375) );
  INV_X1 U87 ( .A(n379), .ZN(n302) );
  OAI21_X1 U88 ( .B1(net185094), .B2(n319), .A(n302), .ZN(net185898) );
  AOI21_X1 U89 ( .B1(n378), .B2(A[20]), .A(B[20]), .ZN(n379) );
  CLKBUF_X1 U90 ( .A(A[20]), .Z(n319) );
  XNOR2_X1 U91 ( .A(n324), .B(net183591), .ZN(SUM[47]) );
  BUF_X1 U92 ( .A(n279), .Z(net183591) );
  OAI22_X1 U93 ( .A1(n325), .A2(net183591), .B1(n312), .B2(B[47]), .ZN(n311)
         );
  AND2_X1 U94 ( .A1(A[47]), .A2(n279), .ZN(n312) );
  XNOR2_X1 U95 ( .A(A[47]), .B(B[47]), .ZN(n324) );
  CLKBUF_X1 U96 ( .A(A[47]), .Z(n325) );
  NAND2_X1 U97 ( .A1(n329), .A2(n339), .ZN(n326) );
  NAND2_X1 U98 ( .A1(n327), .A2(n328), .ZN(n329) );
  NAND2_X1 U99 ( .A1(n329), .A2(n339), .ZN(n337) );
  INV_X1 U100 ( .A(A[32]), .ZN(n327) );
  INV_X1 U103 ( .A(net185161), .ZN(n328) );
  OAI22_X1 U104 ( .A1(n411), .A2(n421), .B1(B[18]), .B2(n273), .ZN(n330) );
  NAND2_X1 U105 ( .A1(n337), .A2(n336), .ZN(n333) );
  OAI21_X1 U106 ( .B1(n336), .B2(n337), .A(n344), .ZN(n335) );
  INV_X1 U107 ( .A(n343), .ZN(n339) );
  INV_X1 U108 ( .A(A[34]), .ZN(n340) );
  XNOR2_X1 U109 ( .A(n326), .B(n350), .ZN(SUM[33]) );
  NAND2_X1 U110 ( .A1(n335), .A2(n333), .ZN(net185453) );
  OAI21_X1 U111 ( .B1(n340), .B2(net185453), .A(n347), .ZN(n348) );
  OAI21_X1 U112 ( .B1(n294), .B2(n340), .A(n347), .ZN(n341) );
  NAND2_X1 U113 ( .A1(net185453), .A2(n340), .ZN(n342) );
  INV_X1 U114 ( .A(B[34]), .ZN(n347) );
  XNOR2_X1 U115 ( .A(A[34]), .B(n347), .ZN(n338) );
  NAND2_X1 U116 ( .A1(n266), .A2(n346), .ZN(net185161) );
  XNOR2_X1 U117 ( .A(n265), .B(net182656), .ZN(SUM[35]) );
  INV_X1 U118 ( .A(n353), .ZN(n344) );
  CLKBUF_X1 U119 ( .A(A[33]), .Z(n353) );
  INV_X1 U120 ( .A(B[33]), .ZN(n336) );
  XNOR2_X1 U121 ( .A(A[33]), .B(n336), .ZN(n350) );
  OAI21_X1 U122 ( .B1(n345), .B2(n268), .A(B[31]), .ZN(n346) );
  AOI21_X1 U123 ( .B1(net185161), .B2(A[32]), .A(B[32]), .ZN(n343) );
  XNOR2_X1 U124 ( .A(A[32]), .B(B[32]), .ZN(net182464) );
  AOI21_X1 U125 ( .B1(n359), .B2(A[30]), .A(B[30]), .ZN(n349) );
  INV_X1 U126 ( .A(n362), .ZN(n359) );
  INV_X1 U127 ( .A(n352), .ZN(n354) );
  AOI21_X1 U128 ( .B1(n357), .B2(n358), .A(n354), .ZN(n362) );
  OAI21_X1 U129 ( .B1(n351), .B2(A[29]), .A(B[29]), .ZN(n352) );
  XNOR2_X1 U130 ( .A(net182434), .B(n357), .ZN(SUM[29]) );
  INV_X1 U131 ( .A(n359), .ZN(n356) );
  XNOR2_X1 U132 ( .A(n359), .B(net183946), .ZN(SUM[30]) );
  NAND2_X1 U133 ( .A1(n365), .A2(n368), .ZN(net185908) );
  INV_X1 U134 ( .A(A[30]), .ZN(net176675) );
  XNOR2_X1 U135 ( .A(A[30]), .B(B[30]), .ZN(net183946) );
  NOR2_X1 U136 ( .A1(n355), .A2(n363), .ZN(n351) );
  AND2_X1 U137 ( .A1(net184622), .A2(net176674), .ZN(n363) );
  XNOR2_X1 U138 ( .A(A[29]), .B(B[29]), .ZN(net182434) );
  CLKBUF_X1 U139 ( .A(A[35]), .Z(net187723) );
  INV_X2 U140 ( .A(B[38]), .ZN(n377) );
  NAND2_X1 U141 ( .A1(A[39]), .A2(B[39]), .ZN(n385) );
  INV_X1 U142 ( .A(n380), .ZN(net176705) );
  OAI21_X1 U143 ( .B1(n371), .B2(n377), .A(n383), .ZN(n380) );
  NAND2_X1 U144 ( .A1(A[38]), .A2(n293), .ZN(n383) );
  XNOR2_X1 U145 ( .A(A[38]), .B(B[38]), .ZN(net182465) );
  NOR2_X1 U146 ( .A1(net185908), .A2(A[38]), .ZN(n371) );
  INV_X1 U147 ( .A(B[39]), .ZN(n374) );
  XNOR2_X1 U148 ( .A(A[39]), .B(n374), .ZN(net190661) );
  NAND2_X1 U149 ( .A1(A[37]), .A2(B[37]), .ZN(n365) );
  OAI21_X1 U150 ( .B1(A[37]), .B2(B[37]), .A(net185452), .ZN(n368) );
  XNOR2_X1 U151 ( .A(A[37]), .B(B[37]), .ZN(net182676) );
  AOI21_X1 U152 ( .B1(net176705), .B2(n385), .A(n392), .ZN(n393) );
  NOR2_X1 U153 ( .A1(A[39]), .A2(B[39]), .ZN(n392) );
  AND2_X1 U154 ( .A1(net176691), .A2(net183664), .ZN(n394) );
  XNOR2_X1 U160 ( .A(net190661), .B(net176705), .ZN(SUM[39]) );
  NAND2_X1 U161 ( .A1(n332), .A2(n394), .ZN(n407) );
  XNOR2_X1 U162 ( .A(n269), .B(net182414), .ZN(SUM[31]) );
  XNOR2_X1 U163 ( .A(net190992), .B(net180768), .ZN(SUM[26]) );
  CLKBUF_X1 U164 ( .A(A[17]), .Z(n395) );
  AND2_X1 U165 ( .A1(net176691), .A2(net183664), .ZN(n396) );
  CLKBUF_X1 U166 ( .A(n420), .Z(n403) );
  XNOR2_X1 U167 ( .A(A[19]), .B(B[19]), .ZN(n397) );
  XNOR2_X1 U168 ( .A(n397), .B(n403), .ZN(SUM[19]) );
  INV_X1 U169 ( .A(n386), .ZN(n398) );
  CLKBUF_X1 U170 ( .A(n395), .Z(n399) );
  CLKBUF_X1 U171 ( .A(n378), .Z(net185094) );
  NOR2_X1 U172 ( .A1(n408), .A2(n400), .ZN(n409) );
  NAND2_X1 U173 ( .A1(net184159), .A2(n334), .ZN(n400) );
  XNOR2_X1 U174 ( .A(n401), .B(A[48]), .ZN(n310) );
  CLKBUF_X1 U175 ( .A(net185898), .Z(net185264) );
  CLKBUF_X1 U176 ( .A(A[16]), .Z(n402) );
  OAI21_X1 U177 ( .B1(n267), .B2(net187723), .A(B[35]), .ZN(n404) );
  XNOR2_X1 U178 ( .A(n421), .B(n405), .ZN(SUM[18]) );
  XNOR2_X1 U179 ( .A(A[18]), .B(B[18]), .ZN(n405) );
  NAND2_X1 U180 ( .A1(n404), .A2(net184159), .ZN(n406) );
  XNOR2_X1 U181 ( .A(n294), .B(n338), .ZN(SUM[34]) );
  NAND2_X1 U182 ( .A1(n364), .A2(n407), .ZN(n360) );
  XNOR2_X1 U183 ( .A(n307), .B(n308), .ZN(SUM[49]) );
  INV_X1 U184 ( .A(n423), .ZN(n408) );
  NOR2_X1 U185 ( .A1(n331), .A2(n409), .ZN(net185452) );
  XNOR2_X1 U186 ( .A(n406), .B(n410), .ZN(SUM[36]) );
  XNOR2_X1 U187 ( .A(A[36]), .B(B[36]), .ZN(n410) );
  INV_X1 U188 ( .A(net185898), .ZN(net183202) );
  CLKBUF_X1 U189 ( .A(A[18]), .Z(n411) );
  OR2_X1 U190 ( .A1(n422), .A2(n330), .ZN(n412) );
  NAND2_X1 U191 ( .A1(n412), .A2(n382), .ZN(n378) );
  BUF_X1 U192 ( .A(n387), .Z(n413) );
  AOI21_X1 U193 ( .B1(n425), .B2(n424), .A(n390), .ZN(n387) );
  CLKBUF_X1 U194 ( .A(A[40]), .Z(n414) );
  XNOR2_X1 U195 ( .A(n415), .B(net184620), .ZN(SUM[40]) );
  XNOR2_X1 U196 ( .A(A[40]), .B(B[40]), .ZN(n415) );
  XNOR2_X1 U197 ( .A(A[22]), .B(B[22]), .ZN(net182726) );
  XNOR2_X1 U198 ( .A(net182676), .B(n295), .ZN(SUM[37]) );
  XNOR2_X1 U199 ( .A(A[24]), .B(B[24]), .ZN(net182664) );
  XNOR2_X1 U200 ( .A(A[35]), .B(B[35]), .ZN(net182656) );
  XNOR2_X1 U201 ( .A(n416), .B(net185094), .ZN(SUM[20]) );
  XNOR2_X1 U202 ( .A(A[20]), .B(B[20]), .ZN(n416) );
  XNOR2_X1 U203 ( .A(net182465), .B(n293), .ZN(SUM[38]) );
  XNOR2_X1 U204 ( .A(net182464), .B(net185161), .ZN(SUM[32]) );
  XNOR2_X1 U205 ( .A(n417), .B(n394), .ZN(SUM[25]) );
  XNOR2_X1 U206 ( .A(A[25]), .B(B[25]), .ZN(n417) );
  XNOR2_X1 U207 ( .A(net182425), .B(net197646), .ZN(SUM[45]) );
  XNOR2_X1 U208 ( .A(n418), .B(net183202), .ZN(SUM[21]) );
  XNOR2_X1 U209 ( .A(A[21]), .B(B[21]), .ZN(n418) );
  OAI22_X1 U210 ( .A1(n411), .A2(n421), .B1(n384), .B2(B[18]), .ZN(n381) );
  AND2_X1 U211 ( .A1(n398), .A2(A[18]), .ZN(n384) );
  INV_X1 U212 ( .A(n311), .ZN(net176708) );
  INV_X1 U213 ( .A(n274), .ZN(n421) );
  OAI22_X1 U214 ( .A1(n395), .A2(n413), .B1(n388), .B2(B[17]), .ZN(n386) );
  AND2_X1 U215 ( .A1(A[17]), .A2(n387), .ZN(n388) );
  INV_X1 U216 ( .A(B[16]), .ZN(n425) );
  INV_X1 U217 ( .A(A[16]), .ZN(n424) );
  AOI21_X1 U218 ( .B1(A[16]), .B2(B[16]), .A(\carry[16] ), .ZN(n390) );
  AND2_X1 U219 ( .A1(A[0]), .A2(B[0]), .ZN(n1) );
  AOI21_X1 U220 ( .B1(n406), .B2(n408), .A(B[36]), .ZN(n331) );
  INV_X1 U221 ( .A(A[36]), .ZN(n423) );
  OAI21_X1 U222 ( .B1(n396), .B2(n332), .A(B[25]), .ZN(n364) );
  INV_X1 U223 ( .A(n304), .ZN(n419) );
  INV_X1 U224 ( .A(n367), .ZN(net176691) );
  INV_X1 U225 ( .A(n381), .ZN(n420) );
  OR2_X1 U226 ( .A1(A[40]), .A2(n393), .ZN(n306) );
  AOI22_X1 U227 ( .A1(net184620), .A2(n414), .B1(n306), .B2(B[40]), .ZN(n304)
         );
  OAI22_X1 U228 ( .A1(n309), .A2(B[48]), .B1(A[48]), .B2(net176708), .ZN(n307)
         );
  AND2_X1 U229 ( .A1(net176708), .A2(A[48]), .ZN(n309) );
  OAI21_X1 U230 ( .B1(n267), .B2(net187723), .A(B[35]), .ZN(n334) );
  OAI21_X1 U231 ( .B1(n420), .B2(A[19]), .A(B[19]), .ZN(n382) );
  INV_X1 U232 ( .A(A[19]), .ZN(n422) );
endmodule


module RCA_NBIT50 ( A, B, Ci, S, Co );
  input [49:0] A;
  input [49:0] B;
  output [49:0] S;
  input Ci;
  output Co;

  assign Co = 1'b0;

  RCA_NBIT50_DW01_add_0 add_95 ( .A(A), .B(B), .CI(1'b0), .SUM(S) );
endmodule


module RCA_NBIT52_DW01_add_0 ( A, B, CI, SUM, CO );
  input [51:0] A;
  input [51:0] B;
  output [51:0] SUM;
  input CI;
  output CO;
  wire   n1, \carry[49] , net79605, n352, n353, n355, n358, n359, n385, n389,
         n400, n403, n404, n406, n407, n410, n412, n413, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, net176742, net176749,
         net182687, net182723, net182728, net183283, net183365, net183876,
         net183884, net184123, net184329, net184328, net184355, net184776,
         net185303, net186814, net187464, net188928, net191198, net193264,
         net194111, n386, n383, n382, n379, net187214, net183460, net182460,
         net182422, n380, n377, n374, n373, net197753, net199641, net199639,
         net199630, net199625, net199623, n401, n398, n397, n395, n394, n365,
         net183362, n341, n339, n338, n336, n335, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n337, n340, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n354, n356, n357, n360,
         n361, n362, n363, n364, n366, n367, n368, n369, n370, n371, n372,
         n375, n376, n378, n381, n384, n387, n388, n390, n391, n392, n393,
         n396, n399, n402, n405, n408, n409, n411, n414, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496;
  wire   [51:1] carry;
  assign net79605 = A[45];

  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U162 ( .A(n488), .B(n417), .Z(SUM[21]) );
  XOR2_X1 U165 ( .A(n466), .B(n423), .Z(SUM[19]) );
  XOR2_X1 U166 ( .A(B[19]), .B(n470), .Z(n423) );
  XOR2_X1 U167 ( .A(n459), .B(n425), .Z(SUM[18]) );
  XOR2_X1 U168 ( .A(carry[18]), .B(B[18]), .Z(n425) );
  XOR2_X1 U169 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U1 ( .A(n321), .Z(net194111) );
  NAND2_X1 U2 ( .A1(n404), .A2(n450), .ZN(n291) );
  CLKBUF_X1 U3 ( .A(A[32]), .Z(n378) );
  OR2_X1 U4 ( .A1(net176742), .A2(net183884), .ZN(n292) );
  OR2_X1 U5 ( .A1(net176742), .A2(net183884), .ZN(n293) );
  OR2_X1 U6 ( .A1(net176742), .A2(net183884), .ZN(n428) );
  OR2_X2 U7 ( .A1(n409), .A2(n414), .ZN(net184328) );
  BUF_X1 U8 ( .A(A[31]), .Z(n294) );
  XNOR2_X1 U9 ( .A(n295), .B(net186814), .ZN(SUM[30]) );
  XOR2_X1 U10 ( .A(A[30]), .B(B[30]), .Z(n295) );
  BUF_X2 U11 ( .A(n373), .Z(n320) );
  INV_X1 U12 ( .A(n335), .ZN(n296) );
  OR2_X1 U13 ( .A1(n465), .A2(n353), .ZN(n330) );
  NOR2_X1 U14 ( .A1(n329), .A2(B[38]), .ZN(n365) );
  INV_X1 U15 ( .A(B[48]), .ZN(n304) );
  INV_X1 U16 ( .A(B[49]), .ZN(n468) );
  NAND2_X1 U17 ( .A1(net199623), .A2(n330), .ZN(n349) );
  AND2_X1 U18 ( .A1(net197753), .A2(n493), .ZN(n461) );
  INV_X1 U19 ( .A(B[37]), .ZN(n314) );
  NAND2_X1 U20 ( .A1(n346), .A2(n345), .ZN(n348) );
  INV_X1 U21 ( .A(B[44]), .ZN(n346) );
  OR2_X1 U22 ( .A1(n299), .A2(n365), .ZN(n297) );
  AND2_X1 U23 ( .A1(net199625), .A2(n349), .ZN(n298) );
  AND2_X1 U24 ( .A1(n319), .A2(n318), .ZN(n299) );
  AND2_X1 U25 ( .A1(B[44]), .A2(A[44]), .ZN(n300) );
  BUF_X1 U26 ( .A(n421), .Z(n466) );
  XNOR2_X1 U27 ( .A(net182460), .B(n325), .ZN(SUM[36]) );
  AOI21_X1 U28 ( .B1(n297), .B2(n308), .A(net182728), .ZN(n301) );
  BUF_X1 U29 ( .A(A[41]), .Z(n430) );
  AOI22_X1 U30 ( .A1(n343), .A2(n334), .B1(n336), .B2(B[47]), .ZN(n302) );
  OR2_X1 U31 ( .A1(n367), .A2(A[29]), .ZN(n375) );
  CLKBUF_X1 U32 ( .A(A[25]), .Z(n303) );
  INV_X1 U33 ( .A(B[39]), .ZN(net182728) );
  INV_X1 U34 ( .A(B[20]), .ZN(n475) );
  INV_X1 U35 ( .A(B[21]), .ZN(n467) );
  INV_X1 U36 ( .A(B[47]), .ZN(n340) );
  OR2_X1 U37 ( .A1(n335), .A2(n304), .ZN(n463) );
  CLKBUF_X1 U38 ( .A(n350), .Z(net183362) );
  NAND2_X1 U39 ( .A1(n361), .A2(n364), .ZN(n305) );
  NAND2_X1 U40 ( .A1(n375), .A2(B[29]), .ZN(n306) );
  NAND2_X1 U41 ( .A1(n305), .A2(n306), .ZN(n307) );
  AOI21_X1 U42 ( .B1(n297), .B2(n308), .A(net182728), .ZN(net176742) );
  INV_X1 U43 ( .A(A[39]), .ZN(n308) );
  OAI21_X1 U44 ( .B1(n313), .B2(n314), .A(n315), .ZN(n312) );
  NOR2_X1 U45 ( .A1(n309), .A2(A[37]), .ZN(n313) );
  OAI21_X1 U46 ( .B1(n322), .B2(n314), .A(n315), .ZN(n321) );
  NAND2_X1 U47 ( .A1(n309), .A2(A[37]), .ZN(n315) );
  INV_X1 U48 ( .A(n321), .ZN(n319) );
  NAND2_X1 U49 ( .A1(n311), .A2(n310), .ZN(n309) );
  NOR2_X1 U50 ( .A1(net188928), .A2(A[37]), .ZN(n322) );
  OAI21_X1 U51 ( .B1(n316), .B2(n328), .A(B[36]), .ZN(n311) );
  NAND2_X1 U52 ( .A1(n323), .A2(n310), .ZN(net188928) );
  OAI21_X1 U53 ( .B1(n316), .B2(n328), .A(B[36]), .ZN(n323) );
  XNOR2_X1 U54 ( .A(net182422), .B(n320), .ZN(SUM[35]) );
  NAND2_X1 U55 ( .A1(n317), .A2(n326), .ZN(n316) );
  NAND2_X1 U56 ( .A1(n327), .A2(n326), .ZN(n324) );
  NAND2_X1 U57 ( .A1(n326), .A2(n327), .ZN(n325) );
  XNOR2_X1 U58 ( .A(A[38]), .B(B[38]), .ZN(net183283) );
  INV_X1 U59 ( .A(A[38]), .ZN(n318) );
  NAND2_X1 U60 ( .A1(n320), .A2(A[35]), .ZN(n326) );
  NAND2_X1 U61 ( .A1(n374), .A2(B[35]), .ZN(n317) );
  NAND2_X1 U62 ( .A1(n374), .A2(B[35]), .ZN(n327) );
  NAND2_X1 U63 ( .A1(n328), .A2(n324), .ZN(n310) );
  BUF_X1 U64 ( .A(A[36]), .Z(n328) );
  AND2_X1 U65 ( .A1(A[38]), .A2(n312), .ZN(n329) );
  OR2_X1 U66 ( .A1(A[43]), .A2(B[43]), .ZN(net199625) );
  BUF_X1 U67 ( .A(n291), .Z(n331) );
  NOR2_X1 U68 ( .A1(B[45]), .A2(net79605), .ZN(net199639) );
  AND2_X1 U69 ( .A1(n495), .A2(n358), .ZN(n332) );
  AND2_X1 U70 ( .A1(n495), .A2(n358), .ZN(n472) );
  AOI22_X1 U71 ( .A1(n343), .A2(n334), .B1(n336), .B2(B[47]), .ZN(n335) );
  INV_X1 U72 ( .A(n302), .ZN(net176749) );
  OR2_X1 U73 ( .A1(n333), .A2(A[47]), .ZN(n336) );
  INV_X1 U74 ( .A(n339), .ZN(n333) );
  INV_X1 U75 ( .A(n333), .ZN(n342) );
  AOI22_X1 U76 ( .A1(n344), .A2(net183362), .B1(n341), .B2(B[46]), .ZN(n339)
         );
  OR2_X1 U77 ( .A1(n350), .A2(A[46]), .ZN(n341) );
  XNOR2_X1 U78 ( .A(n337), .B(net183362), .ZN(SUM[46]) );
  AOI21_X1 U79 ( .B1(n347), .B2(net199630), .A(net199639), .ZN(n350) );
  CLKBUF_X1 U80 ( .A(A[46]), .Z(n344) );
  CLKBUF_X1 U81 ( .A(A[47]), .Z(n334) );
  INV_X1 U82 ( .A(n342), .ZN(n343) );
  XNOR2_X1 U83 ( .A(n338), .B(n342), .ZN(SUM[47]) );
  XNOR2_X1 U84 ( .A(A[47]), .B(n340), .ZN(n338) );
  XNOR2_X1 U85 ( .A(A[46]), .B(B[46]), .ZN(n337) );
  OAI21_X1 U86 ( .B1(n298), .B2(n300), .A(n348), .ZN(n347) );
  INV_X1 U87 ( .A(n347), .ZN(net183365) );
  INV_X1 U88 ( .A(A[44]), .ZN(n345) );
  XNOR2_X1 U89 ( .A(net182723), .B(n298), .ZN(SUM[44]) );
  NAND2_X1 U90 ( .A1(n392), .A2(n391), .ZN(n351) );
  NAND2_X1 U91 ( .A1(n392), .A2(n391), .ZN(n354) );
  AND2_X1 U92 ( .A1(net184123), .A2(A[39]), .ZN(net183884) );
  XNOR2_X1 U93 ( .A(A[39]), .B(B[39]), .ZN(net183876) );
  NOR2_X1 U94 ( .A1(n365), .A2(n299), .ZN(net184123) );
  INV_X1 U95 ( .A(n372), .ZN(n367) );
  INV_X1 U96 ( .A(n395), .ZN(n360) );
  OAI21_X1 U97 ( .B1(n366), .B2(n368), .A(n360), .ZN(n372) );
  AOI21_X1 U98 ( .B1(n394), .B2(A[28]), .A(B[28]), .ZN(n395) );
  CLKBUF_X1 U99 ( .A(A[28]), .Z(n366) );
  BUF_X1 U100 ( .A(n394), .Z(n368) );
  XNOR2_X1 U101 ( .A(n362), .B(n368), .ZN(SUM[28]) );
  CLKBUF_X1 U102 ( .A(A[29]), .Z(n364) );
  AOI22_X1 U103 ( .A1(n361), .A2(n364), .B1(n375), .B2(B[29]), .ZN(net197753)
         );
  AOI22_X1 U104 ( .A1(n361), .A2(n364), .B1(n375), .B2(B[29]), .ZN(net186814)
         );
  INV_X1 U105 ( .A(n372), .ZN(n361) );
  XNOR2_X1 U106 ( .A(n363), .B(n361), .ZN(SUM[29]) );
  XNOR2_X1 U107 ( .A(A[29]), .B(B[29]), .ZN(n363) );
  OAI21_X1 U108 ( .B1(n397), .B2(n356), .A(n398), .ZN(n394) );
  OAI21_X1 U109 ( .B1(n370), .B2(A[27]), .A(B[27]), .ZN(n398) );
  AND2_X1 U110 ( .A1(n357), .A2(n369), .ZN(n370) );
  INV_X1 U111 ( .A(n401), .ZN(n357) );
  AND2_X1 U112 ( .A1(n357), .A2(n369), .ZN(net187464) );
  AOI21_X1 U113 ( .B1(n371), .B2(n400), .A(B[26]), .ZN(n401) );
  BUF_X1 U114 ( .A(A[26]), .Z(n371) );
  OR2_X1 U115 ( .A1(n371), .A2(n291), .ZN(n369) );
  INV_X1 U116 ( .A(A[27]), .ZN(n356) );
  INV_X1 U117 ( .A(net187464), .ZN(n397) );
  XNOR2_X1 U118 ( .A(A[28]), .B(B[28]), .ZN(n362) );
  BUF_X1 U119 ( .A(n432), .Z(n390) );
  CLKBUF_X1 U120 ( .A(A[23]), .Z(n449) );
  NOR2_X1 U121 ( .A1(n384), .A2(n461), .ZN(n376) );
  BUF_X1 U122 ( .A(A[24]), .Z(n453) );
  NOR2_X1 U123 ( .A1(n359), .A2(n332), .ZN(n381) );
  OR2_X1 U124 ( .A1(n409), .A2(n414), .ZN(n426) );
  AOI21_X1 U125 ( .B1(n307), .B2(n476), .A(B[30]), .ZN(n384) );
  AOI21_X1 U126 ( .B1(net184328), .B2(n378), .A(B[32]), .ZN(n387) );
  NAND2_X1 U127 ( .A1(net79605), .A2(B[45]), .ZN(net199630) );
  XNOR2_X1 U128 ( .A(A[44]), .B(B[44]), .ZN(net182723) );
  XNOR2_X1 U129 ( .A(A[43]), .B(B[43]), .ZN(n388) );
  NAND2_X1 U130 ( .A1(A[43]), .A2(B[43]), .ZN(net199623) );
  XNOR2_X1 U131 ( .A(n388), .B(net199641), .ZN(SUM[43]) );
  XNOR2_X1 U132 ( .A(net79605), .B(B[45]), .ZN(net184355) );
  INV_X1 U133 ( .A(n330), .ZN(net199641) );
  NAND2_X1 U134 ( .A1(B[49]), .A2(n443), .ZN(n391) );
  NAND2_X1 U135 ( .A1(\carry[49] ), .A2(n442), .ZN(n392) );
  OAI21_X1 U136 ( .B1(n355), .B2(n430), .A(B[41]), .ZN(n393) );
  XNOR2_X1 U137 ( .A(A[36]), .B(B[36]), .ZN(net182460) );
  OR2_X1 U138 ( .A1(n373), .A2(A[35]), .ZN(n374) );
  XNOR2_X1 U139 ( .A(A[35]), .B(B[35]), .ZN(net182422) );
  NOR2_X1 U140 ( .A1(n377), .A2(n396), .ZN(n373) );
  NOR2_X1 U141 ( .A1(n402), .A2(n405), .ZN(n396) );
  NAND2_X1 U142 ( .A1(n399), .A2(n380), .ZN(n405) );
  OAI21_X1 U143 ( .B1(net187214), .B2(n379), .A(B[33]), .ZN(n380) );
  INV_X1 U144 ( .A(net183460), .ZN(net187214) );
  OAI21_X1 U145 ( .B1(n379), .B2(net187214), .A(B[33]), .ZN(net191198) );
  INV_X1 U146 ( .A(A[33]), .ZN(net183460) );
  OR2_X1 U147 ( .A1(net185303), .A2(net183460), .ZN(net193264) );
  OR2_X1 U148 ( .A1(net183460), .A2(net185303), .ZN(n399) );
  BUF_X1 U149 ( .A(A[34]), .Z(n402) );
  AOI21_X1 U150 ( .B1(net184329), .B2(n402), .A(B[34]), .ZN(n377) );
  NOR2_X1 U151 ( .A1(n387), .A2(n427), .ZN(n379) );
  XNOR2_X1 U152 ( .A(n379), .B(net184776), .ZN(SUM[33]) );
  AND2_X1 U153 ( .A1(n408), .A2(n382), .ZN(n427) );
  INV_X1 U154 ( .A(A[32]), .ZN(n408) );
  AOI21_X1 U155 ( .B1(net184328), .B2(n378), .A(B[32]), .ZN(n383) );
  OR2_X1 U156 ( .A1(n383), .A2(n427), .ZN(net185303) );
  INV_X1 U157 ( .A(n386), .ZN(n409) );
  NOR2_X1 U158 ( .A1(n414), .A2(n409), .ZN(n382) );
  OAI21_X1 U159 ( .B1(n385), .B2(n294), .A(B[31]), .ZN(n386) );
  AND2_X1 U160 ( .A1(n376), .A2(n294), .ZN(n414) );
  XNOR2_X1 U161 ( .A(A[32]), .B(B[32]), .ZN(net182687) );
  XNOR2_X1 U163 ( .A(n411), .B(n376), .ZN(SUM[31]) );
  XNOR2_X1 U164 ( .A(A[31]), .B(B[31]), .ZN(n411) );
  AND2_X1 U170 ( .A1(n486), .A2(n454), .ZN(n429) );
  NAND2_X1 U171 ( .A1(n431), .A2(n449), .ZN(n455) );
  AND2_X1 U172 ( .A1(n448), .A2(n487), .ZN(n431) );
  CLKBUF_X1 U173 ( .A(A[20]), .Z(n441) );
  NAND2_X1 U174 ( .A1(n393), .A2(n452), .ZN(n432) );
  XOR2_X1 U175 ( .A(A[50]), .B(B[50]), .Z(n433) );
  XOR2_X1 U176 ( .A(n354), .B(n433), .Z(SUM[50]) );
  NAND2_X1 U177 ( .A1(n354), .A2(A[50]), .ZN(n434) );
  NAND2_X1 U178 ( .A1(n351), .A2(B[50]), .ZN(n435) );
  NAND2_X1 U179 ( .A1(A[50]), .A2(B[50]), .ZN(n436) );
  NAND3_X1 U180 ( .A1(n434), .A2(n435), .A3(n436), .ZN(carry[51]) );
  INV_X1 U181 ( .A(n491), .ZN(n437) );
  INV_X1 U182 ( .A(n440), .ZN(n438) );
  AOI21_X1 U183 ( .B1(n292), .B2(n457), .A(B[40]), .ZN(n439) );
  OAI22_X1 U184 ( .A1(n441), .A2(n489), .B1(B[20]), .B2(n418), .ZN(n440) );
  XNOR2_X1 U185 ( .A(A[49]), .B(n468), .ZN(n442) );
  CLKBUF_X1 U186 ( .A(A[49]), .Z(n443) );
  NOR2_X1 U187 ( .A1(n359), .A2(n332), .ZN(n444) );
  XNOR2_X1 U188 ( .A(n445), .B(n442), .ZN(SUM[49]) );
  AND3_X1 U189 ( .A1(n462), .A2(n463), .A3(n464), .ZN(n445) );
  AND2_X1 U190 ( .A1(n487), .A2(n448), .ZN(n446) );
  CLKBUF_X1 U191 ( .A(n412), .Z(n447) );
  BUF_X1 U192 ( .A(A[19]), .Z(n470) );
  NOR2_X1 U193 ( .A1(n439), .A2(n472), .ZN(n355) );
  XNOR2_X1 U194 ( .A(A[33]), .B(B[33]), .ZN(net184776) );
  OR2_X1 U195 ( .A1(A[22]), .A2(n412), .ZN(n448) );
  OR2_X1 U196 ( .A1(n403), .A2(n492), .ZN(n450) );
  NAND2_X1 U197 ( .A1(n404), .A2(n450), .ZN(n400) );
  XNOR2_X1 U198 ( .A(n296), .B(n451), .ZN(SUM[48]) );
  XNOR2_X1 U199 ( .A(A[48]), .B(B[48]), .ZN(n451) );
  XNOR2_X1 U200 ( .A(net184355), .B(net183365), .ZN(SUM[45]) );
  NAND2_X1 U201 ( .A1(net191198), .A2(net193264), .ZN(net184329) );
  AND2_X1 U202 ( .A1(n393), .A2(n452), .ZN(n352) );
  NAND2_X1 U203 ( .A1(n444), .A2(n430), .ZN(n452) );
  XNOR2_X1 U204 ( .A(n419), .B(n458), .ZN(SUM[20]) );
  XNOR2_X1 U205 ( .A(A[23]), .B(B[23]), .ZN(n471) );
  OR2_X1 U206 ( .A1(n406), .A2(n453), .ZN(n454) );
  NAND2_X1 U207 ( .A1(n486), .A2(n454), .ZN(n403) );
  NAND2_X1 U208 ( .A1(n410), .A2(n455), .ZN(n406) );
  OR2_X1 U209 ( .A1(n491), .A2(n415), .ZN(n456) );
  NAND2_X1 U210 ( .A1(n416), .A2(n456), .ZN(n412) );
  CLKBUF_X1 U211 ( .A(A[40]), .Z(n457) );
  NOR2_X1 U212 ( .A1(net183884), .A2(n301), .ZN(n358) );
  XNOR2_X1 U213 ( .A(net184123), .B(net183876), .ZN(SUM[39]) );
  OAI22_X1 U214 ( .A1(n470), .A2(n466), .B1(B[19]), .B2(n422), .ZN(n458) );
  INV_X1 U215 ( .A(n490), .ZN(n459) );
  CLKBUF_X1 U216 ( .A(A[48]), .Z(n460) );
  NOR2_X1 U217 ( .A1(n389), .A2(n461), .ZN(n385) );
  NAND2_X1 U218 ( .A1(net176749), .A2(n460), .ZN(n462) );
  NAND2_X1 U219 ( .A1(n460), .A2(B[48]), .ZN(n464) );
  NAND3_X1 U220 ( .A1(n462), .A2(n463), .A3(n464), .ZN(\carry[49] ) );
  AND2_X1 U221 ( .A1(n494), .A2(n352), .ZN(n465) );
  XNOR2_X1 U222 ( .A(A[21]), .B(n467), .ZN(n417) );
  XNOR2_X1 U223 ( .A(net183283), .B(net194111), .ZN(SUM[38]) );
  INV_X1 U224 ( .A(n420), .ZN(n469) );
  AOI21_X1 U225 ( .B1(n496), .B2(n490), .A(n424), .ZN(n421) );
  XNOR2_X1 U226 ( .A(n471), .B(n446), .ZN(SUM[23]) );
  XNOR2_X1 U227 ( .A(n473), .B(n429), .ZN(SUM[25]) );
  XNOR2_X1 U228 ( .A(A[25]), .B(B[25]), .ZN(n473) );
  XNOR2_X1 U229 ( .A(n474), .B(n447), .ZN(SUM[22]) );
  XNOR2_X1 U230 ( .A(A[22]), .B(B[22]), .ZN(n474) );
  XNOR2_X1 U231 ( .A(A[20]), .B(n475), .ZN(n419) );
  INV_X1 U232 ( .A(n493), .ZN(n476) );
  XNOR2_X1 U233 ( .A(n426), .B(net182687), .ZN(SUM[32]) );
  XNOR2_X1 U234 ( .A(net188928), .B(n477), .ZN(SUM[37]) );
  XNOR2_X1 U235 ( .A(A[37]), .B(B[37]), .ZN(n477) );
  XNOR2_X1 U236 ( .A(n478), .B(n406), .ZN(SUM[24]) );
  XNOR2_X1 U237 ( .A(A[24]), .B(B[24]), .ZN(n478) );
  XNOR2_X1 U238 ( .A(n331), .B(n479), .ZN(SUM[26]) );
  XNOR2_X1 U239 ( .A(A[26]), .B(B[26]), .ZN(n479) );
  XNOR2_X1 U240 ( .A(n480), .B(n381), .ZN(SUM[41]) );
  XNOR2_X1 U241 ( .A(A[41]), .B(B[41]), .ZN(n480) );
  XNOR2_X1 U242 ( .A(n293), .B(n481), .ZN(SUM[40]) );
  XNOR2_X1 U243 ( .A(A[40]), .B(B[40]), .ZN(n481) );
  XNOR2_X1 U244 ( .A(n482), .B(n390), .ZN(SUM[42]) );
  XNOR2_X1 U245 ( .A(A[42]), .B(B[42]), .ZN(n482) );
  XNOR2_X1 U246 ( .A(net184329), .B(n483), .ZN(SUM[34]) );
  XNOR2_X1 U247 ( .A(A[34]), .B(B[34]), .ZN(n483) );
  INV_X1 U248 ( .A(A[42]), .ZN(n494) );
  AOI21_X1 U249 ( .B1(A[42]), .B2(n432), .A(B[42]), .ZN(n353) );
  XNOR2_X1 U250 ( .A(n484), .B(net187464), .ZN(SUM[27]) );
  XNOR2_X1 U251 ( .A(A[27]), .B(B[27]), .ZN(n484) );
  XNOR2_X1 U252 ( .A(n485), .B(A[51]), .ZN(SUM[51]) );
  XNOR2_X1 U253 ( .A(carry[51]), .B(B[51]), .ZN(n485) );
  OAI22_X1 U254 ( .A1(n441), .A2(n489), .B1(n418), .B2(B[20]), .ZN(n415) );
  AND2_X1 U255 ( .A1(n469), .A2(A[20]), .ZN(n418) );
  INV_X1 U256 ( .A(B[18]), .ZN(n496) );
  INV_X1 U257 ( .A(A[18]), .ZN(n490) );
  AOI21_X1 U258 ( .B1(A[18]), .B2(B[18]), .A(carry[18]), .ZN(n424) );
  AND2_X1 U259 ( .A1(A[0]), .A2(B[0]), .ZN(n1) );
  INV_X1 U260 ( .A(A[40]), .ZN(n495) );
  OAI21_X1 U261 ( .B1(n446), .B2(n449), .A(B[23]), .ZN(n410) );
  INV_X1 U262 ( .A(A[25]), .ZN(n492) );
  INV_X1 U263 ( .A(A[30]), .ZN(n493) );
  OAI21_X1 U264 ( .B1(n438), .B2(n437), .A(B[21]), .ZN(n416) );
  INV_X1 U265 ( .A(A[21]), .ZN(n491) );
  AOI21_X1 U266 ( .B1(n307), .B2(n476), .A(B[30]), .ZN(n389) );
  OAI21_X1 U267 ( .B1(n429), .B2(n303), .A(B[25]), .ZN(n404) );
  AOI21_X1 U268 ( .B1(n428), .B2(n457), .A(B[40]), .ZN(n359) );
  INV_X1 U269 ( .A(n407), .ZN(n486) );
  INV_X1 U270 ( .A(n413), .ZN(n487) );
  AOI21_X1 U271 ( .B1(n412), .B2(A[22]), .A(B[22]), .ZN(n413) );
  INV_X1 U272 ( .A(n415), .ZN(n488) );
  OAI22_X1 U273 ( .A1(n470), .A2(n466), .B1(n422), .B2(B[19]), .ZN(n420) );
  AND2_X1 U274 ( .A1(A[19]), .A2(n421), .ZN(n422) );
  AOI21_X1 U275 ( .B1(n406), .B2(n453), .A(B[24]), .ZN(n407) );
  INV_X1 U276 ( .A(n458), .ZN(n489) );
endmodule


module RCA_NBIT52 ( A, B, Ci, S, Co );
  input [51:0] A;
  input [51:0] B;
  output [51:0] S;
  input Ci;
  output Co;

  assign Co = 1'b0;

  RCA_NBIT52_DW01_add_0 add_95 ( .A(A), .B(B), .CI(1'b0), .SUM(S) );
endmodule


module RCA_NBIT54_DW01_add_0 ( A, B, CI, SUM, CO );
  input [53:0] A;
  input [53:0] B;
  output [53:0] SUM;
  input CI;
  output CO;
  wire   n1, \carry[49] , \carry[48] , \carry[47] , \carry[46] , n228, n230,
         n231, n232, n235, n236, n238, n249, n260, n261, n268, n269, n271,
         n272, n273, n274, n275, n277, n278, n280, n281, n283, n284, n285,
         n286, n287, n289, n290, n292, n293, n295, n296, n297, n298, n299,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, net176760,
         net182670, net182990, net183126, net184052, net184628, net184627,
         net185339, net185683, net186877, net187258, n243, n241, net183875,
         n256, net186932, net185970, net183577, net193528, net182754,
         net182747, net182702, net176759, n257, n250, net203253, net185306,
         net184333, net183714, net176788, net176757, n251, n248, n245, n244,
         n242, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506;
  wire   [53:1] carry;

  FA_X1 U1_50 ( .A(A[50]), .B(B[50]), .CI(n437), .CO(carry[51]), .S(SUM[50])
         );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  FA_X1 U1_48 ( .A(B[48]), .B(\carry[48] ), .CI(A[48]), .CO(\carry[49] ), .S(
        SUM[48]) );
  FA_X1 U1_47 ( .A(A[47]), .B(B[47]), .CI(\carry[47] ), .CO(\carry[48] ), .S(
        SUM[47]) );
  XOR2_X1 U128 ( .A(n228), .B(carry[51]), .Z(SUM[51]) );
  XOR2_X1 U130 ( .A(n230), .B(\carry[49] ), .Z(SUM[49]) );
  XOR2_X1 U167 ( .A(A[22]), .B(B[22]), .Z(n303) );
  XOR2_X1 U168 ( .A(n474), .B(n306), .Z(SUM[21]) );
  XOR2_X1 U169 ( .A(B[21]), .B(n483), .Z(n306) );
  XOR2_X1 U170 ( .A(B[20]), .B(n427), .Z(n309) );
  XOR2_X1 U171 ( .A(B[19]), .B(A[19]), .Z(n312) );
  XOR2_X1 U172 ( .A(B[18]), .B(A[18]), .Z(n315) );
  XOR2_X1 U173 ( .A(B[17]), .B(A[17]), .Z(n318) );
  XOR2_X1 U174 ( .A(A[16]), .B(n320), .Z(SUM[16]) );
  XOR2_X1 U175 ( .A(carry[16]), .B(B[16]), .Z(n320) );
  XOR2_X1 U176 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  OR2_X1 U1 ( .A1(n235), .A2(n502), .ZN(n472) );
  BUF_X1 U2 ( .A(A[40]), .Z(n386) );
  BUF_X1 U3 ( .A(A[31]), .Z(n414) );
  BUF_X1 U4 ( .A(n467), .Z(n377) );
  OR2_X1 U5 ( .A1(n368), .A2(n493), .ZN(n367) );
  OR2_X2 U6 ( .A1(net184333), .A2(n379), .ZN(net203253) );
  AND2_X1 U7 ( .A1(n474), .A2(n483), .ZN(n368) );
  BUF_X1 U8 ( .A(n304), .Z(n474) );
  BUF_X1 U9 ( .A(A[21]), .Z(n483) );
  INV_X1 U10 ( .A(n251), .ZN(n369) );
  OAI21_X1 U11 ( .B1(n250), .B2(net182702), .A(B[39]), .ZN(n370) );
  INV_X1 U12 ( .A(B[35]), .ZN(n392) );
  INV_X1 U13 ( .A(B[49]), .ZN(n465) );
  BUF_X1 U14 ( .A(A[28]), .Z(n417) );
  CLKBUF_X1 U15 ( .A(n440), .Z(n371) );
  NOR2_X1 U16 ( .A1(net176788), .A2(net183577), .ZN(n372) );
  CLKBUF_X1 U17 ( .A(A[23]), .Z(n430) );
  INV_X1 U18 ( .A(B[36]), .ZN(n396) );
  INV_X1 U19 ( .A(B[40]), .ZN(net185970) );
  INV_X1 U20 ( .A(B[51]), .ZN(n473) );
  INV_X1 U21 ( .A(B[38]), .ZN(n401) );
  INV_X1 U22 ( .A(B[43]), .ZN(n374) );
  INV_X1 U23 ( .A(B[32]), .ZN(n452) );
  NOR2_X1 U24 ( .A1(n375), .A2(n374), .ZN(n373) );
  NOR2_X1 U25 ( .A1(n238), .A2(n482), .ZN(n375) );
  BUF_X1 U26 ( .A(A[43]), .Z(n482) );
  INV_X1 U27 ( .A(B[24]), .ZN(n462) );
  INV_X1 U28 ( .A(B[42]), .ZN(n381) );
  INV_X1 U29 ( .A(B[28]), .ZN(n453) );
  OR2_X1 U30 ( .A1(n488), .A2(n449), .ZN(n412) );
  NAND2_X1 U31 ( .A1(n370), .A2(n376), .ZN(net185306) );
  INV_X1 U32 ( .A(net183577), .ZN(n376) );
  NOR2_X1 U33 ( .A1(n387), .A2(A[35]), .ZN(n391) );
  NOR2_X1 U34 ( .A1(n369), .A2(net183577), .ZN(net184333) );
  NOR2_X1 U35 ( .A1(n380), .A2(n383), .ZN(n241) );
  XNOR2_X1 U36 ( .A(n243), .B(n241), .ZN(SUM[42]) );
  BUF_X1 U37 ( .A(A[39]), .Z(net182702) );
  NOR2_X1 U38 ( .A1(n488), .A2(n449), .ZN(n378) );
  XNOR2_X1 U39 ( .A(net185339), .B(n395), .ZN(SUM[34]) );
  OAI21_X1 U40 ( .B1(n384), .B2(net183714), .A(B[42]), .ZN(n242) );
  NAND2_X1 U41 ( .A1(n242), .A2(net183126), .ZN(n238) );
  INV_X1 U42 ( .A(net176757), .ZN(net183714) );
  OAI21_X1 U43 ( .B1(n385), .B2(net183714), .A(B[42]), .ZN(net184628) );
  INV_X1 U44 ( .A(A[42]), .ZN(net176757) );
  OR2_X1 U45 ( .A1(n241), .A2(net176757), .ZN(net183126) );
  OR2_X1 U46 ( .A1(n380), .A2(n383), .ZN(n384) );
  INV_X1 U47 ( .A(n245), .ZN(n380) );
  OR2_X1 U48 ( .A1(n380), .A2(n383), .ZN(n385) );
  OAI21_X1 U49 ( .B1(n244), .B2(n382), .A(B[41]), .ZN(n245) );
  BUF_X1 U50 ( .A(A[41]), .Z(n382) );
  AND2_X1 U51 ( .A1(n382), .A2(net186877), .ZN(n383) );
  NAND2_X1 U52 ( .A1(n248), .A2(net203253), .ZN(n244) );
  INV_X1 U53 ( .A(A[40]), .ZN(n379) );
  OAI21_X1 U54 ( .B1(net185306), .B2(n386), .A(B[40]), .ZN(n248) );
  OAI21_X1 U55 ( .B1(n386), .B2(net185306), .A(B[40]), .ZN(net186932) );
  XNOR2_X1 U56 ( .A(A[42]), .B(n381), .ZN(n243) );
  XNOR2_X1 U57 ( .A(A[41]), .B(B[41]), .ZN(net182670) );
  XNOR2_X1 U58 ( .A(n249), .B(n372), .ZN(SUM[40]) );
  INV_X1 U59 ( .A(n370), .ZN(net176788) );
  OAI21_X1 U60 ( .B1(n250), .B2(net182702), .A(B[39]), .ZN(n251) );
  INV_X1 U61 ( .A(n390), .ZN(net184052) );
  OAI21_X1 U62 ( .B1(n391), .B2(n392), .A(n393), .ZN(n390) );
  BUF_X1 U63 ( .A(A[37]), .Z(n404) );
  NAND2_X1 U64 ( .A1(n260), .A2(net184627), .ZN(n256) );
  NAND2_X1 U65 ( .A1(n388), .A2(n389), .ZN(n387) );
  OAI21_X1 U66 ( .B1(A[36]), .B2(n390), .A(B[36]), .ZN(n260) );
  INV_X1 U67 ( .A(A[36]), .ZN(net176760) );
  XNOR2_X1 U68 ( .A(A[35]), .B(B[35]), .ZN(n394) );
  NAND2_X1 U69 ( .A1(A[35]), .A2(n387), .ZN(n393) );
  XNOR2_X1 U70 ( .A(A[34]), .B(B[34]), .ZN(n395) );
  NAND2_X1 U71 ( .A1(n397), .A2(B[34]), .ZN(n388) );
  OAI21_X1 U72 ( .B1(B[34]), .B2(n397), .A(net185339), .ZN(n389) );
  XNOR2_X1 U73 ( .A(A[36]), .B(n396), .ZN(n261) );
  XNOR2_X1 U74 ( .A(n394), .B(n387), .ZN(SUM[35]) );
  CLKBUF_X1 U75 ( .A(A[34]), .Z(n397) );
  OR2_X1 U76 ( .A1(net176759), .A2(net193528), .ZN(n398) );
  AND2_X1 U77 ( .A1(n257), .A2(n403), .ZN(n399) );
  OAI21_X1 U78 ( .B1(n402), .B2(A[38]), .A(B[38]), .ZN(n400) );
  AND2_X1 U79 ( .A1(net187258), .A2(net182702), .ZN(net183577) );
  NAND2_X1 U80 ( .A1(net182747), .A2(n400), .ZN(n250) );
  XNOR2_X1 U81 ( .A(A[39]), .B(B[39]), .ZN(net182990) );
  OR2_X1 U82 ( .A1(net176759), .A2(net193528), .ZN(net182747) );
  NAND2_X1 U83 ( .A1(n398), .A2(n400), .ZN(net187258) );
  INV_X1 U84 ( .A(A[38]), .ZN(net176759) );
  NAND2_X1 U85 ( .A1(n405), .A2(n403), .ZN(n402) );
  OAI21_X1 U86 ( .B1(n256), .B2(n404), .A(B[37]), .ZN(n405) );
  OAI21_X1 U87 ( .B1(n256), .B2(n404), .A(B[37]), .ZN(n257) );
  NAND2_X1 U88 ( .A1(net185683), .A2(n404), .ZN(n403) );
  XNOR2_X1 U89 ( .A(net182754), .B(n399), .ZN(SUM[38]) );
  XNOR2_X1 U90 ( .A(A[38]), .B(n401), .ZN(net182754) );
  AND2_X1 U91 ( .A1(n257), .A2(n403), .ZN(net193528) );
  XNOR2_X1 U92 ( .A(A[37]), .B(B[37]), .ZN(net183875) );
  XNOR2_X1 U93 ( .A(A[40]), .B(net185970), .ZN(n249) );
  NAND2_X1 U94 ( .A1(net203253), .A2(net186932), .ZN(net186877) );
  XNOR2_X1 U95 ( .A(net185683), .B(net183875), .ZN(SUM[37]) );
  OR2_X1 U96 ( .A1(n469), .A2(n373), .ZN(n406) );
  NOR2_X1 U97 ( .A1(n492), .A2(n468), .ZN(n289) );
  CLKBUF_X1 U98 ( .A(A[29]), .Z(n486) );
  OR2_X1 U99 ( .A1(n408), .A2(n491), .ZN(n407) );
  BUF_X1 U100 ( .A(A[27]), .Z(n484) );
  AND2_X1 U101 ( .A1(n467), .A2(n484), .ZN(n408) );
  BUF_X1 U102 ( .A(n286), .Z(n467) );
  OR2_X1 U103 ( .A1(n468), .A2(n492), .ZN(n409) );
  AOI22_X1 U104 ( .A1(B[51]), .A2(n464), .B1(n228), .B2(carry[51]), .ZN(n410)
         );
  CLKBUF_X1 U105 ( .A(A[33]), .Z(n411) );
  CLKBUF_X1 U106 ( .A(n475), .Z(n438) );
  OAI21_X1 U107 ( .B1(n448), .B2(n463), .A(B[44]), .ZN(n413) );
  BUF_X1 U108 ( .A(n283), .Z(n476) );
  OAI21_X1 U109 ( .B1(n412), .B2(n429), .A(B[32]), .ZN(n415) );
  OAI21_X1 U110 ( .B1(n301), .B2(n506), .A(n302), .ZN(n298) );
  NAND2_X1 U111 ( .A1(n413), .A2(n472), .ZN(n416) );
  NAND2_X1 U112 ( .A1(n446), .A2(n272), .ZN(n418) );
  XNOR2_X1 U113 ( .A(n410), .B(n419), .ZN(SUM[52]) );
  XOR2_X1 U114 ( .A(A[52]), .B(B[52]), .Z(n419) );
  CLKBUF_X1 U115 ( .A(n232), .Z(n420) );
  BUF_X1 U116 ( .A(n456), .Z(n421) );
  OAI21_X1 U117 ( .B1(n489), .B2(n433), .A(B[30]), .ZN(n422) );
  NAND2_X1 U118 ( .A1(n423), .A2(n424), .ZN(n437) );
  NAND2_X1 U119 ( .A1(n230), .A2(\carry[49] ), .ZN(n423) );
  NAND2_X1 U120 ( .A1(n426), .A2(B[49]), .ZN(n424) );
  BUF_X1 U121 ( .A(A[46]), .Z(n431) );
  OAI21_X1 U122 ( .B1(n420), .B2(n371), .A(B[45]), .ZN(n425) );
  CLKBUF_X1 U123 ( .A(A[49]), .Z(n426) );
  INV_X1 U124 ( .A(n432), .ZN(n295) );
  CLKBUF_X1 U125 ( .A(A[20]), .Z(n427) );
  NAND2_X1 U126 ( .A1(n422), .A2(n454), .ZN(n428) );
  XNOR2_X1 U127 ( .A(A[46]), .B(B[46]), .ZN(n436) );
  BUF_X1 U129 ( .A(n280), .Z(n456) );
  INV_X1 U131 ( .A(n501), .ZN(n429) );
  BUF_X1 U132 ( .A(A[45]), .Z(n440) );
  NAND2_X1 U133 ( .A1(net184627), .A2(n260), .ZN(net185683) );
  XNOR2_X1 U134 ( .A(n460), .B(A[53]), .ZN(SUM[53]) );
  NAND2_X1 U135 ( .A1(n299), .A2(n451), .ZN(n432) );
  INV_X1 U136 ( .A(n500), .ZN(n433) );
  NAND2_X1 U137 ( .A1(n269), .A2(n441), .ZN(net185339) );
  NAND2_X1 U138 ( .A1(n416), .A2(n440), .ZN(n470) );
  XNOR2_X1 U139 ( .A(n406), .B(n435), .ZN(SUM[44]) );
  OR2_X1 U140 ( .A1(n373), .A2(n469), .ZN(n434) );
  XNOR2_X1 U141 ( .A(A[44]), .B(B[44]), .ZN(n435) );
  XNOR2_X1 U142 ( .A(n436), .B(\carry[46] ), .ZN(SUM[46]) );
  XNOR2_X1 U143 ( .A(n439), .B(n289), .ZN(SUM[26]) );
  XOR2_X1 U144 ( .A(A[26]), .B(B[26]), .Z(n439) );
  NAND2_X1 U145 ( .A1(n418), .A2(n411), .ZN(n441) );
  XNOR2_X1 U146 ( .A(n438), .B(n442), .ZN(SUM[25]) );
  XNOR2_X1 U147 ( .A(A[25]), .B(B[25]), .ZN(n442) );
  NAND2_X1 U148 ( .A1(n231), .A2(n470), .ZN(n443) );
  OR2_X1 U149 ( .A1(net176760), .A2(net184052), .ZN(net184627) );
  XNOR2_X1 U150 ( .A(n444), .B(n416), .ZN(SUM[45]) );
  XNOR2_X1 U151 ( .A(A[45]), .B(B[45]), .ZN(n444) );
  XNOR2_X1 U152 ( .A(n445), .B(n447), .ZN(SUM[30]) );
  XOR2_X1 U153 ( .A(A[30]), .B(B[30]), .Z(n445) );
  OR2_X1 U154 ( .A1(n501), .A2(n271), .ZN(n446) );
  NAND2_X1 U155 ( .A1(n415), .A2(n446), .ZN(n268) );
  AOI21_X1 U156 ( .B1(n421), .B2(n486), .A(n490), .ZN(n447) );
  AOI21_X1 U157 ( .B1(n421), .B2(n486), .A(n490), .ZN(n277) );
  OR2_X1 U158 ( .A1(n373), .A2(n469), .ZN(n448) );
  AND2_X1 U159 ( .A1(n428), .A2(n414), .ZN(n449) );
  NOR2_X1 U160 ( .A1(n488), .A2(n449), .ZN(n271) );
  NAND2_X1 U161 ( .A1(net183126), .A2(net184628), .ZN(n450) );
  NAND2_X1 U162 ( .A1(n298), .A2(n430), .ZN(n451) );
  XNOR2_X1 U163 ( .A(A[32]), .B(n452), .ZN(n273) );
  XNOR2_X1 U164 ( .A(A[28]), .B(n453), .ZN(n285) );
  OR2_X1 U165 ( .A1(n447), .A2(n500), .ZN(n454) );
  NAND2_X1 U166 ( .A1(n278), .A2(n454), .ZN(n274) );
  NOR2_X1 U177 ( .A1(n469), .A2(n373), .ZN(n235) );
  XNOR2_X1 U178 ( .A(n428), .B(n455), .ZN(SUM[31]) );
  XNOR2_X1 U179 ( .A(A[31]), .B(B[31]), .ZN(n455) );
  NAND2_X1 U180 ( .A1(n487), .A2(A[52]), .ZN(n457) );
  NAND2_X1 U181 ( .A1(n487), .A2(B[52]), .ZN(n458) );
  NAND2_X1 U182 ( .A1(A[52]), .A2(B[52]), .ZN(n459) );
  NAND3_X1 U183 ( .A1(n457), .A2(n458), .A3(n459), .ZN(carry[53]) );
  XNOR2_X1 U184 ( .A(carry[53]), .B(B[53]), .ZN(n460) );
  XNOR2_X1 U185 ( .A(A[23]), .B(B[23]), .ZN(n461) );
  XNOR2_X1 U186 ( .A(n461), .B(n298), .ZN(SUM[23]) );
  XNOR2_X1 U187 ( .A(A[24]), .B(n462), .ZN(n297) );
  INV_X1 U188 ( .A(n502), .ZN(n463) );
  CLKBUF_X1 U189 ( .A(A[51]), .Z(n464) );
  XNOR2_X1 U190 ( .A(A[49]), .B(n465), .ZN(n230) );
  XNOR2_X1 U191 ( .A(n466), .B(n450), .ZN(SUM[43]) );
  XNOR2_X1 U192 ( .A(A[43]), .B(B[43]), .ZN(n466) );
  AND2_X1 U193 ( .A1(n475), .A2(A[25]), .ZN(n468) );
  BUF_X1 U194 ( .A(n292), .Z(n475) );
  AOI21_X1 U195 ( .B1(n474), .B2(n483), .A(n493), .ZN(n301) );
  AND2_X1 U196 ( .A1(n450), .A2(n482), .ZN(n469) );
  NAND2_X1 U197 ( .A1(n470), .A2(n425), .ZN(\carry[46] ) );
  OR2_X1 U198 ( .A1(n289), .A2(n504), .ZN(n471) );
  NAND2_X1 U199 ( .A1(n290), .A2(n471), .ZN(n286) );
  NAND2_X1 U200 ( .A1(n236), .A2(n472), .ZN(n232) );
  XNOR2_X1 U201 ( .A(A[51]), .B(n473), .ZN(n228) );
  XNOR2_X1 U202 ( .A(net187258), .B(net182990), .ZN(SUM[39]) );
  AOI21_X1 U203 ( .B1(n467), .B2(n484), .A(n491), .ZN(n283) );
  NAND2_X1 U204 ( .A1(n443), .A2(n431), .ZN(n477) );
  NAND2_X1 U205 ( .A1(n443), .A2(B[46]), .ZN(n478) );
  NAND2_X1 U206 ( .A1(n431), .A2(B[46]), .ZN(n479) );
  NAND3_X1 U207 ( .A1(n478), .A2(n477), .A3(n479), .ZN(\carry[47] ) );
  XNOR2_X1 U208 ( .A(n377), .B(n480), .ZN(SUM[27]) );
  XNOR2_X1 U209 ( .A(A[27]), .B(B[27]), .ZN(n480) );
  XNOR2_X1 U210 ( .A(n481), .B(n456), .ZN(SUM[29]) );
  XNOR2_X1 U211 ( .A(A[29]), .B(B[29]), .ZN(n481) );
  XNOR2_X1 U212 ( .A(net182670), .B(net186877), .ZN(SUM[41]) );
  INV_X1 U213 ( .A(A[22]), .ZN(n506) );
  OAI21_X1 U214 ( .B1(n367), .B2(A[22]), .A(B[22]), .ZN(n302) );
  INV_X1 U215 ( .A(n410), .ZN(n487) );
  OAI21_X1 U216 ( .B1(n307), .B2(n499), .A(n308), .ZN(n304) );
  INV_X1 U217 ( .A(n427), .ZN(n499) );
  OAI21_X1 U218 ( .B1(A[20]), .B2(n494), .A(B[20]), .ZN(n308) );
  INV_X1 U219 ( .A(n307), .ZN(n494) );
  AOI22_X1 U220 ( .A1(n495), .A2(A[19]), .B1(n310), .B2(B[19]), .ZN(n307) );
  OR2_X1 U221 ( .A1(A[19]), .A2(n495), .ZN(n310) );
  INV_X1 U222 ( .A(n311), .ZN(n495) );
  AOI22_X1 U223 ( .A1(n497), .A2(A[17]), .B1(n316), .B2(B[17]), .ZN(n314) );
  OR2_X1 U224 ( .A1(A[17]), .A2(n497), .ZN(n316) );
  INV_X1 U225 ( .A(n317), .ZN(n497) );
  AOI22_X1 U226 ( .A1(n496), .A2(A[18]), .B1(n313), .B2(B[18]), .ZN(n311) );
  OR2_X1 U227 ( .A1(A[18]), .A2(n496), .ZN(n313) );
  INV_X1 U228 ( .A(n314), .ZN(n496) );
  AOI21_X1 U229 ( .B1(A[16]), .B2(B[16]), .A(n498), .ZN(n317) );
  INV_X1 U230 ( .A(n319), .ZN(n498) );
  OAI21_X1 U231 ( .B1(A[16]), .B2(B[16]), .A(carry[16]), .ZN(n319) );
  XNOR2_X1 U232 ( .A(n317), .B(n318), .ZN(SUM[17]) );
  XNOR2_X1 U233 ( .A(n314), .B(n315), .ZN(SUM[18]) );
  XNOR2_X1 U234 ( .A(n311), .B(n312), .ZN(SUM[19]) );
  XNOR2_X1 U235 ( .A(n307), .B(n309), .ZN(SUM[20]) );
  AND2_X1 U236 ( .A1(A[0]), .A2(B[0]), .ZN(n1) );
  INV_X1 U237 ( .A(A[44]), .ZN(n502) );
  INV_X1 U238 ( .A(n275), .ZN(n488) );
  XNOR2_X1 U239 ( .A(n418), .B(n485), .ZN(SUM[33]) );
  XNOR2_X1 U240 ( .A(A[33]), .B(B[33]), .ZN(n485) );
  INV_X1 U241 ( .A(A[30]), .ZN(n500) );
  INV_X1 U242 ( .A(A[32]), .ZN(n501) );
  OAI21_X1 U243 ( .B1(n412), .B2(n429), .A(B[32]), .ZN(n272) );
  OAI21_X1 U244 ( .B1(n432), .B2(A[24]), .A(B[24]), .ZN(n296) );
  INV_X1 U245 ( .A(A[24]), .ZN(n505) );
  OAI21_X1 U246 ( .B1(A[21]), .B2(n304), .A(B[21]), .ZN(n305) );
  OAI21_X1 U247 ( .B1(n268), .B2(n411), .A(B[33]), .ZN(n269) );
  INV_X1 U248 ( .A(n287), .ZN(n491) );
  OAI21_X1 U249 ( .B1(n232), .B2(n440), .A(B[45]), .ZN(n231) );
  OAI21_X1 U250 ( .B1(n489), .B2(n433), .A(B[30]), .ZN(n278) );
  INV_X1 U251 ( .A(n293), .ZN(n492) );
  XNOR2_X1 U252 ( .A(n273), .B(n378), .ZN(SUM[32]) );
  OAI21_X1 U253 ( .B1(n274), .B2(n414), .A(B[31]), .ZN(n275) );
  INV_X1 U254 ( .A(n281), .ZN(n490) );
  OAI21_X1 U255 ( .B1(A[27]), .B2(n286), .A(B[27]), .ZN(n287) );
  OAI21_X1 U256 ( .B1(n298), .B2(n430), .A(B[23]), .ZN(n299) );
  INV_X1 U257 ( .A(n305), .ZN(n493) );
  INV_X1 U258 ( .A(A[26]), .ZN(n504) );
  OAI21_X1 U259 ( .B1(n409), .B2(A[26]), .A(B[26]), .ZN(n290) );
  OAI21_X1 U260 ( .B1(n434), .B2(n463), .A(B[44]), .ZN(n236) );
  INV_X1 U261 ( .A(n417), .ZN(n503) );
  OAI21_X1 U262 ( .B1(n407), .B2(n417), .A(B[28]), .ZN(n284) );
  OAI21_X1 U263 ( .B1(n280), .B2(A[29]), .A(B[29]), .ZN(n281) );
  XNOR2_X1 U264 ( .A(net184052), .B(n261), .ZN(SUM[36]) );
  INV_X1 U265 ( .A(n277), .ZN(n489) );
  XNOR2_X1 U266 ( .A(n476), .B(n285), .ZN(SUM[28]) );
  OAI21_X1 U267 ( .B1(n476), .B2(n503), .A(n284), .ZN(n280) );
  OAI21_X1 U268 ( .B1(A[25]), .B2(n292), .A(B[25]), .ZN(n293) );
  XNOR2_X1 U269 ( .A(n297), .B(n295), .ZN(SUM[24]) );
  OAI21_X1 U270 ( .B1(n295), .B2(n505), .A(n296), .ZN(n292) );
  XNOR2_X1 U271 ( .A(n301), .B(n303), .ZN(SUM[22]) );
endmodule


module RCA_NBIT54 ( A, B, Ci, S, Co );
  input [53:0] A;
  input [53:0] B;
  output [53:0] S;
  input Ci;
  output Co;

  assign Co = 1'b0;

  RCA_NBIT54_DW01_add_0 add_95 ( .A(A), .B(B), .CI(1'b0), .SUM(S) );
endmodule


module RCA_NBIT56_DW01_add_0 ( A, B, CI, SUM, CO );
  input [55:0] A;
  input [55:0] B;
  output [55:0] SUM;
  input CI;
  output CO;
  wire   n1, n323, n324, n325, n327, n328, n329, n330, n331, n332, n333, n334,
         n336, n337, n338, n339, n342, n343, n344, n345, n346, n349, n353,
         n355, n357, n358, n359, n361, n363, n364, n381, n382, n384, n385,
         n389, n390, n393, n394, n395, n396, n397, n399, n400, n407, n409,
         n411, n412, n413, n414, n416, n417, net176815, net176817, net176832,
         net182459, net183541, net183568, net183810, net183849, net183848,
         net183944, net184510, net184607, net184677, net184755, net185233,
         net185313, net185701, net186076, net186098, net188923, net190463,
         net191609, net182755, net183811, net183222, net176825, n372, n391,
         n388, n387, n352, n348, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n326, n335, n340, n341, n347, n350, n351,
         n354, n356, n360, n362, n365, n366, n367, n368, n369, n370, n371,
         n373, n374, n375, n376, n377, n378, n379, n380, n383, n386, n392,
         n398, n401, n402, n403, n404, n405, n406, n408, n410, n415, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482;
  wire   [55:1] carry;
  assign net185701 = A[38];

  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(n417), .CO(carry[25]), .S(SUM[24])
         );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U143 ( .A(B[54]), .B(A[54]), .Z(n328) );
  XOR2_X1 U171 ( .A(n454), .B(n323), .Z(SUM[23]) );
  XOR2_X1 U172 ( .A(carry[22]), .B(n416), .Z(SUM[22]) );
  XOR2_X1 U173 ( .A(A[22]), .B(B[22]), .Z(n416) );
  XOR2_X1 U174 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U1 ( .A(n393), .Z(n427) );
  CLKBUF_X1 U2 ( .A(n370), .Z(n281) );
  CLKBUF_X1 U3 ( .A(A[42]), .Z(n279) );
  INV_X1 U4 ( .A(A[32]), .ZN(n280) );
  NOR2_X2 U5 ( .A1(net186098), .A2(n299), .ZN(n406) );
  CLKBUF_X1 U6 ( .A(A[23]), .Z(n282) );
  CLKBUF_X1 U7 ( .A(n432), .Z(n283) );
  OR2_X1 U8 ( .A1(n381), .A2(A[36]), .ZN(n382) );
  INV_X1 U9 ( .A(B[38]), .ZN(net183222) );
  BUF_X1 U10 ( .A(A[47]), .Z(net184677) );
  CLKBUF_X1 U11 ( .A(A[26]), .Z(n458) );
  CLKBUF_X1 U12 ( .A(A[44]), .Z(n423) );
  CLKBUF_X1 U13 ( .A(n408), .Z(n284) );
  CLKBUF_X1 U14 ( .A(A[40]), .Z(n285) );
  AND2_X1 U15 ( .A1(n477), .A2(n345), .ZN(n453) );
  AND2_X1 U16 ( .A1(n474), .A2(n374), .ZN(n286) );
  BUF_X1 U17 ( .A(A[28]), .Z(n403) );
  INV_X1 U18 ( .A(B[26]), .ZN(n425) );
  XNOR2_X1 U19 ( .A(n287), .B(n294), .ZN(SUM[30]) );
  XNOR2_X1 U20 ( .A(A[30]), .B(B[30]), .ZN(n287) );
  BUF_X1 U21 ( .A(A[50]), .Z(n305) );
  INV_X1 U22 ( .A(B[44]), .ZN(n446) );
  NAND2_X1 U23 ( .A1(n406), .A2(n279), .ZN(n288) );
  NAND2_X1 U24 ( .A1(n364), .A2(B[42]), .ZN(n289) );
  NAND2_X1 U25 ( .A1(n288), .A2(n289), .ZN(n290) );
  NAND2_X1 U26 ( .A1(n361), .A2(n291), .ZN(n358) );
  OR2_X1 U27 ( .A1(n479), .A2(n408), .ZN(n291) );
  BUF_X1 U28 ( .A(n402), .Z(n351) );
  INV_X1 U29 ( .A(net183810), .ZN(n292) );
  INV_X1 U30 ( .A(B[46]), .ZN(n302) );
  INV_X1 U31 ( .A(B[29]), .ZN(net183848) );
  XNOR2_X1 U32 ( .A(n293), .B(n426), .ZN(SUM[35]) );
  XNOR2_X1 U33 ( .A(A[35]), .B(B[35]), .ZN(n293) );
  INV_X1 U34 ( .A(B[50]), .ZN(n452) );
  INV_X1 U35 ( .A(B[34]), .ZN(net183944) );
  BUF_X1 U36 ( .A(n387), .Z(net185233) );
  INV_X1 U37 ( .A(B[48]), .ZN(n429) );
  OAI21_X1 U38 ( .B1(n290), .B2(A[43]), .A(B[43]), .ZN(n361) );
  AOI21_X1 U39 ( .B1(n470), .B2(n480), .A(n384), .ZN(n381) );
  NAND2_X1 U40 ( .A1(n294), .A2(A[30]), .ZN(n443) );
  INV_X1 U41 ( .A(n421), .ZN(n294) );
  XNOR2_X1 U42 ( .A(net182755), .B(n298), .ZN(SUM[41]) );
  AOI21_X1 U43 ( .B1(n430), .B2(n305), .A(B[50]), .ZN(n295) );
  CLKBUF_X1 U44 ( .A(A[46]), .Z(n296) );
  BUF_X1 U45 ( .A(A[27]), .Z(n404) );
  CLKBUF_X1 U46 ( .A(n390), .Z(n335) );
  AND2_X1 U47 ( .A1(n298), .A2(n312), .ZN(n299) );
  AOI21_X1 U48 ( .B1(n430), .B2(n305), .A(B[50]), .ZN(n297) );
  AND2_X1 U49 ( .A1(n311), .A2(n310), .ZN(n298) );
  CLKBUF_X1 U50 ( .A(A[51]), .Z(n419) );
  CLKBUF_X1 U51 ( .A(A[39]), .Z(n300) );
  BUF_X1 U52 ( .A(n381), .Z(n444) );
  XNOR2_X1 U53 ( .A(n301), .B(n348), .ZN(SUM[47]) );
  NOR2_X1 U54 ( .A1(n303), .A2(n352), .ZN(n348) );
  XNOR2_X1 U55 ( .A(A[47]), .B(B[47]), .ZN(n301) );
  NOR2_X1 U56 ( .A1(net184755), .A2(n296), .ZN(n303) );
  NOR2_X1 U57 ( .A1(n352), .A2(n303), .ZN(net183568) );
  AOI21_X1 U58 ( .B1(net184755), .B2(n296), .A(B[46]), .ZN(n352) );
  AOI21_X1 U59 ( .B1(net183568), .B2(net184677), .A(B[47]), .ZN(n349) );
  XNOR2_X1 U60 ( .A(A[46]), .B(n302), .ZN(n353) );
  OR2_X1 U61 ( .A1(A[39]), .A2(B[39]), .ZN(n304) );
  NAND2_X1 U62 ( .A1(n304), .A2(n314), .ZN(n308) );
  BUF_X1 U63 ( .A(A[37]), .Z(n354) );
  XNOR2_X1 U64 ( .A(n313), .B(n314), .ZN(SUM[39]) );
  BUF_X1 U65 ( .A(n336), .Z(n455) );
  INV_X1 U66 ( .A(n372), .ZN(n314) );
  NAND2_X1 U67 ( .A1(A[41]), .A2(n309), .ZN(n316) );
  INV_X1 U68 ( .A(A[41]), .ZN(n312) );
  NAND2_X1 U69 ( .A1(n307), .A2(n308), .ZN(n306) );
  NAND2_X1 U70 ( .A1(n317), .A2(n307), .ZN(net190463) );
  OAI21_X1 U71 ( .B1(n300), .B2(B[39]), .A(n314), .ZN(n317) );
  NAND2_X1 U72 ( .A1(net190463), .A2(n285), .ZN(n310) );
  OAI21_X1 U73 ( .B1(n306), .B2(A[40]), .A(B[40]), .ZN(n311) );
  XNOR2_X1 U74 ( .A(A[40]), .B(B[40]), .ZN(net182459) );
  INV_X1 U75 ( .A(B[41]), .ZN(n315) );
  XNOR2_X1 U76 ( .A(A[41]), .B(n315), .ZN(net182755) );
  XNOR2_X1 U77 ( .A(A[39]), .B(B[39]), .ZN(n313) );
  NAND2_X1 U78 ( .A1(B[39]), .A2(A[39]), .ZN(n307) );
  NAND2_X1 U79 ( .A1(n311), .A2(n310), .ZN(n309) );
  AND2_X1 U80 ( .A1(n316), .A2(n315), .ZN(net186098) );
  AND2_X1 U81 ( .A1(n316), .A2(n315), .ZN(n318) );
  NOR2_X1 U82 ( .A1(n318), .A2(n299), .ZN(n363) );
  NOR2_X1 U83 ( .A1(n456), .A2(n297), .ZN(n319) );
  OAI21_X1 U84 ( .B1(n321), .B2(A[34]), .A(B[34]), .ZN(n388) );
  OAI21_X1 U85 ( .B1(net185233), .B2(net183541), .A(n388), .ZN(n385) );
  INV_X1 U86 ( .A(n387), .ZN(n321) );
  OAI21_X1 U87 ( .B1(net188923), .B2(n321), .A(B[34]), .ZN(net185313) );
  BUF_X1 U88 ( .A(A[34]), .Z(net188923) );
  OAI21_X1 U89 ( .B1(n335), .B2(n326), .A(n320), .ZN(n387) );
  INV_X1 U90 ( .A(n391), .ZN(n320) );
  AOI21_X1 U91 ( .B1(n390), .B2(A[33]), .A(B[33]), .ZN(n391) );
  CLKBUF_X1 U92 ( .A(A[33]), .Z(n326) );
  XNOR2_X1 U93 ( .A(n322), .B(n335), .ZN(SUM[33]) );
  XNOR2_X1 U94 ( .A(A[33]), .B(B[33]), .ZN(n322) );
  OR2_X1 U95 ( .A1(n363), .A2(A[42]), .ZN(n340) );
  OR2_X1 U96 ( .A1(n363), .A2(A[42]), .ZN(n364) );
  AOI21_X1 U97 ( .B1(net183811), .B2(n347), .A(net176825), .ZN(n372) );
  AOI21_X1 U98 ( .B1(n350), .B2(net191609), .A(net183222), .ZN(net176825) );
  INV_X1 U99 ( .A(net185701), .ZN(n350) );
  CLKBUF_X1 U100 ( .A(net185701), .Z(n347) );
  INV_X1 U101 ( .A(net191609), .ZN(net183811) );
  XNOR2_X1 U102 ( .A(n341), .B(net183811), .ZN(SUM[38]) );
  XNOR2_X1 U103 ( .A(net185701), .B(B[38]), .ZN(n341) );
  BUF_X1 U104 ( .A(A[36]), .Z(n424) );
  CLKBUF_X1 U105 ( .A(n396), .Z(n438) );
  AOI22_X1 U106 ( .A1(n444), .A2(n424), .B1(n382), .B2(B[36]), .ZN(n356) );
  XNOR2_X1 U107 ( .A(n362), .B(n360), .ZN(SUM[37]) );
  NAND2_X1 U108 ( .A1(A[37]), .A2(B[37]), .ZN(n366) );
  OAI21_X1 U109 ( .B1(n354), .B2(B[37]), .A(n365), .ZN(net191609) );
  INV_X1 U110 ( .A(n354), .ZN(n360) );
  XNOR2_X1 U111 ( .A(net186076), .B(B[37]), .ZN(n362) );
  NAND2_X1 U112 ( .A1(n356), .A2(n366), .ZN(n365) );
  OR2_X1 U113 ( .A1(A[28]), .A2(B[28]), .ZN(n402) );
  AND2_X1 U114 ( .A1(n474), .A2(n374), .ZN(n367) );
  OAI21_X1 U115 ( .B1(n292), .B2(n404), .A(B[27]), .ZN(n368) );
  XNOR2_X1 U116 ( .A(n284), .B(n369), .ZN(SUM[43]) );
  XOR2_X1 U117 ( .A(A[43]), .B(B[43]), .Z(n369) );
  AOI21_X1 U118 ( .B1(n455), .B2(n419), .A(n468), .ZN(n370) );
  NAND2_X1 U119 ( .A1(n351), .A2(n392), .ZN(n371) );
  AND2_X1 U120 ( .A1(n368), .A2(n401), .ZN(n373) );
  OR2_X1 U121 ( .A1(B[25]), .A2(A[25]), .ZN(n374) );
  NAND2_X1 U122 ( .A1(n474), .A2(n374), .ZN(n412) );
  AOI21_X1 U123 ( .B1(n460), .B2(n437), .A(B[48]), .ZN(n375) );
  NOR2_X1 U124 ( .A1(n453), .A2(n375), .ZN(n376) );
  NAND2_X1 U125 ( .A1(n403), .A2(B[28]), .ZN(n378) );
  INV_X1 U126 ( .A(A[28]), .ZN(n383) );
  OAI21_X1 U127 ( .B1(n292), .B2(n404), .A(B[27]), .ZN(n398) );
  XNOR2_X1 U128 ( .A(n292), .B(n386), .ZN(SUM[27]) );
  NAND2_X1 U129 ( .A1(n398), .A2(n401), .ZN(n392) );
  NAND2_X1 U130 ( .A1(A[29]), .A2(n377), .ZN(n380) );
  NAND2_X1 U131 ( .A1(n380), .A2(net183848), .ZN(net176817) );
  XNOR2_X1 U132 ( .A(A[27]), .B(B[27]), .ZN(n386) );
  NAND2_X1 U133 ( .A1(n404), .A2(net176815), .ZN(n401) );
  XNOR2_X1 U134 ( .A(A[29]), .B(B[29]), .ZN(net183849) );
  NAND2_X1 U135 ( .A1(n402), .A2(n392), .ZN(n379) );
  NAND2_X1 U136 ( .A1(n379), .A2(n378), .ZN(n377) );
  NAND2_X1 U137 ( .A1(n371), .A2(n378), .ZN(n405) );
  NAND2_X1 U138 ( .A1(n371), .A2(n378), .ZN(net184607) );
  XNOR2_X1 U139 ( .A(n383), .B(B[28]), .ZN(n407) );
  CLKBUF_X1 U140 ( .A(A[29]), .Z(net184510) );
  AOI22_X1 U141 ( .A1(n406), .A2(n279), .B1(n340), .B2(B[42]), .ZN(n408) );
  BUF_X1 U142 ( .A(n358), .Z(n415) );
  AOI21_X1 U144 ( .B1(n415), .B2(n423), .A(B[44]), .ZN(n410) );
  NOR2_X1 U145 ( .A1(n453), .A2(n346), .ZN(n342) );
  NOR2_X1 U146 ( .A1(n410), .A2(n435), .ZN(n418) );
  AOI22_X1 U147 ( .A1(n444), .A2(n424), .B1(n382), .B2(B[36]), .ZN(net186076)
         );
  CLKBUF_X1 U148 ( .A(A[53]), .Z(n447) );
  CLKBUF_X1 U149 ( .A(A[31]), .Z(n420) );
  OAI21_X1 U150 ( .B1(net184510), .B2(net184607), .A(net176817), .ZN(n421) );
  NOR2_X1 U151 ( .A1(n357), .A2(n435), .ZN(n422) );
  XNOR2_X1 U152 ( .A(n448), .B(n345), .ZN(SUM[48]) );
  XNOR2_X1 U153 ( .A(A[26]), .B(n425), .ZN(n413) );
  OAI21_X1 U154 ( .B1(net185233), .B2(net183541), .A(net185313), .ZN(n426) );
  AOI21_X1 U155 ( .B1(n455), .B2(n419), .A(n468), .ZN(n333) );
  AND2_X1 U156 ( .A1(n451), .A2(n450), .ZN(n428) );
  BUF_X1 U157 ( .A(A[45]), .Z(n432) );
  XNOR2_X1 U158 ( .A(A[48]), .B(n429), .ZN(n448) );
  OR2_X1 U159 ( .A1(n469), .A2(n441), .ZN(n430) );
  BUF_X1 U160 ( .A(A[49]), .Z(n431) );
  CLKBUF_X1 U161 ( .A(n434), .Z(n433) );
  OR2_X1 U162 ( .A1(n466), .A2(n440), .ZN(n434) );
  AND2_X1 U163 ( .A1(n436), .A2(n478), .ZN(n435) );
  INV_X1 U164 ( .A(n358), .ZN(n436) );
  AND2_X1 U165 ( .A1(net176832), .A2(n449), .ZN(n437) );
  NOR2_X1 U166 ( .A1(n440), .A2(n466), .ZN(n329) );
  NAND2_X1 U167 ( .A1(n451), .A2(n450), .ZN(net184755) );
  NOR2_X1 U168 ( .A1(n469), .A2(n441), .ZN(n339) );
  INV_X1 U169 ( .A(n475), .ZN(n439) );
  AND2_X1 U170 ( .A1(n330), .A2(n447), .ZN(n440) );
  AND2_X1 U175 ( .A1(n376), .A2(n431), .ZN(n441) );
  XNOR2_X1 U176 ( .A(n325), .B(n442), .ZN(SUM[55]) );
  XOR2_X1 U177 ( .A(B[55]), .B(A[55]), .Z(n442) );
  NAND2_X1 U178 ( .A1(n443), .A2(n400), .ZN(n396) );
  XNOR2_X1 U179 ( .A(A[34]), .B(net183944), .ZN(n389) );
  XNOR2_X1 U180 ( .A(net183849), .B(n405), .ZN(SUM[29]) );
  OAI22_X1 U181 ( .A1(n458), .A2(n286), .B1(n411), .B2(B[26]), .ZN(net183810)
         );
  XNOR2_X1 U182 ( .A(n370), .B(n445), .ZN(SUM[52]) );
  XOR2_X1 U183 ( .A(A[52]), .B(B[52]), .Z(n445) );
  XNOR2_X1 U184 ( .A(A[44]), .B(n446), .ZN(n359) );
  INV_X1 U185 ( .A(net188923), .ZN(net183541) );
  OR2_X1 U186 ( .A1(net184677), .A2(net183568), .ZN(n449) );
  NAND2_X1 U187 ( .A1(net176832), .A2(n449), .ZN(n345) );
  NAND2_X1 U188 ( .A1(n422), .A2(n283), .ZN(n450) );
  NAND2_X1 U189 ( .A1(n355), .A2(B[45]), .ZN(n451) );
  XNOR2_X1 U190 ( .A(A[50]), .B(n452), .ZN(n457) );
  CLKBUF_X1 U191 ( .A(n324), .Z(n454) );
  AND2_X1 U192 ( .A1(n339), .A2(n476), .ZN(n456) );
  NOR2_X1 U193 ( .A1(n295), .A2(n456), .ZN(n336) );
  XNOR2_X1 U194 ( .A(n330), .B(n332), .ZN(SUM[53]) );
  XNOR2_X1 U195 ( .A(n457), .B(n339), .ZN(SUM[50]) );
  XNOR2_X1 U196 ( .A(n338), .B(n336), .ZN(SUM[51]) );
  XNOR2_X1 U197 ( .A(n329), .B(n328), .ZN(SUM[54]) );
  XNOR2_X1 U198 ( .A(n438), .B(n459), .ZN(SUM[31]) );
  XNOR2_X1 U199 ( .A(A[31]), .B(B[31]), .ZN(n459) );
  INV_X1 U200 ( .A(n477), .ZN(n460) );
  INV_X1 U201 ( .A(A[44]), .ZN(n478) );
  INV_X1 U202 ( .A(n426), .ZN(n470) );
  INV_X1 U203 ( .A(n397), .ZN(n472) );
  XNOR2_X1 U204 ( .A(n422), .B(n461), .ZN(SUM[45]) );
  XNOR2_X1 U205 ( .A(A[45]), .B(B[45]), .ZN(n461) );
  INV_X1 U206 ( .A(n409), .ZN(net176815) );
  XNOR2_X1 U207 ( .A(A[49]), .B(B[49]), .ZN(n344) );
  XNOR2_X1 U208 ( .A(n462), .B(n406), .ZN(SUM[42]) );
  XNOR2_X1 U209 ( .A(A[42]), .B(B[42]), .ZN(n462) );
  XNOR2_X1 U210 ( .A(net182459), .B(net190463), .ZN(SUM[40]) );
  XNOR2_X1 U211 ( .A(n444), .B(n463), .ZN(SUM[36]) );
  XNOR2_X1 U212 ( .A(A[36]), .B(B[36]), .ZN(n463) );
  AOI21_X1 U213 ( .B1(n467), .B2(n439), .A(B[52]), .ZN(n334) );
  AOI21_X1 U214 ( .B1(n415), .B2(n423), .A(B[44]), .ZN(n357) );
  OAI21_X1 U215 ( .B1(n427), .B2(n280), .A(n394), .ZN(n390) );
  INV_X1 U216 ( .A(n393), .ZN(n471) );
  INV_X1 U217 ( .A(n399), .ZN(n473) );
  INV_X1 U218 ( .A(A[50]), .ZN(n476) );
  INV_X1 U219 ( .A(A[52]), .ZN(n475) );
  INV_X1 U220 ( .A(A[48]), .ZN(n477) );
  INV_X1 U221 ( .A(n327), .ZN(n465) );
  INV_X1 U222 ( .A(n337), .ZN(n468) );
  INV_X1 U223 ( .A(B[23]), .ZN(n482) );
  XNOR2_X1 U224 ( .A(n464), .B(A[25]), .ZN(SUM[25]) );
  XNOR2_X1 U225 ( .A(carry[25]), .B(B[25]), .ZN(n464) );
  INV_X1 U226 ( .A(n414), .ZN(n474) );
  AOI22_X1 U227 ( .A1(B[22]), .A2(A[22]), .B1(n416), .B2(carry[22]), .ZN(n323)
         );
  AND2_X1 U228 ( .A1(A[0]), .A2(B[0]), .ZN(n1) );
  XNOR2_X1 U229 ( .A(A[51]), .B(B[51]), .ZN(n338) );
  OAI21_X1 U230 ( .B1(n319), .B2(A[51]), .A(B[51]), .ZN(n337) );
  OAI21_X1 U231 ( .B1(A[54]), .B2(n433), .A(n465), .ZN(n325) );
  AOI21_X1 U232 ( .B1(n434), .B2(A[54]), .A(B[54]), .ZN(n327) );
  XNOR2_X1 U233 ( .A(A[53]), .B(B[53]), .ZN(n332) );
  INV_X1 U234 ( .A(n343), .ZN(n469) );
  AOI21_X1 U235 ( .B1(n437), .B2(n460), .A(B[48]), .ZN(n346) );
  XNOR2_X1 U236 ( .A(n280), .B(B[32]), .ZN(n395) );
  XNOR2_X1 U237 ( .A(n359), .B(n436), .ZN(SUM[44]) );
  XNOR2_X1 U238 ( .A(n395), .B(n427), .ZN(SUM[32]) );
  INV_X1 U239 ( .A(n349), .ZN(net176832) );
  XNOR2_X1 U240 ( .A(n407), .B(n373), .ZN(SUM[28]) );
  OAI21_X1 U241 ( .B1(net184510), .B2(net184607), .A(net176817), .ZN(n399) );
  AOI21_X1 U242 ( .B1(A[25]), .B2(B[25]), .A(carry[25]), .ZN(n414) );
  INV_X1 U243 ( .A(A[43]), .ZN(n479) );
  OAI21_X1 U244 ( .B1(n473), .B2(A[30]), .A(B[30]), .ZN(n400) );
  OAI22_X1 U245 ( .A1(n458), .A2(n286), .B1(B[26]), .B2(n411), .ZN(n409) );
  AND2_X1 U246 ( .A1(A[26]), .A2(n367), .ZN(n411) );
  OAI22_X1 U247 ( .A1(n482), .A2(n481), .B1(n323), .B2(n324), .ZN(n417) );
  AOI21_X1 U248 ( .B1(n385), .B2(A[35]), .A(B[35]), .ZN(n384) );
  INV_X1 U249 ( .A(A[35]), .ZN(n480) );
  XNOR2_X1 U250 ( .A(n389), .B(net185233), .ZN(SUM[34]) );
  OAI21_X1 U251 ( .B1(n471), .B2(A[32]), .A(B[32]), .ZN(n394) );
  AOI21_X1 U252 ( .B1(n281), .B2(n475), .A(n334), .ZN(n330) );
  INV_X1 U253 ( .A(n333), .ZN(n467) );
  OR2_X1 U254 ( .A1(n418), .A2(n432), .ZN(n355) );
  OAI21_X1 U255 ( .B1(n438), .B2(n420), .A(n472), .ZN(n393) );
  AOI21_X1 U256 ( .B1(n396), .B2(A[31]), .A(B[31]), .ZN(n397) );
  INV_X1 U257 ( .A(n282), .ZN(n481) );
  XNOR2_X1 U258 ( .A(A[23]), .B(B[23]), .ZN(n324) );
  INV_X1 U259 ( .A(n331), .ZN(n466) );
  OAI21_X1 U260 ( .B1(n330), .B2(n447), .A(B[53]), .ZN(n331) );
  XNOR2_X1 U261 ( .A(n376), .B(n344), .ZN(SUM[49]) );
  OAI21_X1 U262 ( .B1(n342), .B2(n431), .A(B[49]), .ZN(n343) );
  XNOR2_X1 U263 ( .A(n412), .B(n413), .ZN(SUM[26]) );
  XNOR2_X1 U264 ( .A(n428), .B(n353), .ZN(SUM[46]) );
endmodule


module RCA_NBIT56 ( A, B, Ci, S, Co );
  input [55:0] A;
  input [55:0] B;
  output [55:0] S;
  input Ci;
  output Co;

  assign Co = 1'b0;

  RCA_NBIT56_DW01_add_0 add_95 ( .A(A), .B(B), .CI(1'b0), .SUM(S) );
endmodule


module RCA_NBIT58_DW01_add_0 ( A, B, CI, SUM, CO );
  input [57:0] A;
  input [57:0] B;
  output [57:0] SUM;
  input CI;
  output CO;
  wire   n1, n242, n243, n246, n247, n248, n249, n250, n253, n255, n256, n258,
         n259, n261, n262, n264, n265, n268, n273, n274, n280, n309, n310,
         n320, n321, n324, n325, n326, n327, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, net176843, net176879, net183764, net183763,
         net183827, net183852, net184130, net184494, net184498, net184761,
         net185518, net185538, net185975, net176867, net185857, net191668,
         net191778, net185534, net176848, n279, net193281, n322, n319, n316,
         n315, n313, net182868, net176874, net176873, n284, n283, n282,
         net193299, net186765, net184493, n302, n300, net194076, net194068,
         net193440, net184127, net184089, net183952, net183417, net182384,
         net180710, n292, n289, n285, net197767, net183604, n301, n271, n270,
         n267, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545;
  wire   [57:1] carry;
  assign net193299 = A[37];

  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U174 ( .A(A[27]), .B(B[27]), .Z(n329) );
  XOR2_X1 U175 ( .A(A[26]), .B(B[26]), .Z(n332) );
  XOR2_X1 U176 ( .A(B[25]), .B(n514), .Z(n335) );
  XOR2_X1 U177 ( .A(A[24]), .B(n337), .Z(SUM[24]) );
  XOR2_X1 U178 ( .A(carry[24]), .B(B[24]), .Z(n337) );
  XOR2_X1 U179 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  CLKBUF_X1 U1 ( .A(A[29]), .Z(n385) );
  CLKBUF_X1 U2 ( .A(n536), .Z(n492) );
  OAI21_X1 U3 ( .B1(n431), .B2(n490), .A(B[54]), .ZN(n386) );
  CLKBUF_X1 U4 ( .A(n282), .Z(net182868) );
  AND2_X1 U5 ( .A1(n396), .A2(n395), .ZN(n387) );
  CLKBUF_X1 U6 ( .A(A[42]), .Z(net185534) );
  OR2_X1 U7 ( .A1(n529), .A2(n531), .ZN(n388) );
  CLKBUF_X1 U8 ( .A(n315), .Z(n457) );
  BUF_X1 U9 ( .A(n315), .Z(n453) );
  BUF_X1 U10 ( .A(A[27]), .Z(n498) );
  OR2_X2 U11 ( .A1(n532), .A2(n528), .ZN(n489) );
  CLKBUF_X1 U12 ( .A(n321), .Z(n389) );
  OR2_X1 U13 ( .A1(n529), .A2(n531), .ZN(n431) );
  INV_X1 U14 ( .A(B[38]), .ZN(n437) );
  NAND2_X1 U15 ( .A1(A[26]), .A2(n492), .ZN(n395) );
  OR2_X1 U16 ( .A1(net176843), .A2(n407), .ZN(net191668) );
  AND2_X1 U17 ( .A1(n280), .A2(net184761), .ZN(n475) );
  AND3_X1 U18 ( .A1(n421), .A2(n439), .A3(n442), .ZN(n390) );
  INV_X1 U19 ( .A(B[35]), .ZN(net183763) );
  BUF_X1 U20 ( .A(net185518), .Z(n391) );
  CLKBUF_X1 U21 ( .A(A[30]), .Z(n392) );
  BUF_X1 U22 ( .A(A[53]), .Z(n480) );
  OR2_X1 U23 ( .A1(n403), .A2(n540), .ZN(n393) );
  NAND2_X1 U24 ( .A1(n393), .A2(n242), .ZN(carry[56]) );
  INV_X1 U25 ( .A(B[30]), .ZN(n448) );
  INV_X1 U26 ( .A(B[46]), .ZN(n414) );
  INV_X1 U27 ( .A(B[41]), .ZN(net183952) );
  INV_X1 U28 ( .A(B[48]), .ZN(n473) );
  INV_X1 U29 ( .A(B[50]), .ZN(n519) );
  INV_X1 U30 ( .A(B[42]), .ZN(n444) );
  INV_X1 U31 ( .A(B[44]), .ZN(n523) );
  INV_X1 U32 ( .A(B[36]), .ZN(n423) );
  INV_X1 U33 ( .A(B[40]), .ZN(n429) );
  BUF_X1 U34 ( .A(A[32]), .Z(n449) );
  NAND2_X1 U35 ( .A1(B[26]), .A2(n330), .ZN(n396) );
  BUF_X1 U36 ( .A(A[43]), .Z(n460) );
  NAND2_X1 U37 ( .A1(n396), .A2(n395), .ZN(n394) );
  XNOR2_X1 U38 ( .A(A[33]), .B(B[33]), .ZN(n497) );
  CLKBUF_X1 U39 ( .A(A[34]), .Z(n430) );
  INV_X1 U40 ( .A(B[32]), .ZN(n455) );
  INV_X1 U41 ( .A(B[54]), .ZN(n496) );
  INV_X1 U42 ( .A(B[28]), .ZN(n499) );
  XNOR2_X1 U43 ( .A(n248), .B(n246), .ZN(SUM[54]) );
  AOI21_X1 U44 ( .B1(n397), .B2(n398), .A(net183952), .ZN(net176873) );
  INV_X1 U45 ( .A(n285), .ZN(n397) );
  INV_X1 U46 ( .A(A[41]), .ZN(n398) );
  XNOR2_X1 U47 ( .A(n441), .B(n440), .ZN(SUM[38]) );
  OAI21_X1 U48 ( .B1(B[34]), .B2(A[34]), .A(net183852), .ZN(n468) );
  AOI21_X1 U49 ( .B1(n264), .B2(n543), .A(n473), .ZN(n399) );
  INV_X1 U50 ( .A(n399), .ZN(n265) );
  OR2_X2 U51 ( .A1(net176867), .A2(net193281), .ZN(net184493) );
  BUF_X1 U52 ( .A(n285), .Z(net184127) );
  OAI21_X1 U53 ( .B1(net176874), .B2(net185534), .A(B[42]), .ZN(n400) );
  OAI21_X1 U54 ( .B1(n452), .B2(n449), .A(B[32]), .ZN(n401) );
  OAI21_X1 U55 ( .B1(net176848), .B2(n428), .A(n400), .ZN(n402) );
  AND2_X1 U56 ( .A1(n247), .A2(n522), .ZN(n403) );
  BUF_X1 U57 ( .A(n530), .Z(n404) );
  BUF_X1 U58 ( .A(A[45]), .Z(n491) );
  BUF_X1 U59 ( .A(A[47]), .Z(n412) );
  OR2_X1 U60 ( .A1(n544), .A2(n475), .ZN(n405) );
  NAND2_X1 U61 ( .A1(n405), .A2(n463), .ZN(n273) );
  OAI21_X1 U62 ( .B1(n402), .B2(n460), .A(B[43]), .ZN(n406) );
  AOI21_X1 U63 ( .B1(n453), .B2(n450), .A(n447), .ZN(n407) );
  XNOR2_X1 U64 ( .A(n413), .B(n410), .ZN(SUM[47]) );
  BUF_X1 U65 ( .A(n267), .Z(n410) );
  AND2_X1 U66 ( .A1(n410), .A2(A[47]), .ZN(net197767) );
  AOI21_X1 U67 ( .B1(n410), .B2(n412), .A(net176879), .ZN(net185518) );
  NOR2_X1 U68 ( .A1(n415), .A2(n416), .ZN(n413) );
  NOR2_X1 U69 ( .A1(n412), .A2(n409), .ZN(n416) );
  INV_X1 U70 ( .A(B[47]), .ZN(n409) );
  AND2_X1 U71 ( .A1(A[47]), .A2(n409), .ZN(n415) );
  OAI21_X1 U72 ( .B1(n270), .B2(n408), .A(n271), .ZN(n267) );
  OAI21_X1 U73 ( .B1(A[47]), .B2(n267), .A(B[47]), .ZN(n268) );
  OAI21_X1 U74 ( .B1(net184498), .B2(A[46]), .A(B[46]), .ZN(n271) );
  INV_X1 U75 ( .A(A[46]), .ZN(n408) );
  INV_X1 U76 ( .A(net184498), .ZN(n270) );
  XNOR2_X1 U77 ( .A(n270), .B(n411), .ZN(SUM[46]) );
  XNOR2_X1 U78 ( .A(A[46]), .B(n414), .ZN(n411) );
  CLKBUF_X1 U79 ( .A(A[33]), .Z(n417) );
  OAI21_X1 U80 ( .B1(n390), .B2(n437), .A(n438), .ZN(n418) );
  BUF_X1 U81 ( .A(net193299), .Z(net194076) );
  OAI21_X1 U82 ( .B1(n390), .B2(n437), .A(n438), .ZN(net185857) );
  NOR2_X1 U83 ( .A1(n458), .A2(n446), .ZN(n419) );
  NAND2_X1 U84 ( .A1(n322), .A2(n420), .ZN(n456) );
  NAND2_X1 U85 ( .A1(net184130), .A2(n385), .ZN(n420) );
  OAI21_X1 U86 ( .B1(n426), .B2(net194076), .A(B[37]), .ZN(n421) );
  XNOR2_X1 U87 ( .A(net183604), .B(n426), .ZN(SUM[37]) );
  XNOR2_X1 U88 ( .A(net193299), .B(B[37]), .ZN(net183604) );
  NAND2_X1 U89 ( .A1(n424), .A2(n427), .ZN(n426) );
  OAI21_X1 U90 ( .B1(net194076), .B2(n426), .A(B[37]), .ZN(net194068) );
  OAI21_X1 U91 ( .B1(net184493), .B2(n425), .A(B[36]), .ZN(n301) );
  INV_X1 U92 ( .A(n422), .ZN(n425) );
  OAI21_X1 U93 ( .B1(net184493), .B2(n425), .A(B[36]), .ZN(n427) );
  INV_X1 U94 ( .A(A[36]), .ZN(n422) );
  OR2_X1 U95 ( .A1(n300), .A2(n422), .ZN(n424) );
  NAND2_X1 U96 ( .A1(n301), .A2(n424), .ZN(net186765) );
  XNOR2_X1 U97 ( .A(A[36]), .B(n423), .ZN(n302) );
  NOR2_X1 U98 ( .A1(net197767), .A2(net176879), .ZN(n264) );
  INV_X1 U99 ( .A(net176874), .ZN(n428) );
  XNOR2_X1 U100 ( .A(A[40]), .B(n429), .ZN(n434) );
  XNOR2_X1 U101 ( .A(net184089), .B(net184127), .ZN(SUM[41]) );
  XNOR2_X1 U102 ( .A(A[41]), .B(B[41]), .ZN(net184089) );
  AOI21_X1 U103 ( .B1(net184127), .B2(net183417), .A(net176873), .ZN(n282) );
  CLKBUF_X1 U104 ( .A(A[41]), .Z(net183417) );
  OAI21_X1 U105 ( .B1(n433), .B2(n432), .A(n289), .ZN(n285) );
  OAI21_X1 U106 ( .B1(net180710), .B2(A[40]), .A(B[40]), .ZN(n289) );
  NAND2_X1 U107 ( .A1(n435), .A2(net182384), .ZN(net180710) );
  OAI21_X1 U108 ( .B1(n418), .B2(net193440), .A(B[39]), .ZN(n435) );
  BUF_X1 U109 ( .A(A[39]), .Z(net193440) );
  OAI21_X1 U110 ( .B1(net193440), .B2(net185857), .A(B[39]), .ZN(n292) );
  NAND2_X1 U111 ( .A1(n418), .A2(net193440), .ZN(net182384) );
  INV_X1 U112 ( .A(A[40]), .ZN(n432) );
  XNOR2_X1 U113 ( .A(n434), .B(n433), .ZN(SUM[40]) );
  AND2_X1 U114 ( .A1(n292), .A2(net182384), .ZN(n433) );
  XNOR2_X1 U115 ( .A(n436), .B(net185857), .ZN(SUM[39]) );
  XNOR2_X1 U116 ( .A(A[39]), .B(B[39]), .ZN(n436) );
  XNOR2_X1 U117 ( .A(A[38]), .B(B[38]), .ZN(n440) );
  NAND2_X1 U118 ( .A1(n441), .A2(n443), .ZN(n438) );
  INV_X1 U119 ( .A(A[38]), .ZN(n439) );
  NAND2_X1 U120 ( .A1(net194076), .A2(net186765), .ZN(n442) );
  NAND2_X1 U121 ( .A1(net194068), .A2(n442), .ZN(n441) );
  INV_X1 U122 ( .A(n439), .ZN(n443) );
  NOR2_X1 U123 ( .A1(net193281), .A2(net176867), .ZN(n300) );
  XNOR2_X1 U124 ( .A(n302), .B(n300), .ZN(SUM[36]) );
  XNOR2_X1 U125 ( .A(n284), .B(net182868), .ZN(SUM[42]) );
  XNOR2_X1 U126 ( .A(A[42]), .B(n444), .ZN(n284) );
  OAI21_X1 U127 ( .B1(net176848), .B2(n428), .A(n283), .ZN(n279) );
  OAI21_X1 U128 ( .B1(net176874), .B2(net185534), .A(B[42]), .ZN(n283) );
  INV_X1 U129 ( .A(n282), .ZN(net176874) );
  OAI21_X1 U130 ( .B1(n452), .B2(n449), .A(B[32]), .ZN(n313) );
  NAND2_X1 U131 ( .A1(n401), .A2(net191668), .ZN(n309) );
  NAND2_X1 U132 ( .A1(net191668), .A2(n313), .ZN(net191778) );
  INV_X1 U133 ( .A(n449), .ZN(net176843) );
  OR2_X1 U134 ( .A1(n447), .A2(n451), .ZN(n452) );
  AND2_X1 U135 ( .A1(n453), .A2(n450), .ZN(n451) );
  CLKBUF_X1 U136 ( .A(A[31]), .Z(n450) );
  INV_X1 U137 ( .A(n316), .ZN(n447) );
  OAI21_X1 U138 ( .B1(n315), .B2(A[31]), .A(B[31]), .ZN(n316) );
  XNOR2_X1 U139 ( .A(A[32]), .B(n455), .ZN(net185538) );
  XNOR2_X1 U140 ( .A(A[31]), .B(B[31]), .ZN(net183827) );
  NAND2_X1 U141 ( .A1(n454), .A2(n319), .ZN(n315) );
  OAI21_X1 U142 ( .B1(n456), .B2(n392), .A(B[30]), .ZN(n319) );
  AND2_X1 U143 ( .A1(n389), .A2(n385), .ZN(n458) );
  OAI21_X1 U144 ( .B1(n321), .B2(A[29]), .A(B[29]), .ZN(n322) );
  INV_X1 U145 ( .A(n322), .ZN(n446) );
  NOR2_X1 U146 ( .A1(n446), .A2(n458), .ZN(net185975) );
  OR2_X1 U147 ( .A1(net185975), .A2(n445), .ZN(n454) );
  INV_X1 U148 ( .A(A[30]), .ZN(n445) );
  XNOR2_X1 U149 ( .A(A[30]), .B(n448), .ZN(n320) );
  BUF_X1 U150 ( .A(net184494), .Z(n462) );
  OR2_X1 U151 ( .A1(n479), .A2(n545), .ZN(n459) );
  NAND2_X1 U152 ( .A1(n325), .A2(n459), .ZN(n321) );
  AND2_X1 U153 ( .A1(A[35]), .A2(net184494), .ZN(net193281) );
  BUF_X1 U154 ( .A(n321), .Z(net184130) );
  XNOR2_X1 U155 ( .A(n279), .B(n461), .ZN(SUM[43]) );
  XNOR2_X1 U156 ( .A(A[43]), .B(B[43]), .ZN(n461) );
  OAI21_X1 U157 ( .B1(n402), .B2(n460), .A(B[43]), .ZN(n280) );
  NAND2_X1 U158 ( .A1(n279), .A2(n460), .ZN(net184761) );
  INV_X1 U159 ( .A(net185534), .ZN(net176848) );
  OAI21_X1 U160 ( .B1(n477), .B2(A[44]), .A(B[44]), .ZN(n463) );
  NAND2_X1 U161 ( .A1(n465), .A2(n521), .ZN(n464) );
  OAI21_X1 U162 ( .B1(n489), .B2(n510), .A(B[52]), .ZN(n465) );
  OR2_X1 U163 ( .A1(net185518), .A2(n543), .ZN(n466) );
  NAND2_X1 U164 ( .A1(n265), .A2(n466), .ZN(n261) );
  XNOR2_X1 U165 ( .A(A[34]), .B(B[34]), .ZN(n470) );
  NAND2_X1 U166 ( .A1(n430), .A2(B[34]), .ZN(n467) );
  XNOR2_X1 U167 ( .A(A[35]), .B(B[35]), .ZN(net183764) );
  INV_X1 U168 ( .A(A[35]), .ZN(n469) );
  NAND2_X1 U169 ( .A1(n468), .A2(n467), .ZN(net184494) );
  AOI21_X1 U170 ( .B1(n469), .B2(n471), .A(net183763), .ZN(net176867) );
  AND2_X1 U171 ( .A1(n468), .A2(n467), .ZN(n471) );
  XNOR2_X1 U172 ( .A(n470), .B(net183852), .ZN(SUM[34]) );
  OAI21_X1 U173 ( .B1(n544), .B2(n475), .A(n463), .ZN(n472) );
  XNOR2_X1 U180 ( .A(A[48]), .B(n473), .ZN(n507) );
  CLKBUF_X1 U181 ( .A(A[25]), .Z(n502) );
  OAI21_X1 U182 ( .B1(n511), .B2(n533), .A(B[50]), .ZN(n474) );
  XNOR2_X1 U183 ( .A(n530), .B(n476), .ZN(SUM[49]) );
  XNOR2_X1 U184 ( .A(B[49]), .B(A[49]), .ZN(n476) );
  BUF_X1 U185 ( .A(A[51]), .Z(n508) );
  NAND2_X1 U186 ( .A1(n406), .A2(net184761), .ZN(n477) );
  OR2_X1 U187 ( .A1(n394), .A2(A[27]), .ZN(n478) );
  AOI22_X1 U188 ( .A1(n520), .A2(n498), .B1(n478), .B2(B[27]), .ZN(n479) );
  NAND2_X1 U189 ( .A1(n488), .A2(n474), .ZN(n481) );
  XNOR2_X1 U190 ( .A(carry[57]), .B(B[57]), .ZN(n482) );
  XNOR2_X1 U191 ( .A(n482), .B(A[57]), .ZN(SUM[57]) );
  BUF_X1 U192 ( .A(n261), .Z(n530) );
  INV_X1 U193 ( .A(n487), .ZN(n483) );
  XNOR2_X1 U194 ( .A(net185538), .B(n407), .ZN(SUM[32]) );
  OAI21_X1 U195 ( .B1(n388), .B2(n490), .A(B[54]), .ZN(n484) );
  NAND2_X1 U196 ( .A1(n484), .A2(n522), .ZN(n485) );
  CLKBUF_X1 U197 ( .A(A[49]), .Z(n486) );
  CLKBUF_X1 U198 ( .A(n537), .Z(n487) );
  OR2_X1 U199 ( .A1(n515), .A2(n542), .ZN(n488) );
  NAND2_X1 U200 ( .A1(n259), .A2(n488), .ZN(n255) );
  INV_X1 U201 ( .A(n539), .ZN(n490) );
  NAND2_X1 U202 ( .A1(n274), .A2(n505), .ZN(net184498) );
  XNOR2_X1 U203 ( .A(n493), .B(n481), .ZN(SUM[51]) );
  XNOR2_X1 U204 ( .A(A[51]), .B(B[51]), .ZN(n493) );
  NOR2_X1 U205 ( .A1(n529), .A2(n531), .ZN(n494) );
  NOR2_X1 U206 ( .A1(n529), .A2(n531), .ZN(n246) );
  INV_X1 U207 ( .A(n492), .ZN(n495) );
  XNOR2_X1 U208 ( .A(A[54]), .B(n496), .ZN(n248) );
  XNOR2_X1 U209 ( .A(net191778), .B(n497), .ZN(SUM[33]) );
  XNOR2_X1 U210 ( .A(A[28]), .B(n499), .ZN(n326) );
  NOR2_X1 U211 ( .A1(n532), .A2(n528), .ZN(n500) );
  NOR2_X1 U212 ( .A1(n528), .A2(n532), .ZN(n501) );
  XNOR2_X1 U213 ( .A(n464), .B(n503), .ZN(SUM[53]) );
  XNOR2_X1 U214 ( .A(A[53]), .B(B[53]), .ZN(n503) );
  NAND2_X1 U215 ( .A1(n310), .A2(n504), .ZN(net183852) );
  NAND2_X1 U216 ( .A1(net191778), .A2(n417), .ZN(n504) );
  NAND2_X1 U217 ( .A1(n472), .A2(n491), .ZN(n505) );
  XNOR2_X1 U218 ( .A(carry[56]), .B(n506), .ZN(SUM[56]) );
  XNOR2_X1 U219 ( .A(A[56]), .B(B[56]), .ZN(n506) );
  XNOR2_X1 U220 ( .A(n507), .B(n391), .ZN(SUM[48]) );
  XNOR2_X1 U221 ( .A(n457), .B(net183827), .ZN(SUM[31]) );
  XNOR2_X1 U222 ( .A(net183764), .B(n462), .ZN(SUM[35]) );
  XNOR2_X1 U223 ( .A(n500), .B(n509), .ZN(SUM[52]) );
  XOR2_X1 U224 ( .A(A[52]), .B(B[52]), .Z(n509) );
  INV_X1 U225 ( .A(n541), .ZN(n510) );
  INV_X1 U226 ( .A(n542), .ZN(n511) );
  XNOR2_X1 U227 ( .A(n512), .B(n243), .ZN(SUM[55]) );
  XNOR2_X1 U228 ( .A(A[55]), .B(B[55]), .ZN(n512) );
  XNOR2_X1 U229 ( .A(net184130), .B(n513), .ZN(SUM[29]) );
  XNOR2_X1 U230 ( .A(A[29]), .B(B[29]), .ZN(n513) );
  CLKBUF_X1 U231 ( .A(n502), .Z(n514) );
  AOI21_X1 U232 ( .B1(n404), .B2(n486), .A(n534), .ZN(n515) );
  AOI21_X1 U233 ( .B1(n404), .B2(n486), .A(n534), .ZN(n258) );
  NAND2_X1 U234 ( .A1(carry[56]), .A2(A[56]), .ZN(n516) );
  NAND2_X1 U235 ( .A1(carry[56]), .A2(B[56]), .ZN(n517) );
  NAND2_X1 U236 ( .A1(A[56]), .A2(B[56]), .ZN(n518) );
  NAND3_X1 U237 ( .A1(n517), .A2(n516), .A3(n518), .ZN(carry[57]) );
  XNOR2_X1 U238 ( .A(A[50]), .B(n519), .ZN(n527) );
  INV_X1 U239 ( .A(n387), .ZN(n520) );
  OR2_X1 U240 ( .A1(n501), .A2(n541), .ZN(n521) );
  NAND2_X1 U241 ( .A1(n253), .A2(n521), .ZN(n249) );
  OR2_X1 U242 ( .A1(n494), .A2(n539), .ZN(n522) );
  NAND2_X1 U243 ( .A1(n386), .A2(n522), .ZN(n243) );
  XNOR2_X1 U244 ( .A(A[44]), .B(n523), .ZN(n524) );
  XNOR2_X1 U245 ( .A(n524), .B(n475), .ZN(SUM[44]) );
  XNOR2_X1 U246 ( .A(n525), .B(n472), .ZN(SUM[45]) );
  XNOR2_X1 U247 ( .A(A[45]), .B(B[45]), .ZN(n525) );
  AOI22_X1 U248 ( .A1(n520), .A2(n498), .B1(n327), .B2(B[27]), .ZN(n324) );
  INV_X1 U249 ( .A(n540), .ZN(n526) );
  XNOR2_X1 U250 ( .A(n527), .B(n515), .ZN(SUM[50]) );
  AND2_X1 U251 ( .A1(n481), .A2(n508), .ZN(n528) );
  AND2_X1 U252 ( .A1(n464), .A2(n480), .ZN(n529) );
  XNOR2_X1 U253 ( .A(n320), .B(n419), .ZN(SUM[30]) );
  XNOR2_X1 U254 ( .A(n495), .B(n332), .ZN(SUM[26]) );
  XNOR2_X1 U255 ( .A(n479), .B(n326), .ZN(SUM[28]) );
  AOI22_X1 U256 ( .A1(n487), .A2(n502), .B1(n333), .B2(B[25]), .ZN(n331) );
  INV_X1 U257 ( .A(n336), .ZN(n538) );
  OAI21_X1 U258 ( .B1(A[24]), .B2(B[24]), .A(carry[24]), .ZN(n336) );
  AND2_X1 U259 ( .A1(A[0]), .A2(B[0]), .ZN(n1) );
  INV_X1 U260 ( .A(A[55]), .ZN(n540) );
  INV_X1 U261 ( .A(A[54]), .ZN(n539) );
  XNOR2_X1 U262 ( .A(n483), .B(n335), .ZN(SUM[25]) );
  INV_X1 U263 ( .A(n334), .ZN(n537) );
  AOI21_X1 U264 ( .B1(B[24]), .B2(A[24]), .A(n538), .ZN(n334) );
  INV_X1 U265 ( .A(A[50]), .ZN(n542) );
  INV_X1 U266 ( .A(n258), .ZN(n533) );
  INV_X1 U267 ( .A(A[48]), .ZN(n543) );
  INV_X1 U268 ( .A(A[52]), .ZN(n541) );
  OR2_X1 U269 ( .A1(n394), .A2(A[27]), .ZN(n327) );
  INV_X1 U270 ( .A(A[28]), .ZN(n545) );
  OR2_X1 U271 ( .A1(n536), .A2(A[26]), .ZN(n330) );
  OAI21_X1 U272 ( .B1(n489), .B2(n510), .A(B[52]), .ZN(n253) );
  OAI21_X1 U273 ( .B1(n535), .B2(A[28]), .A(B[28]), .ZN(n325) );
  INV_X1 U274 ( .A(n331), .ZN(n536) );
  OAI21_X1 U275 ( .B1(n431), .B2(n490), .A(B[54]), .ZN(n247) );
  OAI21_X1 U276 ( .B1(n261), .B2(A[49]), .A(B[49]), .ZN(n262) );
  XNOR2_X1 U277 ( .A(n387), .B(n329), .ZN(SUM[27]) );
  OR2_X1 U278 ( .A1(A[25]), .A2(n537), .ZN(n333) );
  OAI21_X1 U279 ( .B1(n309), .B2(n417), .A(B[33]), .ZN(n310) );
  INV_X1 U280 ( .A(n324), .ZN(n535) );
  INV_X1 U281 ( .A(n262), .ZN(n534) );
  INV_X1 U282 ( .A(n250), .ZN(n531) );
  OAI21_X1 U283 ( .B1(n491), .B2(n273), .A(B[45]), .ZN(n274) );
  OAI21_X1 U284 ( .B1(n526), .B2(n485), .A(B[55]), .ZN(n242) );
  OAI21_X1 U285 ( .B1(n249), .B2(n480), .A(B[53]), .ZN(n250) );
  INV_X1 U286 ( .A(n256), .ZN(n532) );
  OAI21_X1 U287 ( .B1(n255), .B2(n508), .A(B[51]), .ZN(n256) );
  INV_X1 U288 ( .A(A[44]), .ZN(n544) );
  OAI21_X1 U289 ( .B1(n533), .B2(n511), .A(B[50]), .ZN(n259) );
  INV_X1 U290 ( .A(n268), .ZN(net176879) );
endmodule


module RCA_NBIT58 ( A, B, Ci, S, Co );
  input [57:0] A;
  input [57:0] B;
  output [57:0] S;
  input Ci;
  output Co;

  assign Co = 1'b0;

  RCA_NBIT58_DW01_add_0 add_95 ( .A(A), .B(B), .CI(1'b0), .SUM(S) );
endmodule


module RCA_NBIT60_DW01_add_0 ( A, B, CI, SUM, CO );
  input [59:0] A;
  input [59:0] B;
  output [59:0] SUM;
  input CI;
  output CO;
  wire   n1, n295, n296, n297, n298, n299, n300, n302, n303, n304, n305, n306,
         n308, n309, n310, n311, n312, n314, n315, n316, n317, n318, n320,
         n321, n329, n340, n356, n359, n360, n362, n363, n365, n366, n369,
         n370, n371, n372, n374, n375, n376, n378, n380, n381, n382, n383,
         net176898, net182615, net182746, net182859, net183396, net184334,
         net184968, net185085, net186806, net197538, net182618, n350, n347,
         net186793, net184798, net183635, net183226, net176894, n348, n345,
         n344, n341, net183653, net176921, n322, net199683, net176919, n326,
         net184500, net184136, net183192, net176897, n327, n324, n323, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n301, n307, n313, n319,
         n325, n328, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n342, n343, n346, n349, n351, n352, n353, n354, n355, n357,
         n358, n361, n364, n367, n368, n373, n377, n379, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436;
  wire   [59:1] carry;

  FA_X1 U1_29 ( .A(B[29]), .B(carry[29]), .CI(A[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XNOR2_X2 U3 ( .A(n297), .B(n298), .ZN(SUM[59]) );
  XOR2_X1 U129 ( .A(B[59]), .B(A[59]), .Z(n298) );
  XOR2_X1 U162 ( .A(carry[26]), .B(n296), .Z(SUM[26]) );
  XOR2_X1 U163 ( .A(A[26]), .B(B[26]), .Z(n296) );
  XOR2_X1 U164 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  CLKBUF_X1 U1 ( .A(A[42]), .Z(n351) );
  NAND2_X1 U2 ( .A1(n313), .A2(n319), .ZN(n254) );
  BUF_X1 U4 ( .A(A[44]), .Z(net183226) );
  AOI21_X2 U5 ( .B1(n436), .B2(n380), .A(n381), .ZN(n263) );
  CLKBUF_X3 U6 ( .A(n341), .Z(net183635) );
  INV_X1 U7 ( .A(n335), .ZN(net185085) );
  INV_X1 U8 ( .A(B[28]), .ZN(n387) );
  AND2_X1 U9 ( .A1(n414), .A2(n429), .ZN(n255) );
  INV_X1 U10 ( .A(B[48]), .ZN(net182859) );
  BUF_X1 U11 ( .A(A[34]), .Z(n257) );
  AOI22_X1 U12 ( .A1(net183635), .A2(net183226), .B1(n294), .B2(B[44]), .ZN(
        n256) );
  BUF_X1 U13 ( .A(A[35]), .Z(n259) );
  BUF_X1 U14 ( .A(A[54]), .Z(n415) );
  BUF_X1 U15 ( .A(A[33]), .Z(n400) );
  CLKBUF_X1 U16 ( .A(A[32]), .Z(n264) );
  CLKBUF_X1 U17 ( .A(A[36]), .Z(n260) );
  CLKBUF_X1 U18 ( .A(A[27]), .Z(n258) );
  NAND2_X1 U19 ( .A1(n336), .A2(n337), .ZN(n335) );
  INV_X1 U20 ( .A(B[53]), .ZN(n404) );
  INV_X1 U21 ( .A(B[57]), .ZN(n417) );
  INV_X1 U22 ( .A(B[55]), .ZN(n395) );
  INV_X1 U23 ( .A(B[31]), .ZN(n293) );
  INV_X1 U24 ( .A(B[47]), .ZN(n279) );
  INV_X1 U25 ( .A(B[37]), .ZN(n262) );
  XNOR2_X1 U26 ( .A(n333), .B(n328), .ZN(SUM[39]) );
  XNOR2_X1 U27 ( .A(A[39]), .B(B[39]), .ZN(n333) );
  XNOR2_X1 U28 ( .A(n422), .B(n371), .ZN(SUM[34]) );
  NAND2_X1 U29 ( .A1(n325), .A2(n356), .ZN(n337) );
  INV_X1 U30 ( .A(B[39]), .ZN(n325) );
  NAND2_X1 U31 ( .A1(net197538), .A2(n268), .ZN(n273) );
  NOR2_X1 U32 ( .A1(n388), .A2(n378), .ZN(n368) );
  NAND2_X1 U33 ( .A1(n330), .A2(n331), .ZN(n313) );
  NAND2_X1 U34 ( .A1(net183635), .A2(net183226), .ZN(n270) );
  OAI21_X1 U35 ( .B1(n379), .B2(n416), .A(B[55]), .ZN(n261) );
  XNOR2_X1 U36 ( .A(A[37]), .B(n262), .ZN(n265) );
  XNOR2_X1 U37 ( .A(n265), .B(n362), .ZN(SUM[37]) );
  OAI21_X1 U38 ( .B1(n266), .B2(n267), .A(net182859), .ZN(net176919) );
  INV_X1 U39 ( .A(n373), .ZN(n380) );
  OAI21_X1 U40 ( .B1(n269), .B2(B[45]), .A(n273), .ZN(n272) );
  INV_X1 U41 ( .A(n272), .ZN(n278) );
  INV_X1 U42 ( .A(A[45]), .ZN(n268) );
  OAI21_X1 U43 ( .B1(n286), .B2(A[46]), .A(B[46]), .ZN(n275) );
  AOI21_X1 U44 ( .B1(n271), .B2(n270), .A(n268), .ZN(n269) );
  NAND2_X1 U45 ( .A1(n284), .A2(n275), .ZN(n274) );
  NAND2_X1 U46 ( .A1(A[47]), .A2(n274), .ZN(n280) );
  XNOR2_X1 U47 ( .A(n282), .B(B[47]), .ZN(n277) );
  OR2_X1 U48 ( .A1(A[47]), .A2(n282), .ZN(n281) );
  XNOR2_X1 U49 ( .A(n277), .B(n285), .ZN(SUM[47]) );
  NAND2_X1 U50 ( .A1(n283), .A2(n284), .ZN(n282) );
  XNOR2_X1 U51 ( .A(A[48]), .B(B[48]), .ZN(net184334) );
  INV_X1 U52 ( .A(net199683), .ZN(n266) );
  OAI21_X1 U53 ( .B1(n278), .B2(A[46]), .A(B[46]), .ZN(n283) );
  XNOR2_X1 U54 ( .A(net182746), .B(n286), .ZN(SUM[46]) );
  NAND2_X1 U55 ( .A1(n278), .A2(A[46]), .ZN(n284) );
  CLKBUF_X1 U56 ( .A(A[47]), .Z(n285) );
  INV_X1 U57 ( .A(n272), .ZN(n286) );
  NAND2_X1 U58 ( .A1(n280), .A2(n279), .ZN(n276) );
  BUF_X1 U59 ( .A(A[48]), .Z(net199683) );
  OAI21_X1 U60 ( .B1(net183226), .B2(net183635), .A(B[44]), .ZN(n271) );
  NAND2_X1 U61 ( .A1(n281), .A2(n276), .ZN(n267) );
  AND2_X1 U62 ( .A1(n281), .A2(n276), .ZN(n329) );
  AOI21_X1 U63 ( .B1(n323), .B2(n288), .A(B[50]), .ZN(n324) );
  INV_X1 U64 ( .A(n324), .ZN(net176921) );
  CLKBUF_X1 U65 ( .A(A[50]), .Z(n288) );
  OR2_X1 U66 ( .A1(n288), .A2(n323), .ZN(net183653) );
  NAND2_X1 U67 ( .A1(n327), .A2(net184136), .ZN(n323) );
  XNOR2_X1 U68 ( .A(n323), .B(n287), .ZN(SUM[50]) );
  OR2_X1 U69 ( .A1(n326), .A2(net176897), .ZN(net184136) );
  INV_X1 U70 ( .A(A[49]), .ZN(net176897) );
  OAI21_X1 U71 ( .B1(net183192), .B2(net184500), .A(B[49]), .ZN(n327) );
  CLKBUF_X1 U72 ( .A(A[49]), .Z(net184500) );
  INV_X1 U73 ( .A(n326), .ZN(net183192) );
  XNOR2_X1 U74 ( .A(A[50]), .B(B[50]), .ZN(n287) );
  XNOR2_X1 U75 ( .A(A[49]), .B(B[49]), .ZN(net182615) );
  CLKBUF_X1 U76 ( .A(n254), .Z(n289) );
  OAI21_X1 U77 ( .B1(net199683), .B2(n329), .A(net176919), .ZN(n326) );
  XNOR2_X1 U78 ( .A(n322), .B(n291), .ZN(SUM[51]) );
  AND2_X1 U79 ( .A1(net176921), .A2(net183653), .ZN(n291) );
  AND2_X1 U80 ( .A1(net176921), .A2(net183653), .ZN(n290) );
  NAND2_X1 U81 ( .A1(net176921), .A2(net183653), .ZN(n320) );
  XNOR2_X1 U82 ( .A(A[51]), .B(B[51]), .ZN(n322) );
  INV_X1 U83 ( .A(A[51]), .ZN(net176898) );
  OAI21_X1 U84 ( .B1(n290), .B2(A[51]), .A(B[51]), .ZN(n321) );
  OAI21_X1 U85 ( .B1(n432), .B2(n308), .A(n261), .ZN(n292) );
  XNOR2_X1 U86 ( .A(A[31]), .B(n293), .ZN(n382) );
  OR2_X1 U87 ( .A1(n341), .A2(A[44]), .ZN(n294) );
  CLKBUF_X1 U88 ( .A(n339), .Z(n301) );
  AND2_X1 U89 ( .A1(n301), .A2(n342), .ZN(n307) );
  NAND2_X1 U90 ( .A1(n350), .A2(n332), .ZN(n342) );
  NAND2_X1 U91 ( .A1(n313), .A2(n319), .ZN(n350) );
  NAND2_X1 U92 ( .A1(n343), .A2(n335), .ZN(n319) );
  NAND2_X1 U93 ( .A1(A[40]), .A2(B[40]), .ZN(n343) );
  INV_X1 U94 ( .A(A[40]), .ZN(n330) );
  INV_X1 U95 ( .A(A[41]), .ZN(n338) );
  INV_X1 U96 ( .A(A[39]), .ZN(n334) );
  OAI21_X1 U97 ( .B1(n254), .B2(n332), .A(n338), .ZN(n339) );
  OAI21_X1 U98 ( .B1(n356), .B2(n325), .A(n334), .ZN(n336) );
  INV_X1 U99 ( .A(n356), .ZN(n328) );
  AND2_X1 U100 ( .A1(n339), .A2(n342), .ZN(n347) );
  INV_X1 U101 ( .A(B[40]), .ZN(n331) );
  INV_X1 U102 ( .A(B[41]), .ZN(n332) );
  XNOR2_X1 U103 ( .A(A[41]), .B(n332), .ZN(net182618) );
  XOR2_X1 U104 ( .A(A[40]), .B(n331), .Z(net183396) );
  BUF_X1 U105 ( .A(n307), .Z(n346) );
  AOI22_X1 U106 ( .A1(net183635), .A2(net183226), .B1(n294), .B2(B[44]), .ZN(
        net197538) );
  XNOR2_X1 U107 ( .A(n354), .B(net183635), .ZN(SUM[44]) );
  XNOR2_X1 U108 ( .A(A[44]), .B(B[44]), .ZN(n354) );
  NOR2_X1 U109 ( .A1(n345), .A2(net184798), .ZN(n341) );
  AND2_X1 U110 ( .A1(net176894), .A2(net186793), .ZN(net184798) );
  AOI22_X1 U111 ( .A1(n346), .A2(n351), .B1(n353), .B2(B[42]), .ZN(net186793)
         );
  OR2_X1 U112 ( .A1(n347), .A2(A[42]), .ZN(n353) );
  AOI22_X1 U113 ( .A1(n307), .A2(n351), .B1(n348), .B2(B[42]), .ZN(n344) );
  XNOR2_X1 U114 ( .A(n346), .B(n352), .ZN(SUM[42]) );
  INV_X1 U115 ( .A(A[43]), .ZN(net176894) );
  AOI21_X1 U116 ( .B1(n349), .B2(A[43]), .A(B[43]), .ZN(n345) );
  INV_X1 U117 ( .A(n344), .ZN(n349) );
  CLKBUF_X1 U118 ( .A(n349), .Z(net184968) );
  OR2_X1 U119 ( .A1(A[42]), .A2(n347), .ZN(n348) );
  XNOR2_X1 U120 ( .A(A[42]), .B(B[42]), .ZN(n352) );
  XNOR2_X1 U121 ( .A(A[43]), .B(B[43]), .ZN(net186806) );
  XNOR2_X1 U122 ( .A(net182618), .B(n289), .ZN(SUM[41]) );
  OR2_X1 U123 ( .A1(n314), .A2(n433), .ZN(n355) );
  BUF_X1 U124 ( .A(A[30]), .Z(n390) );
  NAND2_X1 U125 ( .A1(n259), .A2(n357), .ZN(n384) );
  AND2_X1 U126 ( .A1(n429), .A2(n414), .ZN(n357) );
  XOR2_X1 U127 ( .A(n258), .B(B[27]), .Z(n358) );
  XOR2_X1 U128 ( .A(n430), .B(n358), .Z(SUM[27]) );
  NAND2_X1 U130 ( .A1(n430), .A2(A[27]), .ZN(n361) );
  NAND2_X1 U131 ( .A1(n430), .A2(B[27]), .ZN(n364) );
  NAND2_X1 U132 ( .A1(A[27]), .A2(B[27]), .ZN(n367) );
  NAND3_X1 U133 ( .A1(n361), .A2(n364), .A3(n367), .ZN(carry[28]) );
  NAND2_X1 U134 ( .A1(n383), .A2(n377), .ZN(n373) );
  NAND2_X1 U135 ( .A1(A[30]), .A2(B[30]), .ZN(n377) );
  AND2_X1 U136 ( .A1(n385), .A2(n426), .ZN(n379) );
  NAND2_X1 U137 ( .A1(n369), .A2(n384), .ZN(n365) );
  CLKBUF_X1 U138 ( .A(A[56]), .Z(n393) );
  OR2_X1 U139 ( .A1(n415), .A2(n391), .ZN(n385) );
  NAND2_X1 U140 ( .A1(n385), .A2(n426), .ZN(n308) );
  OAI21_X1 U141 ( .B1(n393), .B2(n389), .A(n425), .ZN(n386) );
  BUF_X1 U142 ( .A(n359), .Z(n403) );
  XNOR2_X1 U143 ( .A(carry[28]), .B(n387), .ZN(n405) );
  OR2_X1 U144 ( .A1(n378), .A2(n388), .ZN(n374) );
  NOR2_X1 U145 ( .A1(n263), .A2(n264), .ZN(n388) );
  XNOR2_X1 U146 ( .A(net184968), .B(net186806), .ZN(SUM[43]) );
  CLKBUF_X1 U147 ( .A(n292), .Z(n389) );
  XOR2_X1 U148 ( .A(A[45]), .B(B[45]), .Z(n340) );
  NAND2_X1 U149 ( .A1(n355), .A2(n315), .ZN(n391) );
  BUF_X1 U150 ( .A(A[55]), .Z(n416) );
  OR2_X1 U151 ( .A1(n399), .A2(n366), .ZN(n362) );
  CLKBUF_X1 U152 ( .A(A[52]), .Z(n392) );
  AND2_X1 U153 ( .A1(n427), .A2(n412), .ZN(n394) );
  XNOR2_X1 U154 ( .A(A[55]), .B(n395), .ZN(n310) );
  XNOR2_X1 U155 ( .A(n300), .B(n396), .ZN(SUM[58]) );
  XNOR2_X1 U156 ( .A(B[58]), .B(A[58]), .ZN(n396) );
  OR2_X1 U157 ( .A1(n320), .A2(net176898), .ZN(n397) );
  NAND2_X1 U158 ( .A1(n397), .A2(n321), .ZN(n317) );
  NOR2_X1 U159 ( .A1(n366), .A2(n399), .ZN(n398) );
  XNOR2_X1 U160 ( .A(A[52]), .B(B[52]), .ZN(n410) );
  NOR2_X1 U161 ( .A1(n365), .A2(n260), .ZN(n399) );
  CLKBUF_X1 U165 ( .A(A[28]), .Z(n401) );
  XNOR2_X1 U166 ( .A(net184334), .B(n329), .ZN(SUM[48]) );
  INV_X1 U167 ( .A(n431), .ZN(n402) );
  XNOR2_X1 U168 ( .A(A[53]), .B(n404), .ZN(n316) );
  XOR2_X1 U169 ( .A(n405), .B(n401), .Z(SUM[28]) );
  NAND2_X1 U170 ( .A1(A[28]), .A2(carry[28]), .ZN(n406) );
  NAND2_X1 U171 ( .A1(A[28]), .A2(B[28]), .ZN(n407) );
  NAND2_X1 U172 ( .A1(carry[28]), .A2(B[28]), .ZN(n408) );
  NAND3_X1 U173 ( .A1(n406), .A2(n407), .A3(n408), .ZN(carry[29]) );
  XNOR2_X1 U174 ( .A(n409), .B(n263), .ZN(SUM[32]) );
  XNOR2_X1 U175 ( .A(A[32]), .B(B[32]), .ZN(n409) );
  XNOR2_X1 U176 ( .A(n410), .B(n317), .ZN(SUM[52]) );
  OR2_X1 U177 ( .A1(n302), .A2(n431), .ZN(n411) );
  NAND2_X1 U178 ( .A1(n303), .A2(n411), .ZN(n300) );
  NAND2_X1 U179 ( .A1(n315), .A2(n355), .ZN(n311) );
  OR2_X1 U180 ( .A1(n392), .A2(n317), .ZN(n412) );
  NAND2_X1 U181 ( .A1(n427), .A2(n412), .ZN(n314) );
  AND2_X1 U182 ( .A1(n429), .A2(n414), .ZN(n413) );
  XNOR2_X1 U183 ( .A(net183396), .B(net185085), .ZN(SUM[40]) );
  OR2_X1 U184 ( .A1(n371), .A2(n257), .ZN(n414) );
  XNOR2_X1 U185 ( .A(A[46]), .B(B[46]), .ZN(net182746) );
  XNOR2_X1 U186 ( .A(A[57]), .B(n417), .ZN(n304) );
  XNOR2_X1 U187 ( .A(net182615), .B(net183192), .ZN(SUM[49]) );
  INV_X1 U188 ( .A(A[31]), .ZN(n436) );
  AND2_X1 U189 ( .A1(n300), .A2(A[58]), .ZN(n299) );
  XNOR2_X1 U190 ( .A(n418), .B(n391), .ZN(SUM[54]) );
  XNOR2_X1 U191 ( .A(A[54]), .B(B[54]), .ZN(n418) );
  XNOR2_X1 U192 ( .A(n419), .B(n390), .ZN(SUM[30]) );
  XNOR2_X1 U193 ( .A(carry[30]), .B(B[30]), .ZN(n419) );
  XNOR2_X1 U194 ( .A(n420), .B(n403), .ZN(SUM[38]) );
  XNOR2_X1 U195 ( .A(A[38]), .B(B[38]), .ZN(n420) );
  XNOR2_X1 U196 ( .A(n421), .B(n365), .ZN(SUM[36]) );
  XNOR2_X1 U197 ( .A(A[36]), .B(B[36]), .ZN(n421) );
  XNOR2_X1 U198 ( .A(A[34]), .B(B[34]), .ZN(n422) );
  AOI21_X1 U199 ( .B1(A[31]), .B2(n373), .A(B[31]), .ZN(n381) );
  XNOR2_X1 U200 ( .A(n423), .B(n305), .ZN(SUM[56]) );
  XNOR2_X1 U201 ( .A(A[56]), .B(B[56]), .ZN(n423) );
  INV_X1 U202 ( .A(n360), .ZN(n428) );
  OAI21_X1 U203 ( .B1(A[30]), .B2(B[30]), .A(carry[30]), .ZN(n383) );
  OAI21_X1 U204 ( .B1(n413), .B2(n259), .A(B[35]), .ZN(n369) );
  AOI21_X1 U205 ( .B1(n365), .B2(n260), .A(B[36]), .ZN(n366) );
  OAI21_X1 U206 ( .B1(n374), .B2(n435), .A(n375), .ZN(n371) );
  INV_X1 U207 ( .A(n400), .ZN(n435) );
  OAI21_X1 U208 ( .B1(n368), .B2(n400), .A(B[33]), .ZN(n375) );
  XNOR2_X1 U209 ( .A(n316), .B(n314), .ZN(SUM[53]) );
  XNOR2_X1 U210 ( .A(n376), .B(n368), .ZN(SUM[33]) );
  XNOR2_X1 U211 ( .A(A[33]), .B(B[33]), .ZN(n376) );
  XNOR2_X1 U212 ( .A(n370), .B(n255), .ZN(SUM[35]) );
  XNOR2_X1 U213 ( .A(A[35]), .B(B[35]), .ZN(n370) );
  XNOR2_X1 U214 ( .A(n382), .B(n380), .ZN(SUM[31]) );
  INV_X1 U215 ( .A(n302), .ZN(n424) );
  AOI21_X1 U216 ( .B1(n292), .B2(n393), .A(B[56]), .ZN(n306) );
  INV_X1 U217 ( .A(A[37]), .ZN(n434) );
  OAI21_X1 U218 ( .B1(n398), .B2(A[37]), .A(B[37]), .ZN(n363) );
  INV_X1 U219 ( .A(A[57]), .ZN(n431) );
  AOI21_X1 U220 ( .B1(n311), .B2(n415), .A(B[54]), .ZN(n312) );
  INV_X1 U221 ( .A(n372), .ZN(n429) );
  INV_X1 U222 ( .A(n295), .ZN(n430) );
  AOI22_X1 U223 ( .A1(B[26]), .A2(A[26]), .B1(n296), .B2(carry[26]), .ZN(n295)
         );
  AND2_X1 U224 ( .A1(A[0]), .A2(B[0]), .ZN(n1) );
  AOI21_X1 U225 ( .B1(n371), .B2(n257), .A(B[34]), .ZN(n372) );
  OAI21_X1 U226 ( .B1(n432), .B2(n308), .A(n309), .ZN(n305) );
  XNOR2_X1 U227 ( .A(n310), .B(n308), .ZN(SUM[55]) );
  AOI21_X1 U228 ( .B1(n264), .B2(n263), .A(B[32]), .ZN(n378) );
  XNOR2_X1 U229 ( .A(n304), .B(n386), .ZN(SUM[57]) );
  XNOR2_X1 U230 ( .A(n256), .B(n340), .ZN(SUM[45]) );
  OAI21_X1 U231 ( .B1(A[38]), .B2(n403), .A(n428), .ZN(n356) );
  AOI21_X1 U232 ( .B1(n359), .B2(A[38]), .A(B[38]), .ZN(n360) );
  OAI21_X1 U233 ( .B1(n362), .B2(n434), .A(n363), .ZN(n359) );
  INV_X1 U234 ( .A(A[53]), .ZN(n433) );
  AOI21_X1 U235 ( .B1(n317), .B2(n392), .A(B[52]), .ZN(n318) );
  OAI21_X1 U236 ( .B1(n394), .B2(A[53]), .A(B[53]), .ZN(n315) );
  OAI21_X1 U237 ( .B1(n393), .B2(n389), .A(n425), .ZN(n302) );
  INV_X1 U238 ( .A(n306), .ZN(n425) );
  INV_X1 U239 ( .A(n312), .ZN(n426) );
  INV_X1 U240 ( .A(n318), .ZN(n427) );
  OAI21_X1 U241 ( .B1(n424), .B2(n402), .A(B[57]), .ZN(n303) );
  OAI22_X1 U242 ( .A1(n299), .A2(B[58]), .B1(n300), .B2(A[58]), .ZN(n297) );
  OAI21_X1 U243 ( .B1(n379), .B2(n416), .A(B[55]), .ZN(n309) );
  INV_X1 U244 ( .A(n416), .ZN(n432) );
endmodule


module RCA_NBIT60 ( A, B, Ci, S, Co );
  input [59:0] A;
  input [59:0] B;
  output [59:0] S;
  input Ci;
  output Co;

  assign Co = 1'b0;

  RCA_NBIT60_DW01_add_0 add_95 ( .A(A), .B(B), .CI(1'b0), .SUM(S) );
endmodule


module RCA_NBIT62_DW01_add_0 ( A, B, CI, SUM, CO );
  input [61:0] A;
  input [61:0] B;
  output [61:0] SUM;
  input CI;
  output CO;
  wire   n1, \carry[59] , \carry[58] , n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n336, n338, n339, n340, n344, n346, n347, n348,
         n350, n351, n353, n354, n360, n367, n370, n371, n373, n374, n375,
         n376, n377, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n394, n395, n397, n398, n400, n401, n405, n411, net176946, net176961,
         net182620, net183453, net183785, net183931, net184000, net184550,
         net184547, net185657, net185823, net186117, net176945, n407, n403,
         net186084, net182688, n357, n356, n355, n352, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n335, n337, n341, n342, n343, n345, n349,
         n358, n359, n361, n362, n363, n364, n365, n366, n368, n369, n372,
         n378, n388, n389, n390, n391, n392, n393, n396, n399, n402, n404,
         n406, n408, n409, n410, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508;
  wire   [61:1] carry;

  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  FA_X1 U1_57 ( .A(A[57]), .B(B[57]), .CI(n492), .CO(\carry[58] ), .S(SUM[57])
         );
  FA_X1 U1_58 ( .A(A[58]), .B(B[58]), .CI(\carry[58] ), .CO(\carry[59] ), .S(
        SUM[58]) );
  XOR2_X1 U131 ( .A(B[61]), .B(A[61]), .Z(n330) );
  XOR2_X1 U132 ( .A(B[60]), .B(A[60]), .Z(n333) );
  XOR2_X1 U135 ( .A(n482), .B(n336), .Z(SUM[56]) );
  XOR2_X1 U136 ( .A(n486), .B(B[56]), .Z(n336) );
  XOR2_X1 U139 ( .A(n292), .B(n348), .Z(SUM[52]) );
  XOR2_X1 U140 ( .A(A[52]), .B(B[52]), .Z(n348) );
  XOR2_X1 U141 ( .A(net184000), .B(n354), .Z(SUM[50]) );
  XOR2_X1 U142 ( .A(A[50]), .B(B[50]), .Z(n354) );
  XOR2_X1 U143 ( .A(net183453), .B(n360), .Z(SUM[48]) );
  XOR2_X1 U149 ( .A(A[43]), .B(B[43]), .Z(n375) );
  XOR2_X1 U152 ( .A(n387), .B(net184547), .Z(SUM[39]) );
  XOR2_X1 U153 ( .A(A[39]), .B(B[39]), .Z(n387) );
  XOR2_X1 U165 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  XOR2_X1 U144 ( .A(net182688), .B(B[48]), .Z(n360) );
  CLKBUF_X1 U1 ( .A(n345), .Z(n285) );
  OAI21_X1 U2 ( .B1(n499), .B2(n469), .A(B[36]), .ZN(n286) );
  INV_X1 U3 ( .A(A[47]), .ZN(n287) );
  BUF_X1 U4 ( .A(n450), .Z(n288) );
  AND2_X1 U5 ( .A1(n395), .A2(n308), .ZN(n289) );
  AND2_X1 U6 ( .A1(n286), .A2(n308), .ZN(n307) );
  OR2_X1 U7 ( .A1(n298), .A2(n297), .ZN(n290) );
  AND2_X1 U8 ( .A1(n428), .A2(n424), .ZN(n291) );
  BUF_X1 U9 ( .A(n397), .Z(n471) );
  NOR2_X1 U10 ( .A1(n298), .A2(n297), .ZN(n292) );
  AND2_X1 U11 ( .A1(n293), .A2(B[38]), .ZN(n444) );
  NAND2_X1 U12 ( .A1(n446), .A2(n445), .ZN(n293) );
  CLKBUF_X1 U13 ( .A(n427), .Z(n294) );
  AND2_X2 U14 ( .A1(n407), .A2(n438), .ZN(n309) );
  NAND2_X1 U15 ( .A1(carry[29]), .A2(B[29]), .ZN(n426) );
  INV_X1 U16 ( .A(B[29]), .ZN(n412) );
  INV_X1 U17 ( .A(B[46]), .ZN(n389) );
  INV_X1 U18 ( .A(B[47]), .ZN(n388) );
  XNOR2_X1 U19 ( .A(n434), .B(n420), .ZN(SUM[29]) );
  XNOR2_X1 U20 ( .A(n433), .B(B[29]), .ZN(n420) );
  NOR2_X1 U21 ( .A1(net185823), .A2(net183785), .ZN(n295) );
  CLKBUF_X1 U22 ( .A(A[59]), .Z(n296) );
  XNOR2_X1 U23 ( .A(n329), .B(n330), .ZN(SUM[61]) );
  NOR2_X1 U24 ( .A1(n463), .A2(A[51]), .ZN(n297) );
  CLKBUF_X1 U25 ( .A(A[44]), .Z(n464) );
  BUF_X1 U26 ( .A(n493), .Z(n460) );
  AOI21_X1 U27 ( .B1(n465), .B2(A[51]), .A(B[51]), .ZN(n298) );
  XNOR2_X1 U28 ( .A(n309), .B(n405), .ZN(SUM[33]) );
  XNOR2_X1 U29 ( .A(n453), .B(n299), .ZN(SUM[54]) );
  XNOR2_X1 U30 ( .A(n337), .B(B[54]), .ZN(n299) );
  CLKBUF_X1 U31 ( .A(A[54]), .Z(n337) );
  OR2_X1 U32 ( .A1(n377), .A2(n480), .ZN(n300) );
  NOR2_X2 U33 ( .A1(n302), .A2(n495), .ZN(n485) );
  AOI21_X1 U34 ( .B1(n453), .B2(n337), .A(n460), .ZN(n301) );
  AND2_X1 U35 ( .A1(A[52]), .A2(n306), .ZN(n302) );
  NAND2_X1 U36 ( .A1(n288), .A2(n303), .ZN(n441) );
  AND2_X1 U37 ( .A1(n293), .A2(n451), .ZN(n303) );
  BUF_X1 U38 ( .A(n327), .Z(n482) );
  BUF_X1 U39 ( .A(A[41]), .Z(n478) );
  OAI21_X1 U40 ( .B1(n346), .B2(A[52]), .A(B[52]), .ZN(n304) );
  INV_X1 U41 ( .A(B[33]), .ZN(n439) );
  AOI21_X1 U42 ( .B1(n503), .B2(n485), .A(n344), .ZN(n305) );
  BUF_X1 U43 ( .A(n441), .Z(net184550) );
  NOR2_X1 U44 ( .A1(n298), .A2(n297), .ZN(n306) );
  NAND2_X1 U45 ( .A1(n499), .A2(n469), .ZN(n308) );
  CLKBUF_X1 U46 ( .A(n394), .Z(n406) );
  INV_X1 U47 ( .A(B[30]), .ZN(n424) );
  INV_X1 U48 ( .A(n309), .ZN(n403) );
  BUF_X1 U49 ( .A(n300), .Z(n408) );
  XNOR2_X1 U50 ( .A(n310), .B(n484), .ZN(SUM[44]) );
  XNOR2_X1 U51 ( .A(B[44]), .B(A[44]), .ZN(n310) );
  XNOR2_X1 U52 ( .A(n294), .B(n431), .ZN(SUM[30]) );
  OAI21_X1 U53 ( .B1(n311), .B2(n290), .A(n304), .ZN(n494) );
  INV_X1 U54 ( .A(A[52]), .ZN(n311) );
  AOI21_X1 U55 ( .B1(n312), .B2(n313), .A(n314), .ZN(n493) );
  INV_X1 U56 ( .A(n305), .ZN(n312) );
  INV_X1 U57 ( .A(A[54]), .ZN(n313) );
  INV_X1 U58 ( .A(B[54]), .ZN(n314) );
  OAI21_X1 U59 ( .B1(n315), .B2(n309), .A(n439), .ZN(net176946) );
  INV_X1 U60 ( .A(A[33]), .ZN(n315) );
  NAND2_X1 U61 ( .A1(n345), .A2(A[46]), .ZN(n316) );
  CLKBUF_X1 U62 ( .A(A[48]), .Z(net182688) );
  XNOR2_X1 U63 ( .A(A[46]), .B(B[46]), .ZN(n369) );
  INV_X1 U64 ( .A(A[46]), .ZN(n366) );
  INV_X1 U65 ( .A(A[36]), .ZN(n317) );
  NAND2_X1 U66 ( .A1(n418), .A2(n419), .ZN(n435) );
  XNOR2_X1 U67 ( .A(A[45]), .B(B[45]), .ZN(n372) );
  AND2_X1 U68 ( .A1(n417), .A2(B[31]), .ZN(n421) );
  NAND2_X1 U69 ( .A1(n392), .A2(n389), .ZN(n318) );
  XOR2_X1 U70 ( .A(A[34]), .B(B[34]), .Z(n487) );
  INV_X1 U71 ( .A(net186117), .ZN(n427) );
  NAND2_X1 U72 ( .A1(n318), .A2(n361), .ZN(n319) );
  CLKBUF_X1 U73 ( .A(n370), .Z(n484) );
  OAI21_X1 U74 ( .B1(n322), .B2(B[45]), .A(A[45]), .ZN(n320) );
  OAI21_X1 U75 ( .B1(n484), .B2(n464), .A(n496), .ZN(n321) );
  INV_X1 U76 ( .A(n367), .ZN(n322) );
  AND2_X1 U77 ( .A1(n318), .A2(n361), .ZN(n323) );
  NAND2_X1 U78 ( .A1(n409), .A2(n410), .ZN(net186117) );
  NAND2_X1 U79 ( .A1(n412), .A2(n413), .ZN(n409) );
  NAND2_X1 U80 ( .A1(n428), .A2(n424), .ZN(n416) );
  AND2_X1 U81 ( .A1(n320), .A2(n349), .ZN(n324) );
  CLKBUF_X1 U82 ( .A(n365), .Z(n325) );
  XNOR2_X1 U83 ( .A(n289), .B(n335), .ZN(SUM[37]) );
  XNOR2_X1 U84 ( .A(A[37]), .B(n445), .ZN(n335) );
  XNOR2_X1 U85 ( .A(n406), .B(n341), .ZN(SUM[36]) );
  XNOR2_X1 U86 ( .A(n317), .B(B[36]), .ZN(n341) );
  NAND2_X1 U87 ( .A1(n426), .A2(n423), .ZN(n410) );
  NAND2_X1 U88 ( .A1(n366), .A2(n324), .ZN(n361) );
  NAND2_X1 U89 ( .A1(n316), .A2(n389), .ZN(n362) );
  AND2_X1 U90 ( .A1(n390), .A2(n391), .ZN(n342) );
  BUF_X1 U91 ( .A(A[56]), .Z(n486) );
  CLKBUF_X1 U92 ( .A(n287), .Z(n343) );
  NAND2_X1 U93 ( .A1(n361), .A2(n362), .ZN(n359) );
  INV_X1 U94 ( .A(n321), .ZN(n365) );
  NAND2_X1 U95 ( .A1(B[45]), .A2(n365), .ZN(n349) );
  OAI21_X1 U96 ( .B1(n322), .B2(B[45]), .A(A[45]), .ZN(n358) );
  XNOR2_X1 U97 ( .A(n372), .B(n325), .ZN(SUM[45]) );
  NAND2_X1 U98 ( .A1(n287), .A2(n359), .ZN(n391) );
  OAI21_X1 U99 ( .B1(n319), .B2(n368), .A(n388), .ZN(n390) );
  XNOR2_X1 U100 ( .A(n378), .B(n343), .ZN(SUM[47]) );
  NAND2_X1 U101 ( .A1(n390), .A2(n391), .ZN(n363) );
  INV_X1 U102 ( .A(A[48]), .ZN(n364) );
  INV_X1 U103 ( .A(A[47]), .ZN(n368) );
  NAND2_X1 U104 ( .A1(n358), .A2(n349), .ZN(n345) );
  NAND2_X1 U105 ( .A1(n363), .A2(n364), .ZN(net186084) );
  XNOR2_X1 U106 ( .A(n323), .B(n388), .ZN(n378) );
  NAND2_X1 U107 ( .A1(n345), .A2(A[46]), .ZN(n392) );
  XNOR2_X1 U108 ( .A(n369), .B(n285), .ZN(SUM[46]) );
  AOI21_X1 U109 ( .B1(n393), .B2(n399), .A(n356), .ZN(n352) );
  CLKBUF_X1 U110 ( .A(n352), .Z(net184000) );
  AND2_X1 U111 ( .A1(n352), .A2(A[50]), .ZN(net183785) );
  OAI21_X1 U112 ( .B1(n352), .B2(A[50]), .A(B[50]), .ZN(n353) );
  AOI21_X1 U113 ( .B1(n396), .B2(A[49]), .A(B[49]), .ZN(n356) );
  INV_X1 U114 ( .A(n402), .ZN(n396) );
  AOI22_X1 U115 ( .A1(n342), .A2(net182688), .B1(net186084), .B2(B[48]), .ZN(
        n402) );
  AOI22_X1 U116 ( .A1(net182688), .A2(n342), .B1(net186084), .B2(B[48]), .ZN(
        n355) );
  CLKBUF_X1 U117 ( .A(n342), .Z(net183453) );
  CLKBUF_X1 U118 ( .A(n355), .Z(n399) );
  XNOR2_X1 U119 ( .A(n357), .B(n399), .ZN(SUM[49]) );
  INV_X1 U120 ( .A(A[49]), .ZN(n393) );
  XNOR2_X1 U121 ( .A(B[49]), .B(n393), .ZN(n357) );
  NAND2_X1 U122 ( .A1(n416), .A2(n417), .ZN(net185657) );
  NAND2_X1 U123 ( .A1(n421), .A2(n416), .ZN(n429) );
  OR2_X1 U124 ( .A1(n291), .A2(n422), .ZN(n404) );
  NAND2_X1 U125 ( .A1(n404), .A2(n425), .ZN(n430) );
  NAND2_X1 U126 ( .A1(n417), .A2(B[31]), .ZN(n422) );
  NAND2_X1 U127 ( .A1(net186117), .A2(n414), .ZN(n417) );
  AOI21_X1 U128 ( .B1(n416), .B2(n417), .A(B[31]), .ZN(n432) );
  INV_X1 U129 ( .A(n432), .ZN(n419) );
  INV_X1 U130 ( .A(A[31]), .ZN(n425) );
  NAND2_X1 U133 ( .A1(n425), .A2(n429), .ZN(n418) );
  XNOR2_X1 U134 ( .A(A[30]), .B(B[30]), .ZN(n431) );
  NAND2_X1 U137 ( .A1(n427), .A2(A[30]), .ZN(n428) );
  INV_X1 U138 ( .A(A[30]), .ZN(n414) );
  INV_X1 U145 ( .A(B[31]), .ZN(n415) );
  XNOR2_X1 U146 ( .A(A[31]), .B(n415), .ZN(n411) );
  INV_X1 U147 ( .A(carry[29]), .ZN(n413) );
  INV_X1 U148 ( .A(n413), .ZN(n433) );
  AND2_X1 U150 ( .A1(n419), .A2(n430), .ZN(net176945) );
  INV_X1 U151 ( .A(A[29]), .ZN(n423) );
  INV_X1 U154 ( .A(n423), .ZN(n434) );
  OR2_X1 U155 ( .A1(n436), .A2(n435), .ZN(n438) );
  INV_X1 U156 ( .A(A[32]), .ZN(n436) );
  OAI21_X1 U157 ( .B1(net176945), .B2(A[32]), .A(B[32]), .ZN(n407) );
  CLKBUF_X1 U158 ( .A(A[33]), .Z(net183931) );
  XNOR2_X1 U159 ( .A(A[33]), .B(n439), .ZN(n405) );
  XNOR2_X1 U160 ( .A(n435), .B(n437), .ZN(SUM[32]) );
  XOR2_X1 U161 ( .A(A[32]), .B(B[32]), .Z(n437) );
  AND2_X1 U162 ( .A1(n449), .A2(n448), .ZN(n440) );
  NAND2_X1 U163 ( .A1(n452), .A2(n447), .ZN(n448) );
  INV_X1 U164 ( .A(A[37]), .ZN(n446) );
  NAND2_X1 U166 ( .A1(n307), .A2(n445), .ZN(n451) );
  NAND2_X1 U167 ( .A1(n289), .A2(n446), .ZN(n450) );
  NAND2_X1 U168 ( .A1(n443), .A2(n444), .ZN(n452) );
  NAND2_X1 U169 ( .A1(n441), .A2(n442), .ZN(n449) );
  INV_X1 U170 ( .A(A[38]), .ZN(n447) );
  AND2_X1 U171 ( .A1(n450), .A2(n451), .ZN(n443) );
  INV_X1 U172 ( .A(B[37]), .ZN(n445) );
  AND2_X1 U173 ( .A1(n449), .A2(n448), .ZN(n385) );
  INV_X1 U174 ( .A(B[38]), .ZN(n442) );
  XNOR2_X1 U175 ( .A(A[38]), .B(n442), .ZN(net182620) );
  CLKBUF_X1 U176 ( .A(n340), .Z(n453) );
  OR2_X1 U177 ( .A1(n493), .A2(n456), .ZN(n454) );
  AND2_X1 U178 ( .A1(n458), .A2(A[60]), .ZN(n455) );
  AND2_X1 U179 ( .A1(A[54]), .A2(n340), .ZN(n456) );
  AND2_X1 U180 ( .A1(n491), .A2(n458), .ZN(n457) );
  OR2_X1 U181 ( .A1(A[59]), .A2(B[59]), .ZN(n458) );
  NAND2_X1 U182 ( .A1(n491), .A2(n458), .ZN(n332) );
  INV_X1 U183 ( .A(n461), .ZN(n459) );
  XOR2_X1 U184 ( .A(A[40]), .B(B[40]), .Z(n384) );
  CLKBUF_X1 U185 ( .A(net176961), .Z(net185823) );
  AOI21_X1 U186 ( .B1(n481), .B2(n478), .A(n498), .ZN(n461) );
  AOI21_X1 U187 ( .B1(n453), .B2(n337), .A(n460), .ZN(n462) );
  CLKBUF_X1 U188 ( .A(n385), .Z(net184547) );
  INV_X1 U189 ( .A(n466), .ZN(n382) );
  NOR2_X1 U190 ( .A1(n463), .A2(A[51]), .ZN(n483) );
  OR2_X1 U191 ( .A1(net176961), .A2(net183785), .ZN(n463) );
  OR2_X1 U192 ( .A1(net176961), .A2(net183785), .ZN(n465) );
  NOR2_X1 U193 ( .A1(n467), .A2(n386), .ZN(n466) );
  NOR2_X1 U194 ( .A1(n385), .A2(A[39]), .ZN(n467) );
  CLKBUF_X1 U195 ( .A(n379), .Z(n481) );
  CLKBUF_X1 U196 ( .A(A[28]), .Z(n468) );
  INV_X1 U197 ( .A(n317), .ZN(n469) );
  CLKBUF_X1 U198 ( .A(A[35]), .Z(n470) );
  INV_X1 U199 ( .A(n501), .ZN(n472) );
  OR2_X1 U200 ( .A1(n508), .A2(n400), .ZN(n473) );
  NAND2_X1 U201 ( .A1(n401), .A2(n473), .ZN(n397) );
  XOR2_X1 U202 ( .A(carry[28]), .B(B[28]), .Z(n474) );
  XOR2_X1 U203 ( .A(n468), .B(n474), .Z(SUM[28]) );
  NAND2_X1 U204 ( .A1(n468), .A2(carry[28]), .ZN(n475) );
  NAND2_X1 U205 ( .A1(A[28]), .A2(B[28]), .ZN(n476) );
  NAND2_X1 U206 ( .A1(carry[28]), .A2(B[28]), .ZN(n477) );
  NAND3_X1 U207 ( .A1(n476), .A2(n475), .A3(n477), .ZN(carry[29]) );
  XNOR2_X1 U208 ( .A(n479), .B(n485), .ZN(SUM[53]) );
  XNOR2_X1 U209 ( .A(B[53]), .B(n503), .ZN(n479) );
  AND2_X1 U210 ( .A1(n506), .A2(n461), .ZN(n480) );
  NOR2_X1 U211 ( .A1(n377), .A2(n480), .ZN(n374) );
  XNOR2_X1 U212 ( .A(n459), .B(n489), .ZN(SUM[42]) );
  NOR2_X1 U213 ( .A1(n350), .A2(n483), .ZN(n346) );
  XNOR2_X1 U214 ( .A(net184550), .B(net182620), .ZN(SUM[38]) );
  XNOR2_X1 U215 ( .A(n487), .B(n472), .ZN(SUM[34]) );
  INV_X1 U216 ( .A(A[34]), .ZN(n508) );
  INV_X1 U217 ( .A(A[53]), .ZN(n503) );
  INV_X1 U218 ( .A(A[51]), .ZN(n504) );
  INV_X1 U219 ( .A(n376), .ZN(n497) );
  OAI21_X1 U220 ( .B1(n501), .B2(A[34]), .A(B[34]), .ZN(n401) );
  XNOR2_X1 U221 ( .A(n504), .B(B[51]), .ZN(n351) );
  XNOR2_X1 U222 ( .A(n471), .B(n488), .ZN(SUM[35]) );
  XNOR2_X1 U223 ( .A(A[35]), .B(B[35]), .ZN(n488) );
  XNOR2_X1 U224 ( .A(A[42]), .B(B[42]), .ZN(n489) );
  INV_X1 U225 ( .A(A[43]), .ZN(n505) );
  XNOR2_X1 U226 ( .A(n490), .B(n296), .ZN(SUM[59]) );
  XNOR2_X1 U227 ( .A(\carry[59] ), .B(B[59]), .ZN(n490) );
  OAI21_X1 U228 ( .B1(n470), .B2(n471), .A(n500), .ZN(n394) );
  INV_X1 U229 ( .A(n398), .ZN(n500) );
  AOI21_X1 U230 ( .B1(n397), .B2(A[35]), .A(B[35]), .ZN(n398) );
  OAI21_X1 U231 ( .B1(n499), .B2(n469), .A(B[36]), .ZN(n395) );
  INV_X1 U232 ( .A(n394), .ZN(n499) );
  AOI21_X1 U233 ( .B1(n481), .B2(n478), .A(n498), .ZN(n376) );
  INV_X1 U234 ( .A(n380), .ZN(n498) );
  XNOR2_X1 U235 ( .A(n332), .B(n333), .ZN(SUM[60]) );
  XNOR2_X1 U236 ( .A(n408), .B(n375), .ZN(SUM[43]) );
  XNOR2_X1 U237 ( .A(B[55]), .B(n502), .ZN(n339) );
  OAI21_X1 U238 ( .B1(net183931), .B2(n403), .A(net176946), .ZN(n400) );
  INV_X1 U239 ( .A(A[42]), .ZN(n506) );
  AOI21_X1 U240 ( .B1(n497), .B2(A[42]), .A(B[42]), .ZN(n377) );
  INV_X1 U241 ( .A(n334), .ZN(n491) );
  AOI21_X1 U242 ( .B1(A[59]), .B2(B[59]), .A(\carry[59] ), .ZN(n334) );
  XNOR2_X1 U243 ( .A(n411), .B(net185657), .ZN(SUM[31]) );
  AND2_X1 U244 ( .A1(A[0]), .A2(B[0]), .ZN(n1) );
  AOI21_X1 U245 ( .B1(n466), .B2(A[40]), .A(B[40]), .ZN(n383) );
  INV_X1 U246 ( .A(A[40]), .ZN(n507) );
  AOI21_X1 U247 ( .B1(n440), .B2(A[39]), .A(B[39]), .ZN(n386) );
  XNOR2_X1 U248 ( .A(n381), .B(n481), .ZN(SUM[41]) );
  XNOR2_X1 U249 ( .A(n384), .B(n382), .ZN(SUM[40]) );
  AOI21_X1 U250 ( .B1(n507), .B2(n382), .A(n383), .ZN(n379) );
  INV_X1 U251 ( .A(n400), .ZN(n501) );
  INV_X1 U252 ( .A(A[55]), .ZN(n502) );
  AOI21_X1 U253 ( .B1(n502), .B2(n462), .A(n338), .ZN(n327) );
  AOI21_X1 U254 ( .B1(A[55]), .B2(n454), .A(B[55]), .ZN(n338) );
  XNOR2_X1 U255 ( .A(n295), .B(n351), .ZN(SUM[51]) );
  OAI21_X1 U256 ( .B1(n300), .B2(n505), .A(n373), .ZN(n370) );
  INV_X1 U257 ( .A(n371), .ZN(n496) );
  AOI21_X1 U258 ( .B1(A[53]), .B2(n494), .A(B[53]), .ZN(n344) );
  OAI22_X1 U259 ( .A1(n331), .A2(B[60]), .B1(n457), .B2(A[60]), .ZN(n329) );
  AND2_X1 U260 ( .A1(n491), .A2(n455), .ZN(n331) );
  XNOR2_X1 U261 ( .A(n339), .B(n301), .ZN(SUM[55]) );
  AOI21_X1 U262 ( .B1(n503), .B2(n485), .A(n344), .ZN(n340) );
  OAI21_X1 U263 ( .B1(n484), .B2(n464), .A(n496), .ZN(n367) );
  AOI21_X1 U264 ( .B1(n370), .B2(A[44]), .A(B[44]), .ZN(n371) );
  OAI21_X1 U265 ( .B1(n374), .B2(A[43]), .A(B[43]), .ZN(n373) );
  XNOR2_X1 U266 ( .A(n478), .B(B[41]), .ZN(n381) );
  OAI21_X1 U267 ( .B1(n379), .B2(A[41]), .A(B[41]), .ZN(n380) );
  INV_X1 U268 ( .A(n326), .ZN(n492) );
  OAI21_X1 U269 ( .B1(n346), .B2(A[52]), .A(B[52]), .ZN(n347) );
  AOI21_X1 U270 ( .B1(n465), .B2(A[51]), .A(B[51]), .ZN(n350) );
  AOI22_X1 U271 ( .A1(n482), .A2(n486), .B1(n328), .B2(B[56]), .ZN(n326) );
  OR2_X1 U272 ( .A1(n327), .A2(A[56]), .ZN(n328) );
  INV_X1 U273 ( .A(n347), .ZN(n495) );
  INV_X1 U274 ( .A(n353), .ZN(net176961) );
endmodule


module RCA_NBIT62 ( A, B, Ci, S, Co );
  input [61:0] A;
  input [61:0] B;
  output [61:0] S;
  input Ci;
  output Co;

  assign Co = 1'b0;

  RCA_NBIT62_DW01_add_0 add_95 ( .A(A), .B(B), .CI(1'b0), .SUM(S) );
endmodule


module RCA_NBIT64_DW01_add_0 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1, net50029, n423, n424, n427, n428, n431, n432, n433, n434, n435,
         n436, n437, n439, n440, n441, n443, n444, n445, n446, n448, n449,
         n451, n452, n454, n455, n457, n458, n460, n461, n463, n464, n466,
         n467, n469, n470, n473, n474, n475, n476, n479, n481, n482, n485,
         n487, n488, n490, n491, n493, n494, n496, n497, n500, n502, n503,
         n505, n506, n508, n509, n510, n511, n512, n514, n515, n516, n517,
         n518, n519, n520, n521, net182739, net183790, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n425, n426,
         n429, n430, n438, n442, n447, n450, n453, n456, n459, n462, n465,
         n468, n471, n472, n477, n478, n480, n483, n484, n486, n489, n492,
         n495, n498, n499, n501, n504, n507, n513, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613;
  wire   [63:1] carry;
  assign net50029 = A[55];

  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U131 ( .A(n410), .B(n423), .Z(SUM[61]) );
  XOR2_X1 U134 ( .A(n432), .B(n545), .Z(SUM[58]) );
  OAI33_X1 U135 ( .A1(n456), .A2(n612), .A3(n613), .B1(n437), .B2(n603), .B3(
        n612), .ZN(n435) );
  XOR2_X1 U136 ( .A(n439), .B(n440), .Z(SUM[57]) );
  XOR2_X1 U137 ( .A(n541), .B(B[57]), .Z(n440) );
  XOR2_X1 U140 ( .A(n456), .B(n444), .Z(SUM[55]) );
  XOR2_X1 U141 ( .A(n603), .B(B[55]), .Z(n444) );
  XOR2_X1 U160 ( .A(n407), .B(n474), .Z(SUM[45]) );
  XOR2_X1 U161 ( .A(B[45]), .B(A[45]), .Z(n474) );
  XOR2_X1 U184 ( .A(n527), .B(n510), .Z(SUM[33]) );
  XOR2_X1 U185 ( .A(B[33]), .B(n535), .Z(n510) );
  XOR2_X1 U187 ( .A(n379), .B(n515), .Z(SUM[31]) );
  XOR2_X1 U188 ( .A(B[31]), .B(n480), .Z(n515) );
  XOR2_X1 U189 ( .A(n597), .B(n518), .Z(SUM[30]) );
  XOR2_X1 U190 ( .A(B[30]), .B(A[30]), .Z(n518) );
  XOR2_X1 U191 ( .A(A[29]), .B(n521), .Z(SUM[29]) );
  XOR2_X1 U192 ( .A(carry[29]), .B(B[29]), .Z(n521) );
  XOR2_X1 U193 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  CLKBUF_X1 U1 ( .A(n443), .Z(n366) );
  CLKBUF_X1 U2 ( .A(n487), .Z(n529) );
  CLKBUF_X1 U3 ( .A(n469), .Z(n550) );
  CLKBUF_X1 U4 ( .A(A[43]), .Z(n367) );
  NAND2_X1 U5 ( .A1(A[38]), .A2(n591), .ZN(n534) );
  NAND2_X1 U6 ( .A1(A[36]), .A2(n368), .ZN(n402) );
  NOR2_X1 U7 ( .A1(n395), .A2(n503), .ZN(n368) );
  NOR2_X1 U8 ( .A1(n395), .A2(n503), .ZN(n369) );
  OR2_X1 U9 ( .A1(n472), .A2(n610), .ZN(n370) );
  INV_X1 U10 ( .A(n421), .ZN(n371) );
  BUF_X1 U11 ( .A(A[40]), .Z(n486) );
  CLKBUF_X1 U12 ( .A(n585), .Z(n372) );
  BUF_X1 U13 ( .A(A[31]), .Z(n480) );
  OR2_X1 U14 ( .A1(n469), .A2(A[46]), .ZN(n373) );
  OR2_X1 U15 ( .A1(n469), .A2(A[46]), .ZN(n470) );
  CLKBUF_X1 U16 ( .A(n529), .Z(n374) );
  INV_X1 U17 ( .A(B[61]), .ZN(n413) );
  INV_X1 U18 ( .A(B[62]), .ZN(n425) );
  XOR2_X1 U19 ( .A(A[62]), .B(B[62]), .Z(n375) );
  XNOR2_X1 U20 ( .A(n409), .B(n376), .ZN(SUM[60]) );
  XOR2_X1 U21 ( .A(B[60]), .B(n450), .Z(n376) );
  BUF_X1 U22 ( .A(A[61]), .Z(n377) );
  CLKBUF_X1 U23 ( .A(n550), .Z(n378) );
  CLKBUF_X1 U24 ( .A(n596), .Z(n379) );
  AND2_X1 U25 ( .A1(n386), .A2(n385), .ZN(n380) );
  CLKBUF_X1 U26 ( .A(A[42]), .Z(n381) );
  CLKBUF_X1 U27 ( .A(A[44]), .Z(n382) );
  CLKBUF_X1 U28 ( .A(A[41]), .Z(n383) );
  OR2_X1 U29 ( .A1(n436), .A2(n613), .ZN(n551) );
  NOR2_X1 U30 ( .A1(n384), .A2(A[43]), .ZN(n539) );
  OR2_X1 U31 ( .A1(n589), .A2(n548), .ZN(n384) );
  NAND2_X1 U32 ( .A1(n529), .A2(n486), .ZN(n385) );
  NAND2_X1 U33 ( .A1(n488), .A2(B[40]), .ZN(n386) );
  NAND2_X1 U34 ( .A1(n386), .A2(n385), .ZN(n387) );
  AND2_X1 U35 ( .A1(n388), .A2(A[56]), .ZN(n434) );
  NAND3_X1 U36 ( .A1(n443), .A2(n551), .A3(n612), .ZN(n388) );
  OR2_X1 U37 ( .A1(n584), .A2(n549), .ZN(n389) );
  OR2_X1 U38 ( .A1(n584), .A2(n549), .ZN(n537) );
  CLKBUF_X1 U39 ( .A(n589), .Z(n390) );
  CLKBUF_X1 U40 ( .A(n586), .Z(n391) );
  OR2_X1 U41 ( .A1(n390), .A2(n548), .ZN(n392) );
  OR2_X1 U42 ( .A1(n372), .A2(n525), .ZN(n393) );
  CLKBUF_X1 U43 ( .A(n496), .Z(n468) );
  CLKBUF_X1 U44 ( .A(n554), .Z(n394) );
  NOR2_X1 U45 ( .A1(n399), .A2(A[35]), .ZN(n395) );
  INV_X1 U46 ( .A(n489), .ZN(n396) );
  INV_X1 U47 ( .A(n472), .ZN(n397) );
  BUF_X1 U48 ( .A(n505), .Z(n472) );
  INV_X1 U49 ( .A(n499), .ZN(n398) );
  NAND2_X1 U50 ( .A1(n370), .A2(n506), .ZN(n399) );
  INV_X1 U51 ( .A(n590), .ZN(n400) );
  OR2_X1 U52 ( .A1(n589), .A2(n548), .ZN(n401) );
  NAND2_X1 U53 ( .A1(n500), .A2(n402), .ZN(n496) );
  AND2_X1 U54 ( .A1(n405), .A2(n420), .ZN(n403) );
  NAND2_X1 U55 ( .A1(n450), .A2(B[60]), .ZN(n404) );
  BUF_X2 U56 ( .A(A[60]), .Z(n450) );
  NAND2_X1 U57 ( .A1(n422), .A2(n429), .ZN(n405) );
  OR2_X1 U58 ( .A1(n513), .A2(n588), .ZN(n406) );
  OR2_X1 U59 ( .A1(n513), .A2(n588), .ZN(n407) );
  CLKBUF_X1 U60 ( .A(n369), .Z(n408) );
  INV_X1 U61 ( .A(n411), .ZN(n421) );
  CLKBUF_X1 U62 ( .A(n422), .Z(n409) );
  CLKBUF_X1 U63 ( .A(net183790), .Z(n410) );
  XNOR2_X1 U64 ( .A(n414), .B(n375), .ZN(SUM[62]) );
  NOR2_X1 U65 ( .A1(n453), .A2(n403), .ZN(n414) );
  INV_X1 U66 ( .A(n424), .ZN(n422) );
  NAND2_X1 U67 ( .A1(n450), .A2(B[60]), .ZN(n429) );
  NAND2_X1 U68 ( .A1(n430), .A2(n377), .ZN(n418) );
  XNOR2_X1 U69 ( .A(A[61]), .B(B[61]), .ZN(n423) );
  INV_X1 U70 ( .A(A[62]), .ZN(n426) );
  NOR2_X1 U71 ( .A1(B[62]), .A2(A[62]), .ZN(n415) );
  AOI21_X1 U72 ( .B1(n417), .B2(n418), .A(n415), .ZN(n416) );
  XNOR2_X1 U73 ( .A(n416), .B(n419), .ZN(SUM[63]) );
  NAND2_X1 U74 ( .A1(n422), .A2(n404), .ZN(n412) );
  NAND2_X1 U75 ( .A1(n405), .A2(n420), .ZN(n438) );
  NAND2_X1 U76 ( .A1(n412), .A2(n371), .ZN(net183790) );
  NAND2_X1 U77 ( .A1(n438), .A2(n426), .ZN(n447) );
  NAND2_X1 U78 ( .A1(n438), .A2(n425), .ZN(n442) );
  NAND2_X1 U79 ( .A1(net183790), .A2(n413), .ZN(n430) );
  AND2_X1 U80 ( .A1(n430), .A2(n377), .ZN(n453) );
  NAND2_X1 U81 ( .A1(n447), .A2(n442), .ZN(n417) );
  NOR2_X1 U82 ( .A1(n413), .A2(n421), .ZN(n420) );
  INV_X1 U83 ( .A(net182739), .ZN(n419) );
  OR2_X1 U84 ( .A1(A[60]), .A2(B[60]), .ZN(n411) );
  INV_X1 U85 ( .A(n582), .ZN(n456) );
  CLKBUF_X1 U86 ( .A(A[36]), .Z(n459) );
  CLKBUF_X1 U87 ( .A(n457), .Z(n462) );
  OR2_X1 U88 ( .A1(n524), .A2(n391), .ZN(n465) );
  OR2_X1 U89 ( .A1(n586), .A2(n524), .ZN(n471) );
  CLKBUF_X1 U90 ( .A(A[38]), .Z(n477) );
  OAI21_X1 U91 ( .B1(n582), .B2(B[55]), .A(net50029), .ZN(n478) );
  OR2_X1 U92 ( .A1(n431), .A2(n546), .ZN(n483) );
  CLKBUF_X1 U93 ( .A(A[37]), .Z(n484) );
  AOI22_X1 U94 ( .A1(n550), .A2(A[46]), .B1(n373), .B2(B[46]), .ZN(n489) );
  CLKBUF_X1 U95 ( .A(n468), .Z(n492) );
  CLKBUF_X1 U96 ( .A(A[34]), .Z(n495) );
  CLKBUF_X1 U97 ( .A(n463), .Z(n498) );
  INV_X1 U98 ( .A(n595), .ZN(n499) );
  NOR2_X1 U99 ( .A1(n441), .A2(B[56]), .ZN(n501) );
  AND2_X1 U100 ( .A1(n583), .A2(n556), .ZN(n504) );
  BUF_X1 U101 ( .A(A[57]), .Z(n522) );
  CLKBUF_X1 U102 ( .A(n399), .Z(n507) );
  AND2_X1 U103 ( .A1(n554), .A2(A[44]), .ZN(n513) );
  BUF_X1 U104 ( .A(n475), .Z(n554) );
  OR2_X1 U105 ( .A1(n585), .A2(n525), .ZN(n523) );
  AND2_X1 U106 ( .A1(n463), .A2(A[48]), .ZN(n524) );
  NOR2_X1 U107 ( .A1(n524), .A2(n586), .ZN(n460) );
  AND2_X1 U108 ( .A1(n457), .A2(A[50]), .ZN(n525) );
  NOR2_X1 U109 ( .A1(n525), .A2(n585), .ZN(n454) );
  INV_X1 U110 ( .A(n407), .ZN(n526) );
  BUF_X1 U111 ( .A(n508), .Z(n527) );
  OR2_X1 U112 ( .A1(n472), .A2(n610), .ZN(n528) );
  NAND2_X1 U113 ( .A1(n528), .A2(n506), .ZN(n502) );
  CLKBUF_X1 U114 ( .A(n451), .Z(n530) );
  CLKBUF_X1 U115 ( .A(n445), .Z(n531) );
  CLKBUF_X1 U116 ( .A(n591), .Z(n532) );
  INV_X1 U117 ( .A(n380), .ZN(n533) );
  NAND2_X1 U118 ( .A1(n534), .A2(n494), .ZN(n491) );
  CLKBUF_X1 U119 ( .A(A[33]), .Z(n535) );
  NAND2_X1 U120 ( .A1(n551), .A2(n478), .ZN(n536) );
  AND2_X1 U121 ( .A1(n607), .A2(n489), .ZN(n538) );
  NOR2_X1 U122 ( .A1(n467), .A2(n538), .ZN(n463) );
  NOR2_X1 U123 ( .A1(n479), .A2(n539), .ZN(n475) );
  INV_X1 U124 ( .A(n609), .ZN(n540) );
  CLKBUF_X1 U125 ( .A(n522), .Z(n541) );
  AND2_X1 U126 ( .A1(n604), .A2(n448), .ZN(n542) );
  NOR2_X1 U127 ( .A1(n449), .A2(n542), .ZN(n445) );
  CLKBUF_X1 U128 ( .A(n481), .Z(n555) );
  CLKBUF_X1 U129 ( .A(A[58]), .Z(n543) );
  OR2_X1 U130 ( .A1(n580), .A2(n547), .ZN(n544) );
  NOR2_X1 U132 ( .A1(n547), .A2(n580), .ZN(n545) );
  AND2_X1 U133 ( .A1(n601), .A2(n545), .ZN(n546) );
  NOR2_X1 U138 ( .A1(n546), .A2(n431), .ZN(n428) );
  AND2_X1 U139 ( .A1(n522), .A2(B[57]), .ZN(n547) );
  AND2_X1 U142 ( .A1(n481), .A2(A[42]), .ZN(n548) );
  AND2_X1 U143 ( .A1(n451), .A2(A[52]), .ZN(n549) );
  NOR2_X1 U144 ( .A1(n549), .A2(n584), .ZN(n448) );
  NAND2_X1 U145 ( .A1(n366), .A2(n551), .ZN(n441) );
  AND2_X1 U146 ( .A1(n605), .A2(n454), .ZN(n552) );
  NOR2_X1 U147 ( .A1(n455), .A2(n552), .ZN(n451) );
  AND2_X1 U148 ( .A1(n460), .A2(n606), .ZN(n553) );
  NOR2_X1 U149 ( .A1(n461), .A2(n553), .ZN(n457) );
  OR2_X1 U150 ( .A1(n445), .A2(A[54]), .ZN(n556) );
  NAND2_X1 U151 ( .A1(n583), .A2(n556), .ZN(n436) );
  XOR2_X1 U152 ( .A(B[63]), .B(A[63]), .Z(net182739) );
  XOR2_X1 U153 ( .A(n530), .B(n557), .Z(SUM[52]) );
  XOR2_X1 U154 ( .A(B[52]), .B(A[52]), .Z(n557) );
  XOR2_X1 U155 ( .A(n462), .B(n558), .Z(SUM[50]) );
  XOR2_X1 U156 ( .A(B[50]), .B(A[50]), .Z(n558) );
  XOR2_X1 U157 ( .A(n378), .B(n559), .Z(SUM[46]) );
  XOR2_X1 U158 ( .A(B[46]), .B(A[46]), .Z(n559) );
  XOR2_X1 U159 ( .A(n507), .B(n560), .Z(SUM[35]) );
  XOR2_X1 U162 ( .A(B[35]), .B(A[35]), .Z(n560) );
  XOR2_X1 U163 ( .A(n397), .B(n561), .Z(SUM[34]) );
  XOR2_X1 U164 ( .A(B[34]), .B(n495), .Z(n561) );
  INV_X1 U165 ( .A(A[32]), .ZN(n611) );
  INV_X1 U166 ( .A(A[56]), .ZN(n602) );
  INV_X1 U167 ( .A(A[59]), .ZN(n600) );
  INV_X1 U168 ( .A(n493), .ZN(n591) );
  INV_X1 U169 ( .A(n505), .ZN(n593) );
  INV_X1 U170 ( .A(A[47]), .ZN(n607) );
  INV_X1 U171 ( .A(A[41]), .ZN(n599) );
  INV_X1 U172 ( .A(A[34]), .ZN(n610) );
  OAI21_X1 U173 ( .B1(n593), .B2(A[34]), .A(B[34]), .ZN(n506) );
  INV_X1 U174 ( .A(n482), .ZN(n589) );
  OAI21_X1 U175 ( .B1(n369), .B2(A[36]), .A(B[36]), .ZN(n500) );
  OAI21_X1 U176 ( .B1(n591), .B2(A[38]), .A(B[38]), .ZN(n494) );
  OAI21_X1 U177 ( .B1(n499), .B2(n611), .A(n512), .ZN(n508) );
  OAI21_X1 U178 ( .B1(n595), .B2(A[32]), .A(B[32]), .ZN(n512) );
  AOI21_X1 U179 ( .B1(n600), .B2(n483), .A(n427), .ZN(n424) );
  OAI21_X1 U180 ( .B1(n484), .B2(n468), .A(n592), .ZN(n493) );
  INV_X1 U181 ( .A(n497), .ZN(n592) );
  AOI21_X1 U182 ( .B1(n496), .B2(A[37]), .A(B[37]), .ZN(n497) );
  AOI21_X1 U183 ( .B1(n609), .B2(n590), .A(n490), .ZN(n487) );
  INV_X1 U186 ( .A(A[39]), .ZN(n609) );
  INV_X1 U194 ( .A(n491), .ZN(n590) );
  AOI21_X1 U195 ( .B1(n491), .B2(A[39]), .A(B[39]), .ZN(n490) );
  OAI21_X1 U196 ( .B1(n535), .B2(n527), .A(n594), .ZN(n505) );
  INV_X1 U197 ( .A(n509), .ZN(n594) );
  AOI21_X1 U198 ( .B1(n508), .B2(A[33]), .A(B[33]), .ZN(n509) );
  INV_X1 U199 ( .A(A[49]), .ZN(n606) );
  INV_X1 U200 ( .A(A[51]), .ZN(n605) );
  INV_X1 U201 ( .A(A[45]), .ZN(n608) );
  AOI21_X1 U202 ( .B1(n406), .B2(A[45]), .A(B[45]), .ZN(n473) );
  XNOR2_X1 U203 ( .A(n562), .B(n483), .ZN(SUM[59]) );
  XNOR2_X1 U204 ( .A(n600), .B(B[59]), .ZN(n562) );
  NOR2_X1 U205 ( .A1(B[55]), .A2(n504), .ZN(n437) );
  INV_X1 U206 ( .A(n511), .ZN(n595) );
  INV_X1 U207 ( .A(A[58]), .ZN(n601) );
  INV_X1 U208 ( .A(n452), .ZN(n584) );
  XNOR2_X1 U209 ( .A(n393), .B(n563), .ZN(SUM[51]) );
  XNOR2_X1 U210 ( .A(B[51]), .B(A[51]), .ZN(n563) );
  XNOR2_X1 U211 ( .A(n389), .B(n564), .ZN(SUM[53]) );
  XNOR2_X1 U212 ( .A(B[53]), .B(A[53]), .ZN(n564) );
  XNOR2_X1 U213 ( .A(n543), .B(B[58]), .ZN(n432) );
  XNOR2_X1 U214 ( .A(n531), .B(n565), .ZN(SUM[54]) );
  XNOR2_X1 U215 ( .A(A[54]), .B(B[54]), .ZN(n565) );
  OAI22_X1 U216 ( .A1(n581), .A2(n612), .B1(n501), .B2(n602), .ZN(n439) );
  XNOR2_X1 U217 ( .A(n536), .B(n566), .ZN(SUM[56]) );
  XNOR2_X1 U218 ( .A(B[56]), .B(A[56]), .ZN(n566) );
  XNOR2_X1 U219 ( .A(n396), .B(n567), .ZN(SUM[47]) );
  XNOR2_X1 U220 ( .A(B[47]), .B(A[47]), .ZN(n567) );
  XNOR2_X1 U221 ( .A(n568), .B(n498), .ZN(SUM[48]) );
  XNOR2_X1 U222 ( .A(B[48]), .B(A[48]), .ZN(n568) );
  XNOR2_X1 U223 ( .A(n465), .B(n569), .ZN(SUM[49]) );
  XNOR2_X1 U224 ( .A(B[49]), .B(A[49]), .ZN(n569) );
  XNOR2_X1 U225 ( .A(n392), .B(n570), .ZN(SUM[43]) );
  XNOR2_X1 U226 ( .A(n367), .B(B[43]), .ZN(n570) );
  XNOR2_X1 U227 ( .A(n394), .B(n571), .ZN(SUM[44]) );
  XNOR2_X1 U228 ( .A(n382), .B(B[44]), .ZN(n571) );
  XNOR2_X1 U229 ( .A(n555), .B(n572), .ZN(SUM[42]) );
  XNOR2_X1 U230 ( .A(n381), .B(B[42]), .ZN(n572) );
  XNOR2_X1 U231 ( .A(n533), .B(n573), .ZN(SUM[41]) );
  XNOR2_X1 U232 ( .A(B[41]), .B(n383), .ZN(n573) );
  XNOR2_X1 U233 ( .A(n408), .B(n574), .ZN(SUM[36]) );
  XNOR2_X1 U234 ( .A(B[36]), .B(n459), .ZN(n574) );
  XNOR2_X1 U235 ( .A(n532), .B(n575), .ZN(SUM[38]) );
  XNOR2_X1 U236 ( .A(B[38]), .B(n477), .ZN(n575) );
  XNOR2_X1 U237 ( .A(n398), .B(n576), .ZN(SUM[32]) );
  XOR2_X1 U238 ( .A(B[32]), .B(n611), .Z(n576) );
  XNOR2_X1 U239 ( .A(n374), .B(n577), .ZN(SUM[40]) );
  XNOR2_X1 U240 ( .A(B[40]), .B(n486), .ZN(n577) );
  XNOR2_X1 U241 ( .A(n400), .B(n578), .ZN(SUM[39]) );
  XNOR2_X1 U242 ( .A(B[39]), .B(n540), .ZN(n578) );
  XNOR2_X1 U243 ( .A(n492), .B(n579), .ZN(SUM[37]) );
  XNOR2_X1 U244 ( .A(B[37]), .B(n484), .ZN(n579) );
  INV_X1 U245 ( .A(B[56]), .ZN(n612) );
  INV_X1 U246 ( .A(B[55]), .ZN(n613) );
  OAI22_X1 U247 ( .A1(n480), .A2(n379), .B1(n514), .B2(B[31]), .ZN(n511) );
  AND2_X1 U248 ( .A1(A[31]), .A2(n596), .ZN(n514) );
  INV_X1 U249 ( .A(n516), .ZN(n596) );
  OAI22_X1 U250 ( .A1(A[30]), .A2(n597), .B1(B[30]), .B2(n517), .ZN(n516) );
  AND2_X1 U251 ( .A1(n597), .A2(A[30]), .ZN(n517) );
  INV_X1 U252 ( .A(n519), .ZN(n597) );
  OAI21_X1 U253 ( .B1(B[29]), .B2(A[29]), .A(n598), .ZN(n519) );
  INV_X1 U254 ( .A(n520), .ZN(n598) );
  AOI21_X1 U255 ( .B1(A[29]), .B2(B[29]), .A(carry[29]), .ZN(n520) );
  AND2_X1 U256 ( .A1(A[0]), .A2(B[0]), .ZN(n1) );
  AOI21_X1 U257 ( .B1(n502), .B2(A[35]), .A(B[35]), .ZN(n503) );
  OAI21_X1 U258 ( .B1(n457), .B2(A[50]), .A(B[50]), .ZN(n458) );
  AOI21_X1 U259 ( .B1(n608), .B2(n526), .A(n473), .ZN(n469) );
  INV_X1 U260 ( .A(n536), .ZN(n581) );
  OAI21_X1 U261 ( .B1(n481), .B2(A[42]), .A(B[42]), .ZN(n482) );
  INV_X1 U262 ( .A(A[53]), .ZN(n604) );
  AOI21_X1 U263 ( .B1(n445), .B2(A[54]), .A(B[54]), .ZN(n446) );
  INV_X1 U264 ( .A(n464), .ZN(n586) );
  INV_X1 U265 ( .A(n466), .ZN(n587) );
  INV_X1 U266 ( .A(n476), .ZN(n588) );
  OAI21_X1 U267 ( .B1(A[44]), .B2(n475), .A(B[44]), .ZN(n476) );
  INV_X1 U268 ( .A(n436), .ZN(n582) );
  OAI21_X1 U269 ( .B1(n451), .B2(A[52]), .A(B[52]), .ZN(n452) );
  OAI21_X1 U270 ( .B1(n463), .B2(A[48]), .A(B[48]), .ZN(n464) );
  INV_X1 U271 ( .A(net50029), .ZN(n603) );
  INV_X1 U272 ( .A(n458), .ZN(n585) );
  OAI21_X1 U273 ( .B1(n504), .B2(B[55]), .A(net50029), .ZN(n443) );
  OR2_X1 U274 ( .A1(n487), .A2(A[40]), .ZN(n488) );
  AOI22_X1 U275 ( .A1(n550), .A2(A[46]), .B1(n470), .B2(B[46]), .ZN(n466) );
  AOI21_X1 U276 ( .B1(n523), .B2(A[51]), .A(B[51]), .ZN(n455) );
  AOI21_X1 U277 ( .B1(n471), .B2(A[49]), .A(B[49]), .ZN(n461) );
  AOI21_X1 U278 ( .B1(n401), .B2(A[43]), .A(B[43]), .ZN(n479) );
  AOI21_X1 U279 ( .B1(n587), .B2(A[47]), .A(B[47]), .ZN(n467) );
  AOI21_X1 U280 ( .B1(n599), .B2(n380), .A(n485), .ZN(n481) );
  AOI21_X1 U281 ( .B1(n387), .B2(A[41]), .A(B[41]), .ZN(n485) );
  AOI21_X1 U282 ( .B1(n537), .B2(A[53]), .A(B[53]), .ZN(n449) );
  INV_X1 U283 ( .A(n446), .ZN(n583) );
  INV_X1 U284 ( .A(n433), .ZN(n580) );
  AOI21_X1 U285 ( .B1(n544), .B2(A[58]), .A(B[58]), .ZN(n431) );
  OAI22_X1 U286 ( .A1(n434), .A2(n435), .B1(A[57]), .B2(B[57]), .ZN(n433) );
  AOI21_X1 U287 ( .B1(n428), .B2(A[59]), .A(B[59]), .ZN(n427) );
endmodule


module RCA_NBIT64 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;

  assign Co = 1'b0;

  RCA_NBIT64_DW01_add_0 add_95 ( .A(A), .B(B), .CI(1'b0), .SUM(S) );
endmodule


module BOOTHMUL_NBIT32_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n96, n97, n98, n100, n102, n103, n104, n106, n107, n108, n110,
         n111, n112, n114, n115, n116, n118, n119, n120, n122, n123, n124, n94,
         n95, n99, n101, n105, n109, n113, n117, n121, n125, n126, n127;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U42 ( .A(n96), .B(B[30]), .Z(DIFF[30]) );
  XOR2_X1 U43 ( .A(n98), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U45 ( .A(n100), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U46 ( .A(n102), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U48 ( .A(n104), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U49 ( .A(n106), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U51 ( .A(n108), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U52 ( .A(n110), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U54 ( .A(n112), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U55 ( .A(n114), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U57 ( .A(n116), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U58 ( .A(n118), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U60 ( .A(n120), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U61 ( .A(n122), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U62 ( .A(\B[0] ), .B(B[1]), .Z(DIFF[1]) );
  NAND3_X1 U1 ( .A1(n94), .A2(n95), .A3(n99), .ZN(n122) );
  INV_X1 U2 ( .A(\B[0] ), .ZN(n94) );
  INV_X1 U3 ( .A(B[2]), .ZN(n95) );
  INV_X1 U4 ( .A(B[1]), .ZN(n99) );
  OR3_X1 U5 ( .A1(B[3]), .A2(B[4]), .A3(n122), .ZN(n120) );
  XOR2_X1 U6 ( .A(n101), .B(B[26]), .Z(DIFF[26]) );
  OR2_X1 U7 ( .A1(n100), .A2(B[25]), .ZN(n101) );
  XOR2_X1 U8 ( .A(n105), .B(B[22]), .Z(DIFF[22]) );
  OR2_X1 U9 ( .A1(n104), .A2(B[21]), .ZN(n105) );
  XOR2_X1 U10 ( .A(B[28]), .B(n109), .Z(DIFF[28]) );
  OR2_X1 U11 ( .A1(B[27]), .A2(n98), .ZN(n109) );
  XOR2_X1 U12 ( .A(n97), .B(n127), .Z(DIFF[29]) );
  NAND2_X1 U13 ( .A1(n97), .A2(n127), .ZN(n96) );
  XNOR2_X1 U14 ( .A(B[4]), .B(n123), .ZN(DIFF[4]) );
  NOR2_X1 U15 ( .A1(B[3]), .A2(n122), .ZN(n123) );
  XNOR2_X1 U16 ( .A(B[8]), .B(n119), .ZN(DIFF[8]) );
  NOR2_X1 U17 ( .A1(B[7]), .A2(n118), .ZN(n119) );
  XNOR2_X1 U18 ( .A(n124), .B(B[2]), .ZN(DIFF[2]) );
  NOR2_X1 U19 ( .A1(\B[0] ), .A2(B[1]), .ZN(n124) );
  OR3_X1 U20 ( .A1(B[5]), .A2(B[6]), .A3(n120), .ZN(n118) );
  OR3_X1 U21 ( .A1(B[7]), .A2(B[8]), .A3(n118), .ZN(n116) );
  XNOR2_X1 U22 ( .A(n113), .B(B[6]), .ZN(DIFF[6]) );
  NOR2_X1 U23 ( .A1(n120), .A2(B[5]), .ZN(n113) );
  XNOR2_X1 U24 ( .A(n117), .B(B[14]), .ZN(DIFF[14]) );
  NOR2_X1 U25 ( .A1(n112), .A2(B[13]), .ZN(n117) );
  XNOR2_X1 U26 ( .A(n121), .B(B[18]), .ZN(DIFF[18]) );
  NOR2_X1 U27 ( .A1(n108), .A2(B[17]), .ZN(n121) );
  XNOR2_X1 U28 ( .A(B[20]), .B(n107), .ZN(DIFF[20]) );
  NOR2_X1 U29 ( .A1(B[19]), .A2(n106), .ZN(n107) );
  XNOR2_X1 U30 ( .A(B[16]), .B(n111), .ZN(DIFF[16]) );
  NOR2_X1 U31 ( .A1(B[15]), .A2(n110), .ZN(n111) );
  XNOR2_X1 U32 ( .A(B[24]), .B(n103), .ZN(DIFF[24]) );
  NOR2_X1 U33 ( .A1(B[23]), .A2(n102), .ZN(n103) );
  XNOR2_X1 U34 ( .A(B[12]), .B(n115), .ZN(DIFF[12]) );
  NOR2_X1 U35 ( .A1(B[11]), .A2(n114), .ZN(n115) );
  OR3_X1 U36 ( .A1(B[21]), .A2(B[22]), .A3(n104), .ZN(n102) );
  OR3_X1 U37 ( .A1(B[17]), .A2(B[18]), .A3(n108), .ZN(n106) );
  OR3_X1 U38 ( .A1(B[13]), .A2(B[14]), .A3(n112), .ZN(n110) );
  OR3_X1 U39 ( .A1(B[10]), .A2(B[9]), .A3(n116), .ZN(n114) );
  OR3_X1 U40 ( .A1(B[19]), .A2(B[20]), .A3(n106), .ZN(n104) );
  OR3_X1 U41 ( .A1(B[15]), .A2(B[16]), .A3(n110), .ZN(n108) );
  OR3_X1 U44 ( .A1(B[11]), .A2(B[12]), .A3(n114), .ZN(n112) );
  XNOR2_X1 U47 ( .A(n125), .B(B[10]), .ZN(DIFF[10]) );
  NOR2_X1 U50 ( .A1(n116), .A2(B[9]), .ZN(n125) );
  NOR3_X1 U53 ( .A1(B[27]), .A2(B[28]), .A3(n98), .ZN(n97) );
  OR3_X1 U56 ( .A1(B[25]), .A2(B[26]), .A3(n100), .ZN(n98) );
  OR3_X1 U59 ( .A1(B[23]), .A2(B[24]), .A3(n102), .ZN(n100) );
  XNOR2_X1 U63 ( .A(n126), .B(B[31]), .ZN(DIFF[31]) );
  NOR2_X1 U64 ( .A1(n96), .A2(B[30]), .ZN(n126) );
  INV_X1 U65 ( .A(B[29]), .ZN(n127) );
endmodule


module BOOTHMUL_NBIT32 ( A, B, S );
  input [31:0] A;
  input [31:0] B;
  output [63:0] S;
  wire   A_n_65, \SHIFT[1][31] , \SHIFT[1][30] , \SHIFT[1][29] ,
         \SHIFT[1][28] , \SHIFT[1][27] , \SHIFT[1][26] , \SHIFT[1][25] ,
         \SHIFT[1][24] , \SHIFT[1][23] , \SHIFT[1][22] , \SHIFT[1][21] ,
         \SHIFT[1][20] , \SHIFT[1][19] , \SHIFT[1][18] , \SHIFT[1][17] ,
         \SHIFT[1][16] , \SHIFT[1][15] , \SHIFT[1][14] , \SHIFT[1][13] ,
         \SHIFT[1][12] , \SHIFT[1][11] , \SHIFT[1][10] , \SHIFT[1][9] ,
         \SHIFT[1][8] , \SHIFT[1][7] , \SHIFT[1][6] , \SHIFT[1][5] ,
         \SHIFT[1][4] , \SHIFT[1][3] , \SHIFT[1][2] , \SHIFT[1][1] ,
         \SHIFT[15][61] , \SHIFT[15][60] , \SHIFT[15][59] , \SHIFT[15][58] ,
         \SHIFT[15][57] , \SHIFT[15][56] , \SHIFT[15][55] , \SHIFT[15][54] ,
         \SHIFT[15][53] , \SHIFT[15][52] , \SHIFT[15][51] , \SHIFT[15][50] ,
         \SHIFT[15][49] , \SHIFT[15][48] , \SHIFT[15][47] , \SHIFT[15][46] ,
         \SHIFT[15][45] , \SHIFT[15][44] , \SHIFT[15][43] , \SHIFT[15][42] ,
         \SHIFT[15][41] , \SHIFT[15][40] , \SHIFT[15][39] , \SHIFT[15][38] ,
         \SHIFT[15][37] , \SHIFT[15][36] , \SHIFT[15][35] , \SHIFT[15][34] ,
         \SHIFT[15][33] , \SHIFT[15][32] , \SHIFT[15][31] , \SHIFT[15][30] ,
         \SHIFT[15][29] , \SHIFT[15][28] , \SHIFT[15][27] , \SHIFT[15][26] ,
         \SHIFT[15][25] , \SHIFT[15][24] , \SHIFT[15][23] , \SHIFT[15][22] ,
         \SHIFT[15][21] , \SHIFT[15][20] , \SHIFT[15][19] , \SHIFT[15][18] ,
         \SHIFT[15][17] , \SHIFT[15][16] , \SHIFT[15][15] , \SHIFT[15][14] ,
         \SHIFT[15][13] , \SHIFT[15][12] , \SHIFT[15][11] , \SHIFT[15][10] ,
         \SHIFT[15][9] , \SHIFT[15][8] , \SHIFT[15][7] , \SHIFT[15][6] ,
         \SHIFT[15][5] , \SHIFT[15][4] , \SHIFT[15][3] , \SHIFT[15][2] ,
         \SHIFT[14][59] , \SHIFT[14][58] , \SHIFT[14][57] , \SHIFT[14][56] ,
         \SHIFT[14][55] , \SHIFT[14][54] , \SHIFT[14][53] , \SHIFT[14][52] ,
         \SHIFT[14][51] , \SHIFT[14][50] , \SHIFT[14][49] , \SHIFT[14][48] ,
         \SHIFT[14][47] , \SHIFT[14][46] , \SHIFT[14][45] , \SHIFT[14][44] ,
         \SHIFT[14][43] , \SHIFT[14][42] , \SHIFT[14][41] , \SHIFT[14][40] ,
         \SHIFT[14][39] , \SHIFT[14][38] , \SHIFT[14][37] , \SHIFT[14][36] ,
         \SHIFT[14][35] , \SHIFT[14][34] , \SHIFT[14][33] , \SHIFT[14][32] ,
         \SHIFT[14][31] , \SHIFT[14][30] , \SHIFT[14][29] , \SHIFT[14][28] ,
         \SHIFT[14][27] , \SHIFT[14][26] , \SHIFT[14][25] , \SHIFT[14][24] ,
         \SHIFT[14][23] , \SHIFT[14][22] , \SHIFT[14][21] , \SHIFT[14][20] ,
         \SHIFT[14][19] , \SHIFT[14][18] , \SHIFT[14][17] , \SHIFT[14][16] ,
         \SHIFT[14][15] , \SHIFT[14][14] , \SHIFT[14][13] , \SHIFT[14][12] ,
         \SHIFT[14][11] , \SHIFT[14][10] , \SHIFT[14][9] , \SHIFT[14][8] ,
         \SHIFT[14][7] , \SHIFT[14][6] , \SHIFT[14][5] , \SHIFT[14][4] ,
         \SHIFT[14][3] , \SHIFT[14][2] , \SHIFT[13][57] , \SHIFT[13][56] ,
         \SHIFT[13][55] , \SHIFT[13][54] , \SHIFT[13][53] , \SHIFT[13][52] ,
         \SHIFT[13][51] , \SHIFT[13][50] , \SHIFT[13][49] , \SHIFT[13][48] ,
         \SHIFT[13][47] , \SHIFT[13][46] , \SHIFT[13][45] , \SHIFT[13][44] ,
         \SHIFT[13][43] , \SHIFT[13][42] , \SHIFT[13][41] , \SHIFT[13][40] ,
         \SHIFT[13][39] , \SHIFT[13][38] , \SHIFT[13][37] , \SHIFT[13][36] ,
         \SHIFT[13][35] , \SHIFT[13][34] , \SHIFT[13][33] , \SHIFT[13][32] ,
         \SHIFT[13][31] , \SHIFT[13][30] , \SHIFT[13][29] , \SHIFT[13][28] ,
         \SHIFT[13][27] , \SHIFT[13][26] , \SHIFT[13][25] , \SHIFT[13][24] ,
         \SHIFT[13][23] , \SHIFT[13][22] , \SHIFT[13][21] , \SHIFT[13][20] ,
         \SHIFT[13][19] , \SHIFT[13][18] , \SHIFT[13][17] , \SHIFT[13][16] ,
         \SHIFT[13][15] , \SHIFT[13][14] , \SHIFT[13][13] , \SHIFT[13][12] ,
         \SHIFT[13][11] , \SHIFT[13][10] , \SHIFT[13][9] , \SHIFT[13][8] ,
         \SHIFT[13][7] , \SHIFT[13][6] , \SHIFT[13][5] , \SHIFT[13][4] ,
         \SHIFT[13][3] , \SHIFT[13][2] , \SHIFT[12][55] , \SHIFT[12][54] ,
         \SHIFT[12][53] , \SHIFT[12][52] , \SHIFT[12][51] , \SHIFT[12][50] ,
         \SHIFT[12][49] , \SHIFT[12][48] , \SHIFT[12][47] , \SHIFT[12][46] ,
         \SHIFT[12][45] , \SHIFT[12][44] , \SHIFT[12][43] , \SHIFT[12][42] ,
         \SHIFT[12][41] , \SHIFT[12][40] , \SHIFT[12][39] , \SHIFT[12][38] ,
         \SHIFT[12][37] , \SHIFT[12][36] , \SHIFT[12][35] , \SHIFT[12][34] ,
         \SHIFT[12][33] , \SHIFT[12][32] , \SHIFT[12][31] , \SHIFT[12][30] ,
         \SHIFT[12][29] , \SHIFT[12][28] , \SHIFT[12][27] , \SHIFT[12][26] ,
         \SHIFT[12][25] , \SHIFT[12][24] , \SHIFT[12][23] , \SHIFT[12][22] ,
         \SHIFT[12][21] , \SHIFT[12][20] , \SHIFT[12][19] , \SHIFT[12][18] ,
         \SHIFT[12][17] , \SHIFT[12][16] , \SHIFT[12][15] , \SHIFT[12][14] ,
         \SHIFT[12][13] , \SHIFT[12][12] , \SHIFT[12][11] , \SHIFT[12][10] ,
         \SHIFT[12][9] , \SHIFT[12][8] , \SHIFT[12][7] , \SHIFT[12][6] ,
         \SHIFT[12][5] , \SHIFT[12][4] , \SHIFT[12][3] , \SHIFT[12][2] ,
         \SHIFT[11][53] , \SHIFT[11][52] , \SHIFT[11][51] , \SHIFT[11][50] ,
         \SHIFT[11][49] , \SHIFT[11][48] , \SHIFT[11][47] , \SHIFT[11][46] ,
         \SHIFT[11][45] , \SHIFT[11][44] , \SHIFT[11][43] , \SHIFT[11][42] ,
         \SHIFT[11][41] , \SHIFT[11][40] , \SHIFT[11][39] , \SHIFT[11][38] ,
         \SHIFT[11][37] , \SHIFT[11][36] , \SHIFT[11][35] , \SHIFT[11][34] ,
         \SHIFT[11][33] , \SHIFT[11][32] , \SHIFT[11][31] , \SHIFT[11][30] ,
         \SHIFT[11][29] , \SHIFT[11][28] , \SHIFT[11][27] , \SHIFT[11][26] ,
         \SHIFT[11][25] , \SHIFT[11][24] , \SHIFT[11][23] , \SHIFT[11][22] ,
         \SHIFT[11][21] , \SHIFT[11][20] , \SHIFT[11][19] , \SHIFT[11][18] ,
         \SHIFT[11][17] , \SHIFT[11][16] , \SHIFT[11][15] , \SHIFT[11][14] ,
         \SHIFT[11][13] , \SHIFT[11][12] , \SHIFT[11][11] , \SHIFT[11][10] ,
         \SHIFT[11][9] , \SHIFT[11][8] , \SHIFT[11][7] , \SHIFT[11][6] ,
         \SHIFT[11][5] , \SHIFT[11][4] , \SHIFT[11][3] , \SHIFT[11][2] ,
         \SHIFT[10][51] , \SHIFT[10][50] , \SHIFT[10][49] , \SHIFT[10][48] ,
         \SHIFT[10][47] , \SHIFT[10][46] , \SHIFT[10][45] , \SHIFT[10][44] ,
         \SHIFT[10][43] , \SHIFT[10][42] , \SHIFT[10][41] , \SHIFT[10][40] ,
         \SHIFT[10][39] , \SHIFT[10][38] , \SHIFT[10][37] , \SHIFT[10][36] ,
         \SHIFT[10][35] , \SHIFT[10][34] , \SHIFT[10][33] , \SHIFT[10][32] ,
         \SHIFT[10][31] , \SHIFT[10][30] , \SHIFT[10][29] , \SHIFT[10][28] ,
         \SHIFT[10][27] , \SHIFT[10][26] , \SHIFT[10][25] , \SHIFT[10][24] ,
         \SHIFT[10][23] , \SHIFT[10][22] , \SHIFT[10][21] , \SHIFT[10][20] ,
         \SHIFT[10][19] , \SHIFT[10][18] , \SHIFT[10][17] , \SHIFT[10][16] ,
         \SHIFT[10][15] , \SHIFT[10][14] , \SHIFT[10][13] , \SHIFT[10][12] ,
         \SHIFT[10][11] , \SHIFT[10][10] , \SHIFT[10][9] , \SHIFT[10][8] ,
         \SHIFT[10][7] , \SHIFT[10][6] , \SHIFT[10][5] , \SHIFT[10][4] ,
         \SHIFT[10][3] , \SHIFT[10][2] , \SHIFT[9][49] , \SHIFT[9][48] ,
         \SHIFT[9][47] , \SHIFT[9][46] , \SHIFT[9][45] , \SHIFT[9][44] ,
         \SHIFT[9][43] , \SHIFT[9][42] , \SHIFT[9][41] , \SHIFT[9][40] ,
         \SHIFT[9][39] , \SHIFT[9][38] , \SHIFT[9][37] , \SHIFT[9][36] ,
         \SHIFT[9][35] , \SHIFT[9][34] , \SHIFT[9][33] , \SHIFT[9][32] ,
         \SHIFT[9][31] , \SHIFT[9][30] , \SHIFT[9][29] , \SHIFT[9][28] ,
         \SHIFT[9][27] , \SHIFT[9][26] , \SHIFT[9][25] , \SHIFT[9][24] ,
         \SHIFT[9][23] , \SHIFT[9][22] , \SHIFT[9][21] , \SHIFT[9][20] ,
         \SHIFT[9][19] , \SHIFT[9][18] , \SHIFT[9][17] , \SHIFT[9][16] ,
         \SHIFT[9][15] , \SHIFT[9][14] , \SHIFT[9][13] , \SHIFT[9][12] ,
         \SHIFT[9][11] , \SHIFT[9][10] , \SHIFT[9][9] , \SHIFT[9][8] ,
         \SHIFT[9][7] , \SHIFT[9][6] , \SHIFT[9][5] , \SHIFT[9][4] ,
         \SHIFT[9][3] , \SHIFT[9][2] , \SHIFT[8][47] , \SHIFT[8][46] ,
         \SHIFT[8][45] , \SHIFT[8][44] , \SHIFT[8][43] , \SHIFT[8][42] ,
         \SHIFT[8][41] , \SHIFT[8][40] , \SHIFT[8][39] , \SHIFT[8][38] ,
         \SHIFT[8][37] , \SHIFT[8][36] , \SHIFT[8][35] , \SHIFT[8][34] ,
         \SHIFT[8][33] , \SHIFT[8][32] , \SHIFT[8][31] , \SHIFT[8][30] ,
         \SHIFT[8][29] , \SHIFT[8][28] , \SHIFT[8][27] , \SHIFT[8][26] ,
         \SHIFT[8][25] , \SHIFT[8][24] , \SHIFT[8][23] , \SHIFT[8][22] ,
         \SHIFT[8][21] , \SHIFT[8][20] , \SHIFT[8][19] , \SHIFT[8][18] ,
         \SHIFT[8][17] , \SHIFT[8][16] , \SHIFT[8][15] , \SHIFT[8][14] ,
         \SHIFT[8][13] , \SHIFT[8][12] , \SHIFT[8][11] , \SHIFT[8][10] ,
         \SHIFT[8][9] , \SHIFT[8][8] , \SHIFT[8][7] , \SHIFT[8][6] ,
         \SHIFT[8][5] , \SHIFT[8][4] , \SHIFT[8][3] , \SHIFT[8][2] ,
         \SHIFT[7][45] , \SHIFT[7][44] , \SHIFT[7][43] , \SHIFT[7][42] ,
         \SHIFT[7][41] , \SHIFT[7][40] , \SHIFT[7][39] , \SHIFT[7][38] ,
         \SHIFT[7][37] , \SHIFT[7][36] , \SHIFT[7][35] , \SHIFT[7][34] ,
         \SHIFT[7][33] , \SHIFT[7][32] , \SHIFT[7][31] , \SHIFT[7][30] ,
         \SHIFT[7][29] , \SHIFT[7][28] , \SHIFT[7][27] , \SHIFT[7][26] ,
         \SHIFT[7][25] , \SHIFT[7][24] , \SHIFT[7][23] , \SHIFT[7][22] ,
         \SHIFT[7][21] , \SHIFT[7][20] , \SHIFT[7][19] , \SHIFT[7][18] ,
         \SHIFT[7][17] , \SHIFT[7][16] , \SHIFT[7][15] , \SHIFT[7][14] ,
         \SHIFT[7][13] , \SHIFT[7][12] , \SHIFT[7][11] , \SHIFT[7][10] ,
         \SHIFT[7][9] , \SHIFT[7][8] , \SHIFT[7][7] , \SHIFT[7][6] ,
         \SHIFT[7][5] , \SHIFT[7][4] , \SHIFT[7][3] , \SHIFT[7][2] ,
         \SHIFT[6][43] , \SHIFT[6][42] , \SHIFT[6][41] , \SHIFT[6][40] ,
         \SHIFT[6][39] , \SHIFT[6][38] , \SHIFT[6][37] , \SHIFT[6][36] ,
         \SHIFT[6][35] , \SHIFT[6][34] , \SHIFT[6][33] , \SHIFT[6][32] ,
         \SHIFT[6][31] , \SHIFT[6][30] , \SHIFT[6][29] , \SHIFT[6][28] ,
         \SHIFT[6][27] , \SHIFT[6][26] , \SHIFT[6][25] , \SHIFT[6][24] ,
         \SHIFT[6][23] , \SHIFT[6][22] , \SHIFT[6][21] , \SHIFT[6][20] ,
         \SHIFT[6][19] , \SHIFT[6][18] , \SHIFT[6][17] , \SHIFT[6][16] ,
         \SHIFT[6][15] , \SHIFT[6][14] , \SHIFT[6][13] , \SHIFT[6][12] ,
         \SHIFT[6][11] , \SHIFT[6][10] , \SHIFT[6][9] , \SHIFT[6][8] ,
         \SHIFT[6][7] , \SHIFT[6][6] , \SHIFT[6][5] , \SHIFT[6][4] ,
         \SHIFT[6][3] , \SHIFT[6][2] , \SHIFT[5][41] , \SHIFT[5][40] ,
         \SHIFT[5][39] , \SHIFT[5][38] , \SHIFT[5][37] , \SHIFT[5][36] ,
         \SHIFT[5][35] , \SHIFT[5][34] , \SHIFT[5][33] , \SHIFT[5][32] ,
         \SHIFT[5][31] , \SHIFT[5][30] , \SHIFT[5][29] , \SHIFT[5][28] ,
         \SHIFT[5][27] , \SHIFT[5][26] , \SHIFT[5][25] , \SHIFT[5][24] ,
         \SHIFT[5][23] , \SHIFT[5][22] , \SHIFT[5][21] , \SHIFT[5][20] ,
         \SHIFT[5][19] , \SHIFT[5][18] , \SHIFT[5][17] , \SHIFT[5][16] ,
         \SHIFT[5][15] , \SHIFT[5][14] , \SHIFT[5][13] , \SHIFT[5][12] ,
         \SHIFT[5][11] , \SHIFT[5][10] , \SHIFT[5][9] , \SHIFT[5][8] ,
         \SHIFT[5][7] , \SHIFT[5][6] , \SHIFT[5][5] , \SHIFT[5][4] ,
         \SHIFT[5][3] , \SHIFT[5][2] , \SHIFT[4][39] , \SHIFT[4][38] ,
         \SHIFT[4][37] , \SHIFT[4][36] , \SHIFT[4][35] , \SHIFT[4][34] ,
         \SHIFT[4][33] , \SHIFT[4][32] , \SHIFT[4][31] , \SHIFT[4][30] ,
         \SHIFT[4][29] , \SHIFT[4][28] , \SHIFT[4][27] , \SHIFT[4][26] ,
         \SHIFT[4][25] , \SHIFT[4][24] , \SHIFT[4][23] , \SHIFT[4][22] ,
         \SHIFT[4][21] , \SHIFT[4][20] , \SHIFT[4][19] , \SHIFT[4][18] ,
         \SHIFT[4][17] , \SHIFT[4][16] , \SHIFT[4][15] , \SHIFT[4][14] ,
         \SHIFT[4][13] , \SHIFT[4][12] , \SHIFT[4][11] , \SHIFT[4][10] ,
         \SHIFT[4][9] , \SHIFT[4][8] , \SHIFT[4][7] , \SHIFT[4][6] ,
         \SHIFT[4][5] , \SHIFT[4][4] , \SHIFT[4][3] , \SHIFT[4][2] ,
         \SHIFT[3][37] , \SHIFT[3][36] , \SHIFT[3][35] , \SHIFT[3][34] ,
         \SHIFT[3][33] , \SHIFT[3][32] , \SHIFT[3][31] , \SHIFT[3][30] ,
         \SHIFT[3][29] , \SHIFT[3][28] , \SHIFT[3][27] , \SHIFT[3][26] ,
         \SHIFT[3][25] , \SHIFT[3][24] , \SHIFT[3][23] , \SHIFT[3][22] ,
         \SHIFT[3][21] , \SHIFT[3][20] , \SHIFT[3][19] , \SHIFT[3][18] ,
         \SHIFT[3][17] , \SHIFT[3][16] , \SHIFT[3][15] , \SHIFT[3][14] ,
         \SHIFT[3][13] , \SHIFT[3][12] , \SHIFT[3][11] , \SHIFT[3][10] ,
         \SHIFT[3][9] , \SHIFT[3][8] , \SHIFT[3][7] , \SHIFT[3][6] ,
         \SHIFT[3][5] , \SHIFT[3][4] , \SHIFT[3][3] , \SHIFT[3][2] ,
         \SHIFT[2][35] , \SHIFT[2][34] , \SHIFT[2][33] , \SHIFT[2][32] ,
         \SHIFT[2][31] , \SHIFT[2][30] , \SHIFT[2][29] , \SHIFT[2][28] ,
         \SHIFT[2][27] , \SHIFT[2][26] , \SHIFT[2][25] , \SHIFT[2][24] ,
         \SHIFT[2][23] , \SHIFT[2][22] , \SHIFT[2][21] , \SHIFT[2][20] ,
         \SHIFT[2][19] , \SHIFT[2][18] , \SHIFT[2][17] , \SHIFT[2][16] ,
         \SHIFT[2][15] , \SHIFT[2][14] , \SHIFT[2][13] , \SHIFT[2][12] ,
         \SHIFT[2][11] , \SHIFT[2][10] , \SHIFT[2][9] , \SHIFT[2][8] ,
         \SHIFT[2][7] , \SHIFT[2][6] , \SHIFT[2][5] , \SHIFT[2][4] ,
         \SHIFT[2][3] , \SHIFT[2][2] , \SHIFT[1][33] , \SHIFT[1][32] ,
         \SHIFT_n[1][31] , \SHIFT_n[1][30] , \SHIFT_n[1][29] ,
         \SHIFT_n[1][28] , \SHIFT_n[1][27] , \SHIFT_n[1][26] ,
         \SHIFT_n[1][25] , \SHIFT_n[1][24] , \SHIFT_n[1][23] ,
         \SHIFT_n[1][22] , \SHIFT_n[1][21] , \SHIFT_n[1][20] ,
         \SHIFT_n[1][19] , \SHIFT_n[1][18] , \SHIFT_n[1][17] ,
         \SHIFT_n[1][16] , \SHIFT_n[1][15] , \SHIFT_n[1][14] ,
         \SHIFT_n[1][13] , \SHIFT_n[1][12] , \SHIFT_n[1][11] ,
         \SHIFT_n[1][10] , \SHIFT_n[1][9] , \SHIFT_n[1][8] , \SHIFT_n[1][7] ,
         \SHIFT_n[1][6] , \SHIFT_n[1][5] , \SHIFT_n[1][4] , \SHIFT_n[1][3] ,
         \SHIFT_n[1][2] , \SHIFT_n[1][1] , \SHIFT_n[15][61] ,
         \SHIFT_n[15][60] , \SHIFT_n[15][59] , \SHIFT_n[15][58] ,
         \SHIFT_n[15][57] , \SHIFT_n[15][56] , \SHIFT_n[15][55] ,
         \SHIFT_n[15][54] , \SHIFT_n[15][53] , \SHIFT_n[15][52] ,
         \SHIFT_n[15][51] , \SHIFT_n[15][50] , \SHIFT_n[15][49] ,
         \SHIFT_n[15][48] , \SHIFT_n[15][47] , \SHIFT_n[15][46] ,
         \SHIFT_n[15][45] , \SHIFT_n[15][44] , \SHIFT_n[15][43] ,
         \SHIFT_n[15][42] , \SHIFT_n[15][41] , \SHIFT_n[15][40] ,
         \SHIFT_n[15][39] , \SHIFT_n[15][38] , \SHIFT_n[15][37] ,
         \SHIFT_n[15][36] , \SHIFT_n[15][35] , \SHIFT_n[15][34] ,
         \SHIFT_n[15][33] , \SHIFT_n[15][32] , \SHIFT_n[15][31] ,
         \SHIFT_n[15][30] , \SHIFT_n[15][29] , \SHIFT_n[15][28] ,
         \SHIFT_n[15][27] , \SHIFT_n[15][26] , \SHIFT_n[15][25] ,
         \SHIFT_n[15][24] , \SHIFT_n[15][23] , \SHIFT_n[15][22] ,
         \SHIFT_n[15][21] , \SHIFT_n[15][20] , \SHIFT_n[15][19] ,
         \SHIFT_n[15][18] , \SHIFT_n[15][17] , \SHIFT_n[15][16] ,
         \SHIFT_n[15][15] , \SHIFT_n[15][14] , \SHIFT_n[15][13] ,
         \SHIFT_n[15][12] , \SHIFT_n[15][11] , \SHIFT_n[15][10] ,
         \SHIFT_n[15][9] , \SHIFT_n[15][8] , \SHIFT_n[15][7] ,
         \SHIFT_n[15][6] , \SHIFT_n[15][5] , \SHIFT_n[15][4] ,
         \SHIFT_n[15][3] , \SHIFT_n[15][2] , \SHIFT_n[14][59] ,
         \SHIFT_n[14][58] , \SHIFT_n[14][57] , \SHIFT_n[14][56] ,
         \SHIFT_n[14][55] , \SHIFT_n[14][54] , \SHIFT_n[14][53] ,
         \SHIFT_n[14][52] , \SHIFT_n[14][51] , \SHIFT_n[14][50] ,
         \SHIFT_n[14][49] , \SHIFT_n[14][48] , \SHIFT_n[14][47] ,
         \SHIFT_n[14][46] , \SHIFT_n[14][45] , \SHIFT_n[14][44] ,
         \SHIFT_n[14][43] , \SHIFT_n[14][42] , \SHIFT_n[14][41] ,
         \SHIFT_n[14][40] , \SHIFT_n[14][39] , \SHIFT_n[14][38] ,
         \SHIFT_n[14][37] , \SHIFT_n[14][36] , \SHIFT_n[14][35] ,
         \SHIFT_n[14][34] , \SHIFT_n[14][33] , \SHIFT_n[14][32] ,
         \SHIFT_n[14][31] , \SHIFT_n[14][30] , \SHIFT_n[14][29] ,
         \SHIFT_n[14][28] , \SHIFT_n[14][27] , \SHIFT_n[14][26] ,
         \SHIFT_n[14][25] , \SHIFT_n[14][24] , \SHIFT_n[14][23] ,
         \SHIFT_n[14][22] , \SHIFT_n[14][21] , \SHIFT_n[14][20] ,
         \SHIFT_n[14][19] , \SHIFT_n[14][18] , \SHIFT_n[14][17] ,
         \SHIFT_n[14][16] , \SHIFT_n[14][15] , \SHIFT_n[14][14] ,
         \SHIFT_n[14][13] , \SHIFT_n[14][12] , \SHIFT_n[14][11] ,
         \SHIFT_n[14][10] , \SHIFT_n[14][9] , \SHIFT_n[14][8] ,
         \SHIFT_n[14][7] , \SHIFT_n[14][6] , \SHIFT_n[14][5] ,
         \SHIFT_n[14][4] , \SHIFT_n[14][3] , \SHIFT_n[14][2] ,
         \SHIFT_n[13][57] , \SHIFT_n[13][56] , \SHIFT_n[13][55] ,
         \SHIFT_n[13][54] , \SHIFT_n[13][53] , \SHIFT_n[13][52] ,
         \SHIFT_n[13][51] , \SHIFT_n[13][50] , \SHIFT_n[13][49] ,
         \SHIFT_n[13][48] , \SHIFT_n[13][47] , \SHIFT_n[13][46] ,
         \SHIFT_n[13][45] , \SHIFT_n[13][44] , \SHIFT_n[13][43] ,
         \SHIFT_n[13][42] , \SHIFT_n[13][41] , \SHIFT_n[13][40] ,
         \SHIFT_n[13][39] , \SHIFT_n[13][38] , \SHIFT_n[13][37] ,
         \SHIFT_n[13][36] , \SHIFT_n[13][35] , \SHIFT_n[13][34] ,
         \SHIFT_n[13][33] , \SHIFT_n[13][32] , \SHIFT_n[13][31] ,
         \SHIFT_n[13][30] , \SHIFT_n[13][29] , \SHIFT_n[13][28] ,
         \SHIFT_n[13][27] , \SHIFT_n[13][26] , \SHIFT_n[13][25] ,
         \SHIFT_n[13][24] , \SHIFT_n[13][23] , \SHIFT_n[13][22] ,
         \SHIFT_n[13][21] , \SHIFT_n[13][20] , \SHIFT_n[13][19] ,
         \SHIFT_n[13][18] , \SHIFT_n[13][17] , \SHIFT_n[13][16] ,
         \SHIFT_n[13][15] , \SHIFT_n[13][14] , \SHIFT_n[13][13] ,
         \SHIFT_n[13][12] , \SHIFT_n[13][11] , \SHIFT_n[13][10] ,
         \SHIFT_n[13][9] , \SHIFT_n[13][8] , \SHIFT_n[13][7] ,
         \SHIFT_n[13][6] , \SHIFT_n[13][5] , \SHIFT_n[13][4] ,
         \SHIFT_n[13][3] , \SHIFT_n[13][2] , \SHIFT_n[12][55] ,
         \SHIFT_n[12][54] , \SHIFT_n[12][53] , \SHIFT_n[12][52] ,
         \SHIFT_n[12][51] , \SHIFT_n[12][50] , \SHIFT_n[12][49] ,
         \SHIFT_n[12][48] , \SHIFT_n[12][47] , \SHIFT_n[12][46] ,
         \SHIFT_n[12][45] , \SHIFT_n[12][44] , \SHIFT_n[12][43] ,
         \SHIFT_n[12][42] , \SHIFT_n[12][41] , \SHIFT_n[12][40] ,
         \SHIFT_n[12][39] , \SHIFT_n[12][38] , \SHIFT_n[12][37] ,
         \SHIFT_n[12][36] , \SHIFT_n[12][35] , \SHIFT_n[12][34] ,
         \SHIFT_n[12][33] , \SHIFT_n[12][32] , \SHIFT_n[12][31] ,
         \SHIFT_n[12][30] , \SHIFT_n[12][29] , \SHIFT_n[12][28] ,
         \SHIFT_n[12][27] , \SHIFT_n[12][26] , \SHIFT_n[12][25] ,
         \SHIFT_n[12][24] , \SHIFT_n[12][23] , \SHIFT_n[12][22] ,
         \SHIFT_n[12][21] , \SHIFT_n[12][20] , \SHIFT_n[12][19] ,
         \SHIFT_n[12][18] , \SHIFT_n[12][17] , \SHIFT_n[12][16] ,
         \SHIFT_n[12][15] , \SHIFT_n[12][14] , \SHIFT_n[12][13] ,
         \SHIFT_n[12][12] , \SHIFT_n[12][11] , \SHIFT_n[12][10] ,
         \SHIFT_n[12][9] , \SHIFT_n[12][8] , \SHIFT_n[12][7] ,
         \SHIFT_n[12][6] , \SHIFT_n[12][5] , \SHIFT_n[12][4] ,
         \SHIFT_n[12][3] , \SHIFT_n[12][2] , \SHIFT_n[11][53] ,
         \SHIFT_n[11][52] , \SHIFT_n[11][51] , \SHIFT_n[11][50] ,
         \SHIFT_n[11][49] , \SHIFT_n[11][48] , \SHIFT_n[11][47] ,
         \SHIFT_n[11][46] , \SHIFT_n[11][45] , \SHIFT_n[11][44] ,
         \SHIFT_n[11][43] , \SHIFT_n[11][42] , \SHIFT_n[11][41] ,
         \SHIFT_n[11][40] , \SHIFT_n[11][39] , \SHIFT_n[11][38] ,
         \SHIFT_n[11][37] , \SHIFT_n[11][36] , \SHIFT_n[11][35] ,
         \SHIFT_n[11][34] , \SHIFT_n[11][33] , \SHIFT_n[11][32] ,
         \SHIFT_n[11][31] , \SHIFT_n[11][30] , \SHIFT_n[11][29] ,
         \SHIFT_n[11][28] , \SHIFT_n[11][27] , \SHIFT_n[11][26] ,
         \SHIFT_n[11][25] , \SHIFT_n[11][24] , \SHIFT_n[11][23] ,
         \SHIFT_n[11][22] , \SHIFT_n[11][21] , \SHIFT_n[11][20] ,
         \SHIFT_n[11][19] , \SHIFT_n[11][18] , \SHIFT_n[11][17] ,
         \SHIFT_n[11][16] , \SHIFT_n[11][15] , \SHIFT_n[11][14] ,
         \SHIFT_n[11][13] , \SHIFT_n[11][12] , \SHIFT_n[11][11] ,
         \SHIFT_n[11][10] , \SHIFT_n[11][9] , \SHIFT_n[11][8] ,
         \SHIFT_n[11][7] , \SHIFT_n[11][6] , \SHIFT_n[11][5] ,
         \SHIFT_n[11][4] , \SHIFT_n[11][3] , \SHIFT_n[11][2] ,
         \SHIFT_n[10][51] , \SHIFT_n[10][50] , \SHIFT_n[10][49] ,
         \SHIFT_n[10][48] , \SHIFT_n[10][47] , \SHIFT_n[10][46] ,
         \SHIFT_n[10][45] , \SHIFT_n[10][44] , \SHIFT_n[10][43] ,
         \SHIFT_n[10][42] , \SHIFT_n[10][41] , \SHIFT_n[10][40] ,
         \SHIFT_n[10][39] , \SHIFT_n[10][38] , \SHIFT_n[10][37] ,
         \SHIFT_n[10][36] , \SHIFT_n[10][35] , \SHIFT_n[10][34] ,
         \SHIFT_n[10][33] , \SHIFT_n[10][32] , \SHIFT_n[10][31] ,
         \SHIFT_n[10][30] , \SHIFT_n[10][29] , \SHIFT_n[10][28] ,
         \SHIFT_n[10][27] , \SHIFT_n[10][26] , \SHIFT_n[10][25] ,
         \SHIFT_n[10][24] , \SHIFT_n[10][23] , \SHIFT_n[10][22] ,
         \SHIFT_n[10][21] , \SHIFT_n[10][20] , \SHIFT_n[10][19] ,
         \SHIFT_n[10][18] , \SHIFT_n[10][17] , \SHIFT_n[10][16] ,
         \SHIFT_n[10][15] , \SHIFT_n[10][14] , \SHIFT_n[10][13] ,
         \SHIFT_n[10][12] , \SHIFT_n[10][11] , \SHIFT_n[10][10] ,
         \SHIFT_n[10][9] , \SHIFT_n[10][8] , \SHIFT_n[10][7] ,
         \SHIFT_n[10][6] , \SHIFT_n[10][5] , \SHIFT_n[10][4] ,
         \SHIFT_n[10][3] , \SHIFT_n[10][2] , \SHIFT_n[9][49] ,
         \SHIFT_n[9][48] , \SHIFT_n[9][47] , \SHIFT_n[9][46] ,
         \SHIFT_n[9][45] , \SHIFT_n[9][44] , \SHIFT_n[9][43] ,
         \SHIFT_n[9][42] , \SHIFT_n[9][41] , \SHIFT_n[9][40] ,
         \SHIFT_n[9][39] , \SHIFT_n[9][38] , \SHIFT_n[9][37] ,
         \SHIFT_n[9][36] , \SHIFT_n[9][35] , \SHIFT_n[9][34] ,
         \SHIFT_n[9][33] , \SHIFT_n[9][32] , \SHIFT_n[9][31] ,
         \SHIFT_n[9][30] , \SHIFT_n[9][29] , \SHIFT_n[9][28] ,
         \SHIFT_n[9][27] , \SHIFT_n[9][26] , \SHIFT_n[9][25] ,
         \SHIFT_n[9][24] , \SHIFT_n[9][23] , \SHIFT_n[9][22] ,
         \SHIFT_n[9][21] , \SHIFT_n[9][20] , \SHIFT_n[9][19] ,
         \SHIFT_n[9][18] , \SHIFT_n[9][17] , \SHIFT_n[9][16] ,
         \SHIFT_n[9][15] , \SHIFT_n[9][14] , \SHIFT_n[9][13] ,
         \SHIFT_n[9][12] , \SHIFT_n[9][11] , \SHIFT_n[9][10] , \SHIFT_n[9][9] ,
         \SHIFT_n[9][8] , \SHIFT_n[9][7] , \SHIFT_n[9][6] , \SHIFT_n[9][5] ,
         \SHIFT_n[9][4] , \SHIFT_n[9][3] , \SHIFT_n[9][2] , \SHIFT_n[8][47] ,
         \SHIFT_n[8][46] , \SHIFT_n[8][45] , \SHIFT_n[8][44] ,
         \SHIFT_n[8][43] , \SHIFT_n[8][42] , \SHIFT_n[8][41] ,
         \SHIFT_n[8][40] , \SHIFT_n[8][39] , \SHIFT_n[8][38] ,
         \SHIFT_n[8][37] , \SHIFT_n[8][36] , \SHIFT_n[8][35] ,
         \SHIFT_n[8][34] , \SHIFT_n[8][33] , \SHIFT_n[8][32] ,
         \SHIFT_n[8][31] , \SHIFT_n[8][30] , \SHIFT_n[8][29] ,
         \SHIFT_n[8][28] , \SHIFT_n[8][27] , \SHIFT_n[8][26] ,
         \SHIFT_n[8][25] , \SHIFT_n[8][24] , \SHIFT_n[8][23] ,
         \SHIFT_n[8][22] , \SHIFT_n[8][21] , \SHIFT_n[8][20] ,
         \SHIFT_n[8][19] , \SHIFT_n[8][18] , \SHIFT_n[8][17] ,
         \SHIFT_n[8][16] , \SHIFT_n[8][15] , \SHIFT_n[8][14] ,
         \SHIFT_n[8][13] , \SHIFT_n[8][12] , \SHIFT_n[8][11] ,
         \SHIFT_n[8][10] , \SHIFT_n[8][9] , \SHIFT_n[8][8] , \SHIFT_n[8][7] ,
         \SHIFT_n[8][6] , \SHIFT_n[8][5] , \SHIFT_n[8][4] , \SHIFT_n[8][3] ,
         \SHIFT_n[8][2] , \SHIFT_n[7][45] , \SHIFT_n[7][44] , \SHIFT_n[7][43] ,
         \SHIFT_n[7][42] , \SHIFT_n[7][41] , \SHIFT_n[7][40] ,
         \SHIFT_n[7][39] , \SHIFT_n[7][38] , \SHIFT_n[7][37] ,
         \SHIFT_n[7][36] , \SHIFT_n[7][35] , \SHIFT_n[7][34] ,
         \SHIFT_n[7][33] , \SHIFT_n[7][32] , \SHIFT_n[7][31] ,
         \SHIFT_n[7][30] , \SHIFT_n[7][29] , \SHIFT_n[7][28] ,
         \SHIFT_n[7][27] , \SHIFT_n[7][26] , \SHIFT_n[7][25] ,
         \SHIFT_n[7][24] , \SHIFT_n[7][23] , \SHIFT_n[7][22] ,
         \SHIFT_n[7][21] , \SHIFT_n[7][20] , \SHIFT_n[7][19] ,
         \SHIFT_n[7][18] , \SHIFT_n[7][17] , \SHIFT_n[7][16] ,
         \SHIFT_n[7][15] , \SHIFT_n[7][14] , \SHIFT_n[7][13] ,
         \SHIFT_n[7][12] , \SHIFT_n[7][11] , \SHIFT_n[7][10] , \SHIFT_n[7][9] ,
         \SHIFT_n[7][8] , \SHIFT_n[7][7] , \SHIFT_n[7][6] , \SHIFT_n[7][5] ,
         \SHIFT_n[7][4] , \SHIFT_n[7][3] , \SHIFT_n[7][2] , \SHIFT_n[6][43] ,
         \SHIFT_n[6][42] , \SHIFT_n[6][41] , \SHIFT_n[6][40] ,
         \SHIFT_n[6][39] , \SHIFT_n[6][38] , \SHIFT_n[6][37] ,
         \SHIFT_n[6][36] , \SHIFT_n[6][35] , \SHIFT_n[6][34] ,
         \SHIFT_n[6][33] , \SHIFT_n[6][32] , \SHIFT_n[6][31] ,
         \SHIFT_n[6][30] , \SHIFT_n[6][29] , \SHIFT_n[6][28] ,
         \SHIFT_n[6][27] , \SHIFT_n[6][26] , \SHIFT_n[6][25] ,
         \SHIFT_n[6][24] , \SHIFT_n[6][23] , \SHIFT_n[6][22] ,
         \SHIFT_n[6][21] , \SHIFT_n[6][20] , \SHIFT_n[6][19] ,
         \SHIFT_n[6][18] , \SHIFT_n[6][17] , \SHIFT_n[6][16] ,
         \SHIFT_n[6][15] , \SHIFT_n[6][14] , \SHIFT_n[6][13] ,
         \SHIFT_n[6][12] , \SHIFT_n[6][11] , \SHIFT_n[6][10] , \SHIFT_n[6][9] ,
         \SHIFT_n[6][8] , \SHIFT_n[6][7] , \SHIFT_n[6][6] , \SHIFT_n[6][5] ,
         \SHIFT_n[6][4] , \SHIFT_n[6][3] , \SHIFT_n[6][2] , \SHIFT_n[5][41] ,
         \SHIFT_n[5][40] , \SHIFT_n[5][39] , \SHIFT_n[5][38] ,
         \SHIFT_n[5][37] , \SHIFT_n[5][36] , \SHIFT_n[5][35] ,
         \SHIFT_n[5][34] , \SHIFT_n[5][33] , \SHIFT_n[5][32] ,
         \SHIFT_n[5][31] , \SHIFT_n[5][30] , \SHIFT_n[5][29] ,
         \SHIFT_n[5][28] , \SHIFT_n[5][27] , \SHIFT_n[5][26] ,
         \SHIFT_n[5][25] , \SHIFT_n[5][24] , \SHIFT_n[5][23] ,
         \SHIFT_n[5][22] , \SHIFT_n[5][21] , \SHIFT_n[5][20] ,
         \SHIFT_n[5][19] , \SHIFT_n[5][18] , \SHIFT_n[5][17] ,
         \SHIFT_n[5][16] , \SHIFT_n[5][15] , \SHIFT_n[5][14] ,
         \SHIFT_n[5][13] , \SHIFT_n[5][12] , \SHIFT_n[5][11] ,
         \SHIFT_n[5][10] , \SHIFT_n[5][9] , \SHIFT_n[5][8] , \SHIFT_n[5][7] ,
         \SHIFT_n[5][6] , \SHIFT_n[5][5] , \SHIFT_n[5][4] , \SHIFT_n[5][3] ,
         \SHIFT_n[5][2] , \SHIFT_n[4][39] , \SHIFT_n[4][38] , \SHIFT_n[4][37] ,
         \SHIFT_n[4][36] , \SHIFT_n[4][35] , \SHIFT_n[4][34] ,
         \SHIFT_n[4][33] , \SHIFT_n[4][32] , \SHIFT_n[4][31] ,
         \SHIFT_n[4][30] , \SHIFT_n[4][29] , \SHIFT_n[4][28] ,
         \SHIFT_n[4][27] , \SHIFT_n[4][26] , \SHIFT_n[4][25] ,
         \SHIFT_n[4][24] , \SHIFT_n[4][23] , \SHIFT_n[4][22] ,
         \SHIFT_n[4][21] , \SHIFT_n[4][20] , \SHIFT_n[4][19] ,
         \SHIFT_n[4][18] , \SHIFT_n[4][17] , \SHIFT_n[4][16] ,
         \SHIFT_n[4][15] , \SHIFT_n[4][14] , \SHIFT_n[4][13] ,
         \SHIFT_n[4][12] , \SHIFT_n[4][11] , \SHIFT_n[4][10] , \SHIFT_n[4][9] ,
         \SHIFT_n[4][8] , \SHIFT_n[4][7] , \SHIFT_n[4][6] , \SHIFT_n[4][5] ,
         \SHIFT_n[4][4] , \SHIFT_n[4][3] , \SHIFT_n[4][2] , \SHIFT_n[3][37] ,
         \SHIFT_n[3][36] , \SHIFT_n[3][35] , \SHIFT_n[3][34] ,
         \SHIFT_n[3][33] , \SHIFT_n[3][32] , \SHIFT_n[3][31] ,
         \SHIFT_n[3][30] , \SHIFT_n[3][29] , \SHIFT_n[3][28] ,
         \SHIFT_n[3][27] , \SHIFT_n[3][26] , \SHIFT_n[3][25] ,
         \SHIFT_n[3][24] , \SHIFT_n[3][23] , \SHIFT_n[3][22] ,
         \SHIFT_n[3][21] , \SHIFT_n[3][20] , \SHIFT_n[3][19] ,
         \SHIFT_n[3][18] , \SHIFT_n[3][17] , \SHIFT_n[3][16] ,
         \SHIFT_n[3][15] , \SHIFT_n[3][14] , \SHIFT_n[3][13] ,
         \SHIFT_n[3][12] , \SHIFT_n[3][11] , \SHIFT_n[3][10] , \SHIFT_n[3][9] ,
         \SHIFT_n[3][8] , \SHIFT_n[3][7] , \SHIFT_n[3][6] , \SHIFT_n[3][5] ,
         \SHIFT_n[3][4] , \SHIFT_n[3][3] , \SHIFT_n[3][2] , \SHIFT_n[2][35] ,
         \SHIFT_n[2][34] , \SHIFT_n[2][33] , \SHIFT_n[2][32] ,
         \SHIFT_n[2][31] , \SHIFT_n[2][30] , \SHIFT_n[2][29] ,
         \SHIFT_n[2][28] , \SHIFT_n[2][27] , \SHIFT_n[2][26] ,
         \SHIFT_n[2][25] , \SHIFT_n[2][24] , \SHIFT_n[2][23] ,
         \SHIFT_n[2][22] , \SHIFT_n[2][21] , \SHIFT_n[2][20] ,
         \SHIFT_n[2][19] , \SHIFT_n[2][18] , \SHIFT_n[2][17] ,
         \SHIFT_n[2][16] , \SHIFT_n[2][15] , \SHIFT_n[2][14] ,
         \SHIFT_n[2][13] , \SHIFT_n[2][12] , \SHIFT_n[2][11] ,
         \SHIFT_n[2][10] , \SHIFT_n[2][9] , \SHIFT_n[2][8] , \SHIFT_n[2][7] ,
         \SHIFT_n[2][6] , \SHIFT_n[2][5] , \SHIFT_n[2][4] , \SHIFT_n[2][3] ,
         \SHIFT_n[2][2] , \SHIFT_n[1][33] , \SHIFT_n[1][32] , \OTMP[8][15] ,
         \OTMP[8][14] , \OTMP[8][13] , \OTMP[8][12] , \OTMP[8][11] ,
         \OTMP[8][10] , \OTMP[8][9] , \OTMP[8][8] , \OTMP[8][7] , \OTMP[8][6] ,
         \OTMP[8][5] , \OTMP[8][4] , \OTMP[8][3] , \OTMP[8][2] , \OTMP[8][1] ,
         \OTMP[7][47] , \OTMP[7][46] , \OTMP[7][45] , \OTMP[7][44] ,
         \OTMP[7][43] , \OTMP[7][42] , \OTMP[7][41] , \OTMP[7][40] ,
         \OTMP[7][39] , \OTMP[7][38] , \OTMP[7][37] , \OTMP[7][36] ,
         \OTMP[7][35] , \OTMP[7][34] , \OTMP[7][33] , \OTMP[7][32] ,
         \OTMP[7][31] , \OTMP[7][30] , \OTMP[7][29] , \OTMP[7][28] ,
         \OTMP[7][27] , \OTMP[7][26] , \OTMP[7][25] , \OTMP[7][24] ,
         \OTMP[7][23] , \OTMP[7][22] , \OTMP[7][21] , \OTMP[7][20] ,
         \OTMP[7][19] , \OTMP[7][18] , \OTMP[7][17] , \OTMP[7][16] ,
         \OTMP[7][15] , \OTMP[7][14] , \OTMP[7][13] , \OTMP[7][12] ,
         \OTMP[7][11] , \OTMP[7][10] , \OTMP[7][9] , \OTMP[7][8] ,
         \OTMP[7][7] , \OTMP[7][6] , \OTMP[7][5] , \OTMP[7][4] , \OTMP[7][3] ,
         \OTMP[7][2] , \OTMP[7][1] , \OTMP[6][45] , \OTMP[6][44] ,
         \OTMP[6][43] , \OTMP[6][42] , \OTMP[6][41] , \OTMP[6][40] ,
         \OTMP[6][39] , \OTMP[6][38] , \OTMP[6][37] , \OTMP[6][36] ,
         \OTMP[6][35] , \OTMP[6][34] , \OTMP[6][33] , \OTMP[6][32] ,
         \OTMP[6][31] , \OTMP[6][30] , \OTMP[6][29] , \OTMP[6][28] ,
         \OTMP[6][27] , \OTMP[6][26] , \OTMP[6][25] , \OTMP[6][24] ,
         \OTMP[6][23] , \OTMP[6][22] , \OTMP[6][21] , \OTMP[6][20] ,
         \OTMP[6][19] , \OTMP[6][18] , \OTMP[6][17] , \OTMP[6][16] ,
         \OTMP[6][15] , \OTMP[6][14] , \OTMP[6][13] , \OTMP[6][12] ,
         \OTMP[6][11] , \OTMP[6][10] , \OTMP[6][9] , \OTMP[6][8] ,
         \OTMP[6][7] , \OTMP[6][6] , \OTMP[6][5] , \OTMP[6][4] , \OTMP[6][3] ,
         \OTMP[6][2] , \OTMP[6][1] , \OTMP[5][43] , \OTMP[5][42] ,
         \OTMP[5][41] , \OTMP[5][40] , \OTMP[5][39] , \OTMP[5][38] ,
         \OTMP[5][37] , \OTMP[5][36] , \OTMP[5][35] , \OTMP[5][34] ,
         \OTMP[5][33] , \OTMP[5][32] , \OTMP[5][31] , \OTMP[5][30] ,
         \OTMP[5][29] , \OTMP[5][28] , \OTMP[5][27] , \OTMP[5][26] ,
         \OTMP[5][25] , \OTMP[5][24] , \OTMP[5][23] , \OTMP[5][22] ,
         \OTMP[5][21] , \OTMP[5][20] , \OTMP[5][19] , \OTMP[5][18] ,
         \OTMP[5][17] , \OTMP[5][16] , \OTMP[5][15] , \OTMP[5][14] ,
         \OTMP[5][13] , \OTMP[5][12] , \OTMP[5][11] , \OTMP[5][10] ,
         \OTMP[5][9] , \OTMP[5][8] , \OTMP[5][7] , \OTMP[5][6] , \OTMP[5][5] ,
         \OTMP[5][4] , \OTMP[5][3] , \OTMP[5][2] , \OTMP[5][1] , \OTMP[4][41] ,
         \OTMP[4][40] , \OTMP[4][39] , \OTMP[4][38] , \OTMP[4][37] ,
         \OTMP[4][36] , \OTMP[4][35] , \OTMP[4][34] , \OTMP[4][33] ,
         \OTMP[4][32] , \OTMP[4][31] , \OTMP[4][30] , \OTMP[4][29] ,
         \OTMP[4][28] , \OTMP[4][27] , \OTMP[4][26] , \OTMP[4][25] ,
         \OTMP[4][24] , \OTMP[4][23] , \OTMP[4][22] , \OTMP[4][21] ,
         \OTMP[4][20] , \OTMP[4][19] , \OTMP[4][18] , \OTMP[4][17] ,
         \OTMP[4][16] , \OTMP[4][15] , \OTMP[4][14] , \OTMP[4][13] ,
         \OTMP[4][12] , \OTMP[4][11] , \OTMP[4][10] , \OTMP[4][9] ,
         \OTMP[4][8] , \OTMP[4][7] , \OTMP[4][6] , \OTMP[4][5] , \OTMP[4][4] ,
         \OTMP[4][3] , \OTMP[4][2] , \OTMP[4][1] , \OTMP[3][39] ,
         \OTMP[3][38] , \OTMP[3][37] , \OTMP[3][36] , \OTMP[3][35] ,
         \OTMP[3][34] , \OTMP[3][33] , \OTMP[3][32] , \OTMP[3][31] ,
         \OTMP[3][30] , \OTMP[3][29] , \OTMP[3][28] , \OTMP[3][27] ,
         \OTMP[3][26] , \OTMP[3][25] , \OTMP[3][24] , \OTMP[3][23] ,
         \OTMP[3][22] , \OTMP[3][21] , \OTMP[3][20] , \OTMP[3][19] ,
         \OTMP[3][18] , \OTMP[3][17] , \OTMP[3][16] , \OTMP[3][15] ,
         \OTMP[3][14] , \OTMP[3][13] , \OTMP[3][12] , \OTMP[3][11] ,
         \OTMP[3][10] , \OTMP[3][9] , \OTMP[3][8] , \OTMP[3][7] , \OTMP[3][6] ,
         \OTMP[3][5] , \OTMP[3][4] , \OTMP[3][3] , \OTMP[3][2] , \OTMP[3][1] ,
         \OTMP[2][37] , \OTMP[2][36] , \OTMP[2][35] , \OTMP[2][34] ,
         \OTMP[2][33] , \OTMP[2][32] , \OTMP[2][31] , \OTMP[2][30] ,
         \OTMP[2][29] , \OTMP[2][28] , \OTMP[2][27] , \OTMP[2][26] ,
         \OTMP[2][25] , \OTMP[2][24] , \OTMP[2][23] , \OTMP[2][22] ,
         \OTMP[2][21] , \OTMP[2][20] , \OTMP[2][19] , \OTMP[2][18] ,
         \OTMP[2][17] , \OTMP[2][16] , \OTMP[2][15] , \OTMP[2][14] ,
         \OTMP[2][13] , \OTMP[2][12] , \OTMP[2][11] , \OTMP[2][10] ,
         \OTMP[2][9] , \OTMP[2][8] , \OTMP[2][7] , \OTMP[2][6] , \OTMP[2][5] ,
         \OTMP[2][4] , \OTMP[2][3] , \OTMP[2][2] , \OTMP[2][1] , \OTMP[1][35] ,
         \OTMP[1][34] , \OTMP[1][33] , \OTMP[1][32] , \OTMP[1][31] ,
         \OTMP[1][30] , \OTMP[1][29] , \OTMP[1][28] , \OTMP[1][27] ,
         \OTMP[1][26] , \OTMP[1][25] , \OTMP[1][24] , \OTMP[1][23] ,
         \OTMP[1][22] , \OTMP[1][21] , \OTMP[1][20] , \OTMP[1][19] ,
         \OTMP[1][18] , \OTMP[1][17] , \OTMP[1][16] , \OTMP[1][15] ,
         \OTMP[1][14] , \OTMP[1][13] , \OTMP[1][12] , \OTMP[1][11] ,
         \OTMP[1][10] , \OTMP[1][9] , \OTMP[1][8] , \OTMP[1][7] , \OTMP[1][6] ,
         \OTMP[1][5] , \OTMP[1][4] , \OTMP[1][3] , \OTMP[1][2] , \OTMP[1][1] ,
         \OTMP[0][34] , \OTMP[0][32] , \OTMP[0][31] , \OTMP[0][30] ,
         \OTMP[0][29] , \OTMP[0][28] , \OTMP[0][27] , \OTMP[0][26] ,
         \OTMP[0][25] , \OTMP[0][24] , \OTMP[0][23] , \OTMP[0][22] ,
         \OTMP[0][21] , \OTMP[0][20] , \OTMP[0][19] , \OTMP[0][18] ,
         \OTMP[0][17] , \OTMP[0][16] , \OTMP[0][15] , \OTMP[0][14] ,
         \OTMP[0][13] , \OTMP[0][12] , \OTMP[0][11] , \OTMP[0][10] ,
         \OTMP[0][9] , \OTMP[0][8] , \OTMP[0][7] , \OTMP[0][6] , \OTMP[0][5] ,
         \OTMP[0][4] , \OTMP[0][3] , \OTMP[0][2] , \OTMP[0][1] , \OTMP[0][0] ,
         \OTMP[15][63] , \OTMP[15][62] , \OTMP[15][61] , \OTMP[15][60] ,
         \OTMP[15][59] , \OTMP[15][58] , \OTMP[15][57] , \OTMP[15][56] ,
         \OTMP[15][55] , \OTMP[15][54] , \OTMP[15][53] , \OTMP[15][52] ,
         \OTMP[15][51] , \OTMP[15][50] , \OTMP[15][49] , \OTMP[15][48] ,
         \OTMP[15][47] , \OTMP[15][46] , \OTMP[15][45] , \OTMP[15][44] ,
         \OTMP[15][43] , \OTMP[15][42] , \OTMP[15][41] , \OTMP[15][40] ,
         \OTMP[15][39] , \OTMP[15][38] , \OTMP[15][37] , \OTMP[15][36] ,
         \OTMP[15][35] , \OTMP[15][34] , \OTMP[15][33] , \OTMP[15][32] ,
         \OTMP[15][31] , \OTMP[15][30] , \OTMP[15][29] , \OTMP[15][28] ,
         \OTMP[15][27] , \OTMP[15][26] , \OTMP[15][25] , \OTMP[15][24] ,
         \OTMP[15][23] , \OTMP[15][22] , \OTMP[15][21] , \OTMP[15][20] ,
         \OTMP[15][19] , \OTMP[15][18] , \OTMP[15][17] , \OTMP[15][16] ,
         \OTMP[15][15] , \OTMP[15][14] , \OTMP[15][13] , \OTMP[15][12] ,
         \OTMP[15][11] , \OTMP[15][10] , \OTMP[15][9] , \OTMP[15][8] ,
         \OTMP[15][7] , \OTMP[15][6] , \OTMP[15][5] , \OTMP[15][4] ,
         \OTMP[15][3] , \OTMP[15][2] , \OTMP[15][1] , \OTMP[14][61] ,
         \OTMP[14][60] , \OTMP[14][59] , \OTMP[14][58] , \OTMP[14][57] ,
         \OTMP[14][56] , \OTMP[14][55] , \OTMP[14][54] , \OTMP[14][53] ,
         \OTMP[14][52] , \OTMP[14][51] , \OTMP[14][50] , \OTMP[14][49] ,
         \OTMP[14][48] , \OTMP[14][47] , \OTMP[14][46] , \OTMP[14][45] ,
         \OTMP[14][44] , \OTMP[14][43] , \OTMP[14][42] , \OTMP[14][41] ,
         \OTMP[14][40] , \OTMP[14][39] , \OTMP[14][38] , \OTMP[14][37] ,
         \OTMP[14][36] , \OTMP[14][35] , \OTMP[14][34] , \OTMP[14][33] ,
         \OTMP[14][32] , \OTMP[14][31] , \OTMP[14][30] , \OTMP[14][29] ,
         \OTMP[14][28] , \OTMP[14][27] , \OTMP[14][26] , \OTMP[14][25] ,
         \OTMP[14][24] , \OTMP[14][23] , \OTMP[14][22] , \OTMP[14][21] ,
         \OTMP[14][20] , \OTMP[14][19] , \OTMP[14][18] , \OTMP[14][17] ,
         \OTMP[14][16] , \OTMP[14][15] , \OTMP[14][14] , \OTMP[14][13] ,
         \OTMP[14][12] , \OTMP[14][11] , \OTMP[14][10] , \OTMP[14][9] ,
         \OTMP[14][8] , \OTMP[14][7] , \OTMP[14][6] , \OTMP[14][5] ,
         \OTMP[14][4] , \OTMP[14][3] , \OTMP[14][2] , \OTMP[14][1] ,
         \OTMP[13][59] , \OTMP[13][58] , \OTMP[13][57] , \OTMP[13][56] ,
         \OTMP[13][55] , \OTMP[13][54] , \OTMP[13][53] , \OTMP[13][52] ,
         \OTMP[13][51] , \OTMP[13][50] , \OTMP[13][49] , \OTMP[13][48] ,
         \OTMP[13][47] , \OTMP[13][46] , \OTMP[13][45] , \OTMP[13][44] ,
         \OTMP[13][43] , \OTMP[13][42] , \OTMP[13][41] , \OTMP[13][40] ,
         \OTMP[13][39] , \OTMP[13][38] , \OTMP[13][37] , \OTMP[13][36] ,
         \OTMP[13][35] , \OTMP[13][34] , \OTMP[13][33] , \OTMP[13][32] ,
         \OTMP[13][31] , \OTMP[13][30] , \OTMP[13][29] , \OTMP[13][28] ,
         \OTMP[13][27] , \OTMP[13][26] , \OTMP[13][25] , \OTMP[13][24] ,
         \OTMP[13][23] , \OTMP[13][22] , \OTMP[13][21] , \OTMP[13][20] ,
         \OTMP[13][19] , \OTMP[13][18] , \OTMP[13][17] , \OTMP[13][16] ,
         \OTMP[13][15] , \OTMP[13][14] , \OTMP[13][13] , \OTMP[13][12] ,
         \OTMP[13][11] , \OTMP[13][10] , \OTMP[13][9] , \OTMP[13][8] ,
         \OTMP[13][7] , \OTMP[13][6] , \OTMP[13][5] , \OTMP[13][4] ,
         \OTMP[13][3] , \OTMP[13][2] , \OTMP[13][1] , \OTMP[12][57] ,
         \OTMP[12][56] , \OTMP[12][55] , \OTMP[12][54] , \OTMP[12][53] ,
         \OTMP[12][52] , \OTMP[12][51] , \OTMP[12][50] , \OTMP[12][49] ,
         \OTMP[12][48] , \OTMP[12][47] , \OTMP[12][46] , \OTMP[12][45] ,
         \OTMP[12][44] , \OTMP[12][43] , \OTMP[12][42] , \OTMP[12][41] ,
         \OTMP[12][40] , \OTMP[12][39] , \OTMP[12][38] , \OTMP[12][37] ,
         \OTMP[12][36] , \OTMP[12][35] , \OTMP[12][34] , \OTMP[12][33] ,
         \OTMP[12][32] , \OTMP[12][31] , \OTMP[12][30] , \OTMP[12][29] ,
         \OTMP[12][28] , \OTMP[12][27] , \OTMP[12][26] , \OTMP[12][25] ,
         \OTMP[12][24] , \OTMP[12][23] , \OTMP[12][22] , \OTMP[12][21] ,
         \OTMP[12][20] , \OTMP[12][19] , \OTMP[12][18] , \OTMP[12][17] ,
         \OTMP[12][16] , \OTMP[12][15] , \OTMP[12][14] , \OTMP[12][13] ,
         \OTMP[12][12] , \OTMP[12][11] , \OTMP[12][10] , \OTMP[12][9] ,
         \OTMP[12][8] , \OTMP[12][7] , \OTMP[12][6] , \OTMP[12][5] ,
         \OTMP[12][4] , \OTMP[12][3] , \OTMP[12][2] , \OTMP[12][1] ,
         \OTMP[11][55] , \OTMP[11][54] , \OTMP[11][53] , \OTMP[11][52] ,
         \OTMP[11][51] , \OTMP[11][50] , \OTMP[11][49] , \OTMP[11][48] ,
         \OTMP[11][47] , \OTMP[11][46] , \OTMP[11][45] , \OTMP[11][44] ,
         \OTMP[11][43] , \OTMP[11][42] , \OTMP[11][41] , \OTMP[11][40] ,
         \OTMP[11][39] , \OTMP[11][38] , \OTMP[11][37] , \OTMP[11][36] ,
         \OTMP[11][35] , \OTMP[11][34] , \OTMP[11][33] , \OTMP[11][32] ,
         \OTMP[11][31] , \OTMP[11][30] , \OTMP[11][29] , \OTMP[11][28] ,
         \OTMP[11][27] , \OTMP[11][26] , \OTMP[11][25] , \OTMP[11][24] ,
         \OTMP[11][23] , \OTMP[11][22] , \OTMP[11][21] , \OTMP[11][20] ,
         \OTMP[11][19] , \OTMP[11][18] , \OTMP[11][17] , \OTMP[11][16] ,
         \OTMP[11][15] , \OTMP[11][14] , \OTMP[11][13] , \OTMP[11][12] ,
         \OTMP[11][11] , \OTMP[11][10] , \OTMP[11][9] , \OTMP[11][8] ,
         \OTMP[11][7] , \OTMP[11][6] , \OTMP[11][5] , \OTMP[11][4] ,
         \OTMP[11][3] , \OTMP[11][2] , \OTMP[11][1] , \OTMP[10][53] ,
         \OTMP[10][52] , \OTMP[10][51] , \OTMP[10][50] , \OTMP[10][49] ,
         \OTMP[10][48] , \OTMP[10][47] , \OTMP[10][46] , \OTMP[10][45] ,
         \OTMP[10][44] , \OTMP[10][43] , \OTMP[10][42] , \OTMP[10][41] ,
         \OTMP[10][40] , \OTMP[10][39] , \OTMP[10][38] , \OTMP[10][37] ,
         \OTMP[10][36] , \OTMP[10][35] , \OTMP[10][34] , \OTMP[10][33] ,
         \OTMP[10][32] , \OTMP[10][31] , \OTMP[10][30] , \OTMP[10][29] ,
         \OTMP[10][28] , \OTMP[10][27] , \OTMP[10][26] , \OTMP[10][25] ,
         \OTMP[10][24] , \OTMP[10][23] , \OTMP[10][22] , \OTMP[10][21] ,
         \OTMP[10][20] , \OTMP[10][19] , \OTMP[10][18] , \OTMP[10][17] ,
         \OTMP[10][16] , \OTMP[10][15] , \OTMP[10][14] , \OTMP[10][13] ,
         \OTMP[10][12] , \OTMP[10][11] , \OTMP[10][10] , \OTMP[10][9] ,
         \OTMP[10][8] , \OTMP[10][7] , \OTMP[10][6] , \OTMP[10][5] ,
         \OTMP[10][4] , \OTMP[10][3] , \OTMP[10][2] , \OTMP[10][1] ,
         \OTMP[9][51] , \OTMP[9][50] , \OTMP[9][49] , \OTMP[9][48] ,
         \OTMP[9][47] , \OTMP[9][46] , \OTMP[9][45] , \OTMP[9][44] ,
         \OTMP[9][43] , \OTMP[9][42] , \OTMP[9][41] , \OTMP[9][40] ,
         \OTMP[9][39] , \OTMP[9][38] , \OTMP[9][37] , \OTMP[9][36] ,
         \OTMP[9][35] , \OTMP[9][34] , \OTMP[9][33] , \OTMP[9][32] ,
         \OTMP[9][31] , \OTMP[9][30] , \OTMP[9][29] , \OTMP[9][28] ,
         \OTMP[9][27] , \OTMP[9][26] , \OTMP[9][25] , \OTMP[9][24] ,
         \OTMP[9][23] , \OTMP[9][22] , \OTMP[9][21] , \OTMP[9][20] ,
         \OTMP[9][19] , \OTMP[9][18] , \OTMP[9][17] , \OTMP[9][16] ,
         \OTMP[9][15] , \OTMP[9][14] , \OTMP[9][13] , \OTMP[9][12] ,
         \OTMP[9][11] , \OTMP[9][10] , \OTMP[9][9] , \OTMP[9][8] ,
         \OTMP[9][7] , \OTMP[9][6] , \OTMP[9][5] , \OTMP[9][4] , \OTMP[9][3] ,
         \OTMP[9][2] , \OTMP[9][1] , \OTMP[8][49] , \OTMP[8][48] ,
         \OTMP[8][47] , \OTMP[8][46] , \OTMP[8][45] , \OTMP[8][44] ,
         \OTMP[8][43] , \OTMP[8][42] , \OTMP[8][41] , \OTMP[8][40] ,
         \OTMP[8][39] , \OTMP[8][38] , \OTMP[8][37] , \OTMP[8][36] ,
         \OTMP[8][35] , \OTMP[8][34] , \OTMP[8][33] , \OTMP[8][32] ,
         \OTMP[8][31] , \OTMP[8][30] , \OTMP[8][29] , \OTMP[8][28] ,
         \OTMP[8][27] , \OTMP[8][26] , \OTMP[8][25] , \OTMP[8][24] ,
         \OTMP[8][23] , \OTMP[8][22] , \OTMP[8][21] , \OTMP[8][20] ,
         \OTMP[8][19] , \OTMP[8][18] , \OTMP[8][17] , \OTMP[8][16] ,
         \PTMP[8][15] , \PTMP[8][14] , \PTMP[8][13] , \PTMP[8][12] ,
         \PTMP[8][11] , \PTMP[8][10] , \PTMP[8][9] , \PTMP[8][8] ,
         \PTMP[8][7] , \PTMP[8][6] , \PTMP[8][5] , \PTMP[8][4] , \PTMP[8][3] ,
         \PTMP[8][2] , \PTMP[8][1] , \PTMP[8][0] , \PTMP[7][49] ,
         \PTMP[7][48] , \PTMP[7][47] , \PTMP[7][46] , \PTMP[7][45] ,
         \PTMP[7][44] , \PTMP[7][43] , \PTMP[7][42] , \PTMP[7][41] ,
         \PTMP[7][40] , \PTMP[7][39] , \PTMP[7][38] , \PTMP[7][37] ,
         \PTMP[7][36] , \PTMP[7][35] , \PTMP[7][34] , \PTMP[7][33] ,
         \PTMP[7][32] , \PTMP[7][31] , \PTMP[7][30] , \PTMP[7][29] ,
         \PTMP[7][28] , \PTMP[7][27] , \PTMP[7][26] , \PTMP[7][25] ,
         \PTMP[7][24] , \PTMP[7][23] , \PTMP[7][22] , \PTMP[7][21] ,
         \PTMP[7][20] , \PTMP[7][19] , \PTMP[7][18] , \PTMP[7][17] ,
         \PTMP[7][16] , \PTMP[7][15] , \PTMP[7][14] , \PTMP[7][13] ,
         \PTMP[7][12] , \PTMP[7][11] , \PTMP[7][10] , \PTMP[7][9] ,
         \PTMP[7][8] , \PTMP[7][7] , \PTMP[7][6] , \PTMP[7][5] , \PTMP[7][4] ,
         \PTMP[7][3] , \PTMP[7][2] , \PTMP[7][1] , \PTMP[7][0] , \PTMP[6][47] ,
         \PTMP[6][46] , \PTMP[6][45] , \PTMP[6][44] , \PTMP[6][43] ,
         \PTMP[6][42] , \PTMP[6][41] , \PTMP[6][40] , \PTMP[6][39] ,
         \PTMP[6][38] , \PTMP[6][37] , \PTMP[6][36] , \PTMP[6][35] ,
         \PTMP[6][34] , \PTMP[6][33] , \PTMP[6][32] , \PTMP[6][31] ,
         \PTMP[6][30] , \PTMP[6][29] , \PTMP[6][28] , \PTMP[6][27] ,
         \PTMP[6][26] , \PTMP[6][25] , \PTMP[6][24] , \PTMP[6][23] ,
         \PTMP[6][22] , \PTMP[6][21] , \PTMP[6][20] , \PTMP[6][19] ,
         \PTMP[6][18] , \PTMP[6][17] , \PTMP[6][16] , \PTMP[6][15] ,
         \PTMP[6][14] , \PTMP[6][13] , \PTMP[6][12] , \PTMP[6][11] ,
         \PTMP[6][10] , \PTMP[6][9] , \PTMP[6][8] , \PTMP[6][7] , \PTMP[6][6] ,
         \PTMP[6][5] , \PTMP[6][4] , \PTMP[6][3] , \PTMP[6][2] , \PTMP[6][1] ,
         \PTMP[6][0] , \PTMP[5][45] , \PTMP[5][44] , \PTMP[5][43] ,
         \PTMP[5][42] , \PTMP[5][41] , \PTMP[5][40] , \PTMP[5][39] ,
         \PTMP[5][38] , \PTMP[5][37] , \PTMP[5][36] , \PTMP[5][35] ,
         \PTMP[5][34] , \PTMP[5][33] , \PTMP[5][32] , \PTMP[5][31] ,
         \PTMP[5][30] , \PTMP[5][29] , \PTMP[5][28] , \PTMP[5][27] ,
         \PTMP[5][26] , \PTMP[5][25] , \PTMP[5][24] , \PTMP[5][23] ,
         \PTMP[5][22] , \PTMP[5][21] , \PTMP[5][20] , \PTMP[5][19] ,
         \PTMP[5][18] , \PTMP[5][17] , \PTMP[5][16] , \PTMP[5][15] ,
         \PTMP[5][14] , \PTMP[5][13] , \PTMP[5][12] , \PTMP[5][11] ,
         \PTMP[5][10] , \PTMP[5][9] , \PTMP[5][8] , \PTMP[5][7] , \PTMP[5][6] ,
         \PTMP[5][5] , \PTMP[5][4] , \PTMP[5][3] , \PTMP[5][2] , \PTMP[5][1] ,
         \PTMP[5][0] , \PTMP[4][43] , \PTMP[4][42] , \PTMP[4][41] ,
         \PTMP[4][40] , \PTMP[4][39] , \PTMP[4][38] , \PTMP[4][37] ,
         \PTMP[4][36] , \PTMP[4][35] , \PTMP[4][34] , \PTMP[4][33] ,
         \PTMP[4][32] , \PTMP[4][31] , \PTMP[4][30] , \PTMP[4][29] ,
         \PTMP[4][28] , \PTMP[4][27] , \PTMP[4][26] , \PTMP[4][25] ,
         \PTMP[4][24] , \PTMP[4][23] , \PTMP[4][22] , \PTMP[4][21] ,
         \PTMP[4][20] , \PTMP[4][19] , \PTMP[4][18] , \PTMP[4][17] ,
         \PTMP[4][16] , \PTMP[4][15] , \PTMP[4][14] , \PTMP[4][13] ,
         \PTMP[4][12] , \PTMP[4][11] , \PTMP[4][10] , \PTMP[4][9] ,
         \PTMP[4][8] , \PTMP[4][7] , \PTMP[4][6] , \PTMP[4][5] , \PTMP[4][4] ,
         \PTMP[4][3] , \PTMP[4][2] , \PTMP[4][1] , \PTMP[4][0] , \PTMP[3][41] ,
         \PTMP[3][40] , \PTMP[3][39] , \PTMP[3][38] , \PTMP[3][37] ,
         \PTMP[3][36] , \PTMP[3][35] , \PTMP[3][34] , \PTMP[3][33] ,
         \PTMP[3][32] , \PTMP[3][31] , \PTMP[3][30] , \PTMP[3][29] ,
         \PTMP[3][28] , \PTMP[3][27] , \PTMP[3][26] , \PTMP[3][25] ,
         \PTMP[3][24] , \PTMP[3][23] , \PTMP[3][22] , \PTMP[3][21] ,
         \PTMP[3][20] , \PTMP[3][19] , \PTMP[3][18] , \PTMP[3][17] ,
         \PTMP[3][16] , \PTMP[3][15] , \PTMP[3][14] , \PTMP[3][13] ,
         \PTMP[3][12] , \PTMP[3][11] , \PTMP[3][10] , \PTMP[3][9] ,
         \PTMP[3][8] , \PTMP[3][7] , \PTMP[3][6] , \PTMP[3][5] , \PTMP[3][4] ,
         \PTMP[3][3] , \PTMP[3][2] , \PTMP[3][1] , \PTMP[3][0] , \PTMP[2][39] ,
         \PTMP[2][38] , \PTMP[2][37] , \PTMP[2][36] , \PTMP[2][35] ,
         \PTMP[2][34] , \PTMP[2][33] , \PTMP[2][32] , \PTMP[2][31] ,
         \PTMP[2][30] , \PTMP[2][29] , \PTMP[2][28] , \PTMP[2][27] ,
         \PTMP[2][26] , \PTMP[2][25] , \PTMP[2][24] , \PTMP[2][23] ,
         \PTMP[2][22] , \PTMP[2][21] , \PTMP[2][20] , \PTMP[2][19] ,
         \PTMP[2][18] , \PTMP[2][17] , \PTMP[2][16] , \PTMP[2][15] ,
         \PTMP[2][14] , \PTMP[2][13] , \PTMP[2][12] , \PTMP[2][11] ,
         \PTMP[2][10] , \PTMP[2][9] , \PTMP[2][8] , \PTMP[2][7] , \PTMP[2][6] ,
         \PTMP[2][5] , \PTMP[2][4] , \PTMP[2][3] , \PTMP[2][2] , \PTMP[2][1] ,
         \PTMP[2][0] , \PTMP[1][37] , \PTMP[1][36] , \PTMP[1][35] ,
         \PTMP[1][34] , \PTMP[1][33] , \PTMP[1][32] , \PTMP[1][31] ,
         \PTMP[1][30] , \PTMP[1][29] , \PTMP[1][28] , \PTMP[1][27] ,
         \PTMP[1][26] , \PTMP[1][25] , \PTMP[1][24] , \PTMP[1][23] ,
         \PTMP[1][22] , \PTMP[1][21] , \PTMP[1][20] , \PTMP[1][19] ,
         \PTMP[1][18] , \PTMP[1][17] , \PTMP[1][16] , \PTMP[1][15] ,
         \PTMP[1][14] , \PTMP[1][13] , \PTMP[1][12] , \PTMP[1][11] ,
         \PTMP[1][10] , \PTMP[1][9] , \PTMP[1][8] , \PTMP[1][7] , \PTMP[1][6] ,
         \PTMP[1][5] , \PTMP[1][4] , \PTMP[1][3] , \PTMP[1][2] , \PTMP[1][1] ,
         \PTMP[1][0] , \PTMP[0][36] , \PTMP[0][34] , \PTMP[0][33] ,
         \PTMP[0][32] , \PTMP[0][31] , \PTMP[0][30] , \PTMP[0][29] ,
         \PTMP[0][28] , \PTMP[0][27] , \PTMP[0][26] , \PTMP[0][25] ,
         \PTMP[0][24] , \PTMP[0][23] , \PTMP[0][22] , \PTMP[0][21] ,
         \PTMP[0][20] , \PTMP[0][19] , \PTMP[0][18] , \PTMP[0][17] ,
         \PTMP[0][16] , \PTMP[0][15] , \PTMP[0][14] , \PTMP[0][13] ,
         \PTMP[0][12] , \PTMP[0][11] , \PTMP[0][10] , \PTMP[0][9] ,
         \PTMP[0][8] , \PTMP[0][7] , \PTMP[0][6] , \PTMP[0][5] , \PTMP[0][4] ,
         \PTMP[0][3] , \PTMP[0][2] , \PTMP[0][1] , \PTMP[0][0] ,
         \PTMP[13][61] , \PTMP[13][60] , \PTMP[13][59] , \PTMP[13][58] ,
         \PTMP[13][57] , \PTMP[13][56] , \PTMP[13][55] , \PTMP[13][54] ,
         \PTMP[13][53] , \PTMP[13][52] , \PTMP[13][51] , \PTMP[13][50] ,
         \PTMP[13][49] , \PTMP[13][48] , \PTMP[13][47] , \PTMP[13][46] ,
         \PTMP[13][45] , \PTMP[13][44] , \PTMP[13][43] , \PTMP[13][42] ,
         \PTMP[13][41] , \PTMP[13][40] , \PTMP[13][39] , \PTMP[13][38] ,
         \PTMP[13][37] , \PTMP[13][36] , \PTMP[13][35] , \PTMP[13][34] ,
         \PTMP[13][33] , \PTMP[13][32] , \PTMP[13][31] , \PTMP[13][30] ,
         \PTMP[13][29] , \PTMP[13][28] , \PTMP[13][27] , \PTMP[13][26] ,
         \PTMP[13][25] , \PTMP[13][24] , \PTMP[13][23] , \PTMP[13][22] ,
         \PTMP[13][21] , \PTMP[13][20] , \PTMP[13][19] , \PTMP[13][18] ,
         \PTMP[13][17] , \PTMP[13][16] , \PTMP[13][15] , \PTMP[13][14] ,
         \PTMP[13][13] , \PTMP[13][12] , \PTMP[13][11] , \PTMP[13][10] ,
         \PTMP[13][9] , \PTMP[13][8] , \PTMP[13][7] , \PTMP[13][6] ,
         \PTMP[13][5] , \PTMP[13][4] , \PTMP[13][3] , \PTMP[13][2] ,
         \PTMP[13][1] , \PTMP[13][0] , \PTMP[12][59] , \PTMP[12][58] ,
         \PTMP[12][57] , \PTMP[12][56] , \PTMP[12][55] , \PTMP[12][54] ,
         \PTMP[12][53] , \PTMP[12][52] , \PTMP[12][51] , \PTMP[12][50] ,
         \PTMP[12][49] , \PTMP[12][48] , \PTMP[12][47] , \PTMP[12][46] ,
         \PTMP[12][45] , \PTMP[12][44] , \PTMP[12][43] , \PTMP[12][42] ,
         \PTMP[12][41] , \PTMP[12][40] , \PTMP[12][39] , \PTMP[12][38] ,
         \PTMP[12][37] , \PTMP[12][36] , \PTMP[12][35] , \PTMP[12][34] ,
         \PTMP[12][33] , \PTMP[12][32] , \PTMP[12][31] , \PTMP[12][30] ,
         \PTMP[12][29] , \PTMP[12][28] , \PTMP[12][27] , \PTMP[12][26] ,
         \PTMP[12][25] , \PTMP[12][24] , \PTMP[12][23] , \PTMP[12][22] ,
         \PTMP[12][21] , \PTMP[12][20] , \PTMP[12][19] , \PTMP[12][18] ,
         \PTMP[12][17] , \PTMP[12][16] , \PTMP[12][15] , \PTMP[12][14] ,
         \PTMP[12][13] , \PTMP[12][12] , \PTMP[12][11] , \PTMP[12][10] ,
         \PTMP[12][9] , \PTMP[12][8] , \PTMP[12][7] , \PTMP[12][6] ,
         \PTMP[12][5] , \PTMP[12][4] , \PTMP[12][3] , \PTMP[12][2] ,
         \PTMP[12][1] , \PTMP[12][0] , \PTMP[11][57] , \PTMP[11][56] ,
         \PTMP[11][55] , \PTMP[11][54] , \PTMP[11][53] , \PTMP[11][52] ,
         \PTMP[11][51] , \PTMP[11][50] , \PTMP[11][49] , \PTMP[11][48] ,
         \PTMP[11][47] , \PTMP[11][46] , \PTMP[11][45] , \PTMP[11][44] ,
         \PTMP[11][43] , \PTMP[11][42] , \PTMP[11][41] , \PTMP[11][40] ,
         \PTMP[11][39] , \PTMP[11][38] , \PTMP[11][37] , \PTMP[11][36] ,
         \PTMP[11][35] , \PTMP[11][34] , \PTMP[11][33] , \PTMP[11][32] ,
         \PTMP[11][31] , \PTMP[11][30] , \PTMP[11][29] , \PTMP[11][28] ,
         \PTMP[11][27] , \PTMP[11][26] , \PTMP[11][25] , \PTMP[11][24] ,
         \PTMP[11][23] , \PTMP[11][22] , \PTMP[11][21] , \PTMP[11][20] ,
         \PTMP[11][19] , \PTMP[11][18] , \PTMP[11][17] , \PTMP[11][16] ,
         \PTMP[11][15] , \PTMP[11][14] , \PTMP[11][13] , \PTMP[11][12] ,
         \PTMP[11][11] , \PTMP[11][10] , \PTMP[11][9] , \PTMP[11][8] ,
         \PTMP[11][7] , \PTMP[11][6] , \PTMP[11][5] , \PTMP[11][4] ,
         \PTMP[11][3] , \PTMP[11][2] , \PTMP[11][1] , \PTMP[11][0] ,
         \PTMP[10][55] , \PTMP[10][54] , \PTMP[10][53] , \PTMP[10][52] ,
         \PTMP[10][51] , \PTMP[10][50] , \PTMP[10][49] , \PTMP[10][48] ,
         \PTMP[10][47] , \PTMP[10][46] , \PTMP[10][45] , \PTMP[10][44] ,
         \PTMP[10][43] , \PTMP[10][42] , \PTMP[10][41] , \PTMP[10][40] ,
         \PTMP[10][39] , \PTMP[10][38] , \PTMP[10][37] , \PTMP[10][36] ,
         \PTMP[10][35] , \PTMP[10][34] , \PTMP[10][33] , \PTMP[10][32] ,
         \PTMP[10][31] , \PTMP[10][30] , \PTMP[10][29] , \PTMP[10][28] ,
         \PTMP[10][27] , \PTMP[10][26] , \PTMP[10][25] , \PTMP[10][24] ,
         \PTMP[10][23] , \PTMP[10][22] , \PTMP[10][21] , \PTMP[10][20] ,
         \PTMP[10][19] , \PTMP[10][18] , \PTMP[10][17] , \PTMP[10][16] ,
         \PTMP[10][15] , \PTMP[10][14] , \PTMP[10][13] , \PTMP[10][12] ,
         \PTMP[10][11] , \PTMP[10][10] , \PTMP[10][9] , \PTMP[10][8] ,
         \PTMP[10][7] , \PTMP[10][6] , \PTMP[10][5] , \PTMP[10][4] ,
         \PTMP[10][3] , \PTMP[10][2] , \PTMP[10][1] , \PTMP[10][0] ,
         \PTMP[9][53] , \PTMP[9][52] , \PTMP[9][51] , \PTMP[9][50] ,
         \PTMP[9][49] , \PTMP[9][48] , \PTMP[9][47] , \PTMP[9][46] ,
         \PTMP[9][45] , \PTMP[9][44] , \PTMP[9][43] , \PTMP[9][42] ,
         \PTMP[9][41] , \PTMP[9][40] , \PTMP[9][39] , \PTMP[9][38] ,
         \PTMP[9][37] , \PTMP[9][36] , \PTMP[9][35] , \PTMP[9][34] ,
         \PTMP[9][33] , \PTMP[9][32] , \PTMP[9][31] , \PTMP[9][30] ,
         \PTMP[9][29] , \PTMP[9][28] , \PTMP[9][27] , \PTMP[9][26] ,
         \PTMP[9][25] , \PTMP[9][24] , \PTMP[9][23] , \PTMP[9][22] ,
         \PTMP[9][21] , \PTMP[9][20] , \PTMP[9][19] , \PTMP[9][18] ,
         \PTMP[9][17] , \PTMP[9][16] , \PTMP[9][15] , \PTMP[9][14] ,
         \PTMP[9][13] , \PTMP[9][12] , \PTMP[9][11] , \PTMP[9][10] ,
         \PTMP[9][9] , \PTMP[9][8] , \PTMP[9][7] , \PTMP[9][6] , \PTMP[9][5] ,
         \PTMP[9][4] , \PTMP[9][3] , \PTMP[9][2] , \PTMP[9][1] , \PTMP[9][0] ,
         \PTMP[8][51] , \PTMP[8][50] , \PTMP[8][49] , \PTMP[8][48] ,
         \PTMP[8][47] , \PTMP[8][46] , \PTMP[8][45] , \PTMP[8][44] ,
         \PTMP[8][43] , \PTMP[8][42] , \PTMP[8][41] , \PTMP[8][40] ,
         \PTMP[8][39] , \PTMP[8][38] , \PTMP[8][37] , \PTMP[8][36] ,
         \PTMP[8][35] , \PTMP[8][34] , \PTMP[8][33] , \PTMP[8][32] ,
         \PTMP[8][31] , \PTMP[8][30] , \PTMP[8][29] , \PTMP[8][28] ,
         \PTMP[8][27] , \PTMP[8][26] , \PTMP[8][25] , \PTMP[8][24] ,
         \PTMP[8][23] , \PTMP[8][22] , \PTMP[8][21] , \PTMP[8][20] ,
         \PTMP[8][19] , \PTMP[8][18] , \PTMP[8][17] , \PTMP[8][16] , n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22;
  wire   [30:0] A_n;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72;

  BOOTHENC_NBIT34_i0 ENC1 ( .A_s({A[31], A[31], A[31:2], n11, A[0]}), .A_ns({
        A_n_65, A_n_65, A_n_65, A_n}), .B({B[31], B[31], B}), .O({
        \OTMP[0][34] , \OTMP[0][32] , \OTMP[0][31] , \OTMP[0][30] , 
        \OTMP[0][29] , \OTMP[0][28] , \OTMP[0][27] , \OTMP[0][26] , 
        \OTMP[0][25] , \OTMP[0][24] , \OTMP[0][23] , \OTMP[0][22] , 
        \OTMP[0][21] , \OTMP[0][20] , \OTMP[0][19] , \OTMP[0][18] , 
        \OTMP[0][17] , \OTMP[0][16] , \OTMP[0][15] , \OTMP[0][14] , 
        \OTMP[0][13] , \OTMP[0][12] , \OTMP[0][11] , \OTMP[0][10] , 
        \OTMP[0][9] , \OTMP[0][8] , \OTMP[0][7] , \OTMP[0][6] , \OTMP[0][5] , 
        \OTMP[0][4] , \OTMP[0][3] , \OTMP[0][2] , \OTMP[0][1] , \OTMP[0][0] }), 
        .A_so({\SHIFT[1][33] , \SHIFT[1][32] , \SHIFT[1][31] , \SHIFT[1][30] , 
        \SHIFT[1][29] , \SHIFT[1][28] , \SHIFT[1][27] , \SHIFT[1][26] , 
        \SHIFT[1][25] , \SHIFT[1][24] , \SHIFT[1][23] , \SHIFT[1][22] , 
        \SHIFT[1][21] , \SHIFT[1][20] , \SHIFT[1][19] , \SHIFT[1][18] , 
        \SHIFT[1][17] , \SHIFT[1][16] , \SHIFT[1][15] , \SHIFT[1][14] , 
        \SHIFT[1][13] , \SHIFT[1][12] , \SHIFT[1][11] , \SHIFT[1][10] , 
        \SHIFT[1][9] , \SHIFT[1][8] , \SHIFT[1][7] , \SHIFT[1][6] , 
        \SHIFT[1][5] , \SHIFT[1][4] , \SHIFT[1][3] , \SHIFT[1][2] , 
        \SHIFT[1][1] , SYNOPSYS_UNCONNECTED__0}), .A_nso({\SHIFT_n[1][33] , 
        \SHIFT_n[1][32] , \SHIFT_n[1][31] , \SHIFT_n[1][30] , \SHIFT_n[1][29] , 
        \SHIFT_n[1][28] , \SHIFT_n[1][27] , \SHIFT_n[1][26] , \SHIFT_n[1][25] , 
        \SHIFT_n[1][24] , \SHIFT_n[1][23] , \SHIFT_n[1][22] , \SHIFT_n[1][21] , 
        \SHIFT_n[1][20] , \SHIFT_n[1][19] , \SHIFT_n[1][18] , \SHIFT_n[1][17] , 
        \SHIFT_n[1][16] , \SHIFT_n[1][15] , \SHIFT_n[1][14] , \SHIFT_n[1][13] , 
        \SHIFT_n[1][12] , \SHIFT_n[1][11] , \SHIFT_n[1][10] , \SHIFT_n[1][9] , 
        \SHIFT_n[1][8] , \SHIFT_n[1][7] , \SHIFT_n[1][6] , \SHIFT_n[1][5] , 
        \SHIFT_n[1][4] , \SHIFT_n[1][3] , \SHIFT_n[1][2] , \SHIFT_n[1][1] , 
        SYNOPSYS_UNCONNECTED__1}) );
  BOOTHENC_NBIT36_i2 ENC_1 ( .A_s({\SHIFT[1][33] , \SHIFT[1][33] , 
        \SHIFT[1][33] , \SHIFT[1][32] , \SHIFT[1][31] , \SHIFT[1][30] , 
        \SHIFT[1][29] , \SHIFT[1][28] , \SHIFT[1][27] , \SHIFT[1][26] , 
        \SHIFT[1][25] , \SHIFT[1][24] , \SHIFT[1][23] , \SHIFT[1][22] , 
        \SHIFT[1][21] , \SHIFT[1][20] , \SHIFT[1][19] , \SHIFT[1][18] , 
        \SHIFT[1][17] , \SHIFT[1][16] , \SHIFT[1][15] , \SHIFT[1][14] , 
        \SHIFT[1][13] , \SHIFT[1][12] , \SHIFT[1][11] , \SHIFT[1][10] , 
        \SHIFT[1][9] , \SHIFT[1][8] , \SHIFT[1][7] , \SHIFT[1][6] , 
        \SHIFT[1][5] , \SHIFT[1][4] , \SHIFT[1][3] , \SHIFT[1][2] , 
        \SHIFT[1][1] , 1'b0}), .A_ns({\SHIFT_n[1][33] , \SHIFT_n[1][33] , 
        \SHIFT_n[1][33] , \SHIFT_n[1][32] , \SHIFT_n[1][31] , \SHIFT_n[1][30] , 
        \SHIFT_n[1][29] , \SHIFT_n[1][28] , \SHIFT_n[1][27] , \SHIFT_n[1][26] , 
        \SHIFT_n[1][25] , \SHIFT_n[1][24] , \SHIFT_n[1][23] , \SHIFT_n[1][22] , 
        \SHIFT_n[1][21] , \SHIFT_n[1][20] , \SHIFT_n[1][19] , \SHIFT_n[1][18] , 
        \SHIFT_n[1][17] , \SHIFT_n[1][16] , \SHIFT_n[1][15] , \SHIFT_n[1][14] , 
        \SHIFT_n[1][13] , \SHIFT_n[1][12] , \SHIFT_n[1][11] , \SHIFT_n[1][10] , 
        \SHIFT_n[1][9] , \SHIFT_n[1][8] , \SHIFT_n[1][7] , \SHIFT_n[1][6] , 
        \SHIFT_n[1][5] , \SHIFT_n[1][4] , \SHIFT_n[1][3] , \SHIFT_n[1][2] , 
        \SHIFT_n[1][1] , 1'b0}), .B({B[31], B[31], B[31], B[31], B}), .O({
        \OTMP[1][35] , \OTMP[1][34] , \OTMP[1][33] , \OTMP[1][32] , 
        \OTMP[1][31] , \OTMP[1][30] , \OTMP[1][29] , \OTMP[1][28] , 
        \OTMP[1][27] , \OTMP[1][26] , \OTMP[1][25] , \OTMP[1][24] , 
        \OTMP[1][23] , \OTMP[1][22] , \OTMP[1][21] , \OTMP[1][20] , 
        \OTMP[1][19] , \OTMP[1][18] , \OTMP[1][17] , \OTMP[1][16] , 
        \OTMP[1][15] , \OTMP[1][14] , \OTMP[1][13] , \OTMP[1][12] , 
        \OTMP[1][11] , \OTMP[1][10] , \OTMP[1][9] , \OTMP[1][8] , \OTMP[1][7] , 
        \OTMP[1][6] , \OTMP[1][5] , \OTMP[1][4] , \OTMP[1][3] , \OTMP[1][2] , 
        \OTMP[1][1] , SYNOPSYS_UNCONNECTED__2}), .A_so({\SHIFT[2][35] , 
        \SHIFT[2][34] , \SHIFT[2][33] , \SHIFT[2][32] , \SHIFT[2][31] , 
        \SHIFT[2][30] , \SHIFT[2][29] , \SHIFT[2][28] , \SHIFT[2][27] , 
        \SHIFT[2][26] , \SHIFT[2][25] , \SHIFT[2][24] , \SHIFT[2][23] , 
        \SHIFT[2][22] , \SHIFT[2][21] , \SHIFT[2][20] , \SHIFT[2][19] , 
        \SHIFT[2][18] , \SHIFT[2][17] , \SHIFT[2][16] , \SHIFT[2][15] , 
        \SHIFT[2][14] , \SHIFT[2][13] , \SHIFT[2][12] , \SHIFT[2][11] , 
        \SHIFT[2][10] , \SHIFT[2][9] , \SHIFT[2][8] , \SHIFT[2][7] , 
        \SHIFT[2][6] , \SHIFT[2][5] , \SHIFT[2][4] , \SHIFT[2][3] , 
        \SHIFT[2][2] , SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4}), 
        .A_nso({\SHIFT_n[2][35] , \SHIFT_n[2][34] , \SHIFT_n[2][33] , 
        \SHIFT_n[2][32] , \SHIFT_n[2][31] , \SHIFT_n[2][30] , \SHIFT_n[2][29] , 
        \SHIFT_n[2][28] , \SHIFT_n[2][27] , \SHIFT_n[2][26] , \SHIFT_n[2][25] , 
        \SHIFT_n[2][24] , \SHIFT_n[2][23] , \SHIFT_n[2][22] , \SHIFT_n[2][21] , 
        \SHIFT_n[2][20] , \SHIFT_n[2][19] , \SHIFT_n[2][18] , \SHIFT_n[2][17] , 
        \SHIFT_n[2][16] , \SHIFT_n[2][15] , \SHIFT_n[2][14] , \SHIFT_n[2][13] , 
        \SHIFT_n[2][12] , \SHIFT_n[2][11] , \SHIFT_n[2][10] , \SHIFT_n[2][9] , 
        \SHIFT_n[2][8] , \SHIFT_n[2][7] , \SHIFT_n[2][6] , \SHIFT_n[2][5] , 
        \SHIFT_n[2][4] , \SHIFT_n[2][3] , \SHIFT_n[2][2] , 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6}) );
  BOOTHENC_NBIT38_i4 ENC_2 ( .A_s({\SHIFT[2][35] , \SHIFT[2][35] , 
        \SHIFT[2][35] , \SHIFT[2][34] , \SHIFT[2][33] , \SHIFT[2][32] , 
        \SHIFT[2][31] , \SHIFT[2][30] , \SHIFT[2][29] , \SHIFT[2][28] , 
        \SHIFT[2][27] , \SHIFT[2][26] , \SHIFT[2][25] , \SHIFT[2][24] , 
        \SHIFT[2][23] , \SHIFT[2][22] , \SHIFT[2][21] , \SHIFT[2][20] , 
        \SHIFT[2][19] , \SHIFT[2][18] , \SHIFT[2][17] , \SHIFT[2][16] , 
        \SHIFT[2][15] , \SHIFT[2][14] , \SHIFT[2][13] , \SHIFT[2][12] , 
        \SHIFT[2][11] , \SHIFT[2][10] , \SHIFT[2][9] , \SHIFT[2][8] , 
        \SHIFT[2][7] , \SHIFT[2][6] , \SHIFT[2][5] , \SHIFT[2][4] , 
        \SHIFT[2][3] , \SHIFT[2][2] , 1'b0, 1'b0}), .A_ns({\SHIFT_n[2][35] , 
        \SHIFT_n[2][35] , \SHIFT_n[2][35] , \SHIFT_n[2][34] , \SHIFT_n[2][33] , 
        \SHIFT_n[2][32] , \SHIFT_n[2][31] , \SHIFT_n[2][30] , \SHIFT_n[2][29] , 
        \SHIFT_n[2][28] , \SHIFT_n[2][27] , \SHIFT_n[2][26] , \SHIFT_n[2][25] , 
        \SHIFT_n[2][24] , \SHIFT_n[2][23] , \SHIFT_n[2][22] , \SHIFT_n[2][21] , 
        \SHIFT_n[2][20] , \SHIFT_n[2][19] , \SHIFT_n[2][18] , \SHIFT_n[2][17] , 
        \SHIFT_n[2][16] , \SHIFT_n[2][15] , \SHIFT_n[2][14] , \SHIFT_n[2][13] , 
        \SHIFT_n[2][12] , \SHIFT_n[2][11] , \SHIFT_n[2][10] , \SHIFT_n[2][9] , 
        \SHIFT_n[2][8] , \SHIFT_n[2][7] , \SHIFT_n[2][6] , \SHIFT_n[2][5] , 
        \SHIFT_n[2][4] , \SHIFT_n[2][3] , \SHIFT_n[2][2] , 1'b0, 1'b0}), .B({
        B[31], B[31], B[31], B[31], B[31], B[31], B}), .O({\OTMP[2][37] , 
        \OTMP[2][36] , \OTMP[2][35] , \OTMP[2][34] , \OTMP[2][33] , 
        \OTMP[2][32] , \OTMP[2][31] , \OTMP[2][30] , \OTMP[2][29] , 
        \OTMP[2][28] , \OTMP[2][27] , \OTMP[2][26] , \OTMP[2][25] , 
        \OTMP[2][24] , \OTMP[2][23] , \OTMP[2][22] , \OTMP[2][21] , 
        \OTMP[2][20] , \OTMP[2][19] , \OTMP[2][18] , \OTMP[2][17] , 
        \OTMP[2][16] , \OTMP[2][15] , \OTMP[2][14] , \OTMP[2][13] , 
        \OTMP[2][12] , \OTMP[2][11] , \OTMP[2][10] , \OTMP[2][9] , 
        \OTMP[2][8] , \OTMP[2][7] , \OTMP[2][6] , \OTMP[2][5] , \OTMP[2][4] , 
        \OTMP[2][3] , \OTMP[2][2] , \OTMP[2][1] , SYNOPSYS_UNCONNECTED__7}), 
        .A_so({\SHIFT[3][37] , \SHIFT[3][36] , \SHIFT[3][35] , \SHIFT[3][34] , 
        \SHIFT[3][33] , \SHIFT[3][32] , \SHIFT[3][31] , \SHIFT[3][30] , 
        \SHIFT[3][29] , \SHIFT[3][28] , \SHIFT[3][27] , \SHIFT[3][26] , 
        \SHIFT[3][25] , \SHIFT[3][24] , \SHIFT[3][23] , \SHIFT[3][22] , 
        \SHIFT[3][21] , \SHIFT[3][20] , \SHIFT[3][19] , \SHIFT[3][18] , 
        \SHIFT[3][17] , \SHIFT[3][16] , \SHIFT[3][15] , \SHIFT[3][14] , 
        \SHIFT[3][13] , \SHIFT[3][12] , \SHIFT[3][11] , \SHIFT[3][10] , 
        \SHIFT[3][9] , \SHIFT[3][8] , \SHIFT[3][7] , \SHIFT[3][6] , 
        \SHIFT[3][5] , \SHIFT[3][4] , \SHIFT[3][3] , \SHIFT[3][2] , 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9}), .A_nso({
        \SHIFT_n[3][37] , \SHIFT_n[3][36] , \SHIFT_n[3][35] , \SHIFT_n[3][34] , 
        \SHIFT_n[3][33] , \SHIFT_n[3][32] , \SHIFT_n[3][31] , \SHIFT_n[3][30] , 
        \SHIFT_n[3][29] , \SHIFT_n[3][28] , \SHIFT_n[3][27] , \SHIFT_n[3][26] , 
        \SHIFT_n[3][25] , \SHIFT_n[3][24] , \SHIFT_n[3][23] , \SHIFT_n[3][22] , 
        \SHIFT_n[3][21] , \SHIFT_n[3][20] , \SHIFT_n[3][19] , \SHIFT_n[3][18] , 
        \SHIFT_n[3][17] , \SHIFT_n[3][16] , \SHIFT_n[3][15] , \SHIFT_n[3][14] , 
        \SHIFT_n[3][13] , \SHIFT_n[3][12] , \SHIFT_n[3][11] , \SHIFT_n[3][10] , 
        \SHIFT_n[3][9] , \SHIFT_n[3][8] , \SHIFT_n[3][7] , \SHIFT_n[3][6] , 
        \SHIFT_n[3][5] , \SHIFT_n[3][4] , \SHIFT_n[3][3] , \SHIFT_n[3][2] , 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11}) );
  BOOTHENC_NBIT40_i6 ENC_3 ( .A_s({\SHIFT[3][37] , \SHIFT[3][37] , 
        \SHIFT[3][37] , \SHIFT[3][36] , \SHIFT[3][35] , \SHIFT[3][34] , 
        \SHIFT[3][33] , \SHIFT[3][32] , \SHIFT[3][31] , \SHIFT[3][30] , 
        \SHIFT[3][29] , \SHIFT[3][28] , \SHIFT[3][27] , \SHIFT[3][26] , 
        \SHIFT[3][25] , \SHIFT[3][24] , \SHIFT[3][23] , \SHIFT[3][22] , 
        \SHIFT[3][21] , \SHIFT[3][20] , \SHIFT[3][19] , \SHIFT[3][18] , 
        \SHIFT[3][17] , \SHIFT[3][16] , \SHIFT[3][15] , \SHIFT[3][14] , 
        \SHIFT[3][13] , \SHIFT[3][12] , \SHIFT[3][11] , \SHIFT[3][10] , 
        \SHIFT[3][9] , \SHIFT[3][8] , \SHIFT[3][7] , \SHIFT[3][6] , 
        \SHIFT[3][5] , \SHIFT[3][4] , \SHIFT[3][3] , \SHIFT[3][2] , 1'b0, 1'b0}), .A_ns({\SHIFT_n[3][37] , \SHIFT_n[3][37] , \SHIFT_n[3][37] , 
        \SHIFT_n[3][36] , \SHIFT_n[3][35] , \SHIFT_n[3][34] , \SHIFT_n[3][33] , 
        \SHIFT_n[3][32] , \SHIFT_n[3][31] , \SHIFT_n[3][30] , \SHIFT_n[3][29] , 
        \SHIFT_n[3][28] , \SHIFT_n[3][27] , \SHIFT_n[3][26] , \SHIFT_n[3][25] , 
        \SHIFT_n[3][24] , \SHIFT_n[3][23] , \SHIFT_n[3][22] , \SHIFT_n[3][21] , 
        \SHIFT_n[3][20] , \SHIFT_n[3][19] , \SHIFT_n[3][18] , \SHIFT_n[3][17] , 
        \SHIFT_n[3][16] , \SHIFT_n[3][15] , \SHIFT_n[3][14] , \SHIFT_n[3][13] , 
        \SHIFT_n[3][12] , \SHIFT_n[3][11] , \SHIFT_n[3][10] , \SHIFT_n[3][9] , 
        \SHIFT_n[3][8] , \SHIFT_n[3][7] , \SHIFT_n[3][6] , \SHIFT_n[3][5] , 
        \SHIFT_n[3][4] , \SHIFT_n[3][3] , \SHIFT_n[3][2] , 1'b0, 1'b0}), .B({
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B}), .O({
        \OTMP[3][39] , \OTMP[3][38] , \OTMP[3][37] , \OTMP[3][36] , 
        \OTMP[3][35] , \OTMP[3][34] , \OTMP[3][33] , \OTMP[3][32] , 
        \OTMP[3][31] , \OTMP[3][30] , \OTMP[3][29] , \OTMP[3][28] , 
        \OTMP[3][27] , \OTMP[3][26] , \OTMP[3][25] , \OTMP[3][24] , 
        \OTMP[3][23] , \OTMP[3][22] , \OTMP[3][21] , \OTMP[3][20] , 
        \OTMP[3][19] , \OTMP[3][18] , \OTMP[3][17] , \OTMP[3][16] , 
        \OTMP[3][15] , \OTMP[3][14] , \OTMP[3][13] , \OTMP[3][12] , 
        \OTMP[3][11] , \OTMP[3][10] , \OTMP[3][9] , \OTMP[3][8] , \OTMP[3][7] , 
        \OTMP[3][6] , \OTMP[3][5] , \OTMP[3][4] , \OTMP[3][3] , \OTMP[3][2] , 
        \OTMP[3][1] , SYNOPSYS_UNCONNECTED__12}), .A_so({\SHIFT[4][39] , 
        \SHIFT[4][38] , \SHIFT[4][37] , \SHIFT[4][36] , \SHIFT[4][35] , 
        \SHIFT[4][34] , \SHIFT[4][33] , \SHIFT[4][32] , \SHIFT[4][31] , 
        \SHIFT[4][30] , \SHIFT[4][29] , \SHIFT[4][28] , \SHIFT[4][27] , 
        \SHIFT[4][26] , \SHIFT[4][25] , \SHIFT[4][24] , \SHIFT[4][23] , 
        \SHIFT[4][22] , \SHIFT[4][21] , \SHIFT[4][20] , \SHIFT[4][19] , 
        \SHIFT[4][18] , \SHIFT[4][17] , \SHIFT[4][16] , \SHIFT[4][15] , 
        \SHIFT[4][14] , \SHIFT[4][13] , \SHIFT[4][12] , \SHIFT[4][11] , 
        \SHIFT[4][10] , \SHIFT[4][9] , \SHIFT[4][8] , \SHIFT[4][7] , 
        \SHIFT[4][6] , \SHIFT[4][5] , \SHIFT[4][4] , \SHIFT[4][3] , 
        \SHIFT[4][2] , SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14}), 
        .A_nso({\SHIFT_n[4][39] , \SHIFT_n[4][38] , \SHIFT_n[4][37] , 
        \SHIFT_n[4][36] , \SHIFT_n[4][35] , \SHIFT_n[4][34] , \SHIFT_n[4][33] , 
        \SHIFT_n[4][32] , \SHIFT_n[4][31] , \SHIFT_n[4][30] , \SHIFT_n[4][29] , 
        \SHIFT_n[4][28] , \SHIFT_n[4][27] , \SHIFT_n[4][26] , \SHIFT_n[4][25] , 
        \SHIFT_n[4][24] , \SHIFT_n[4][23] , \SHIFT_n[4][22] , \SHIFT_n[4][21] , 
        \SHIFT_n[4][20] , \SHIFT_n[4][19] , \SHIFT_n[4][18] , \SHIFT_n[4][17] , 
        \SHIFT_n[4][16] , \SHIFT_n[4][15] , \SHIFT_n[4][14] , \SHIFT_n[4][13] , 
        \SHIFT_n[4][12] , \SHIFT_n[4][11] , \SHIFT_n[4][10] , \SHIFT_n[4][9] , 
        \SHIFT_n[4][8] , \SHIFT_n[4][7] , \SHIFT_n[4][6] , \SHIFT_n[4][5] , 
        \SHIFT_n[4][4] , \SHIFT_n[4][3] , \SHIFT_n[4][2] , 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16}) );
  BOOTHENC_NBIT42_i8 ENC_4 ( .A_s({\SHIFT[4][39] , \SHIFT[4][39] , 
        \SHIFT[4][39] , \SHIFT[4][38] , \SHIFT[4][37] , \SHIFT[4][36] , 
        \SHIFT[4][35] , \SHIFT[4][34] , \SHIFT[4][33] , \SHIFT[4][32] , 
        \SHIFT[4][31] , \SHIFT[4][30] , \SHIFT[4][29] , \SHIFT[4][28] , 
        \SHIFT[4][27] , \SHIFT[4][26] , \SHIFT[4][25] , \SHIFT[4][24] , 
        \SHIFT[4][23] , \SHIFT[4][22] , \SHIFT[4][21] , \SHIFT[4][20] , 
        \SHIFT[4][19] , \SHIFT[4][18] , \SHIFT[4][17] , \SHIFT[4][16] , 
        \SHIFT[4][15] , \SHIFT[4][14] , \SHIFT[4][13] , \SHIFT[4][12] , 
        \SHIFT[4][11] , \SHIFT[4][10] , \SHIFT[4][9] , \SHIFT[4][8] , 
        \SHIFT[4][7] , \SHIFT[4][6] , \SHIFT[4][5] , \SHIFT[4][4] , 
        \SHIFT[4][3] , \SHIFT[4][2] , 1'b0, 1'b0}), .A_ns({\SHIFT_n[4][39] , 
        \SHIFT_n[4][39] , \SHIFT_n[4][39] , \SHIFT_n[4][38] , \SHIFT_n[4][37] , 
        \SHIFT_n[4][36] , \SHIFT_n[4][35] , \SHIFT_n[4][34] , \SHIFT_n[4][33] , 
        \SHIFT_n[4][32] , \SHIFT_n[4][31] , \SHIFT_n[4][30] , \SHIFT_n[4][29] , 
        \SHIFT_n[4][28] , \SHIFT_n[4][27] , \SHIFT_n[4][26] , \SHIFT_n[4][25] , 
        \SHIFT_n[4][24] , \SHIFT_n[4][23] , \SHIFT_n[4][22] , \SHIFT_n[4][21] , 
        \SHIFT_n[4][20] , \SHIFT_n[4][19] , \SHIFT_n[4][18] , \SHIFT_n[4][17] , 
        \SHIFT_n[4][16] , \SHIFT_n[4][15] , \SHIFT_n[4][14] , \SHIFT_n[4][13] , 
        \SHIFT_n[4][12] , \SHIFT_n[4][11] , \SHIFT_n[4][10] , \SHIFT_n[4][9] , 
        \SHIFT_n[4][8] , \SHIFT_n[4][7] , \SHIFT_n[4][6] , \SHIFT_n[4][5] , 
        \SHIFT_n[4][4] , \SHIFT_n[4][3] , \SHIFT_n[4][2] , 1'b0, 1'b0}), .B({
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B}), .O({\OTMP[4][41] , \OTMP[4][40] , \OTMP[4][39] , \OTMP[4][38] , 
        \OTMP[4][37] , \OTMP[4][36] , \OTMP[4][35] , \OTMP[4][34] , 
        \OTMP[4][33] , \OTMP[4][32] , \OTMP[4][31] , \OTMP[4][30] , 
        \OTMP[4][29] , \OTMP[4][28] , \OTMP[4][27] , \OTMP[4][26] , 
        \OTMP[4][25] , \OTMP[4][24] , \OTMP[4][23] , \OTMP[4][22] , 
        \OTMP[4][21] , \OTMP[4][20] , \OTMP[4][19] , \OTMP[4][18] , 
        \OTMP[4][17] , \OTMP[4][16] , \OTMP[4][15] , \OTMP[4][14] , 
        \OTMP[4][13] , \OTMP[4][12] , \OTMP[4][11] , \OTMP[4][10] , 
        \OTMP[4][9] , \OTMP[4][8] , \OTMP[4][7] , \OTMP[4][6] , \OTMP[4][5] , 
        \OTMP[4][4] , \OTMP[4][3] , \OTMP[4][2] , \OTMP[4][1] , 
        SYNOPSYS_UNCONNECTED__17}), .A_so({\SHIFT[5][41] , \SHIFT[5][40] , 
        \SHIFT[5][39] , \SHIFT[5][38] , \SHIFT[5][37] , \SHIFT[5][36] , 
        \SHIFT[5][35] , \SHIFT[5][34] , \SHIFT[5][33] , \SHIFT[5][32] , 
        \SHIFT[5][31] , \SHIFT[5][30] , \SHIFT[5][29] , \SHIFT[5][28] , 
        \SHIFT[5][27] , \SHIFT[5][26] , \SHIFT[5][25] , \SHIFT[5][24] , 
        \SHIFT[5][23] , \SHIFT[5][22] , \SHIFT[5][21] , \SHIFT[5][20] , 
        \SHIFT[5][19] , \SHIFT[5][18] , \SHIFT[5][17] , \SHIFT[5][16] , 
        \SHIFT[5][15] , \SHIFT[5][14] , \SHIFT[5][13] , \SHIFT[5][12] , 
        \SHIFT[5][11] , \SHIFT[5][10] , \SHIFT[5][9] , \SHIFT[5][8] , 
        \SHIFT[5][7] , \SHIFT[5][6] , \SHIFT[5][5] , \SHIFT[5][4] , 
        \SHIFT[5][3] , \SHIFT[5][2] , SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19}), .A_nso({\SHIFT_n[5][41] , \SHIFT_n[5][40] , 
        \SHIFT_n[5][39] , \SHIFT_n[5][38] , \SHIFT_n[5][37] , \SHIFT_n[5][36] , 
        \SHIFT_n[5][35] , \SHIFT_n[5][34] , \SHIFT_n[5][33] , \SHIFT_n[5][32] , 
        \SHIFT_n[5][31] , \SHIFT_n[5][30] , \SHIFT_n[5][29] , \SHIFT_n[5][28] , 
        \SHIFT_n[5][27] , \SHIFT_n[5][26] , \SHIFT_n[5][25] , \SHIFT_n[5][24] , 
        \SHIFT_n[5][23] , \SHIFT_n[5][22] , \SHIFT_n[5][21] , \SHIFT_n[5][20] , 
        \SHIFT_n[5][19] , \SHIFT_n[5][18] , \SHIFT_n[5][17] , \SHIFT_n[5][16] , 
        \SHIFT_n[5][15] , \SHIFT_n[5][14] , \SHIFT_n[5][13] , \SHIFT_n[5][12] , 
        \SHIFT_n[5][11] , \SHIFT_n[5][10] , \SHIFT_n[5][9] , \SHIFT_n[5][8] , 
        \SHIFT_n[5][7] , \SHIFT_n[5][6] , \SHIFT_n[5][5] , \SHIFT_n[5][4] , 
        \SHIFT_n[5][3] , \SHIFT_n[5][2] , SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21}) );
  BOOTHENC_NBIT44_i10 ENC_5 ( .A_s({\SHIFT[5][41] , \SHIFT[5][41] , 
        \SHIFT[5][41] , \SHIFT[5][40] , \SHIFT[5][39] , \SHIFT[5][38] , 
        \SHIFT[5][37] , \SHIFT[5][36] , \SHIFT[5][35] , \SHIFT[5][34] , 
        \SHIFT[5][33] , \SHIFT[5][32] , \SHIFT[5][31] , \SHIFT[5][30] , 
        \SHIFT[5][29] , \SHIFT[5][28] , \SHIFT[5][27] , \SHIFT[5][26] , 
        \SHIFT[5][25] , \SHIFT[5][24] , \SHIFT[5][23] , \SHIFT[5][22] , 
        \SHIFT[5][21] , \SHIFT[5][20] , \SHIFT[5][19] , \SHIFT[5][18] , 
        \SHIFT[5][17] , \SHIFT[5][16] , \SHIFT[5][15] , \SHIFT[5][14] , 
        \SHIFT[5][13] , \SHIFT[5][12] , \SHIFT[5][11] , \SHIFT[5][10] , 
        \SHIFT[5][9] , \SHIFT[5][8] , \SHIFT[5][7] , \SHIFT[5][6] , 
        \SHIFT[5][5] , \SHIFT[5][4] , \SHIFT[5][3] , \SHIFT[5][2] , 1'b0, 1'b0}), .A_ns({\SHIFT_n[5][41] , \SHIFT_n[5][41] , \SHIFT_n[5][41] , 
        \SHIFT_n[5][40] , \SHIFT_n[5][39] , \SHIFT_n[5][38] , \SHIFT_n[5][37] , 
        \SHIFT_n[5][36] , \SHIFT_n[5][35] , \SHIFT_n[5][34] , \SHIFT_n[5][33] , 
        \SHIFT_n[5][32] , \SHIFT_n[5][31] , \SHIFT_n[5][30] , \SHIFT_n[5][29] , 
        \SHIFT_n[5][28] , \SHIFT_n[5][27] , \SHIFT_n[5][26] , \SHIFT_n[5][25] , 
        \SHIFT_n[5][24] , \SHIFT_n[5][23] , \SHIFT_n[5][22] , \SHIFT_n[5][21] , 
        \SHIFT_n[5][20] , \SHIFT_n[5][19] , \SHIFT_n[5][18] , \SHIFT_n[5][17] , 
        \SHIFT_n[5][16] , \SHIFT_n[5][15] , \SHIFT_n[5][14] , \SHIFT_n[5][13] , 
        \SHIFT_n[5][12] , \SHIFT_n[5][11] , \SHIFT_n[5][10] , \SHIFT_n[5][9] , 
        \SHIFT_n[5][8] , \SHIFT_n[5][7] , \SHIFT_n[5][6] , \SHIFT_n[5][5] , 
        \SHIFT_n[5][4] , \SHIFT_n[5][3] , \SHIFT_n[5][2] , 1'b0, 1'b0}), .B({
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31:3], n10, B[1:0]}), .O({\OTMP[5][43] , \OTMP[5][42] , 
        \OTMP[5][41] , \OTMP[5][40] , \OTMP[5][39] , \OTMP[5][38] , 
        \OTMP[5][37] , \OTMP[5][36] , \OTMP[5][35] , \OTMP[5][34] , 
        \OTMP[5][33] , \OTMP[5][32] , \OTMP[5][31] , \OTMP[5][30] , 
        \OTMP[5][29] , \OTMP[5][28] , \OTMP[5][27] , \OTMP[5][26] , 
        \OTMP[5][25] , \OTMP[5][24] , \OTMP[5][23] , \OTMP[5][22] , 
        \OTMP[5][21] , \OTMP[5][20] , \OTMP[5][19] , \OTMP[5][18] , 
        \OTMP[5][17] , \OTMP[5][16] , \OTMP[5][15] , \OTMP[5][14] , 
        \OTMP[5][13] , \OTMP[5][12] , \OTMP[5][11] , \OTMP[5][10] , 
        \OTMP[5][9] , \OTMP[5][8] , \OTMP[5][7] , \OTMP[5][6] , \OTMP[5][5] , 
        \OTMP[5][4] , \OTMP[5][3] , \OTMP[5][2] , \OTMP[5][1] , 
        SYNOPSYS_UNCONNECTED__22}), .A_so({\SHIFT[6][43] , \SHIFT[6][42] , 
        \SHIFT[6][41] , \SHIFT[6][40] , \SHIFT[6][39] , \SHIFT[6][38] , 
        \SHIFT[6][37] , \SHIFT[6][36] , \SHIFT[6][35] , \SHIFT[6][34] , 
        \SHIFT[6][33] , \SHIFT[6][32] , \SHIFT[6][31] , \SHIFT[6][30] , 
        \SHIFT[6][29] , \SHIFT[6][28] , \SHIFT[6][27] , \SHIFT[6][26] , 
        \SHIFT[6][25] , \SHIFT[6][24] , \SHIFT[6][23] , \SHIFT[6][22] , 
        \SHIFT[6][21] , \SHIFT[6][20] , \SHIFT[6][19] , \SHIFT[6][18] , 
        \SHIFT[6][17] , \SHIFT[6][16] , \SHIFT[6][15] , \SHIFT[6][14] , 
        \SHIFT[6][13] , \SHIFT[6][12] , \SHIFT[6][11] , \SHIFT[6][10] , 
        \SHIFT[6][9] , \SHIFT[6][8] , \SHIFT[6][7] , \SHIFT[6][6] , 
        \SHIFT[6][5] , \SHIFT[6][4] , \SHIFT[6][3] , \SHIFT[6][2] , 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24}), .A_nso({
        \SHIFT_n[6][43] , \SHIFT_n[6][42] , \SHIFT_n[6][41] , \SHIFT_n[6][40] , 
        \SHIFT_n[6][39] , \SHIFT_n[6][38] , \SHIFT_n[6][37] , \SHIFT_n[6][36] , 
        \SHIFT_n[6][35] , \SHIFT_n[6][34] , \SHIFT_n[6][33] , \SHIFT_n[6][32] , 
        \SHIFT_n[6][31] , \SHIFT_n[6][30] , \SHIFT_n[6][29] , \SHIFT_n[6][28] , 
        \SHIFT_n[6][27] , \SHIFT_n[6][26] , \SHIFT_n[6][25] , \SHIFT_n[6][24] , 
        \SHIFT_n[6][23] , \SHIFT_n[6][22] , \SHIFT_n[6][21] , \SHIFT_n[6][20] , 
        \SHIFT_n[6][19] , \SHIFT_n[6][18] , \SHIFT_n[6][17] , \SHIFT_n[6][16] , 
        \SHIFT_n[6][15] , \SHIFT_n[6][14] , \SHIFT_n[6][13] , \SHIFT_n[6][12] , 
        \SHIFT_n[6][11] , \SHIFT_n[6][10] , \SHIFT_n[6][9] , \SHIFT_n[6][8] , 
        \SHIFT_n[6][7] , \SHIFT_n[6][6] , \SHIFT_n[6][5] , \SHIFT_n[6][4] , 
        \SHIFT_n[6][3] , \SHIFT_n[6][2] , SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26}) );
  BOOTHENC_NBIT46_i12 ENC_6 ( .A_s({\SHIFT[6][43] , \SHIFT[6][43] , 
        \SHIFT[6][43] , \SHIFT[6][42] , \SHIFT[6][41] , \SHIFT[6][40] , 
        \SHIFT[6][39] , \SHIFT[6][38] , \SHIFT[6][37] , \SHIFT[6][36] , 
        \SHIFT[6][35] , \SHIFT[6][34] , \SHIFT[6][33] , \SHIFT[6][32] , 
        \SHIFT[6][31] , \SHIFT[6][30] , \SHIFT[6][29] , \SHIFT[6][28] , 
        \SHIFT[6][27] , \SHIFT[6][26] , \SHIFT[6][25] , \SHIFT[6][24] , 
        \SHIFT[6][23] , \SHIFT[6][22] , \SHIFT[6][21] , \SHIFT[6][20] , 
        \SHIFT[6][19] , \SHIFT[6][18] , \SHIFT[6][17] , \SHIFT[6][16] , 
        \SHIFT[6][15] , \SHIFT[6][14] , \SHIFT[6][13] , \SHIFT[6][12] , 
        \SHIFT[6][11] , \SHIFT[6][10] , \SHIFT[6][9] , \SHIFT[6][8] , 
        \SHIFT[6][7] , \SHIFT[6][6] , \SHIFT[6][5] , \SHIFT[6][4] , 
        \SHIFT[6][3] , \SHIFT[6][2] , 1'b0, 1'b0}), .A_ns({\SHIFT_n[6][43] , 
        \SHIFT_n[6][43] , \SHIFT_n[6][43] , \SHIFT_n[6][42] , \SHIFT_n[6][41] , 
        \SHIFT_n[6][40] , \SHIFT_n[6][39] , \SHIFT_n[6][38] , \SHIFT_n[6][37] , 
        \SHIFT_n[6][36] , \SHIFT_n[6][35] , \SHIFT_n[6][34] , \SHIFT_n[6][33] , 
        \SHIFT_n[6][32] , \SHIFT_n[6][31] , \SHIFT_n[6][30] , \SHIFT_n[6][29] , 
        \SHIFT_n[6][28] , \SHIFT_n[6][27] , \SHIFT_n[6][26] , \SHIFT_n[6][25] , 
        \SHIFT_n[6][24] , \SHIFT_n[6][23] , \SHIFT_n[6][22] , \SHIFT_n[6][21] , 
        \SHIFT_n[6][20] , \SHIFT_n[6][19] , \SHIFT_n[6][18] , \SHIFT_n[6][17] , 
        \SHIFT_n[6][16] , \SHIFT_n[6][15] , \SHIFT_n[6][14] , \SHIFT_n[6][13] , 
        \SHIFT_n[6][12] , \SHIFT_n[6][11] , \SHIFT_n[6][10] , \SHIFT_n[6][9] , 
        \SHIFT_n[6][8] , \SHIFT_n[6][7] , \SHIFT_n[6][6] , \SHIFT_n[6][5] , 
        \SHIFT_n[6][4] , \SHIFT_n[6][3] , \SHIFT_n[6][2] , 1'b0, 1'b0}), .B({
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31:3], n9, B[1:0]}), .O({\OTMP[6][45] , 
        \OTMP[6][44] , \OTMP[6][43] , \OTMP[6][42] , \OTMP[6][41] , 
        \OTMP[6][40] , \OTMP[6][39] , \OTMP[6][38] , \OTMP[6][37] , 
        \OTMP[6][36] , \OTMP[6][35] , \OTMP[6][34] , \OTMP[6][33] , 
        \OTMP[6][32] , \OTMP[6][31] , \OTMP[6][30] , \OTMP[6][29] , 
        \OTMP[6][28] , \OTMP[6][27] , \OTMP[6][26] , \OTMP[6][25] , 
        \OTMP[6][24] , \OTMP[6][23] , \OTMP[6][22] , \OTMP[6][21] , 
        \OTMP[6][20] , \OTMP[6][19] , \OTMP[6][18] , \OTMP[6][17] , 
        \OTMP[6][16] , \OTMP[6][15] , \OTMP[6][14] , \OTMP[6][13] , 
        \OTMP[6][12] , \OTMP[6][11] , \OTMP[6][10] , \OTMP[6][9] , 
        \OTMP[6][8] , \OTMP[6][7] , \OTMP[6][6] , \OTMP[6][5] , \OTMP[6][4] , 
        \OTMP[6][3] , \OTMP[6][2] , \OTMP[6][1] , SYNOPSYS_UNCONNECTED__27}), 
        .A_so({\SHIFT[7][45] , \SHIFT[7][44] , \SHIFT[7][43] , \SHIFT[7][42] , 
        \SHIFT[7][41] , \SHIFT[7][40] , \SHIFT[7][39] , \SHIFT[7][38] , 
        \SHIFT[7][37] , \SHIFT[7][36] , \SHIFT[7][35] , \SHIFT[7][34] , 
        \SHIFT[7][33] , \SHIFT[7][32] , \SHIFT[7][31] , \SHIFT[7][30] , 
        \SHIFT[7][29] , \SHIFT[7][28] , \SHIFT[7][27] , \SHIFT[7][26] , 
        \SHIFT[7][25] , \SHIFT[7][24] , \SHIFT[7][23] , \SHIFT[7][22] , 
        \SHIFT[7][21] , \SHIFT[7][20] , \SHIFT[7][19] , \SHIFT[7][18] , 
        \SHIFT[7][17] , \SHIFT[7][16] , \SHIFT[7][15] , \SHIFT[7][14] , 
        \SHIFT[7][13] , \SHIFT[7][12] , \SHIFT[7][11] , \SHIFT[7][10] , 
        \SHIFT[7][9] , \SHIFT[7][8] , \SHIFT[7][7] , \SHIFT[7][6] , 
        \SHIFT[7][5] , \SHIFT[7][4] , \SHIFT[7][3] , \SHIFT[7][2] , 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29}), .A_nso({
        \SHIFT_n[7][45] , \SHIFT_n[7][44] , \SHIFT_n[7][43] , \SHIFT_n[7][42] , 
        \SHIFT_n[7][41] , \SHIFT_n[7][40] , \SHIFT_n[7][39] , \SHIFT_n[7][38] , 
        \SHIFT_n[7][37] , \SHIFT_n[7][36] , \SHIFT_n[7][35] , \SHIFT_n[7][34] , 
        \SHIFT_n[7][33] , \SHIFT_n[7][32] , \SHIFT_n[7][31] , \SHIFT_n[7][30] , 
        \SHIFT_n[7][29] , \SHIFT_n[7][28] , \SHIFT_n[7][27] , \SHIFT_n[7][26] , 
        \SHIFT_n[7][25] , \SHIFT_n[7][24] , \SHIFT_n[7][23] , \SHIFT_n[7][22] , 
        \SHIFT_n[7][21] , \SHIFT_n[7][20] , \SHIFT_n[7][19] , \SHIFT_n[7][18] , 
        \SHIFT_n[7][17] , \SHIFT_n[7][16] , \SHIFT_n[7][15] , \SHIFT_n[7][14] , 
        \SHIFT_n[7][13] , \SHIFT_n[7][12] , \SHIFT_n[7][11] , \SHIFT_n[7][10] , 
        \SHIFT_n[7][9] , \SHIFT_n[7][8] , \SHIFT_n[7][7] , \SHIFT_n[7][6] , 
        \SHIFT_n[7][5] , \SHIFT_n[7][4] , \SHIFT_n[7][3] , \SHIFT_n[7][2] , 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31}) );
  BOOTHENC_NBIT48_i14 ENC_7 ( .A_s({\SHIFT[7][45] , \SHIFT[7][45] , 
        \SHIFT[7][45] , \SHIFT[7][44] , \SHIFT[7][43] , \SHIFT[7][42] , 
        \SHIFT[7][41] , \SHIFT[7][40] , \SHIFT[7][39] , \SHIFT[7][38] , 
        \SHIFT[7][37] , \SHIFT[7][36] , \SHIFT[7][35] , \SHIFT[7][34] , 
        \SHIFT[7][33] , \SHIFT[7][32] , \SHIFT[7][31] , \SHIFT[7][30] , 
        \SHIFT[7][29] , \SHIFT[7][28] , \SHIFT[7][27] , \SHIFT[7][26] , 
        \SHIFT[7][25] , \SHIFT[7][24] , \SHIFT[7][23] , \SHIFT[7][22] , 
        \SHIFT[7][21] , \SHIFT[7][20] , \SHIFT[7][19] , \SHIFT[7][18] , 
        \SHIFT[7][17] , \SHIFT[7][16] , \SHIFT[7][15] , \SHIFT[7][14] , 
        \SHIFT[7][13] , \SHIFT[7][12] , \SHIFT[7][11] , \SHIFT[7][10] , 
        \SHIFT[7][9] , \SHIFT[7][8] , \SHIFT[7][7] , \SHIFT[7][6] , 
        \SHIFT[7][5] , \SHIFT[7][4] , \SHIFT[7][3] , \SHIFT[7][2] , 1'b0, 1'b0}), .A_ns({\SHIFT_n[7][45] , \SHIFT_n[7][45] , \SHIFT_n[7][45] , 
        \SHIFT_n[7][44] , \SHIFT_n[7][43] , \SHIFT_n[7][42] , \SHIFT_n[7][41] , 
        \SHIFT_n[7][40] , \SHIFT_n[7][39] , \SHIFT_n[7][38] , \SHIFT_n[7][37] , 
        \SHIFT_n[7][36] , \SHIFT_n[7][35] , \SHIFT_n[7][34] , \SHIFT_n[7][33] , 
        \SHIFT_n[7][32] , \SHIFT_n[7][31] , \SHIFT_n[7][30] , \SHIFT_n[7][29] , 
        \SHIFT_n[7][28] , \SHIFT_n[7][27] , \SHIFT_n[7][26] , \SHIFT_n[7][25] , 
        \SHIFT_n[7][24] , \SHIFT_n[7][23] , \SHIFT_n[7][22] , \SHIFT_n[7][21] , 
        \SHIFT_n[7][20] , \SHIFT_n[7][19] , \SHIFT_n[7][18] , \SHIFT_n[7][17] , 
        \SHIFT_n[7][16] , \SHIFT_n[7][15] , \SHIFT_n[7][14] , \SHIFT_n[7][13] , 
        \SHIFT_n[7][12] , \SHIFT_n[7][11] , \SHIFT_n[7][10] , \SHIFT_n[7][9] , 
        \SHIFT_n[7][8] , \SHIFT_n[7][7] , \SHIFT_n[7][6] , \SHIFT_n[7][5] , 
        \SHIFT_n[7][4] , \SHIFT_n[7][3] , \SHIFT_n[7][2] , 1'b0, 1'b0}), .B({
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B}), .O({\OTMP[7][47] , 
        \OTMP[7][46] , \OTMP[7][45] , \OTMP[7][44] , \OTMP[7][43] , 
        \OTMP[7][42] , \OTMP[7][41] , \OTMP[7][40] , \OTMP[7][39] , 
        \OTMP[7][38] , \OTMP[7][37] , \OTMP[7][36] , \OTMP[7][35] , 
        \OTMP[7][34] , \OTMP[7][33] , \OTMP[7][32] , \OTMP[7][31] , 
        \OTMP[7][30] , \OTMP[7][29] , \OTMP[7][28] , \OTMP[7][27] , 
        \OTMP[7][26] , \OTMP[7][25] , \OTMP[7][24] , \OTMP[7][23] , 
        \OTMP[7][22] , \OTMP[7][21] , \OTMP[7][20] , \OTMP[7][19] , 
        \OTMP[7][18] , \OTMP[7][17] , \OTMP[7][16] , \OTMP[7][15] , 
        \OTMP[7][14] , \OTMP[7][13] , \OTMP[7][12] , \OTMP[7][11] , 
        \OTMP[7][10] , \OTMP[7][9] , \OTMP[7][8] , \OTMP[7][7] , \OTMP[7][6] , 
        \OTMP[7][5] , \OTMP[7][4] , \OTMP[7][3] , \OTMP[7][2] , \OTMP[7][1] , 
        SYNOPSYS_UNCONNECTED__32}), .A_so({\SHIFT[8][47] , \SHIFT[8][46] , 
        \SHIFT[8][45] , \SHIFT[8][44] , \SHIFT[8][43] , \SHIFT[8][42] , 
        \SHIFT[8][41] , \SHIFT[8][40] , \SHIFT[8][39] , \SHIFT[8][38] , 
        \SHIFT[8][37] , \SHIFT[8][36] , \SHIFT[8][35] , \SHIFT[8][34] , 
        \SHIFT[8][33] , \SHIFT[8][32] , \SHIFT[8][31] , \SHIFT[8][30] , 
        \SHIFT[8][29] , \SHIFT[8][28] , \SHIFT[8][27] , \SHIFT[8][26] , 
        \SHIFT[8][25] , \SHIFT[8][24] , \SHIFT[8][23] , \SHIFT[8][22] , 
        \SHIFT[8][21] , \SHIFT[8][20] , \SHIFT[8][19] , \SHIFT[8][18] , 
        \SHIFT[8][17] , \SHIFT[8][16] , \SHIFT[8][15] , \SHIFT[8][14] , 
        \SHIFT[8][13] , \SHIFT[8][12] , \SHIFT[8][11] , \SHIFT[8][10] , 
        \SHIFT[8][9] , \SHIFT[8][8] , \SHIFT[8][7] , \SHIFT[8][6] , 
        \SHIFT[8][5] , \SHIFT[8][4] , \SHIFT[8][3] , \SHIFT[8][2] , 
        SYNOPSYS_UNCONNECTED__33, SYNOPSYS_UNCONNECTED__34}), .A_nso({
        \SHIFT_n[8][47] , \SHIFT_n[8][46] , \SHIFT_n[8][45] , \SHIFT_n[8][44] , 
        \SHIFT_n[8][43] , \SHIFT_n[8][42] , \SHIFT_n[8][41] , \SHIFT_n[8][40] , 
        \SHIFT_n[8][39] , \SHIFT_n[8][38] , \SHIFT_n[8][37] , \SHIFT_n[8][36] , 
        \SHIFT_n[8][35] , \SHIFT_n[8][34] , \SHIFT_n[8][33] , \SHIFT_n[8][32] , 
        \SHIFT_n[8][31] , \SHIFT_n[8][30] , \SHIFT_n[8][29] , \SHIFT_n[8][28] , 
        \SHIFT_n[8][27] , \SHIFT_n[8][26] , \SHIFT_n[8][25] , \SHIFT_n[8][24] , 
        \SHIFT_n[8][23] , \SHIFT_n[8][22] , \SHIFT_n[8][21] , \SHIFT_n[8][20] , 
        \SHIFT_n[8][19] , \SHIFT_n[8][18] , \SHIFT_n[8][17] , \SHIFT_n[8][16] , 
        \SHIFT_n[8][15] , \SHIFT_n[8][14] , \SHIFT_n[8][13] , \SHIFT_n[8][12] , 
        \SHIFT_n[8][11] , \SHIFT_n[8][10] , \SHIFT_n[8][9] , \SHIFT_n[8][8] , 
        \SHIFT_n[8][7] , \SHIFT_n[8][6] , \SHIFT_n[8][5] , \SHIFT_n[8][4] , 
        \SHIFT_n[8][3] , \SHIFT_n[8][2] , SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36}) );
  BOOTHENC_NBIT50_i16 ENC_8 ( .A_s({\SHIFT[8][47] , \SHIFT[8][47] , 
        \SHIFT[8][47] , \SHIFT[8][46] , \SHIFT[8][45] , \SHIFT[8][44] , 
        \SHIFT[8][43] , \SHIFT[8][42] , \SHIFT[8][41] , \SHIFT[8][40] , 
        \SHIFT[8][39] , \SHIFT[8][38] , \SHIFT[8][37] , \SHIFT[8][36] , 
        \SHIFT[8][35] , \SHIFT[8][34] , \SHIFT[8][33] , \SHIFT[8][32] , 
        \SHIFT[8][31] , \SHIFT[8][30] , \SHIFT[8][29] , \SHIFT[8][28] , 
        \SHIFT[8][27] , \SHIFT[8][26] , \SHIFT[8][25] , \SHIFT[8][24] , 
        \SHIFT[8][23] , \SHIFT[8][22] , \SHIFT[8][21] , \SHIFT[8][20] , 
        \SHIFT[8][19] , \SHIFT[8][18] , \SHIFT[8][17] , \SHIFT[8][16] , 
        \SHIFT[8][15] , \SHIFT[8][14] , \SHIFT[8][13] , \SHIFT[8][12] , 
        \SHIFT[8][11] , \SHIFT[8][10] , \SHIFT[8][9] , \SHIFT[8][8] , 
        \SHIFT[8][7] , \SHIFT[8][6] , \SHIFT[8][5] , \SHIFT[8][4] , 
        \SHIFT[8][3] , \SHIFT[8][2] , 1'b0, 1'b0}), .A_ns({\SHIFT_n[8][47] , 
        \SHIFT_n[8][47] , \SHIFT_n[8][47] , \SHIFT_n[8][46] , \SHIFT_n[8][45] , 
        \SHIFT_n[8][44] , \SHIFT_n[8][43] , \SHIFT_n[8][42] , \SHIFT_n[8][41] , 
        \SHIFT_n[8][40] , \SHIFT_n[8][39] , \SHIFT_n[8][38] , \SHIFT_n[8][37] , 
        \SHIFT_n[8][36] , \SHIFT_n[8][35] , \SHIFT_n[8][34] , \SHIFT_n[8][33] , 
        \SHIFT_n[8][32] , \SHIFT_n[8][31] , \SHIFT_n[8][30] , \SHIFT_n[8][29] , 
        \SHIFT_n[8][28] , \SHIFT_n[8][27] , \SHIFT_n[8][26] , \SHIFT_n[8][25] , 
        \SHIFT_n[8][24] , \SHIFT_n[8][23] , \SHIFT_n[8][22] , \SHIFT_n[8][21] , 
        \SHIFT_n[8][20] , \SHIFT_n[8][19] , \SHIFT_n[8][18] , \SHIFT_n[8][17] , 
        \SHIFT_n[8][16] , \SHIFT_n[8][15] , \SHIFT_n[8][14] , \SHIFT_n[8][13] , 
        \SHIFT_n[8][12] , \SHIFT_n[8][11] , \SHIFT_n[8][10] , \SHIFT_n[8][9] , 
        \SHIFT_n[8][8] , \SHIFT_n[8][7] , \SHIFT_n[8][6] , \SHIFT_n[8][5] , 
        \SHIFT_n[8][4] , \SHIFT_n[8][3] , \SHIFT_n[8][2] , 1'b0, 1'b0}), .B({
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B}), .O({
        \OTMP[8][49] , \OTMP[8][48] , \OTMP[8][47] , \OTMP[8][46] , 
        \OTMP[8][45] , \OTMP[8][44] , \OTMP[8][43] , \OTMP[8][42] , 
        \OTMP[8][41] , \OTMP[8][40] , \OTMP[8][39] , \OTMP[8][38] , 
        \OTMP[8][37] , \OTMP[8][36] , \OTMP[8][35] , \OTMP[8][34] , 
        \OTMP[8][33] , \OTMP[8][32] , \OTMP[8][31] , \OTMP[8][30] , 
        \OTMP[8][29] , \OTMP[8][28] , \OTMP[8][27] , \OTMP[8][26] , 
        \OTMP[8][25] , \OTMP[8][24] , \OTMP[8][23] , \OTMP[8][22] , 
        \OTMP[8][21] , \OTMP[8][20] , \OTMP[8][19] , \OTMP[8][18] , 
        \OTMP[8][17] , \OTMP[8][16] , \OTMP[8][15] , \OTMP[8][14] , 
        \OTMP[8][13] , \OTMP[8][12] , \OTMP[8][11] , \OTMP[8][10] , 
        \OTMP[8][9] , \OTMP[8][8] , \OTMP[8][7] , \OTMP[8][6] , \OTMP[8][5] , 
        \OTMP[8][4] , \OTMP[8][3] , \OTMP[8][2] , \OTMP[8][1] , 
        SYNOPSYS_UNCONNECTED__37}), .A_so({\SHIFT[9][49] , \SHIFT[9][48] , 
        \SHIFT[9][47] , \SHIFT[9][46] , \SHIFT[9][45] , \SHIFT[9][44] , 
        \SHIFT[9][43] , \SHIFT[9][42] , \SHIFT[9][41] , \SHIFT[9][40] , 
        \SHIFT[9][39] , \SHIFT[9][38] , \SHIFT[9][37] , \SHIFT[9][36] , 
        \SHIFT[9][35] , \SHIFT[9][34] , \SHIFT[9][33] , \SHIFT[9][32] , 
        \SHIFT[9][31] , \SHIFT[9][30] , \SHIFT[9][29] , \SHIFT[9][28] , 
        \SHIFT[9][27] , \SHIFT[9][26] , \SHIFT[9][25] , \SHIFT[9][24] , 
        \SHIFT[9][23] , \SHIFT[9][22] , \SHIFT[9][21] , \SHIFT[9][20] , 
        \SHIFT[9][19] , \SHIFT[9][18] , \SHIFT[9][17] , \SHIFT[9][16] , 
        \SHIFT[9][15] , \SHIFT[9][14] , \SHIFT[9][13] , \SHIFT[9][12] , 
        \SHIFT[9][11] , \SHIFT[9][10] , \SHIFT[9][9] , \SHIFT[9][8] , 
        \SHIFT[9][7] , \SHIFT[9][6] , \SHIFT[9][5] , \SHIFT[9][4] , 
        \SHIFT[9][3] , \SHIFT[9][2] , SYNOPSYS_UNCONNECTED__38, 
        SYNOPSYS_UNCONNECTED__39}), .A_nso({\SHIFT_n[9][49] , \SHIFT_n[9][48] , 
        \SHIFT_n[9][47] , \SHIFT_n[9][46] , \SHIFT_n[9][45] , \SHIFT_n[9][44] , 
        \SHIFT_n[9][43] , \SHIFT_n[9][42] , \SHIFT_n[9][41] , \SHIFT_n[9][40] , 
        \SHIFT_n[9][39] , \SHIFT_n[9][38] , \SHIFT_n[9][37] , \SHIFT_n[9][36] , 
        \SHIFT_n[9][35] , \SHIFT_n[9][34] , \SHIFT_n[9][33] , \SHIFT_n[9][32] , 
        \SHIFT_n[9][31] , \SHIFT_n[9][30] , \SHIFT_n[9][29] , \SHIFT_n[9][28] , 
        \SHIFT_n[9][27] , \SHIFT_n[9][26] , \SHIFT_n[9][25] , \SHIFT_n[9][24] , 
        \SHIFT_n[9][23] , \SHIFT_n[9][22] , \SHIFT_n[9][21] , \SHIFT_n[9][20] , 
        \SHIFT_n[9][19] , \SHIFT_n[9][18] , \SHIFT_n[9][17] , \SHIFT_n[9][16] , 
        \SHIFT_n[9][15] , \SHIFT_n[9][14] , \SHIFT_n[9][13] , \SHIFT_n[9][12] , 
        \SHIFT_n[9][11] , \SHIFT_n[9][10] , \SHIFT_n[9][9] , \SHIFT_n[9][8] , 
        \SHIFT_n[9][7] , \SHIFT_n[9][6] , \SHIFT_n[9][5] , \SHIFT_n[9][4] , 
        \SHIFT_n[9][3] , \SHIFT_n[9][2] , SYNOPSYS_UNCONNECTED__40, 
        SYNOPSYS_UNCONNECTED__41}) );
  BOOTHENC_NBIT52_i18 ENC_9 ( .A_s({\SHIFT[9][49] , \SHIFT[9][49] , 
        \SHIFT[9][49] , \SHIFT[9][48] , \SHIFT[9][47] , \SHIFT[9][46] , 
        \SHIFT[9][45] , \SHIFT[9][44] , \SHIFT[9][43] , \SHIFT[9][42] , 
        \SHIFT[9][41] , \SHIFT[9][40] , \SHIFT[9][39] , \SHIFT[9][38] , 
        \SHIFT[9][37] , \SHIFT[9][36] , \SHIFT[9][35] , \SHIFT[9][34] , 
        \SHIFT[9][33] , \SHIFT[9][32] , \SHIFT[9][31] , \SHIFT[9][30] , 
        \SHIFT[9][29] , \SHIFT[9][28] , \SHIFT[9][27] , \SHIFT[9][26] , 
        \SHIFT[9][25] , \SHIFT[9][24] , \SHIFT[9][23] , \SHIFT[9][22] , 
        \SHIFT[9][21] , \SHIFT[9][20] , \SHIFT[9][19] , \SHIFT[9][18] , 
        \SHIFT[9][17] , \SHIFT[9][16] , \SHIFT[9][15] , \SHIFT[9][14] , 
        \SHIFT[9][13] , \SHIFT[9][12] , \SHIFT[9][11] , \SHIFT[9][10] , 
        \SHIFT[9][9] , \SHIFT[9][8] , \SHIFT[9][7] , \SHIFT[9][6] , 
        \SHIFT[9][5] , \SHIFT[9][4] , \SHIFT[9][3] , \SHIFT[9][2] , 1'b0, 1'b0}), .A_ns({\SHIFT_n[9][49] , \SHIFT_n[9][49] , \SHIFT_n[9][49] , 
        \SHIFT_n[9][48] , \SHIFT_n[9][47] , \SHIFT_n[9][46] , \SHIFT_n[9][45] , 
        \SHIFT_n[9][44] , \SHIFT_n[9][43] , \SHIFT_n[9][42] , \SHIFT_n[9][41] , 
        \SHIFT_n[9][40] , \SHIFT_n[9][39] , \SHIFT_n[9][38] , \SHIFT_n[9][37] , 
        \SHIFT_n[9][36] , \SHIFT_n[9][35] , \SHIFT_n[9][34] , \SHIFT_n[9][33] , 
        \SHIFT_n[9][32] , \SHIFT_n[9][31] , \SHIFT_n[9][30] , \SHIFT_n[9][29] , 
        \SHIFT_n[9][28] , \SHIFT_n[9][27] , \SHIFT_n[9][26] , \SHIFT_n[9][25] , 
        \SHIFT_n[9][24] , \SHIFT_n[9][23] , \SHIFT_n[9][22] , \SHIFT_n[9][21] , 
        \SHIFT_n[9][20] , \SHIFT_n[9][19] , \SHIFT_n[9][18] , \SHIFT_n[9][17] , 
        \SHIFT_n[9][16] , \SHIFT_n[9][15] , \SHIFT_n[9][14] , \SHIFT_n[9][13] , 
        \SHIFT_n[9][12] , \SHIFT_n[9][11] , \SHIFT_n[9][10] , \SHIFT_n[9][9] , 
        \SHIFT_n[9][8] , \SHIFT_n[9][7] , \SHIFT_n[9][6] , \SHIFT_n[9][5] , 
        \SHIFT_n[9][4] , \SHIFT_n[9][3] , \SHIFT_n[9][2] , 1'b0, 1'b0}), .B({
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B}), .O({\OTMP[9][51] , \OTMP[9][50] , \OTMP[9][49] , \OTMP[9][48] , 
        \OTMP[9][47] , \OTMP[9][46] , \OTMP[9][45] , \OTMP[9][44] , 
        \OTMP[9][43] , \OTMP[9][42] , \OTMP[9][41] , \OTMP[9][40] , 
        \OTMP[9][39] , \OTMP[9][38] , \OTMP[9][37] , \OTMP[9][36] , 
        \OTMP[9][35] , \OTMP[9][34] , \OTMP[9][33] , \OTMP[9][32] , 
        \OTMP[9][31] , \OTMP[9][30] , \OTMP[9][29] , \OTMP[9][28] , 
        \OTMP[9][27] , \OTMP[9][26] , \OTMP[9][25] , \OTMP[9][24] , 
        \OTMP[9][23] , \OTMP[9][22] , \OTMP[9][21] , \OTMP[9][20] , 
        \OTMP[9][19] , \OTMP[9][18] , \OTMP[9][17] , \OTMP[9][16] , 
        \OTMP[9][15] , \OTMP[9][14] , \OTMP[9][13] , \OTMP[9][12] , 
        \OTMP[9][11] , \OTMP[9][10] , \OTMP[9][9] , \OTMP[9][8] , \OTMP[9][7] , 
        \OTMP[9][6] , \OTMP[9][5] , \OTMP[9][4] , \OTMP[9][3] , \OTMP[9][2] , 
        \OTMP[9][1] , SYNOPSYS_UNCONNECTED__42}), .A_so({\SHIFT[10][51] , 
        \SHIFT[10][50] , \SHIFT[10][49] , \SHIFT[10][48] , \SHIFT[10][47] , 
        \SHIFT[10][46] , \SHIFT[10][45] , \SHIFT[10][44] , \SHIFT[10][43] , 
        \SHIFT[10][42] , \SHIFT[10][41] , \SHIFT[10][40] , \SHIFT[10][39] , 
        \SHIFT[10][38] , \SHIFT[10][37] , \SHIFT[10][36] , \SHIFT[10][35] , 
        \SHIFT[10][34] , \SHIFT[10][33] , \SHIFT[10][32] , \SHIFT[10][31] , 
        \SHIFT[10][30] , \SHIFT[10][29] , \SHIFT[10][28] , \SHIFT[10][27] , 
        \SHIFT[10][26] , \SHIFT[10][25] , \SHIFT[10][24] , \SHIFT[10][23] , 
        \SHIFT[10][22] , \SHIFT[10][21] , \SHIFT[10][20] , \SHIFT[10][19] , 
        \SHIFT[10][18] , \SHIFT[10][17] , \SHIFT[10][16] , \SHIFT[10][15] , 
        \SHIFT[10][14] , \SHIFT[10][13] , \SHIFT[10][12] , \SHIFT[10][11] , 
        \SHIFT[10][10] , \SHIFT[10][9] , \SHIFT[10][8] , \SHIFT[10][7] , 
        \SHIFT[10][6] , \SHIFT[10][5] , \SHIFT[10][4] , \SHIFT[10][3] , 
        \SHIFT[10][2] , SYNOPSYS_UNCONNECTED__43, SYNOPSYS_UNCONNECTED__44}), 
        .A_nso({\SHIFT_n[10][51] , \SHIFT_n[10][50] , \SHIFT_n[10][49] , 
        \SHIFT_n[10][48] , \SHIFT_n[10][47] , \SHIFT_n[10][46] , 
        \SHIFT_n[10][45] , \SHIFT_n[10][44] , \SHIFT_n[10][43] , 
        \SHIFT_n[10][42] , \SHIFT_n[10][41] , \SHIFT_n[10][40] , 
        \SHIFT_n[10][39] , \SHIFT_n[10][38] , \SHIFT_n[10][37] , 
        \SHIFT_n[10][36] , \SHIFT_n[10][35] , \SHIFT_n[10][34] , 
        \SHIFT_n[10][33] , \SHIFT_n[10][32] , \SHIFT_n[10][31] , 
        \SHIFT_n[10][30] , \SHIFT_n[10][29] , \SHIFT_n[10][28] , 
        \SHIFT_n[10][27] , \SHIFT_n[10][26] , \SHIFT_n[10][25] , 
        \SHIFT_n[10][24] , \SHIFT_n[10][23] , \SHIFT_n[10][22] , 
        \SHIFT_n[10][21] , \SHIFT_n[10][20] , \SHIFT_n[10][19] , 
        \SHIFT_n[10][18] , \SHIFT_n[10][17] , \SHIFT_n[10][16] , 
        \SHIFT_n[10][15] , \SHIFT_n[10][14] , \SHIFT_n[10][13] , 
        \SHIFT_n[10][12] , \SHIFT_n[10][11] , \SHIFT_n[10][10] , 
        \SHIFT_n[10][9] , \SHIFT_n[10][8] , \SHIFT_n[10][7] , \SHIFT_n[10][6] , 
        \SHIFT_n[10][5] , \SHIFT_n[10][4] , \SHIFT_n[10][3] , \SHIFT_n[10][2] , 
        SYNOPSYS_UNCONNECTED__45, SYNOPSYS_UNCONNECTED__46}) );
  BOOTHENC_NBIT54_i20 ENC_10 ( .A_s({\SHIFT[10][51] , \SHIFT[10][51] , 
        \SHIFT[10][51] , \SHIFT[10][50] , \SHIFT[10][49] , \SHIFT[10][48] , 
        \SHIFT[10][47] , \SHIFT[10][46] , \SHIFT[10][45] , \SHIFT[10][44] , 
        \SHIFT[10][43] , \SHIFT[10][42] , \SHIFT[10][41] , \SHIFT[10][40] , 
        \SHIFT[10][39] , \SHIFT[10][38] , \SHIFT[10][37] , \SHIFT[10][36] , 
        \SHIFT[10][35] , \SHIFT[10][34] , \SHIFT[10][33] , \SHIFT[10][32] , 
        \SHIFT[10][31] , \SHIFT[10][30] , \SHIFT[10][29] , \SHIFT[10][28] , 
        \SHIFT[10][27] , \SHIFT[10][26] , \SHIFT[10][25] , \SHIFT[10][24] , 
        \SHIFT[10][23] , \SHIFT[10][22] , \SHIFT[10][21] , \SHIFT[10][20] , 
        \SHIFT[10][19] , \SHIFT[10][18] , \SHIFT[10][17] , \SHIFT[10][16] , 
        \SHIFT[10][15] , \SHIFT[10][14] , \SHIFT[10][13] , \SHIFT[10][12] , 
        \SHIFT[10][11] , \SHIFT[10][10] , \SHIFT[10][9] , \SHIFT[10][8] , 
        \SHIFT[10][7] , \SHIFT[10][6] , \SHIFT[10][5] , \SHIFT[10][4] , 
        \SHIFT[10][3] , \SHIFT[10][2] , 1'b0, 1'b0}), .A_ns({\SHIFT_n[10][51] , 
        \SHIFT_n[10][51] , \SHIFT_n[10][51] , \SHIFT_n[10][50] , 
        \SHIFT_n[10][49] , \SHIFT_n[10][48] , \SHIFT_n[10][47] , 
        \SHIFT_n[10][46] , \SHIFT_n[10][45] , \SHIFT_n[10][44] , 
        \SHIFT_n[10][43] , \SHIFT_n[10][42] , \SHIFT_n[10][41] , 
        \SHIFT_n[10][40] , \SHIFT_n[10][39] , \SHIFT_n[10][38] , 
        \SHIFT_n[10][37] , \SHIFT_n[10][36] , \SHIFT_n[10][35] , 
        \SHIFT_n[10][34] , \SHIFT_n[10][33] , \SHIFT_n[10][32] , 
        \SHIFT_n[10][31] , \SHIFT_n[10][30] , \SHIFT_n[10][29] , 
        \SHIFT_n[10][28] , \SHIFT_n[10][27] , \SHIFT_n[10][26] , 
        \SHIFT_n[10][25] , \SHIFT_n[10][24] , \SHIFT_n[10][23] , 
        \SHIFT_n[10][22] , \SHIFT_n[10][21] , \SHIFT_n[10][20] , 
        \SHIFT_n[10][19] , \SHIFT_n[10][18] , \SHIFT_n[10][17] , 
        \SHIFT_n[10][16] , \SHIFT_n[10][15] , \SHIFT_n[10][14] , 
        \SHIFT_n[10][13] , \SHIFT_n[10][12] , \SHIFT_n[10][11] , 
        \SHIFT_n[10][10] , \SHIFT_n[10][9] , \SHIFT_n[10][8] , 
        \SHIFT_n[10][7] , \SHIFT_n[10][6] , \SHIFT_n[10][5] , \SHIFT_n[10][4] , 
        \SHIFT_n[10][3] , \SHIFT_n[10][2] , 1'b0, 1'b0}), .B({B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B}), .O({\OTMP[10][53] , \OTMP[10][52] , \OTMP[10][51] , 
        \OTMP[10][50] , \OTMP[10][49] , \OTMP[10][48] , \OTMP[10][47] , 
        \OTMP[10][46] , \OTMP[10][45] , \OTMP[10][44] , \OTMP[10][43] , 
        \OTMP[10][42] , \OTMP[10][41] , \OTMP[10][40] , \OTMP[10][39] , 
        \OTMP[10][38] , \OTMP[10][37] , \OTMP[10][36] , \OTMP[10][35] , 
        \OTMP[10][34] , \OTMP[10][33] , \OTMP[10][32] , \OTMP[10][31] , 
        \OTMP[10][30] , \OTMP[10][29] , \OTMP[10][28] , \OTMP[10][27] , 
        \OTMP[10][26] , \OTMP[10][25] , \OTMP[10][24] , \OTMP[10][23] , 
        \OTMP[10][22] , \OTMP[10][21] , \OTMP[10][20] , \OTMP[10][19] , 
        \OTMP[10][18] , \OTMP[10][17] , \OTMP[10][16] , \OTMP[10][15] , 
        \OTMP[10][14] , \OTMP[10][13] , \OTMP[10][12] , \OTMP[10][11] , 
        \OTMP[10][10] , \OTMP[10][9] , \OTMP[10][8] , \OTMP[10][7] , 
        \OTMP[10][6] , \OTMP[10][5] , \OTMP[10][4] , \OTMP[10][3] , 
        \OTMP[10][2] , \OTMP[10][1] , SYNOPSYS_UNCONNECTED__47}), .A_so({
        \SHIFT[11][53] , \SHIFT[11][52] , \SHIFT[11][51] , \SHIFT[11][50] , 
        \SHIFT[11][49] , \SHIFT[11][48] , \SHIFT[11][47] , \SHIFT[11][46] , 
        \SHIFT[11][45] , \SHIFT[11][44] , \SHIFT[11][43] , \SHIFT[11][42] , 
        \SHIFT[11][41] , \SHIFT[11][40] , \SHIFT[11][39] , \SHIFT[11][38] , 
        \SHIFT[11][37] , \SHIFT[11][36] , \SHIFT[11][35] , \SHIFT[11][34] , 
        \SHIFT[11][33] , \SHIFT[11][32] , \SHIFT[11][31] , \SHIFT[11][30] , 
        \SHIFT[11][29] , \SHIFT[11][28] , \SHIFT[11][27] , \SHIFT[11][26] , 
        \SHIFT[11][25] , \SHIFT[11][24] , \SHIFT[11][23] , \SHIFT[11][22] , 
        \SHIFT[11][21] , \SHIFT[11][20] , \SHIFT[11][19] , \SHIFT[11][18] , 
        \SHIFT[11][17] , \SHIFT[11][16] , \SHIFT[11][15] , \SHIFT[11][14] , 
        \SHIFT[11][13] , \SHIFT[11][12] , \SHIFT[11][11] , \SHIFT[11][10] , 
        \SHIFT[11][9] , \SHIFT[11][8] , \SHIFT[11][7] , \SHIFT[11][6] , 
        \SHIFT[11][5] , \SHIFT[11][4] , \SHIFT[11][3] , \SHIFT[11][2] , 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49}), .A_nso({
        \SHIFT_n[11][53] , \SHIFT_n[11][52] , \SHIFT_n[11][51] , 
        \SHIFT_n[11][50] , \SHIFT_n[11][49] , \SHIFT_n[11][48] , 
        \SHIFT_n[11][47] , \SHIFT_n[11][46] , \SHIFT_n[11][45] , 
        \SHIFT_n[11][44] , \SHIFT_n[11][43] , \SHIFT_n[11][42] , 
        \SHIFT_n[11][41] , \SHIFT_n[11][40] , \SHIFT_n[11][39] , 
        \SHIFT_n[11][38] , \SHIFT_n[11][37] , \SHIFT_n[11][36] , 
        \SHIFT_n[11][35] , \SHIFT_n[11][34] , \SHIFT_n[11][33] , 
        \SHIFT_n[11][32] , \SHIFT_n[11][31] , \SHIFT_n[11][30] , 
        \SHIFT_n[11][29] , \SHIFT_n[11][28] , \SHIFT_n[11][27] , 
        \SHIFT_n[11][26] , \SHIFT_n[11][25] , \SHIFT_n[11][24] , 
        \SHIFT_n[11][23] , \SHIFT_n[11][22] , \SHIFT_n[11][21] , 
        \SHIFT_n[11][20] , \SHIFT_n[11][19] , \SHIFT_n[11][18] , 
        \SHIFT_n[11][17] , \SHIFT_n[11][16] , \SHIFT_n[11][15] , 
        \SHIFT_n[11][14] , \SHIFT_n[11][13] , \SHIFT_n[11][12] , 
        \SHIFT_n[11][11] , \SHIFT_n[11][10] , \SHIFT_n[11][9] , 
        \SHIFT_n[11][8] , \SHIFT_n[11][7] , \SHIFT_n[11][6] , \SHIFT_n[11][5] , 
        \SHIFT_n[11][4] , \SHIFT_n[11][3] , \SHIFT_n[11][2] , 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51}) );
  BOOTHENC_NBIT56_i22 ENC_11 ( .A_s({\SHIFT[11][53] , \SHIFT[11][53] , 
        \SHIFT[11][53] , \SHIFT[11][52] , \SHIFT[11][51] , \SHIFT[11][50] , 
        \SHIFT[11][49] , \SHIFT[11][48] , \SHIFT[11][47] , \SHIFT[11][46] , 
        \SHIFT[11][45] , \SHIFT[11][44] , \SHIFT[11][43] , \SHIFT[11][42] , 
        \SHIFT[11][41] , \SHIFT[11][40] , \SHIFT[11][39] , \SHIFT[11][38] , 
        \SHIFT[11][37] , \SHIFT[11][36] , \SHIFT[11][35] , \SHIFT[11][34] , 
        \SHIFT[11][33] , \SHIFT[11][32] , \SHIFT[11][31] , \SHIFT[11][30] , 
        \SHIFT[11][29] , \SHIFT[11][28] , \SHIFT[11][27] , \SHIFT[11][26] , 
        \SHIFT[11][25] , \SHIFT[11][24] , \SHIFT[11][23] , \SHIFT[11][22] , 
        \SHIFT[11][21] , \SHIFT[11][20] , \SHIFT[11][19] , \SHIFT[11][18] , 
        \SHIFT[11][17] , \SHIFT[11][16] , \SHIFT[11][15] , \SHIFT[11][14] , 
        \SHIFT[11][13] , \SHIFT[11][12] , \SHIFT[11][11] , \SHIFT[11][10] , 
        \SHIFT[11][9] , \SHIFT[11][8] , \SHIFT[11][7] , \SHIFT[11][6] , 
        \SHIFT[11][5] , \SHIFT[11][4] , \SHIFT[11][3] , \SHIFT[11][2] , 1'b0, 
        1'b0}), .A_ns({\SHIFT_n[11][53] , \SHIFT_n[11][53] , \SHIFT_n[11][53] , 
        \SHIFT_n[11][52] , \SHIFT_n[11][51] , \SHIFT_n[11][50] , 
        \SHIFT_n[11][49] , \SHIFT_n[11][48] , \SHIFT_n[11][47] , 
        \SHIFT_n[11][46] , \SHIFT_n[11][45] , \SHIFT_n[11][44] , 
        \SHIFT_n[11][43] , \SHIFT_n[11][42] , \SHIFT_n[11][41] , 
        \SHIFT_n[11][40] , \SHIFT_n[11][39] , \SHIFT_n[11][38] , 
        \SHIFT_n[11][37] , \SHIFT_n[11][36] , \SHIFT_n[11][35] , 
        \SHIFT_n[11][34] , \SHIFT_n[11][33] , \SHIFT_n[11][32] , 
        \SHIFT_n[11][31] , \SHIFT_n[11][30] , \SHIFT_n[11][29] , 
        \SHIFT_n[11][28] , \SHIFT_n[11][27] , \SHIFT_n[11][26] , 
        \SHIFT_n[11][25] , \SHIFT_n[11][24] , \SHIFT_n[11][23] , 
        \SHIFT_n[11][22] , \SHIFT_n[11][21] , \SHIFT_n[11][20] , 
        \SHIFT_n[11][19] , \SHIFT_n[11][18] , \SHIFT_n[11][17] , 
        \SHIFT_n[11][16] , \SHIFT_n[11][15] , \SHIFT_n[11][14] , 
        \SHIFT_n[11][13] , \SHIFT_n[11][12] , \SHIFT_n[11][11] , 
        \SHIFT_n[11][10] , \SHIFT_n[11][9] , \SHIFT_n[11][8] , 
        \SHIFT_n[11][7] , \SHIFT_n[11][6] , \SHIFT_n[11][5] , \SHIFT_n[11][4] , 
        \SHIFT_n[11][3] , \SHIFT_n[11][2] , 1'b0, 1'b0}), .B({B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B}), .O({\OTMP[11][55] , \OTMP[11][54] , \OTMP[11][53] , 
        \OTMP[11][52] , \OTMP[11][51] , \OTMP[11][50] , \OTMP[11][49] , 
        \OTMP[11][48] , \OTMP[11][47] , \OTMP[11][46] , \OTMP[11][45] , 
        \OTMP[11][44] , \OTMP[11][43] , \OTMP[11][42] , \OTMP[11][41] , 
        \OTMP[11][40] , \OTMP[11][39] , \OTMP[11][38] , \OTMP[11][37] , 
        \OTMP[11][36] , \OTMP[11][35] , \OTMP[11][34] , \OTMP[11][33] , 
        \OTMP[11][32] , \OTMP[11][31] , \OTMP[11][30] , \OTMP[11][29] , 
        \OTMP[11][28] , \OTMP[11][27] , \OTMP[11][26] , \OTMP[11][25] , 
        \OTMP[11][24] , \OTMP[11][23] , \OTMP[11][22] , \OTMP[11][21] , 
        \OTMP[11][20] , \OTMP[11][19] , \OTMP[11][18] , \OTMP[11][17] , 
        \OTMP[11][16] , \OTMP[11][15] , \OTMP[11][14] , \OTMP[11][13] , 
        \OTMP[11][12] , \OTMP[11][11] , \OTMP[11][10] , \OTMP[11][9] , 
        \OTMP[11][8] , \OTMP[11][7] , \OTMP[11][6] , \OTMP[11][5] , 
        \OTMP[11][4] , \OTMP[11][3] , \OTMP[11][2] , \OTMP[11][1] , 
        SYNOPSYS_UNCONNECTED__52}), .A_so({\SHIFT[12][55] , \SHIFT[12][54] , 
        \SHIFT[12][53] , \SHIFT[12][52] , \SHIFT[12][51] , \SHIFT[12][50] , 
        \SHIFT[12][49] , \SHIFT[12][48] , \SHIFT[12][47] , \SHIFT[12][46] , 
        \SHIFT[12][45] , \SHIFT[12][44] , \SHIFT[12][43] , \SHIFT[12][42] , 
        \SHIFT[12][41] , \SHIFT[12][40] , \SHIFT[12][39] , \SHIFT[12][38] , 
        \SHIFT[12][37] , \SHIFT[12][36] , \SHIFT[12][35] , \SHIFT[12][34] , 
        \SHIFT[12][33] , \SHIFT[12][32] , \SHIFT[12][31] , \SHIFT[12][30] , 
        \SHIFT[12][29] , \SHIFT[12][28] , \SHIFT[12][27] , \SHIFT[12][26] , 
        \SHIFT[12][25] , \SHIFT[12][24] , \SHIFT[12][23] , \SHIFT[12][22] , 
        \SHIFT[12][21] , \SHIFT[12][20] , \SHIFT[12][19] , \SHIFT[12][18] , 
        \SHIFT[12][17] , \SHIFT[12][16] , \SHIFT[12][15] , \SHIFT[12][14] , 
        \SHIFT[12][13] , \SHIFT[12][12] , \SHIFT[12][11] , \SHIFT[12][10] , 
        \SHIFT[12][9] , \SHIFT[12][8] , \SHIFT[12][7] , \SHIFT[12][6] , 
        \SHIFT[12][5] , \SHIFT[12][4] , \SHIFT[12][3] , \SHIFT[12][2] , 
        SYNOPSYS_UNCONNECTED__53, SYNOPSYS_UNCONNECTED__54}), .A_nso({
        \SHIFT_n[12][55] , \SHIFT_n[12][54] , \SHIFT_n[12][53] , 
        \SHIFT_n[12][52] , \SHIFT_n[12][51] , \SHIFT_n[12][50] , 
        \SHIFT_n[12][49] , \SHIFT_n[12][48] , \SHIFT_n[12][47] , 
        \SHIFT_n[12][46] , \SHIFT_n[12][45] , \SHIFT_n[12][44] , 
        \SHIFT_n[12][43] , \SHIFT_n[12][42] , \SHIFT_n[12][41] , 
        \SHIFT_n[12][40] , \SHIFT_n[12][39] , \SHIFT_n[12][38] , 
        \SHIFT_n[12][37] , \SHIFT_n[12][36] , \SHIFT_n[12][35] , 
        \SHIFT_n[12][34] , \SHIFT_n[12][33] , \SHIFT_n[12][32] , 
        \SHIFT_n[12][31] , \SHIFT_n[12][30] , \SHIFT_n[12][29] , 
        \SHIFT_n[12][28] , \SHIFT_n[12][27] , \SHIFT_n[12][26] , 
        \SHIFT_n[12][25] , \SHIFT_n[12][24] , \SHIFT_n[12][23] , 
        \SHIFT_n[12][22] , \SHIFT_n[12][21] , \SHIFT_n[12][20] , 
        \SHIFT_n[12][19] , \SHIFT_n[12][18] , \SHIFT_n[12][17] , 
        \SHIFT_n[12][16] , \SHIFT_n[12][15] , \SHIFT_n[12][14] , 
        \SHIFT_n[12][13] , \SHIFT_n[12][12] , \SHIFT_n[12][11] , 
        \SHIFT_n[12][10] , \SHIFT_n[12][9] , \SHIFT_n[12][8] , 
        \SHIFT_n[12][7] , \SHIFT_n[12][6] , \SHIFT_n[12][5] , \SHIFT_n[12][4] , 
        \SHIFT_n[12][3] , \SHIFT_n[12][2] , SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56}) );
  BOOTHENC_NBIT58_i24 ENC_12 ( .A_s({\SHIFT[12][55] , \SHIFT[12][55] , 
        \SHIFT[12][55] , \SHIFT[12][54] , \SHIFT[12][53] , \SHIFT[12][52] , 
        \SHIFT[12][51] , \SHIFT[12][50] , \SHIFT[12][49] , \SHIFT[12][48] , 
        \SHIFT[12][47] , \SHIFT[12][46] , \SHIFT[12][45] , \SHIFT[12][44] , 
        \SHIFT[12][43] , \SHIFT[12][42] , \SHIFT[12][41] , \SHIFT[12][40] , 
        \SHIFT[12][39] , \SHIFT[12][38] , \SHIFT[12][37] , \SHIFT[12][36] , 
        \SHIFT[12][35] , \SHIFT[12][34] , \SHIFT[12][33] , \SHIFT[12][32] , 
        \SHIFT[12][31] , \SHIFT[12][30] , \SHIFT[12][29] , \SHIFT[12][28] , 
        \SHIFT[12][27] , \SHIFT[12][26] , \SHIFT[12][25] , \SHIFT[12][24] , 
        \SHIFT[12][23] , \SHIFT[12][22] , \SHIFT[12][21] , \SHIFT[12][20] , 
        \SHIFT[12][19] , \SHIFT[12][18] , \SHIFT[12][17] , \SHIFT[12][16] , 
        \SHIFT[12][15] , \SHIFT[12][14] , \SHIFT[12][13] , \SHIFT[12][12] , 
        \SHIFT[12][11] , \SHIFT[12][10] , \SHIFT[12][9] , \SHIFT[12][8] , 
        \SHIFT[12][7] , \SHIFT[12][6] , \SHIFT[12][5] , \SHIFT[12][4] , 
        \SHIFT[12][3] , \SHIFT[12][2] , 1'b0, 1'b0}), .A_ns({\SHIFT_n[12][55] , 
        \SHIFT_n[12][55] , \SHIFT_n[12][55] , \SHIFT_n[12][54] , 
        \SHIFT_n[12][53] , \SHIFT_n[12][52] , \SHIFT_n[12][51] , 
        \SHIFT_n[12][50] , \SHIFT_n[12][49] , \SHIFT_n[12][48] , 
        \SHIFT_n[12][47] , \SHIFT_n[12][46] , \SHIFT_n[12][45] , 
        \SHIFT_n[12][44] , \SHIFT_n[12][43] , \SHIFT_n[12][42] , 
        \SHIFT_n[12][41] , \SHIFT_n[12][40] , \SHIFT_n[12][39] , 
        \SHIFT_n[12][38] , \SHIFT_n[12][37] , \SHIFT_n[12][36] , 
        \SHIFT_n[12][35] , \SHIFT_n[12][34] , \SHIFT_n[12][33] , 
        \SHIFT_n[12][32] , \SHIFT_n[12][31] , \SHIFT_n[12][30] , 
        \SHIFT_n[12][29] , \SHIFT_n[12][28] , \SHIFT_n[12][27] , 
        \SHIFT_n[12][26] , \SHIFT_n[12][25] , \SHIFT_n[12][24] , 
        \SHIFT_n[12][23] , \SHIFT_n[12][22] , \SHIFT_n[12][21] , 
        \SHIFT_n[12][20] , \SHIFT_n[12][19] , \SHIFT_n[12][18] , 
        \SHIFT_n[12][17] , \SHIFT_n[12][16] , \SHIFT_n[12][15] , 
        \SHIFT_n[12][14] , \SHIFT_n[12][13] , \SHIFT_n[12][12] , 
        \SHIFT_n[12][11] , \SHIFT_n[12][10] , \SHIFT_n[12][9] , 
        \SHIFT_n[12][8] , \SHIFT_n[12][7] , \SHIFT_n[12][6] , \SHIFT_n[12][5] , 
        \SHIFT_n[12][4] , \SHIFT_n[12][3] , \SHIFT_n[12][2] , 1'b0, 1'b0}), 
        .B({B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B}), .O({
        \OTMP[12][57] , \OTMP[12][56] , \OTMP[12][55] , \OTMP[12][54] , 
        \OTMP[12][53] , \OTMP[12][52] , \OTMP[12][51] , \OTMP[12][50] , 
        \OTMP[12][49] , \OTMP[12][48] , \OTMP[12][47] , \OTMP[12][46] , 
        \OTMP[12][45] , \OTMP[12][44] , \OTMP[12][43] , \OTMP[12][42] , 
        \OTMP[12][41] , \OTMP[12][40] , \OTMP[12][39] , \OTMP[12][38] , 
        \OTMP[12][37] , \OTMP[12][36] , \OTMP[12][35] , \OTMP[12][34] , 
        \OTMP[12][33] , \OTMP[12][32] , \OTMP[12][31] , \OTMP[12][30] , 
        \OTMP[12][29] , \OTMP[12][28] , \OTMP[12][27] , \OTMP[12][26] , 
        \OTMP[12][25] , \OTMP[12][24] , \OTMP[12][23] , \OTMP[12][22] , 
        \OTMP[12][21] , \OTMP[12][20] , \OTMP[12][19] , \OTMP[12][18] , 
        \OTMP[12][17] , \OTMP[12][16] , \OTMP[12][15] , \OTMP[12][14] , 
        \OTMP[12][13] , \OTMP[12][12] , \OTMP[12][11] , \OTMP[12][10] , 
        \OTMP[12][9] , \OTMP[12][8] , \OTMP[12][7] , \OTMP[12][6] , 
        \OTMP[12][5] , \OTMP[12][4] , \OTMP[12][3] , \OTMP[12][2] , 
        \OTMP[12][1] , SYNOPSYS_UNCONNECTED__57}), .A_so({\SHIFT[13][57] , 
        \SHIFT[13][56] , \SHIFT[13][55] , \SHIFT[13][54] , \SHIFT[13][53] , 
        \SHIFT[13][52] , \SHIFT[13][51] , \SHIFT[13][50] , \SHIFT[13][49] , 
        \SHIFT[13][48] , \SHIFT[13][47] , \SHIFT[13][46] , \SHIFT[13][45] , 
        \SHIFT[13][44] , \SHIFT[13][43] , \SHIFT[13][42] , \SHIFT[13][41] , 
        \SHIFT[13][40] , \SHIFT[13][39] , \SHIFT[13][38] , \SHIFT[13][37] , 
        \SHIFT[13][36] , \SHIFT[13][35] , \SHIFT[13][34] , \SHIFT[13][33] , 
        \SHIFT[13][32] , \SHIFT[13][31] , \SHIFT[13][30] , \SHIFT[13][29] , 
        \SHIFT[13][28] , \SHIFT[13][27] , \SHIFT[13][26] , \SHIFT[13][25] , 
        \SHIFT[13][24] , \SHIFT[13][23] , \SHIFT[13][22] , \SHIFT[13][21] , 
        \SHIFT[13][20] , \SHIFT[13][19] , \SHIFT[13][18] , \SHIFT[13][17] , 
        \SHIFT[13][16] , \SHIFT[13][15] , \SHIFT[13][14] , \SHIFT[13][13] , 
        \SHIFT[13][12] , \SHIFT[13][11] , \SHIFT[13][10] , \SHIFT[13][9] , 
        \SHIFT[13][8] , \SHIFT[13][7] , \SHIFT[13][6] , \SHIFT[13][5] , 
        \SHIFT[13][4] , \SHIFT[13][3] , \SHIFT[13][2] , 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59}), .A_nso({
        \SHIFT_n[13][57] , \SHIFT_n[13][56] , \SHIFT_n[13][55] , 
        \SHIFT_n[13][54] , \SHIFT_n[13][53] , \SHIFT_n[13][52] , 
        \SHIFT_n[13][51] , \SHIFT_n[13][50] , \SHIFT_n[13][49] , 
        \SHIFT_n[13][48] , \SHIFT_n[13][47] , \SHIFT_n[13][46] , 
        \SHIFT_n[13][45] , \SHIFT_n[13][44] , \SHIFT_n[13][43] , 
        \SHIFT_n[13][42] , \SHIFT_n[13][41] , \SHIFT_n[13][40] , 
        \SHIFT_n[13][39] , \SHIFT_n[13][38] , \SHIFT_n[13][37] , 
        \SHIFT_n[13][36] , \SHIFT_n[13][35] , \SHIFT_n[13][34] , 
        \SHIFT_n[13][33] , \SHIFT_n[13][32] , \SHIFT_n[13][31] , 
        \SHIFT_n[13][30] , \SHIFT_n[13][29] , \SHIFT_n[13][28] , 
        \SHIFT_n[13][27] , \SHIFT_n[13][26] , \SHIFT_n[13][25] , 
        \SHIFT_n[13][24] , \SHIFT_n[13][23] , \SHIFT_n[13][22] , 
        \SHIFT_n[13][21] , \SHIFT_n[13][20] , \SHIFT_n[13][19] , 
        \SHIFT_n[13][18] , \SHIFT_n[13][17] , \SHIFT_n[13][16] , 
        \SHIFT_n[13][15] , \SHIFT_n[13][14] , \SHIFT_n[13][13] , 
        \SHIFT_n[13][12] , \SHIFT_n[13][11] , \SHIFT_n[13][10] , 
        \SHIFT_n[13][9] , \SHIFT_n[13][8] , \SHIFT_n[13][7] , \SHIFT_n[13][6] , 
        \SHIFT_n[13][5] , \SHIFT_n[13][4] , \SHIFT_n[13][3] , \SHIFT_n[13][2] , 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61}) );
  BOOTHENC_NBIT60_i26 ENC_13 ( .A_s({\SHIFT[13][57] , \SHIFT[13][57] , 
        \SHIFT[13][57] , \SHIFT[13][56] , \SHIFT[13][55] , \SHIFT[13][54] , 
        \SHIFT[13][53] , \SHIFT[13][52] , \SHIFT[13][51] , \SHIFT[13][50] , 
        \SHIFT[13][49] , \SHIFT[13][48] , \SHIFT[13][47] , \SHIFT[13][46] , 
        \SHIFT[13][45] , \SHIFT[13][44] , \SHIFT[13][43] , \SHIFT[13][42] , 
        \SHIFT[13][41] , \SHIFT[13][40] , \SHIFT[13][39] , \SHIFT[13][38] , 
        \SHIFT[13][37] , \SHIFT[13][36] , \SHIFT[13][35] , \SHIFT[13][34] , 
        \SHIFT[13][33] , \SHIFT[13][32] , \SHIFT[13][31] , \SHIFT[13][30] , 
        \SHIFT[13][29] , \SHIFT[13][28] , \SHIFT[13][27] , \SHIFT[13][26] , 
        \SHIFT[13][25] , \SHIFT[13][24] , \SHIFT[13][23] , \SHIFT[13][22] , 
        \SHIFT[13][21] , \SHIFT[13][20] , \SHIFT[13][19] , \SHIFT[13][18] , 
        \SHIFT[13][17] , \SHIFT[13][16] , \SHIFT[13][15] , \SHIFT[13][14] , 
        \SHIFT[13][13] , \SHIFT[13][12] , \SHIFT[13][11] , \SHIFT[13][10] , 
        \SHIFT[13][9] , \SHIFT[13][8] , \SHIFT[13][7] , \SHIFT[13][6] , 
        \SHIFT[13][5] , \SHIFT[13][4] , \SHIFT[13][3] , \SHIFT[13][2] , 1'b0, 
        1'b0}), .A_ns({\SHIFT_n[13][57] , \SHIFT_n[13][57] , \SHIFT_n[13][57] , 
        \SHIFT_n[13][56] , \SHIFT_n[13][55] , \SHIFT_n[13][54] , 
        \SHIFT_n[13][53] , \SHIFT_n[13][52] , \SHIFT_n[13][51] , 
        \SHIFT_n[13][50] , \SHIFT_n[13][49] , \SHIFT_n[13][48] , 
        \SHIFT_n[13][47] , \SHIFT_n[13][46] , \SHIFT_n[13][45] , 
        \SHIFT_n[13][44] , \SHIFT_n[13][43] , \SHIFT_n[13][42] , 
        \SHIFT_n[13][41] , \SHIFT_n[13][40] , \SHIFT_n[13][39] , 
        \SHIFT_n[13][38] , \SHIFT_n[13][37] , \SHIFT_n[13][36] , 
        \SHIFT_n[13][35] , \SHIFT_n[13][34] , \SHIFT_n[13][33] , 
        \SHIFT_n[13][32] , \SHIFT_n[13][31] , \SHIFT_n[13][30] , 
        \SHIFT_n[13][29] , \SHIFT_n[13][28] , \SHIFT_n[13][27] , 
        \SHIFT_n[13][26] , \SHIFT_n[13][25] , \SHIFT_n[13][24] , 
        \SHIFT_n[13][23] , \SHIFT_n[13][22] , \SHIFT_n[13][21] , 
        \SHIFT_n[13][20] , \SHIFT_n[13][19] , \SHIFT_n[13][18] , 
        \SHIFT_n[13][17] , \SHIFT_n[13][16] , \SHIFT_n[13][15] , 
        \SHIFT_n[13][14] , \SHIFT_n[13][13] , \SHIFT_n[13][12] , 
        \SHIFT_n[13][11] , \SHIFT_n[13][10] , \SHIFT_n[13][9] , 
        \SHIFT_n[13][8] , \SHIFT_n[13][7] , \SHIFT_n[13][6] , \SHIFT_n[13][5] , 
        \SHIFT_n[13][4] , \SHIFT_n[13][3] , \SHIFT_n[13][2] , 1'b0, 1'b0}), 
        .B({B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B}), 
        .O({\OTMP[13][59] , \OTMP[13][58] , \OTMP[13][57] , \OTMP[13][56] , 
        \OTMP[13][55] , \OTMP[13][54] , \OTMP[13][53] , \OTMP[13][52] , 
        \OTMP[13][51] , \OTMP[13][50] , \OTMP[13][49] , \OTMP[13][48] , 
        \OTMP[13][47] , \OTMP[13][46] , \OTMP[13][45] , \OTMP[13][44] , 
        \OTMP[13][43] , \OTMP[13][42] , \OTMP[13][41] , \OTMP[13][40] , 
        \OTMP[13][39] , \OTMP[13][38] , \OTMP[13][37] , \OTMP[13][36] , 
        \OTMP[13][35] , \OTMP[13][34] , \OTMP[13][33] , \OTMP[13][32] , 
        \OTMP[13][31] , \OTMP[13][30] , \OTMP[13][29] , \OTMP[13][28] , 
        \OTMP[13][27] , \OTMP[13][26] , \OTMP[13][25] , \OTMP[13][24] , 
        \OTMP[13][23] , \OTMP[13][22] , \OTMP[13][21] , \OTMP[13][20] , 
        \OTMP[13][19] , \OTMP[13][18] , \OTMP[13][17] , \OTMP[13][16] , 
        \OTMP[13][15] , \OTMP[13][14] , \OTMP[13][13] , \OTMP[13][12] , 
        \OTMP[13][11] , \OTMP[13][10] , \OTMP[13][9] , \OTMP[13][8] , 
        \OTMP[13][7] , \OTMP[13][6] , \OTMP[13][5] , \OTMP[13][4] , 
        \OTMP[13][3] , \OTMP[13][2] , \OTMP[13][1] , SYNOPSYS_UNCONNECTED__62}), .A_so({\SHIFT[14][59] , \SHIFT[14][58] , \SHIFT[14][57] , \SHIFT[14][56] , 
        \SHIFT[14][55] , \SHIFT[14][54] , \SHIFT[14][53] , \SHIFT[14][52] , 
        \SHIFT[14][51] , \SHIFT[14][50] , \SHIFT[14][49] , \SHIFT[14][48] , 
        \SHIFT[14][47] , \SHIFT[14][46] , \SHIFT[14][45] , \SHIFT[14][44] , 
        \SHIFT[14][43] , \SHIFT[14][42] , \SHIFT[14][41] , \SHIFT[14][40] , 
        \SHIFT[14][39] , \SHIFT[14][38] , \SHIFT[14][37] , \SHIFT[14][36] , 
        \SHIFT[14][35] , \SHIFT[14][34] , \SHIFT[14][33] , \SHIFT[14][32] , 
        \SHIFT[14][31] , \SHIFT[14][30] , \SHIFT[14][29] , \SHIFT[14][28] , 
        \SHIFT[14][27] , \SHIFT[14][26] , \SHIFT[14][25] , \SHIFT[14][24] , 
        \SHIFT[14][23] , \SHIFT[14][22] , \SHIFT[14][21] , \SHIFT[14][20] , 
        \SHIFT[14][19] , \SHIFT[14][18] , \SHIFT[14][17] , \SHIFT[14][16] , 
        \SHIFT[14][15] , \SHIFT[14][14] , \SHIFT[14][13] , \SHIFT[14][12] , 
        \SHIFT[14][11] , \SHIFT[14][10] , \SHIFT[14][9] , \SHIFT[14][8] , 
        \SHIFT[14][7] , \SHIFT[14][6] , \SHIFT[14][5] , \SHIFT[14][4] , 
        \SHIFT[14][3] , \SHIFT[14][2] , SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64}), .A_nso({\SHIFT_n[14][59] , 
        \SHIFT_n[14][58] , \SHIFT_n[14][57] , \SHIFT_n[14][56] , 
        \SHIFT_n[14][55] , \SHIFT_n[14][54] , \SHIFT_n[14][53] , 
        \SHIFT_n[14][52] , \SHIFT_n[14][51] , \SHIFT_n[14][50] , 
        \SHIFT_n[14][49] , \SHIFT_n[14][48] , \SHIFT_n[14][47] , 
        \SHIFT_n[14][46] , \SHIFT_n[14][45] , \SHIFT_n[14][44] , 
        \SHIFT_n[14][43] , \SHIFT_n[14][42] , \SHIFT_n[14][41] , 
        \SHIFT_n[14][40] , \SHIFT_n[14][39] , \SHIFT_n[14][38] , 
        \SHIFT_n[14][37] , \SHIFT_n[14][36] , \SHIFT_n[14][35] , 
        \SHIFT_n[14][34] , \SHIFT_n[14][33] , \SHIFT_n[14][32] , 
        \SHIFT_n[14][31] , \SHIFT_n[14][30] , \SHIFT_n[14][29] , 
        \SHIFT_n[14][28] , \SHIFT_n[14][27] , \SHIFT_n[14][26] , 
        \SHIFT_n[14][25] , \SHIFT_n[14][24] , \SHIFT_n[14][23] , 
        \SHIFT_n[14][22] , \SHIFT_n[14][21] , \SHIFT_n[14][20] , 
        \SHIFT_n[14][19] , \SHIFT_n[14][18] , \SHIFT_n[14][17] , 
        \SHIFT_n[14][16] , \SHIFT_n[14][15] , \SHIFT_n[14][14] , 
        \SHIFT_n[14][13] , \SHIFT_n[14][12] , \SHIFT_n[14][11] , 
        \SHIFT_n[14][10] , \SHIFT_n[14][9] , \SHIFT_n[14][8] , 
        \SHIFT_n[14][7] , \SHIFT_n[14][6] , \SHIFT_n[14][5] , \SHIFT_n[14][4] , 
        \SHIFT_n[14][3] , \SHIFT_n[14][2] , SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66}) );
  BOOTHENC_NBIT62_i28 ENC_14 ( .A_s({\SHIFT[14][59] , \SHIFT[14][59] , 
        \SHIFT[14][59] , \SHIFT[14][58] , \SHIFT[14][57] , \SHIFT[14][56] , 
        \SHIFT[14][55] , \SHIFT[14][54] , \SHIFT[14][53] , \SHIFT[14][52] , 
        \SHIFT[14][51] , \SHIFT[14][50] , \SHIFT[14][49] , \SHIFT[14][48] , 
        \SHIFT[14][47] , \SHIFT[14][46] , \SHIFT[14][45] , \SHIFT[14][44] , 
        \SHIFT[14][43] , \SHIFT[14][42] , \SHIFT[14][41] , \SHIFT[14][40] , 
        \SHIFT[14][39] , \SHIFT[14][38] , \SHIFT[14][37] , \SHIFT[14][36] , 
        \SHIFT[14][35] , \SHIFT[14][34] , \SHIFT[14][33] , \SHIFT[14][32] , 
        \SHIFT[14][31] , \SHIFT[14][30] , \SHIFT[14][29] , \SHIFT[14][28] , 
        \SHIFT[14][27] , \SHIFT[14][26] , \SHIFT[14][25] , \SHIFT[14][24] , 
        \SHIFT[14][23] , \SHIFT[14][22] , \SHIFT[14][21] , \SHIFT[14][20] , 
        \SHIFT[14][19] , \SHIFT[14][18] , \SHIFT[14][17] , \SHIFT[14][16] , 
        \SHIFT[14][15] , \SHIFT[14][14] , \SHIFT[14][13] , \SHIFT[14][12] , 
        \SHIFT[14][11] , \SHIFT[14][10] , \SHIFT[14][9] , \SHIFT[14][8] , 
        \SHIFT[14][7] , \SHIFT[14][6] , \SHIFT[14][5] , \SHIFT[14][4] , 
        \SHIFT[14][3] , \SHIFT[14][2] , 1'b0, 1'b0}), .A_ns({\SHIFT_n[14][59] , 
        \SHIFT_n[14][59] , \SHIFT_n[14][59] , \SHIFT_n[14][58] , 
        \SHIFT_n[14][57] , \SHIFT_n[14][56] , \SHIFT_n[14][55] , 
        \SHIFT_n[14][54] , \SHIFT_n[14][53] , \SHIFT_n[14][52] , 
        \SHIFT_n[14][51] , \SHIFT_n[14][50] , \SHIFT_n[14][49] , 
        \SHIFT_n[14][48] , \SHIFT_n[14][47] , \SHIFT_n[14][46] , 
        \SHIFT_n[14][45] , \SHIFT_n[14][44] , \SHIFT_n[14][43] , 
        \SHIFT_n[14][42] , \SHIFT_n[14][41] , \SHIFT_n[14][40] , 
        \SHIFT_n[14][39] , \SHIFT_n[14][38] , \SHIFT_n[14][37] , 
        \SHIFT_n[14][36] , \SHIFT_n[14][35] , \SHIFT_n[14][34] , 
        \SHIFT_n[14][33] , \SHIFT_n[14][32] , \SHIFT_n[14][31] , 
        \SHIFT_n[14][30] , \SHIFT_n[14][29] , \SHIFT_n[14][28] , 
        \SHIFT_n[14][27] , \SHIFT_n[14][26] , \SHIFT_n[14][25] , 
        \SHIFT_n[14][24] , \SHIFT_n[14][23] , \SHIFT_n[14][22] , 
        \SHIFT_n[14][21] , \SHIFT_n[14][20] , \SHIFT_n[14][19] , 
        \SHIFT_n[14][18] , \SHIFT_n[14][17] , \SHIFT_n[14][16] , 
        \SHIFT_n[14][15] , \SHIFT_n[14][14] , \SHIFT_n[14][13] , 
        \SHIFT_n[14][12] , \SHIFT_n[14][11] , \SHIFT_n[14][10] , 
        \SHIFT_n[14][9] , \SHIFT_n[14][8] , \SHIFT_n[14][7] , \SHIFT_n[14][6] , 
        \SHIFT_n[14][5] , \SHIFT_n[14][4] , \SHIFT_n[14][3] , \SHIFT_n[14][2] , 
        1'b0, 1'b0}), .B({B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B}), .O({\OTMP[14][61] , \OTMP[14][60] , 
        \OTMP[14][59] , \OTMP[14][58] , \OTMP[14][57] , \OTMP[14][56] , 
        \OTMP[14][55] , \OTMP[14][54] , \OTMP[14][53] , \OTMP[14][52] , 
        \OTMP[14][51] , \OTMP[14][50] , \OTMP[14][49] , \OTMP[14][48] , 
        \OTMP[14][47] , \OTMP[14][46] , \OTMP[14][45] , \OTMP[14][44] , 
        \OTMP[14][43] , \OTMP[14][42] , \OTMP[14][41] , \OTMP[14][40] , 
        \OTMP[14][39] , \OTMP[14][38] , \OTMP[14][37] , \OTMP[14][36] , 
        \OTMP[14][35] , \OTMP[14][34] , \OTMP[14][33] , \OTMP[14][32] , 
        \OTMP[14][31] , \OTMP[14][30] , \OTMP[14][29] , \OTMP[14][28] , 
        \OTMP[14][27] , \OTMP[14][26] , \OTMP[14][25] , \OTMP[14][24] , 
        \OTMP[14][23] , \OTMP[14][22] , \OTMP[14][21] , \OTMP[14][20] , 
        \OTMP[14][19] , \OTMP[14][18] , \OTMP[14][17] , \OTMP[14][16] , 
        \OTMP[14][15] , \OTMP[14][14] , \OTMP[14][13] , \OTMP[14][12] , 
        \OTMP[14][11] , \OTMP[14][10] , \OTMP[14][9] , \OTMP[14][8] , 
        \OTMP[14][7] , \OTMP[14][6] , \OTMP[14][5] , \OTMP[14][4] , 
        \OTMP[14][3] , \OTMP[14][2] , \OTMP[14][1] , SYNOPSYS_UNCONNECTED__67}), .A_so({\SHIFT[15][61] , \SHIFT[15][60] , \SHIFT[15][59] , \SHIFT[15][58] , 
        \SHIFT[15][57] , \SHIFT[15][56] , \SHIFT[15][55] , \SHIFT[15][54] , 
        \SHIFT[15][53] , \SHIFT[15][52] , \SHIFT[15][51] , \SHIFT[15][50] , 
        \SHIFT[15][49] , \SHIFT[15][48] , \SHIFT[15][47] , \SHIFT[15][46] , 
        \SHIFT[15][45] , \SHIFT[15][44] , \SHIFT[15][43] , \SHIFT[15][42] , 
        \SHIFT[15][41] , \SHIFT[15][40] , \SHIFT[15][39] , \SHIFT[15][38] , 
        \SHIFT[15][37] , \SHIFT[15][36] , \SHIFT[15][35] , \SHIFT[15][34] , 
        \SHIFT[15][33] , \SHIFT[15][32] , \SHIFT[15][31] , \SHIFT[15][30] , 
        \SHIFT[15][29] , \SHIFT[15][28] , \SHIFT[15][27] , \SHIFT[15][26] , 
        \SHIFT[15][25] , \SHIFT[15][24] , \SHIFT[15][23] , \SHIFT[15][22] , 
        \SHIFT[15][21] , \SHIFT[15][20] , \SHIFT[15][19] , \SHIFT[15][18] , 
        \SHIFT[15][17] , \SHIFT[15][16] , \SHIFT[15][15] , \SHIFT[15][14] , 
        \SHIFT[15][13] , \SHIFT[15][12] , \SHIFT[15][11] , \SHIFT[15][10] , 
        \SHIFT[15][9] , \SHIFT[15][8] , \SHIFT[15][7] , \SHIFT[15][6] , 
        \SHIFT[15][5] , \SHIFT[15][4] , \SHIFT[15][3] , \SHIFT[15][2] , 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69}), .A_nso({
        \SHIFT_n[15][61] , \SHIFT_n[15][60] , \SHIFT_n[15][59] , 
        \SHIFT_n[15][58] , \SHIFT_n[15][57] , \SHIFT_n[15][56] , 
        \SHIFT_n[15][55] , \SHIFT_n[15][54] , \SHIFT_n[15][53] , 
        \SHIFT_n[15][52] , \SHIFT_n[15][51] , \SHIFT_n[15][50] , 
        \SHIFT_n[15][49] , \SHIFT_n[15][48] , \SHIFT_n[15][47] , 
        \SHIFT_n[15][46] , \SHIFT_n[15][45] , \SHIFT_n[15][44] , 
        \SHIFT_n[15][43] , \SHIFT_n[15][42] , \SHIFT_n[15][41] , 
        \SHIFT_n[15][40] , \SHIFT_n[15][39] , \SHIFT_n[15][38] , 
        \SHIFT_n[15][37] , \SHIFT_n[15][36] , \SHIFT_n[15][35] , 
        \SHIFT_n[15][34] , \SHIFT_n[15][33] , \SHIFT_n[15][32] , 
        \SHIFT_n[15][31] , \SHIFT_n[15][30] , \SHIFT_n[15][29] , 
        \SHIFT_n[15][28] , \SHIFT_n[15][27] , \SHIFT_n[15][26] , 
        \SHIFT_n[15][25] , \SHIFT_n[15][24] , \SHIFT_n[15][23] , 
        \SHIFT_n[15][22] , \SHIFT_n[15][21] , \SHIFT_n[15][20] , 
        \SHIFT_n[15][19] , \SHIFT_n[15][18] , \SHIFT_n[15][17] , 
        \SHIFT_n[15][16] , \SHIFT_n[15][15] , \SHIFT_n[15][14] , 
        \SHIFT_n[15][13] , \SHIFT_n[15][12] , \SHIFT_n[15][11] , 
        \SHIFT_n[15][10] , \SHIFT_n[15][9] , \SHIFT_n[15][8] , 
        \SHIFT_n[15][7] , \SHIFT_n[15][6] , \SHIFT_n[15][5] , \SHIFT_n[15][4] , 
        \SHIFT_n[15][3] , \SHIFT_n[15][2] , SYNOPSYS_UNCONNECTED__70, 
        SYNOPSYS_UNCONNECTED__71}) );
  BOOTHENC_NBIT64_i30 ENC_15 ( .A_s({\SHIFT[15][61] , \SHIFT[15][61] , 
        \SHIFT[15][61] , \SHIFT[15][60] , \SHIFT[15][59] , \SHIFT[15][58] , 
        \SHIFT[15][57] , \SHIFT[15][56] , \SHIFT[15][55] , \SHIFT[15][54] , 
        \SHIFT[15][53] , \SHIFT[15][52] , \SHIFT[15][51] , \SHIFT[15][50] , 
        \SHIFT[15][49] , \SHIFT[15][48] , \SHIFT[15][47] , \SHIFT[15][46] , 
        \SHIFT[15][45] , \SHIFT[15][44] , \SHIFT[15][43] , \SHIFT[15][42] , 
        \SHIFT[15][41] , \SHIFT[15][40] , \SHIFT[15][39] , \SHIFT[15][38] , 
        \SHIFT[15][37] , \SHIFT[15][36] , \SHIFT[15][35] , \SHIFT[15][34] , 
        \SHIFT[15][33] , \SHIFT[15][32] , \SHIFT[15][31] , \SHIFT[15][30] , 
        \SHIFT[15][29] , \SHIFT[15][28] , \SHIFT[15][27] , \SHIFT[15][26] , 
        \SHIFT[15][25] , \SHIFT[15][24] , \SHIFT[15][23] , \SHIFT[15][22] , 
        \SHIFT[15][21] , \SHIFT[15][20] , \SHIFT[15][19] , \SHIFT[15][18] , 
        \SHIFT[15][17] , \SHIFT[15][16] , \SHIFT[15][15] , \SHIFT[15][14] , 
        \SHIFT[15][13] , \SHIFT[15][12] , \SHIFT[15][11] , \SHIFT[15][10] , 
        \SHIFT[15][9] , \SHIFT[15][8] , \SHIFT[15][7] , \SHIFT[15][6] , 
        \SHIFT[15][5] , \SHIFT[15][4] , \SHIFT[15][3] , \SHIFT[15][2] , 1'b0, 
        1'b0}), .A_ns({\SHIFT_n[15][61] , \SHIFT_n[15][61] , \SHIFT_n[15][61] , 
        \SHIFT_n[15][60] , \SHIFT_n[15][59] , \SHIFT_n[15][58] , 
        \SHIFT_n[15][57] , \SHIFT_n[15][56] , \SHIFT_n[15][55] , 
        \SHIFT_n[15][54] , \SHIFT_n[15][53] , \SHIFT_n[15][52] , 
        \SHIFT_n[15][51] , \SHIFT_n[15][50] , \SHIFT_n[15][49] , 
        \SHIFT_n[15][48] , \SHIFT_n[15][47] , \SHIFT_n[15][46] , 
        \SHIFT_n[15][45] , \SHIFT_n[15][44] , \SHIFT_n[15][43] , 
        \SHIFT_n[15][42] , \SHIFT_n[15][41] , \SHIFT_n[15][40] , 
        \SHIFT_n[15][39] , \SHIFT_n[15][38] , \SHIFT_n[15][37] , 
        \SHIFT_n[15][36] , \SHIFT_n[15][35] , \SHIFT_n[15][34] , 
        \SHIFT_n[15][33] , \SHIFT_n[15][32] , \SHIFT_n[15][31] , 
        \SHIFT_n[15][30] , \SHIFT_n[15][29] , \SHIFT_n[15][28] , 
        \SHIFT_n[15][27] , \SHIFT_n[15][26] , \SHIFT_n[15][25] , 
        \SHIFT_n[15][24] , \SHIFT_n[15][23] , \SHIFT_n[15][22] , 
        \SHIFT_n[15][21] , \SHIFT_n[15][20] , \SHIFT_n[15][19] , 
        \SHIFT_n[15][18] , \SHIFT_n[15][17] , \SHIFT_n[15][16] , 
        \SHIFT_n[15][15] , \SHIFT_n[15][14] , \SHIFT_n[15][13] , 
        \SHIFT_n[15][12] , \SHIFT_n[15][11] , \SHIFT_n[15][10] , 
        \SHIFT_n[15][9] , \SHIFT_n[15][8] , \SHIFT_n[15][7] , \SHIFT_n[15][6] , 
        \SHIFT_n[15][5] , \SHIFT_n[15][4] , \SHIFT_n[15][3] , \SHIFT_n[15][2] , 
        1'b0, 1'b0}), .B({B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B}), .O({\OTMP[15][63] , 
        \OTMP[15][62] , \OTMP[15][61] , \OTMP[15][60] , \OTMP[15][59] , 
        \OTMP[15][58] , \OTMP[15][57] , \OTMP[15][56] , \OTMP[15][55] , 
        \OTMP[15][54] , \OTMP[15][53] , \OTMP[15][52] , \OTMP[15][51] , 
        \OTMP[15][50] , \OTMP[15][49] , \OTMP[15][48] , \OTMP[15][47] , 
        \OTMP[15][46] , \OTMP[15][45] , \OTMP[15][44] , \OTMP[15][43] , 
        \OTMP[15][42] , \OTMP[15][41] , \OTMP[15][40] , \OTMP[15][39] , 
        \OTMP[15][38] , \OTMP[15][37] , \OTMP[15][36] , \OTMP[15][35] , 
        \OTMP[15][34] , \OTMP[15][33] , \OTMP[15][32] , \OTMP[15][31] , 
        \OTMP[15][30] , \OTMP[15][29] , \OTMP[15][28] , \OTMP[15][27] , 
        \OTMP[15][26] , \OTMP[15][25] , \OTMP[15][24] , \OTMP[15][23] , 
        \OTMP[15][22] , \OTMP[15][21] , \OTMP[15][20] , \OTMP[15][19] , 
        \OTMP[15][18] , \OTMP[15][17] , \OTMP[15][16] , \OTMP[15][15] , 
        \OTMP[15][14] , \OTMP[15][13] , \OTMP[15][12] , \OTMP[15][11] , 
        \OTMP[15][10] , \OTMP[15][9] , \OTMP[15][8] , \OTMP[15][7] , 
        \OTMP[15][6] , \OTMP[15][5] , \OTMP[15][4] , \OTMP[15][3] , 
        \OTMP[15][2] , \OTMP[15][1] , SYNOPSYS_UNCONNECTED__72}) );
  RCA_NBIT36 ADDER1 ( .A({\OTMP[0][34] , \OTMP[0][34] , \OTMP[0][34] , 
        \OTMP[0][32] , \OTMP[0][31] , \OTMP[0][30] , \OTMP[0][29] , 
        \OTMP[0][28] , \OTMP[0][27] , \OTMP[0][26] , \OTMP[0][25] , 
        \OTMP[0][24] , \OTMP[0][23] , \OTMP[0][22] , \OTMP[0][21] , 
        \OTMP[0][20] , \OTMP[0][19] , \OTMP[0][18] , \OTMP[0][17] , 
        \OTMP[0][16] , \OTMP[0][15] , \OTMP[0][14] , \OTMP[0][13] , 
        \OTMP[0][12] , \OTMP[0][11] , \OTMP[0][10] , \OTMP[0][9] , 
        \OTMP[0][8] , \OTMP[0][7] , \OTMP[0][6] , \OTMP[0][5] , \OTMP[0][4] , 
        \OTMP[0][3] , \OTMP[0][2] , \OTMP[0][1] , \OTMP[0][0] }), .B({
        \OTMP[1][35] , \OTMP[1][34] , \OTMP[1][33] , \OTMP[1][32] , 
        \OTMP[1][31] , \OTMP[1][30] , \OTMP[1][29] , \OTMP[1][28] , 
        \OTMP[1][27] , \OTMP[1][26] , \OTMP[1][25] , \OTMP[1][24] , 
        \OTMP[1][23] , \OTMP[1][22] , \OTMP[1][21] , \OTMP[1][20] , 
        \OTMP[1][19] , \OTMP[1][18] , \OTMP[1][17] , \OTMP[1][16] , 
        \OTMP[1][15] , \OTMP[1][14] , \OTMP[1][13] , \OTMP[1][12] , 
        \OTMP[1][11] , \OTMP[1][10] , \OTMP[1][9] , \OTMP[1][8] , \OTMP[1][7] , 
        \OTMP[1][6] , \OTMP[1][5] , \OTMP[1][4] , \OTMP[1][3] , \OTMP[1][2] , 
        \OTMP[1][1] , 1'b0}), .Ci(1'b0), .S({\PTMP[0][36] , \PTMP[0][34] , 
        \PTMP[0][33] , \PTMP[0][32] , \PTMP[0][31] , \PTMP[0][30] , 
        \PTMP[0][29] , \PTMP[0][28] , \PTMP[0][27] , \PTMP[0][26] , 
        \PTMP[0][25] , \PTMP[0][24] , \PTMP[0][23] , \PTMP[0][22] , 
        \PTMP[0][21] , \PTMP[0][20] , \PTMP[0][19] , \PTMP[0][18] , 
        \PTMP[0][17] , \PTMP[0][16] , \PTMP[0][15] , \PTMP[0][14] , 
        \PTMP[0][13] , \PTMP[0][12] , \PTMP[0][11] , \PTMP[0][10] , 
        \PTMP[0][9] , \PTMP[0][8] , \PTMP[0][7] , \PTMP[0][6] , \PTMP[0][5] , 
        \PTMP[0][4] , \PTMP[0][3] , \PTMP[0][2] , \PTMP[0][1] , \PTMP[0][0] })
         );
  RCA_NBIT38 ADDER_2 ( .A({\PTMP[0][36] , \PTMP[0][36] , \PTMP[0][36] , 
        \PTMP[0][34] , \PTMP[0][33] , \PTMP[0][32] , \PTMP[0][31] , 
        \PTMP[0][30] , \PTMP[0][29] , \PTMP[0][28] , \PTMP[0][27] , 
        \PTMP[0][26] , \PTMP[0][25] , \PTMP[0][24] , \PTMP[0][23] , 
        \PTMP[0][22] , \PTMP[0][21] , \PTMP[0][20] , \PTMP[0][19] , 
        \PTMP[0][18] , \PTMP[0][17] , \PTMP[0][16] , \PTMP[0][15] , 
        \PTMP[0][14] , \PTMP[0][13] , \PTMP[0][12] , \PTMP[0][11] , 
        \PTMP[0][10] , \PTMP[0][9] , \PTMP[0][8] , \PTMP[0][7] , \PTMP[0][6] , 
        \PTMP[0][5] , \PTMP[0][4] , \PTMP[0][3] , \PTMP[0][2] , \PTMP[0][1] , 
        \PTMP[0][0] }), .B({\OTMP[2][37] , \OTMP[2][36] , \OTMP[2][35] , 
        \OTMP[2][34] , \OTMP[2][33] , \OTMP[2][32] , \OTMP[2][31] , 
        \OTMP[2][30] , \OTMP[2][29] , \OTMP[2][28] , \OTMP[2][27] , 
        \OTMP[2][26] , \OTMP[2][25] , \OTMP[2][24] , \OTMP[2][23] , 
        \OTMP[2][22] , \OTMP[2][21] , \OTMP[2][20] , \OTMP[2][19] , 
        \OTMP[2][18] , \OTMP[2][17] , \OTMP[2][16] , \OTMP[2][15] , 
        \OTMP[2][14] , \OTMP[2][13] , \OTMP[2][12] , \OTMP[2][11] , 
        \OTMP[2][10] , \OTMP[2][9] , \OTMP[2][8] , \OTMP[2][7] , \OTMP[2][6] , 
        \OTMP[2][5] , \OTMP[2][4] , \OTMP[2][3] , \OTMP[2][2] , \OTMP[2][1] , 
        1'b0}), .Ci(1'b0), .S({\PTMP[1][37] , \PTMP[1][36] , \PTMP[1][35] , 
        \PTMP[1][34] , \PTMP[1][33] , \PTMP[1][32] , \PTMP[1][31] , 
        \PTMP[1][30] , \PTMP[1][29] , \PTMP[1][28] , \PTMP[1][27] , 
        \PTMP[1][26] , \PTMP[1][25] , \PTMP[1][24] , \PTMP[1][23] , 
        \PTMP[1][22] , \PTMP[1][21] , \PTMP[1][20] , \PTMP[1][19] , 
        \PTMP[1][18] , \PTMP[1][17] , \PTMP[1][16] , \PTMP[1][15] , 
        \PTMP[1][14] , \PTMP[1][13] , \PTMP[1][12] , \PTMP[1][11] , 
        \PTMP[1][10] , \PTMP[1][9] , \PTMP[1][8] , \PTMP[1][7] , \PTMP[1][6] , 
        \PTMP[1][5] , \PTMP[1][4] , \PTMP[1][3] , \PTMP[1][2] , \PTMP[1][1] , 
        \PTMP[1][0] }) );
  RCA_NBIT40 ADDER_3 ( .A({\PTMP[1][37] , \PTMP[1][37] , \PTMP[1][37] , 
        \PTMP[1][36] , \PTMP[1][35] , \PTMP[1][34] , \PTMP[1][33] , 
        \PTMP[1][32] , \PTMP[1][31] , \PTMP[1][30] , \PTMP[1][29] , 
        \PTMP[1][28] , \PTMP[1][27] , \PTMP[1][26] , \PTMP[1][25] , 
        \PTMP[1][24] , \PTMP[1][23] , \PTMP[1][22] , \PTMP[1][21] , 
        \PTMP[1][20] , \PTMP[1][19] , \PTMP[1][18] , \PTMP[1][17] , 
        \PTMP[1][16] , \PTMP[1][15] , \PTMP[1][14] , \PTMP[1][13] , 
        \PTMP[1][12] , \PTMP[1][11] , \PTMP[1][10] , \PTMP[1][9] , 
        \PTMP[1][8] , \PTMP[1][7] , \PTMP[1][6] , \PTMP[1][5] , \PTMP[1][4] , 
        \PTMP[1][3] , \PTMP[1][2] , \PTMP[1][1] , \PTMP[1][0] }), .B({
        \OTMP[3][39] , \OTMP[3][38] , \OTMP[3][37] , \OTMP[3][36] , 
        \OTMP[3][35] , \OTMP[3][34] , \OTMP[3][33] , \OTMP[3][32] , 
        \OTMP[3][31] , \OTMP[3][30] , \OTMP[3][29] , \OTMP[3][28] , 
        \OTMP[3][27] , \OTMP[3][26] , \OTMP[3][25] , \OTMP[3][24] , 
        \OTMP[3][23] , \OTMP[3][22] , \OTMP[3][21] , \OTMP[3][20] , 
        \OTMP[3][19] , \OTMP[3][18] , \OTMP[3][17] , \OTMP[3][16] , 
        \OTMP[3][15] , \OTMP[3][14] , \OTMP[3][13] , \OTMP[3][12] , 
        \OTMP[3][11] , \OTMP[3][10] , \OTMP[3][9] , \OTMP[3][8] , \OTMP[3][7] , 
        \OTMP[3][6] , \OTMP[3][5] , \OTMP[3][4] , \OTMP[3][3] , \OTMP[3][2] , 
        \OTMP[3][1] , 1'b0}), .Ci(1'b0), .S({\PTMP[2][39] , \PTMP[2][38] , 
        \PTMP[2][37] , \PTMP[2][36] , \PTMP[2][35] , \PTMP[2][34] , 
        \PTMP[2][33] , \PTMP[2][32] , \PTMP[2][31] , \PTMP[2][30] , 
        \PTMP[2][29] , \PTMP[2][28] , \PTMP[2][27] , \PTMP[2][26] , 
        \PTMP[2][25] , \PTMP[2][24] , \PTMP[2][23] , \PTMP[2][22] , 
        \PTMP[2][21] , \PTMP[2][20] , \PTMP[2][19] , \PTMP[2][18] , 
        \PTMP[2][17] , \PTMP[2][16] , \PTMP[2][15] , \PTMP[2][14] , 
        \PTMP[2][13] , \PTMP[2][12] , \PTMP[2][11] , \PTMP[2][10] , 
        \PTMP[2][9] , \PTMP[2][8] , \PTMP[2][7] , \PTMP[2][6] , \PTMP[2][5] , 
        \PTMP[2][4] , \PTMP[2][3] , \PTMP[2][2] , \PTMP[2][1] , \PTMP[2][0] })
         );
  RCA_NBIT42 ADDER_4 ( .A({n7, n7, \PTMP[2][39] , \PTMP[2][38] , \PTMP[2][37] , 
        \PTMP[2][36] , \PTMP[2][35] , \PTMP[2][34] , \PTMP[2][33] , 
        \PTMP[2][32] , \PTMP[2][31] , \PTMP[2][30] , \PTMP[2][29] , 
        \PTMP[2][28] , \PTMP[2][27] , \PTMP[2][26] , \PTMP[2][25] , 
        \PTMP[2][24] , \PTMP[2][23] , \PTMP[2][22] , \PTMP[2][21] , 
        \PTMP[2][20] , \PTMP[2][19] , \PTMP[2][18] , \PTMP[2][17] , 
        \PTMP[2][16] , \PTMP[2][15] , \PTMP[2][14] , \PTMP[2][13] , 
        \PTMP[2][12] , \PTMP[2][11] , \PTMP[2][10] , \PTMP[2][9] , 
        \PTMP[2][8] , \PTMP[2][7] , \PTMP[2][6] , \PTMP[2][5] , \PTMP[2][4] , 
        \PTMP[2][3] , \PTMP[2][2] , \PTMP[2][1] , \PTMP[2][0] }), .B({
        \OTMP[4][41] , \OTMP[4][40] , \OTMP[4][39] , \OTMP[4][38] , 
        \OTMP[4][37] , \OTMP[4][36] , \OTMP[4][35] , \OTMP[4][34] , 
        \OTMP[4][33] , \OTMP[4][32] , \OTMP[4][31] , \OTMP[4][30] , 
        \OTMP[4][29] , \OTMP[4][28] , \OTMP[4][27] , \OTMP[4][26] , 
        \OTMP[4][25] , \OTMP[4][24] , \OTMP[4][23] , \OTMP[4][22] , 
        \OTMP[4][21] , \OTMP[4][20] , \OTMP[4][19] , \OTMP[4][18] , 
        \OTMP[4][17] , \OTMP[4][16] , \OTMP[4][15] , \OTMP[4][14] , 
        \OTMP[4][13] , \OTMP[4][12] , \OTMP[4][11] , \OTMP[4][10] , 
        \OTMP[4][9] , \OTMP[4][8] , \OTMP[4][7] , \OTMP[4][6] , \OTMP[4][5] , 
        \OTMP[4][4] , \OTMP[4][3] , \OTMP[4][2] , \OTMP[4][1] , 1'b0}), .Ci(
        1'b0), .S({\PTMP[3][41] , \PTMP[3][40] , \PTMP[3][39] , \PTMP[3][38] , 
        \PTMP[3][37] , \PTMP[3][36] , \PTMP[3][35] , \PTMP[3][34] , 
        \PTMP[3][33] , \PTMP[3][32] , \PTMP[3][31] , \PTMP[3][30] , 
        \PTMP[3][29] , \PTMP[3][28] , \PTMP[3][27] , \PTMP[3][26] , 
        \PTMP[3][25] , \PTMP[3][24] , \PTMP[3][23] , \PTMP[3][22] , 
        \PTMP[3][21] , \PTMP[3][20] , \PTMP[3][19] , \PTMP[3][18] , 
        \PTMP[3][17] , \PTMP[3][16] , \PTMP[3][15] , \PTMP[3][14] , 
        \PTMP[3][13] , \PTMP[3][12] , \PTMP[3][11] , \PTMP[3][10] , 
        \PTMP[3][9] , \PTMP[3][8] , \PTMP[3][7] , \PTMP[3][6] , \PTMP[3][5] , 
        \PTMP[3][4] , \PTMP[3][3] , \PTMP[3][2] , \PTMP[3][1] , \PTMP[3][0] })
         );
  RCA_NBIT44 ADDER_5 ( .A({\PTMP[3][41] , \PTMP[3][41] , \PTMP[3][41] , 
        \PTMP[3][40] , \PTMP[3][39] , \PTMP[3][38] , \PTMP[3][37] , 
        \PTMP[3][36] , \PTMP[3][35] , \PTMP[3][34] , \PTMP[3][33] , 
        \PTMP[3][32] , \PTMP[3][31] , \PTMP[3][30] , \PTMP[3][29] , 
        \PTMP[3][28] , \PTMP[3][27] , \PTMP[3][26] , \PTMP[3][25] , 
        \PTMP[3][24] , \PTMP[3][23] , \PTMP[3][22] , \PTMP[3][21] , 
        \PTMP[3][20] , \PTMP[3][19] , \PTMP[3][18] , \PTMP[3][17] , 
        \PTMP[3][16] , \PTMP[3][15] , \PTMP[3][14] , \PTMP[3][13] , 
        \PTMP[3][12] , \PTMP[3][11] , \PTMP[3][10] , \PTMP[3][9] , 
        \PTMP[3][8] , \PTMP[3][7] , \PTMP[3][6] , \PTMP[3][5] , \PTMP[3][4] , 
        \PTMP[3][3] , \PTMP[3][2] , \PTMP[3][1] , \PTMP[3][0] }), .B({
        \OTMP[5][43] , \OTMP[5][42] , \OTMP[5][41] , \OTMP[5][40] , 
        \OTMP[5][39] , \OTMP[5][38] , \OTMP[5][37] , \OTMP[5][36] , 
        \OTMP[5][35] , \OTMP[5][34] , \OTMP[5][33] , \OTMP[5][32] , 
        \OTMP[5][31] , \OTMP[5][30] , \OTMP[5][29] , \OTMP[5][28] , 
        \OTMP[5][27] , \OTMP[5][26] , \OTMP[5][25] , \OTMP[5][24] , 
        \OTMP[5][23] , \OTMP[5][22] , \OTMP[5][21] , \OTMP[5][20] , 
        \OTMP[5][19] , \OTMP[5][18] , \OTMP[5][17] , \OTMP[5][16] , 
        \OTMP[5][15] , \OTMP[5][14] , \OTMP[5][13] , \OTMP[5][12] , 
        \OTMP[5][11] , \OTMP[5][10] , \OTMP[5][9] , \OTMP[5][8] , \OTMP[5][7] , 
        \OTMP[5][6] , \OTMP[5][5] , \OTMP[5][4] , \OTMP[5][3] , \OTMP[5][2] , 
        \OTMP[5][1] , 1'b0}), .Ci(1'b0), .S({\PTMP[4][43] , \PTMP[4][42] , 
        \PTMP[4][41] , \PTMP[4][40] , \PTMP[4][39] , \PTMP[4][38] , 
        \PTMP[4][37] , \PTMP[4][36] , \PTMP[4][35] , \PTMP[4][34] , 
        \PTMP[4][33] , \PTMP[4][32] , \PTMP[4][31] , \PTMP[4][30] , 
        \PTMP[4][29] , \PTMP[4][28] , \PTMP[4][27] , \PTMP[4][26] , 
        \PTMP[4][25] , \PTMP[4][24] , \PTMP[4][23] , \PTMP[4][22] , 
        \PTMP[4][21] , \PTMP[4][20] , \PTMP[4][19] , \PTMP[4][18] , 
        \PTMP[4][17] , \PTMP[4][16] , \PTMP[4][15] , \PTMP[4][14] , 
        \PTMP[4][13] , \PTMP[4][12] , \PTMP[4][11] , \PTMP[4][10] , 
        \PTMP[4][9] , \PTMP[4][8] , \PTMP[4][7] , \PTMP[4][6] , \PTMP[4][5] , 
        \PTMP[4][4] , \PTMP[4][3] , \PTMP[4][2] , \PTMP[4][1] , \PTMP[4][0] })
         );
  RCA_NBIT46 ADDER_6 ( .A({n13, n13, \PTMP[4][43] , \PTMP[4][42] , 
        \PTMP[4][41] , \PTMP[4][40] , \PTMP[4][39] , \PTMP[4][38] , 
        \PTMP[4][37] , \PTMP[4][36] , \PTMP[4][35] , \PTMP[4][34] , 
        \PTMP[4][33] , \PTMP[4][32] , \PTMP[4][31] , \PTMP[4][30] , 
        \PTMP[4][29] , \PTMP[4][28] , \PTMP[4][27] , \PTMP[4][26] , 
        \PTMP[4][25] , \PTMP[4][24] , \PTMP[4][23] , \PTMP[4][22] , 
        \PTMP[4][21] , \PTMP[4][20] , \PTMP[4][19] , \PTMP[4][18] , 
        \PTMP[4][17] , \PTMP[4][16] , \PTMP[4][15] , \PTMP[4][14] , 
        \PTMP[4][13] , \PTMP[4][12] , \PTMP[4][11] , \PTMP[4][10] , 
        \PTMP[4][9] , \PTMP[4][8] , \PTMP[4][7] , \PTMP[4][6] , \PTMP[4][5] , 
        \PTMP[4][4] , \PTMP[4][3] , \PTMP[4][2] , \PTMP[4][1] , \PTMP[4][0] }), 
        .B({\OTMP[6][45] , \OTMP[6][44] , \OTMP[6][43] , \OTMP[6][42] , 
        \OTMP[6][41] , \OTMP[6][40] , \OTMP[6][39] , \OTMP[6][38] , 
        \OTMP[6][37] , \OTMP[6][36] , \OTMP[6][35] , \OTMP[6][34] , 
        \OTMP[6][33] , \OTMP[6][32] , \OTMP[6][31] , \OTMP[6][30] , 
        \OTMP[6][29] , \OTMP[6][28] , \OTMP[6][27] , \OTMP[6][26] , 
        \OTMP[6][25] , \OTMP[6][24] , \OTMP[6][23] , \OTMP[6][22] , 
        \OTMP[6][21] , \OTMP[6][20] , \OTMP[6][19] , \OTMP[6][18] , 
        \OTMP[6][17] , \OTMP[6][16] , \OTMP[6][15] , \OTMP[6][14] , 
        \OTMP[6][13] , \OTMP[6][12] , \OTMP[6][11] , \OTMP[6][10] , 
        \OTMP[6][9] , \OTMP[6][8] , \OTMP[6][7] , \OTMP[6][6] , \OTMP[6][5] , 
        \OTMP[6][4] , \OTMP[6][3] , \OTMP[6][2] , \OTMP[6][1] , 1'b0}), .Ci(
        1'b0), .S({\PTMP[5][45] , \PTMP[5][44] , \PTMP[5][43] , \PTMP[5][42] , 
        \PTMP[5][41] , \PTMP[5][40] , \PTMP[5][39] , \PTMP[5][38] , 
        \PTMP[5][37] , \PTMP[5][36] , \PTMP[5][35] , \PTMP[5][34] , 
        \PTMP[5][33] , \PTMP[5][32] , \PTMP[5][31] , \PTMP[5][30] , 
        \PTMP[5][29] , \PTMP[5][28] , \PTMP[5][27] , \PTMP[5][26] , 
        \PTMP[5][25] , \PTMP[5][24] , \PTMP[5][23] , \PTMP[5][22] , 
        \PTMP[5][21] , \PTMP[5][20] , \PTMP[5][19] , \PTMP[5][18] , 
        \PTMP[5][17] , \PTMP[5][16] , \PTMP[5][15] , \PTMP[5][14] , 
        \PTMP[5][13] , \PTMP[5][12] , \PTMP[5][11] , \PTMP[5][10] , 
        \PTMP[5][9] , \PTMP[5][8] , \PTMP[5][7] , \PTMP[5][6] , \PTMP[5][5] , 
        \PTMP[5][4] , \PTMP[5][3] , \PTMP[5][2] , \PTMP[5][1] , \PTMP[5][0] })
         );
  RCA_NBIT48 ADDER_7 ( .A({n6, n15, \PTMP[5][45] , \PTMP[5][44] , 
        \PTMP[5][43] , \PTMP[5][42] , \PTMP[5][41] , \PTMP[5][40] , 
        \PTMP[5][39] , \PTMP[5][38] , \PTMP[5][37] , \PTMP[5][36] , 
        \PTMP[5][35] , \PTMP[5][34] , \PTMP[5][33] , \PTMP[5][32] , 
        \PTMP[5][31] , \PTMP[5][30] , \PTMP[5][29] , \PTMP[5][28] , 
        \PTMP[5][27] , \PTMP[5][26] , \PTMP[5][25] , \PTMP[5][24] , 
        \PTMP[5][23] , \PTMP[5][22] , \PTMP[5][21] , \PTMP[5][20] , 
        \PTMP[5][19] , \PTMP[5][18] , \PTMP[5][17] , \PTMP[5][16] , 
        \PTMP[5][15] , \PTMP[5][14] , \PTMP[5][13] , \PTMP[5][12] , 
        \PTMP[5][11] , \PTMP[5][10] , \PTMP[5][9] , \PTMP[5][8] , \PTMP[5][7] , 
        \PTMP[5][6] , \PTMP[5][5] , \PTMP[5][4] , \PTMP[5][3] , \PTMP[5][2] , 
        \PTMP[5][1] , \PTMP[5][0] }), .B({\OTMP[7][47] , \OTMP[7][46] , 
        \OTMP[7][45] , \OTMP[7][44] , \OTMP[7][43] , \OTMP[7][42] , 
        \OTMP[7][41] , \OTMP[7][40] , \OTMP[7][39] , \OTMP[7][38] , 
        \OTMP[7][37] , \OTMP[7][36] , \OTMP[7][35] , \OTMP[7][34] , 
        \OTMP[7][33] , \OTMP[7][32] , \OTMP[7][31] , \OTMP[7][30] , 
        \OTMP[7][29] , \OTMP[7][28] , \OTMP[7][27] , \OTMP[7][26] , 
        \OTMP[7][25] , \OTMP[7][24] , \OTMP[7][23] , \OTMP[7][22] , 
        \OTMP[7][21] , \OTMP[7][20] , \OTMP[7][19] , \OTMP[7][18] , 
        \OTMP[7][17] , \OTMP[7][16] , \OTMP[7][15] , \OTMP[7][14] , 
        \OTMP[7][13] , \OTMP[7][12] , \OTMP[7][11] , \OTMP[7][10] , 
        \OTMP[7][9] , \OTMP[7][8] , \OTMP[7][7] , \OTMP[7][6] , \OTMP[7][5] , 
        \OTMP[7][4] , \OTMP[7][3] , \OTMP[7][2] , \OTMP[7][1] , 1'b0}), .Ci(
        1'b0), .S({\PTMP[6][47] , \PTMP[6][46] , \PTMP[6][45] , \PTMP[6][44] , 
        \PTMP[6][43] , \PTMP[6][42] , \PTMP[6][41] , \PTMP[6][40] , 
        \PTMP[6][39] , \PTMP[6][38] , \PTMP[6][37] , \PTMP[6][36] , 
        \PTMP[6][35] , \PTMP[6][34] , \PTMP[6][33] , \PTMP[6][32] , 
        \PTMP[6][31] , \PTMP[6][30] , \PTMP[6][29] , \PTMP[6][28] , 
        \PTMP[6][27] , \PTMP[6][26] , \PTMP[6][25] , \PTMP[6][24] , 
        \PTMP[6][23] , \PTMP[6][22] , \PTMP[6][21] , \PTMP[6][20] , 
        \PTMP[6][19] , \PTMP[6][18] , \PTMP[6][17] , \PTMP[6][16] , 
        \PTMP[6][15] , \PTMP[6][14] , \PTMP[6][13] , \PTMP[6][12] , 
        \PTMP[6][11] , \PTMP[6][10] , \PTMP[6][9] , \PTMP[6][8] , \PTMP[6][7] , 
        \PTMP[6][6] , \PTMP[6][5] , \PTMP[6][4] , \PTMP[6][3] , \PTMP[6][2] , 
        \PTMP[6][1] , \PTMP[6][0] }) );
  RCA_NBIT50 ADDER_8 ( .A({n21, n17, \PTMP[6][47] , \PTMP[6][46] , 
        \PTMP[6][45] , \PTMP[6][44] , \PTMP[6][43] , \PTMP[6][42] , 
        \PTMP[6][41] , \PTMP[6][40] , \PTMP[6][39] , \PTMP[6][38] , 
        \PTMP[6][37] , \PTMP[6][36] , \PTMP[6][35] , \PTMP[6][34] , 
        \PTMP[6][33] , \PTMP[6][32] , \PTMP[6][31] , \PTMP[6][30] , 
        \PTMP[6][29] , \PTMP[6][28] , \PTMP[6][27] , \PTMP[6][26] , 
        \PTMP[6][25] , \PTMP[6][24] , \PTMP[6][23] , \PTMP[6][22] , 
        \PTMP[6][21] , \PTMP[6][20] , \PTMP[6][19] , \PTMP[6][18] , 
        \PTMP[6][17] , \PTMP[6][16] , \PTMP[6][15] , \PTMP[6][14] , 
        \PTMP[6][13] , \PTMP[6][12] , \PTMP[6][11] , \PTMP[6][10] , 
        \PTMP[6][9] , \PTMP[6][8] , \PTMP[6][7] , \PTMP[6][6] , \PTMP[6][5] , 
        \PTMP[6][4] , \PTMP[6][3] , \PTMP[6][2] , \PTMP[6][1] , \PTMP[6][0] }), 
        .B({\OTMP[8][49] , \OTMP[8][48] , \OTMP[8][47] , \OTMP[8][46] , 
        \OTMP[8][45] , \OTMP[8][44] , \OTMP[8][43] , \OTMP[8][42] , 
        \OTMP[8][41] , \OTMP[8][40] , \OTMP[8][39] , \OTMP[8][38] , 
        \OTMP[8][37] , \OTMP[8][36] , \OTMP[8][35] , \OTMP[8][34] , 
        \OTMP[8][33] , \OTMP[8][32] , \OTMP[8][31] , \OTMP[8][30] , 
        \OTMP[8][29] , \OTMP[8][28] , \OTMP[8][27] , \OTMP[8][26] , 
        \OTMP[8][25] , \OTMP[8][24] , \OTMP[8][23] , \OTMP[8][22] , 
        \OTMP[8][21] , \OTMP[8][20] , \OTMP[8][19] , \OTMP[8][18] , 
        \OTMP[8][17] , \OTMP[8][16] , \OTMP[8][15] , \OTMP[8][14] , 
        \OTMP[8][13] , \OTMP[8][12] , \OTMP[8][11] , \OTMP[8][10] , 
        \OTMP[8][9] , \OTMP[8][8] , \OTMP[8][7] , \OTMP[8][6] , \OTMP[8][5] , 
        \OTMP[8][4] , \OTMP[8][3] , \OTMP[8][2] , \OTMP[8][1] , 1'b0}), .Ci(
        1'b0), .S({\PTMP[7][49] , \PTMP[7][48] , \PTMP[7][47] , \PTMP[7][46] , 
        \PTMP[7][45] , \PTMP[7][44] , \PTMP[7][43] , \PTMP[7][42] , 
        \PTMP[7][41] , \PTMP[7][40] , \PTMP[7][39] , \PTMP[7][38] , 
        \PTMP[7][37] , \PTMP[7][36] , \PTMP[7][35] , \PTMP[7][34] , 
        \PTMP[7][33] , \PTMP[7][32] , \PTMP[7][31] , \PTMP[7][30] , 
        \PTMP[7][29] , \PTMP[7][28] , \PTMP[7][27] , \PTMP[7][26] , 
        \PTMP[7][25] , \PTMP[7][24] , \PTMP[7][23] , \PTMP[7][22] , 
        \PTMP[7][21] , \PTMP[7][20] , \PTMP[7][19] , \PTMP[7][18] , 
        \PTMP[7][17] , \PTMP[7][16] , \PTMP[7][15] , \PTMP[7][14] , 
        \PTMP[7][13] , \PTMP[7][12] , \PTMP[7][11] , \PTMP[7][10] , 
        \PTMP[7][9] , \PTMP[7][8] , \PTMP[7][7] , \PTMP[7][6] , \PTMP[7][5] , 
        \PTMP[7][4] , \PTMP[7][3] , \PTMP[7][2] , \PTMP[7][1] , \PTMP[7][0] })
         );
  RCA_NBIT52 ADDER_9 ( .A({n16, n16, \PTMP[7][49] , \PTMP[7][48] , 
        \PTMP[7][47] , \PTMP[7][46] , \PTMP[7][45] , \PTMP[7][44] , 
        \PTMP[7][43] , \PTMP[7][42] , \PTMP[7][41] , \PTMP[7][40] , 
        \PTMP[7][39] , \PTMP[7][38] , \PTMP[7][37] , \PTMP[7][36] , 
        \PTMP[7][35] , \PTMP[7][34] , \PTMP[7][33] , \PTMP[7][32] , 
        \PTMP[7][31] , \PTMP[7][30] , \PTMP[7][29] , \PTMP[7][28] , 
        \PTMP[7][27] , \PTMP[7][26] , \PTMP[7][25] , \PTMP[7][24] , 
        \PTMP[7][23] , \PTMP[7][22] , \PTMP[7][21] , \PTMP[7][20] , 
        \PTMP[7][19] , \PTMP[7][18] , \PTMP[7][17] , \PTMP[7][16] , 
        \PTMP[7][15] , \PTMP[7][14] , \PTMP[7][13] , \PTMP[7][12] , 
        \PTMP[7][11] , \PTMP[7][10] , \PTMP[7][9] , \PTMP[7][8] , \PTMP[7][7] , 
        \PTMP[7][6] , \PTMP[7][5] , \PTMP[7][4] , \PTMP[7][3] , \PTMP[7][2] , 
        \PTMP[7][1] , \PTMP[7][0] }), .B({\OTMP[9][51] , \OTMP[9][50] , 
        \OTMP[9][49] , \OTMP[9][48] , \OTMP[9][47] , \OTMP[9][46] , 
        \OTMP[9][45] , \OTMP[9][44] , \OTMP[9][43] , \OTMP[9][42] , 
        \OTMP[9][41] , \OTMP[9][40] , \OTMP[9][39] , \OTMP[9][38] , 
        \OTMP[9][37] , \OTMP[9][36] , \OTMP[9][35] , \OTMP[9][34] , 
        \OTMP[9][33] , \OTMP[9][32] , \OTMP[9][31] , \OTMP[9][30] , 
        \OTMP[9][29] , \OTMP[9][28] , \OTMP[9][27] , \OTMP[9][26] , 
        \OTMP[9][25] , \OTMP[9][24] , \OTMP[9][23] , \OTMP[9][22] , 
        \OTMP[9][21] , \OTMP[9][20] , \OTMP[9][19] , \OTMP[9][18] , 
        \OTMP[9][17] , \OTMP[9][16] , \OTMP[9][15] , \OTMP[9][14] , 
        \OTMP[9][13] , \OTMP[9][12] , \OTMP[9][11] , \OTMP[9][10] , 
        \OTMP[9][9] , \OTMP[9][8] , \OTMP[9][7] , \OTMP[9][6] , \OTMP[9][5] , 
        \OTMP[9][4] , \OTMP[9][3] , \OTMP[9][2] , \OTMP[9][1] , 1'b0}), .Ci(
        1'b0), .S({\PTMP[8][51] , \PTMP[8][50] , \PTMP[8][49] , \PTMP[8][48] , 
        \PTMP[8][47] , \PTMP[8][46] , \PTMP[8][45] , \PTMP[8][44] , 
        \PTMP[8][43] , \PTMP[8][42] , \PTMP[8][41] , \PTMP[8][40] , 
        \PTMP[8][39] , \PTMP[8][38] , \PTMP[8][37] , \PTMP[8][36] , 
        \PTMP[8][35] , \PTMP[8][34] , \PTMP[8][33] , \PTMP[8][32] , 
        \PTMP[8][31] , \PTMP[8][30] , \PTMP[8][29] , \PTMP[8][28] , 
        \PTMP[8][27] , \PTMP[8][26] , \PTMP[8][25] , \PTMP[8][24] , 
        \PTMP[8][23] , \PTMP[8][22] , \PTMP[8][21] , \PTMP[8][20] , 
        \PTMP[8][19] , \PTMP[8][18] , \PTMP[8][17] , \PTMP[8][16] , 
        \PTMP[8][15] , \PTMP[8][14] , \PTMP[8][13] , \PTMP[8][12] , 
        \PTMP[8][11] , \PTMP[8][10] , \PTMP[8][9] , \PTMP[8][8] , \PTMP[8][7] , 
        \PTMP[8][6] , \PTMP[8][5] , \PTMP[8][4] , \PTMP[8][3] , \PTMP[8][2] , 
        \PTMP[8][1] , \PTMP[8][0] }) );
  RCA_NBIT54 ADDER_10 ( .A({n18, n18, \PTMP[8][51] , \PTMP[8][50] , 
        \PTMP[8][49] , \PTMP[8][48] , \PTMP[8][47] , \PTMP[8][46] , 
        \PTMP[8][45] , \PTMP[8][44] , \PTMP[8][43] , \PTMP[8][42] , 
        \PTMP[8][41] , \PTMP[8][40] , \PTMP[8][39] , \PTMP[8][38] , 
        \PTMP[8][37] , \PTMP[8][36] , \PTMP[8][35] , \PTMP[8][34] , 
        \PTMP[8][33] , \PTMP[8][32] , \PTMP[8][31] , \PTMP[8][30] , 
        \PTMP[8][29] , \PTMP[8][28] , \PTMP[8][27] , \PTMP[8][26] , 
        \PTMP[8][25] , \PTMP[8][24] , \PTMP[8][23] , \PTMP[8][22] , 
        \PTMP[8][21] , \PTMP[8][20] , \PTMP[8][19] , \PTMP[8][18] , 
        \PTMP[8][17] , \PTMP[8][16] , \PTMP[8][15] , \PTMP[8][14] , 
        \PTMP[8][13] , \PTMP[8][12] , \PTMP[8][11] , \PTMP[8][10] , 
        \PTMP[8][9] , \PTMP[8][8] , \PTMP[8][7] , \PTMP[8][6] , \PTMP[8][5] , 
        \PTMP[8][4] , \PTMP[8][3] , \PTMP[8][2] , \PTMP[8][1] , \PTMP[8][0] }), 
        .B({\OTMP[10][53] , \OTMP[10][52] , \OTMP[10][51] , \OTMP[10][50] , 
        \OTMP[10][49] , \OTMP[10][48] , \OTMP[10][47] , \OTMP[10][46] , 
        \OTMP[10][45] , \OTMP[10][44] , \OTMP[10][43] , \OTMP[10][42] , 
        \OTMP[10][41] , \OTMP[10][40] , \OTMP[10][39] , \OTMP[10][38] , 
        \OTMP[10][37] , \OTMP[10][36] , \OTMP[10][35] , \OTMP[10][34] , 
        \OTMP[10][33] , \OTMP[10][32] , \OTMP[10][31] , \OTMP[10][30] , 
        \OTMP[10][29] , \OTMP[10][28] , \OTMP[10][27] , \OTMP[10][26] , 
        \OTMP[10][25] , \OTMP[10][24] , \OTMP[10][23] , \OTMP[10][22] , 
        \OTMP[10][21] , \OTMP[10][20] , \OTMP[10][19] , \OTMP[10][18] , 
        \OTMP[10][17] , \OTMP[10][16] , \OTMP[10][15] , \OTMP[10][14] , 
        \OTMP[10][13] , \OTMP[10][12] , \OTMP[10][11] , \OTMP[10][10] , 
        \OTMP[10][9] , \OTMP[10][8] , \OTMP[10][7] , \OTMP[10][6] , 
        \OTMP[10][5] , \OTMP[10][4] , \OTMP[10][3] , \OTMP[10][2] , 
        \OTMP[10][1] , 1'b0}), .Ci(1'b0), .S({\PTMP[9][53] , \PTMP[9][52] , 
        \PTMP[9][51] , \PTMP[9][50] , \PTMP[9][49] , \PTMP[9][48] , 
        \PTMP[9][47] , \PTMP[9][46] , \PTMP[9][45] , \PTMP[9][44] , 
        \PTMP[9][43] , \PTMP[9][42] , \PTMP[9][41] , \PTMP[9][40] , 
        \PTMP[9][39] , \PTMP[9][38] , \PTMP[9][37] , \PTMP[9][36] , 
        \PTMP[9][35] , \PTMP[9][34] , \PTMP[9][33] , \PTMP[9][32] , 
        \PTMP[9][31] , \PTMP[9][30] , \PTMP[9][29] , \PTMP[9][28] , 
        \PTMP[9][27] , \PTMP[9][26] , \PTMP[9][25] , \PTMP[9][24] , 
        \PTMP[9][23] , \PTMP[9][22] , \PTMP[9][21] , \PTMP[9][20] , 
        \PTMP[9][19] , \PTMP[9][18] , \PTMP[9][17] , \PTMP[9][16] , 
        \PTMP[9][15] , \PTMP[9][14] , \PTMP[9][13] , \PTMP[9][12] , 
        \PTMP[9][11] , \PTMP[9][10] , \PTMP[9][9] , \PTMP[9][8] , \PTMP[9][7] , 
        \PTMP[9][6] , \PTMP[9][5] , \PTMP[9][4] , \PTMP[9][3] , \PTMP[9][2] , 
        \PTMP[9][1] , \PTMP[9][0] }) );
  RCA_NBIT56 ADDER_11 ( .A({n14, n14, \PTMP[9][53] , \PTMP[9][52] , 
        \PTMP[9][51] , \PTMP[9][50] , \PTMP[9][49] , \PTMP[9][48] , 
        \PTMP[9][47] , \PTMP[9][46] , \PTMP[9][45] , \PTMP[9][44] , 
        \PTMP[9][43] , \PTMP[9][42] , \PTMP[9][41] , \PTMP[9][40] , 
        \PTMP[9][39] , \PTMP[9][38] , \PTMP[9][37] , \PTMP[9][36] , 
        \PTMP[9][35] , \PTMP[9][34] , \PTMP[9][33] , \PTMP[9][32] , 
        \PTMP[9][31] , \PTMP[9][30] , \PTMP[9][29] , \PTMP[9][28] , 
        \PTMP[9][27] , \PTMP[9][26] , \PTMP[9][25] , \PTMP[9][24] , 
        \PTMP[9][23] , \PTMP[9][22] , \PTMP[9][21] , \PTMP[9][20] , 
        \PTMP[9][19] , \PTMP[9][18] , \PTMP[9][17] , \PTMP[9][16] , 
        \PTMP[9][15] , \PTMP[9][14] , \PTMP[9][13] , \PTMP[9][12] , 
        \PTMP[9][11] , \PTMP[9][10] , \PTMP[9][9] , \PTMP[9][8] , \PTMP[9][7] , 
        \PTMP[9][6] , \PTMP[9][5] , \PTMP[9][4] , \PTMP[9][3] , \PTMP[9][2] , 
        \PTMP[9][1] , \PTMP[9][0] }), .B({\OTMP[11][55] , \OTMP[11][54] , 
        \OTMP[11][53] , \OTMP[11][52] , \OTMP[11][51] , \OTMP[11][50] , 
        \OTMP[11][49] , \OTMP[11][48] , \OTMP[11][47] , \OTMP[11][46] , 
        \OTMP[11][45] , \OTMP[11][44] , \OTMP[11][43] , \OTMP[11][42] , 
        \OTMP[11][41] , \OTMP[11][40] , \OTMP[11][39] , \OTMP[11][38] , 
        \OTMP[11][37] , \OTMP[11][36] , \OTMP[11][35] , \OTMP[11][34] , 
        \OTMP[11][33] , \OTMP[11][32] , \OTMP[11][31] , \OTMP[11][30] , 
        \OTMP[11][29] , \OTMP[11][28] , \OTMP[11][27] , \OTMP[11][26] , 
        \OTMP[11][25] , \OTMP[11][24] , \OTMP[11][23] , \OTMP[11][22] , 
        \OTMP[11][21] , \OTMP[11][20] , \OTMP[11][19] , \OTMP[11][18] , 
        \OTMP[11][17] , \OTMP[11][16] , \OTMP[11][15] , \OTMP[11][14] , 
        \OTMP[11][13] , \OTMP[11][12] , \OTMP[11][11] , \OTMP[11][10] , 
        \OTMP[11][9] , \OTMP[11][8] , \OTMP[11][7] , \OTMP[11][6] , 
        \OTMP[11][5] , \OTMP[11][4] , \OTMP[11][3] , \OTMP[11][2] , 
        \OTMP[11][1] , 1'b0}), .Ci(1'b0), .S({\PTMP[10][55] , \PTMP[10][54] , 
        \PTMP[10][53] , \PTMP[10][52] , \PTMP[10][51] , \PTMP[10][50] , 
        \PTMP[10][49] , \PTMP[10][48] , \PTMP[10][47] , \PTMP[10][46] , 
        \PTMP[10][45] , \PTMP[10][44] , \PTMP[10][43] , \PTMP[10][42] , 
        \PTMP[10][41] , \PTMP[10][40] , \PTMP[10][39] , \PTMP[10][38] , 
        \PTMP[10][37] , \PTMP[10][36] , \PTMP[10][35] , \PTMP[10][34] , 
        \PTMP[10][33] , \PTMP[10][32] , \PTMP[10][31] , \PTMP[10][30] , 
        \PTMP[10][29] , \PTMP[10][28] , \PTMP[10][27] , \PTMP[10][26] , 
        \PTMP[10][25] , \PTMP[10][24] , \PTMP[10][23] , \PTMP[10][22] , 
        \PTMP[10][21] , \PTMP[10][20] , \PTMP[10][19] , \PTMP[10][18] , 
        \PTMP[10][17] , \PTMP[10][16] , \PTMP[10][15] , \PTMP[10][14] , 
        \PTMP[10][13] , \PTMP[10][12] , \PTMP[10][11] , \PTMP[10][10] , 
        \PTMP[10][9] , \PTMP[10][8] , \PTMP[10][7] , \PTMP[10][6] , 
        \PTMP[10][5] , \PTMP[10][4] , \PTMP[10][3] , \PTMP[10][2] , 
        \PTMP[10][1] , \PTMP[10][0] }) );
  RCA_NBIT58 ADDER_12 ( .A({n19, n19, \PTMP[10][55] , \PTMP[10][54] , 
        \PTMP[10][53] , \PTMP[10][52] , \PTMP[10][51] , \PTMP[10][50] , 
        \PTMP[10][49] , \PTMP[10][48] , \PTMP[10][47] , \PTMP[10][46] , 
        \PTMP[10][45] , \PTMP[10][44] , \PTMP[10][43] , \PTMP[10][42] , 
        \PTMP[10][41] , \PTMP[10][40] , \PTMP[10][39] , \PTMP[10][38] , 
        \PTMP[10][37] , \PTMP[10][36] , \PTMP[10][35] , \PTMP[10][34] , 
        \PTMP[10][33] , \PTMP[10][32] , \PTMP[10][31] , \PTMP[10][30] , 
        \PTMP[10][29] , \PTMP[10][28] , \PTMP[10][27] , \PTMP[10][26] , 
        \PTMP[10][25] , \PTMP[10][24] , \PTMP[10][23] , \PTMP[10][22] , 
        \PTMP[10][21] , \PTMP[10][20] , \PTMP[10][19] , \PTMP[10][18] , 
        \PTMP[10][17] , \PTMP[10][16] , \PTMP[10][15] , \PTMP[10][14] , 
        \PTMP[10][13] , \PTMP[10][12] , \PTMP[10][11] , \PTMP[10][10] , 
        \PTMP[10][9] , \PTMP[10][8] , \PTMP[10][7] , \PTMP[10][6] , 
        \PTMP[10][5] , \PTMP[10][4] , \PTMP[10][3] , \PTMP[10][2] , 
        \PTMP[10][1] , \PTMP[10][0] }), .B({\OTMP[12][57] , \OTMP[12][56] , 
        \OTMP[12][55] , \OTMP[12][54] , \OTMP[12][53] , \OTMP[12][52] , 
        \OTMP[12][51] , \OTMP[12][50] , \OTMP[12][49] , \OTMP[12][48] , 
        \OTMP[12][47] , \OTMP[12][46] , \OTMP[12][45] , \OTMP[12][44] , 
        \OTMP[12][43] , \OTMP[12][42] , \OTMP[12][41] , \OTMP[12][40] , 
        \OTMP[12][39] , \OTMP[12][38] , \OTMP[12][37] , \OTMP[12][36] , 
        \OTMP[12][35] , \OTMP[12][34] , \OTMP[12][33] , \OTMP[12][32] , 
        \OTMP[12][31] , \OTMP[12][30] , \OTMP[12][29] , \OTMP[12][28] , 
        \OTMP[12][27] , \OTMP[12][26] , \OTMP[12][25] , \OTMP[12][24] , 
        \OTMP[12][23] , \OTMP[12][22] , \OTMP[12][21] , \OTMP[12][20] , 
        \OTMP[12][19] , \OTMP[12][18] , \OTMP[12][17] , \OTMP[12][16] , 
        \OTMP[12][15] , \OTMP[12][14] , \OTMP[12][13] , \OTMP[12][12] , 
        \OTMP[12][11] , \OTMP[12][10] , \OTMP[12][9] , \OTMP[12][8] , 
        \OTMP[12][7] , \OTMP[12][6] , \OTMP[12][5] , \OTMP[12][4] , 
        \OTMP[12][3] , \OTMP[12][2] , \OTMP[12][1] , 1'b0}), .Ci(1'b0), .S({
        \PTMP[11][57] , \PTMP[11][56] , \PTMP[11][55] , \PTMP[11][54] , 
        \PTMP[11][53] , \PTMP[11][52] , \PTMP[11][51] , \PTMP[11][50] , 
        \PTMP[11][49] , \PTMP[11][48] , \PTMP[11][47] , \PTMP[11][46] , 
        \PTMP[11][45] , \PTMP[11][44] , \PTMP[11][43] , \PTMP[11][42] , 
        \PTMP[11][41] , \PTMP[11][40] , \PTMP[11][39] , \PTMP[11][38] , 
        \PTMP[11][37] , \PTMP[11][36] , \PTMP[11][35] , \PTMP[11][34] , 
        \PTMP[11][33] , \PTMP[11][32] , \PTMP[11][31] , \PTMP[11][30] , 
        \PTMP[11][29] , \PTMP[11][28] , \PTMP[11][27] , \PTMP[11][26] , 
        \PTMP[11][25] , \PTMP[11][24] , \PTMP[11][23] , \PTMP[11][22] , 
        \PTMP[11][21] , \PTMP[11][20] , \PTMP[11][19] , \PTMP[11][18] , 
        \PTMP[11][17] , \PTMP[11][16] , \PTMP[11][15] , \PTMP[11][14] , 
        \PTMP[11][13] , \PTMP[11][12] , \PTMP[11][11] , \PTMP[11][10] , 
        \PTMP[11][9] , \PTMP[11][8] , \PTMP[11][7] , \PTMP[11][6] , 
        \PTMP[11][5] , \PTMP[11][4] , \PTMP[11][3] , \PTMP[11][2] , 
        \PTMP[11][1] , \PTMP[11][0] }) );
  RCA_NBIT60 ADDER_13 ( .A({n22, n22, \PTMP[11][57] , \PTMP[11][56] , 
        \PTMP[11][55] , \PTMP[11][54] , \PTMP[11][53] , \PTMP[11][52] , 
        \PTMP[11][51] , \PTMP[11][50] , \PTMP[11][49] , \PTMP[11][48] , 
        \PTMP[11][47] , \PTMP[11][46] , \PTMP[11][45] , \PTMP[11][44] , 
        \PTMP[11][43] , \PTMP[11][42] , \PTMP[11][41] , \PTMP[11][40] , 
        \PTMP[11][39] , \PTMP[11][38] , \PTMP[11][37] , \PTMP[11][36] , 
        \PTMP[11][35] , \PTMP[11][34] , \PTMP[11][33] , \PTMP[11][32] , 
        \PTMP[11][31] , \PTMP[11][30] , \PTMP[11][29] , \PTMP[11][28] , 
        \PTMP[11][27] , \PTMP[11][26] , \PTMP[11][25] , \PTMP[11][24] , 
        \PTMP[11][23] , \PTMP[11][22] , \PTMP[11][21] , \PTMP[11][20] , 
        \PTMP[11][19] , \PTMP[11][18] , \PTMP[11][17] , \PTMP[11][16] , 
        \PTMP[11][15] , \PTMP[11][14] , \PTMP[11][13] , \PTMP[11][12] , 
        \PTMP[11][11] , \PTMP[11][10] , \PTMP[11][9] , \PTMP[11][8] , 
        \PTMP[11][7] , \PTMP[11][6] , \PTMP[11][5] , \PTMP[11][4] , 
        \PTMP[11][3] , \PTMP[11][2] , \PTMP[11][1] , \PTMP[11][0] }), .B({
        \OTMP[13][59] , \OTMP[13][58] , \OTMP[13][57] , \OTMP[13][56] , 
        \OTMP[13][55] , \OTMP[13][54] , \OTMP[13][53] , \OTMP[13][52] , 
        \OTMP[13][51] , \OTMP[13][50] , \OTMP[13][49] , \OTMP[13][48] , 
        \OTMP[13][47] , \OTMP[13][46] , \OTMP[13][45] , \OTMP[13][44] , 
        \OTMP[13][43] , \OTMP[13][42] , \OTMP[13][41] , \OTMP[13][40] , 
        \OTMP[13][39] , \OTMP[13][38] , \OTMP[13][37] , \OTMP[13][36] , 
        \OTMP[13][35] , \OTMP[13][34] , \OTMP[13][33] , \OTMP[13][32] , 
        \OTMP[13][31] , \OTMP[13][30] , \OTMP[13][29] , \OTMP[13][28] , 
        \OTMP[13][27] , \OTMP[13][26] , \OTMP[13][25] , \OTMP[13][24] , 
        \OTMP[13][23] , \OTMP[13][22] , \OTMP[13][21] , \OTMP[13][20] , 
        \OTMP[13][19] , \OTMP[13][18] , \OTMP[13][17] , \OTMP[13][16] , 
        \OTMP[13][15] , \OTMP[13][14] , \OTMP[13][13] , \OTMP[13][12] , 
        \OTMP[13][11] , \OTMP[13][10] , \OTMP[13][9] , \OTMP[13][8] , 
        \OTMP[13][7] , \OTMP[13][6] , \OTMP[13][5] , \OTMP[13][4] , 
        \OTMP[13][3] , \OTMP[13][2] , \OTMP[13][1] , 1'b0}), .Ci(1'b0), .S({
        \PTMP[12][59] , \PTMP[12][58] , \PTMP[12][57] , \PTMP[12][56] , 
        \PTMP[12][55] , \PTMP[12][54] , \PTMP[12][53] , \PTMP[12][52] , 
        \PTMP[12][51] , \PTMP[12][50] , \PTMP[12][49] , \PTMP[12][48] , 
        \PTMP[12][47] , \PTMP[12][46] , \PTMP[12][45] , \PTMP[12][44] , 
        \PTMP[12][43] , \PTMP[12][42] , \PTMP[12][41] , \PTMP[12][40] , 
        \PTMP[12][39] , \PTMP[12][38] , \PTMP[12][37] , \PTMP[12][36] , 
        \PTMP[12][35] , \PTMP[12][34] , \PTMP[12][33] , \PTMP[12][32] , 
        \PTMP[12][31] , \PTMP[12][30] , \PTMP[12][29] , \PTMP[12][28] , 
        \PTMP[12][27] , \PTMP[12][26] , \PTMP[12][25] , \PTMP[12][24] , 
        \PTMP[12][23] , \PTMP[12][22] , \PTMP[12][21] , \PTMP[12][20] , 
        \PTMP[12][19] , \PTMP[12][18] , \PTMP[12][17] , \PTMP[12][16] , 
        \PTMP[12][15] , \PTMP[12][14] , \PTMP[12][13] , \PTMP[12][12] , 
        \PTMP[12][11] , \PTMP[12][10] , \PTMP[12][9] , \PTMP[12][8] , 
        \PTMP[12][7] , \PTMP[12][6] , \PTMP[12][5] , \PTMP[12][4] , 
        \PTMP[12][3] , \PTMP[12][2] , \PTMP[12][1] , \PTMP[12][0] }) );
  RCA_NBIT62 ADDER_14 ( .A({n12, \PTMP[12][59] , \PTMP[12][59] , 
        \PTMP[12][58] , \PTMP[12][57] , \PTMP[12][56] , \PTMP[12][55] , 
        \PTMP[12][54] , \PTMP[12][53] , \PTMP[12][52] , \PTMP[12][51] , 
        \PTMP[12][50] , \PTMP[12][49] , \PTMP[12][48] , \PTMP[12][47] , 
        \PTMP[12][46] , \PTMP[12][45] , \PTMP[12][44] , \PTMP[12][43] , 
        \PTMP[12][42] , \PTMP[12][41] , \PTMP[12][40] , \PTMP[12][39] , 
        \PTMP[12][38] , \PTMP[12][37] , \PTMP[12][36] , \PTMP[12][35] , 
        \PTMP[12][34] , \PTMP[12][33] , \PTMP[12][32] , \PTMP[12][31] , 
        \PTMP[12][30] , \PTMP[12][29] , \PTMP[12][28] , \PTMP[12][27] , 
        \PTMP[12][26] , \PTMP[12][25] , \PTMP[12][24] , \PTMP[12][23] , 
        \PTMP[12][22] , \PTMP[12][21] , \PTMP[12][20] , \PTMP[12][19] , 
        \PTMP[12][18] , \PTMP[12][17] , \PTMP[12][16] , \PTMP[12][15] , 
        \PTMP[12][14] , \PTMP[12][13] , \PTMP[12][12] , \PTMP[12][11] , 
        \PTMP[12][10] , \PTMP[12][9] , \PTMP[12][8] , \PTMP[12][7] , 
        \PTMP[12][6] , \PTMP[12][5] , \PTMP[12][4] , \PTMP[12][3] , 
        \PTMP[12][2] , \PTMP[12][1] , \PTMP[12][0] }), .B({\OTMP[14][61] , 
        \OTMP[14][60] , \OTMP[14][59] , \OTMP[14][58] , \OTMP[14][57] , 
        \OTMP[14][56] , \OTMP[14][55] , \OTMP[14][54] , \OTMP[14][53] , 
        \OTMP[14][52] , \OTMP[14][51] , \OTMP[14][50] , \OTMP[14][49] , 
        \OTMP[14][48] , \OTMP[14][47] , \OTMP[14][46] , \OTMP[14][45] , 
        \OTMP[14][44] , \OTMP[14][43] , \OTMP[14][42] , \OTMP[14][41] , 
        \OTMP[14][40] , \OTMP[14][39] , \OTMP[14][38] , \OTMP[14][37] , 
        \OTMP[14][36] , \OTMP[14][35] , \OTMP[14][34] , \OTMP[14][33] , 
        \OTMP[14][32] , \OTMP[14][31] , \OTMP[14][30] , \OTMP[14][29] , 
        \OTMP[14][28] , \OTMP[14][27] , \OTMP[14][26] , \OTMP[14][25] , 
        \OTMP[14][24] , \OTMP[14][23] , \OTMP[14][22] , \OTMP[14][21] , 
        \OTMP[14][20] , \OTMP[14][19] , \OTMP[14][18] , \OTMP[14][17] , 
        \OTMP[14][16] , \OTMP[14][15] , \OTMP[14][14] , \OTMP[14][13] , 
        \OTMP[14][12] , \OTMP[14][11] , \OTMP[14][10] , \OTMP[14][9] , 
        \OTMP[14][8] , \OTMP[14][7] , \OTMP[14][6] , \OTMP[14][5] , 
        \OTMP[14][4] , \OTMP[14][3] , \OTMP[14][2] , \OTMP[14][1] , 1'b0}), 
        .Ci(1'b0), .S({\PTMP[13][61] , \PTMP[13][60] , \PTMP[13][59] , 
        \PTMP[13][58] , \PTMP[13][57] , \PTMP[13][56] , \PTMP[13][55] , 
        \PTMP[13][54] , \PTMP[13][53] , \PTMP[13][52] , \PTMP[13][51] , 
        \PTMP[13][50] , \PTMP[13][49] , \PTMP[13][48] , \PTMP[13][47] , 
        \PTMP[13][46] , \PTMP[13][45] , \PTMP[13][44] , \PTMP[13][43] , 
        \PTMP[13][42] , \PTMP[13][41] , \PTMP[13][40] , \PTMP[13][39] , 
        \PTMP[13][38] , \PTMP[13][37] , \PTMP[13][36] , \PTMP[13][35] , 
        \PTMP[13][34] , \PTMP[13][33] , \PTMP[13][32] , \PTMP[13][31] , 
        \PTMP[13][30] , \PTMP[13][29] , \PTMP[13][28] , \PTMP[13][27] , 
        \PTMP[13][26] , \PTMP[13][25] , \PTMP[13][24] , \PTMP[13][23] , 
        \PTMP[13][22] , \PTMP[13][21] , \PTMP[13][20] , \PTMP[13][19] , 
        \PTMP[13][18] , \PTMP[13][17] , \PTMP[13][16] , \PTMP[13][15] , 
        \PTMP[13][14] , \PTMP[13][13] , \PTMP[13][12] , \PTMP[13][11] , 
        \PTMP[13][10] , \PTMP[13][9] , \PTMP[13][8] , \PTMP[13][7] , 
        \PTMP[13][6] , \PTMP[13][5] , \PTMP[13][4] , \PTMP[13][3] , 
        \PTMP[13][2] , \PTMP[13][1] , \PTMP[13][0] }) );
  RCA_NBIT64 ADDER_15 ( .A({\PTMP[13][61] , \PTMP[13][61] , \PTMP[13][61] , 
        \PTMP[13][60] , \PTMP[13][59] , \PTMP[13][58] , \PTMP[13][57] , 
        \PTMP[13][56] , \PTMP[13][55] , \PTMP[13][54] , \PTMP[13][53] , 
        \PTMP[13][52] , \PTMP[13][51] , \PTMP[13][50] , \PTMP[13][49] , 
        \PTMP[13][48] , \PTMP[13][47] , \PTMP[13][46] , \PTMP[13][45] , 
        \PTMP[13][44] , \PTMP[13][43] , \PTMP[13][42] , \PTMP[13][41] , 
        \PTMP[13][40] , \PTMP[13][39] , \PTMP[13][38] , \PTMP[13][37] , 
        \PTMP[13][36] , \PTMP[13][35] , \PTMP[13][34] , \PTMP[13][33] , 
        \PTMP[13][32] , \PTMP[13][31] , \PTMP[13][30] , \PTMP[13][29] , 
        \PTMP[13][28] , \PTMP[13][27] , \PTMP[13][26] , \PTMP[13][25] , 
        \PTMP[13][24] , \PTMP[13][23] , \PTMP[13][22] , \PTMP[13][21] , 
        \PTMP[13][20] , \PTMP[13][19] , \PTMP[13][18] , \PTMP[13][17] , 
        \PTMP[13][16] , \PTMP[13][15] , \PTMP[13][14] , \PTMP[13][13] , 
        \PTMP[13][12] , \PTMP[13][11] , \PTMP[13][10] , \PTMP[13][9] , 
        \PTMP[13][8] , \PTMP[13][7] , \PTMP[13][6] , \PTMP[13][5] , 
        \PTMP[13][4] , \PTMP[13][3] , \PTMP[13][2] , \PTMP[13][1] , 
        \PTMP[13][0] }), .B({\OTMP[15][63] , \OTMP[15][62] , \OTMP[15][61] , 
        \OTMP[15][60] , \OTMP[15][59] , \OTMP[15][58] , \OTMP[15][57] , 
        \OTMP[15][56] , \OTMP[15][55] , \OTMP[15][54] , \OTMP[15][53] , 
        \OTMP[15][52] , \OTMP[15][51] , \OTMP[15][50] , \OTMP[15][49] , 
        \OTMP[15][48] , \OTMP[15][47] , \OTMP[15][46] , \OTMP[15][45] , 
        \OTMP[15][44] , \OTMP[15][43] , \OTMP[15][42] , \OTMP[15][41] , 
        \OTMP[15][40] , \OTMP[15][39] , \OTMP[15][38] , \OTMP[15][37] , 
        \OTMP[15][36] , \OTMP[15][35] , \OTMP[15][34] , \OTMP[15][33] , 
        \OTMP[15][32] , \OTMP[15][31] , \OTMP[15][30] , \OTMP[15][29] , 
        \OTMP[15][28] , \OTMP[15][27] , \OTMP[15][26] , \OTMP[15][25] , 
        \OTMP[15][24] , \OTMP[15][23] , \OTMP[15][22] , \OTMP[15][21] , 
        \OTMP[15][20] , \OTMP[15][19] , \OTMP[15][18] , \OTMP[15][17] , 
        \OTMP[15][16] , \OTMP[15][15] , \OTMP[15][14] , \OTMP[15][13] , 
        \OTMP[15][12] , \OTMP[15][11] , \OTMP[15][10] , \OTMP[15][9] , 
        \OTMP[15][8] , \OTMP[15][7] , \OTMP[15][6] , \OTMP[15][5] , 
        \OTMP[15][4] , \OTMP[15][3] , \OTMP[15][2] , \OTMP[15][1] , 1'b0}), 
        .Ci(1'b0), .S(S) );
  BOOTHMUL_NBIT32_DW01_sub_0 sub_101 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF({A_n_65, A_n}) );
  CLKBUF_X1 U80 ( .A(n15), .Z(n6) );
  BUF_X1 U81 ( .A(\PTMP[5][45] ), .Z(n15) );
  BUF_X1 U82 ( .A(\PTMP[9][53] ), .Z(n14) );
  BUF_X1 U83 ( .A(\PTMP[4][43] ), .Z(n13) );
  BUF_X1 U84 ( .A(\PTMP[2][39] ), .Z(n7) );
  BUF_X2 U85 ( .A(n8), .Z(n16) );
  CLKBUF_X1 U86 ( .A(\PTMP[8][51] ), .Z(n18) );
  CLKBUF_X1 U87 ( .A(\PTMP[7][49] ), .Z(n8) );
  CLKBUF_X1 U88 ( .A(\PTMP[6][47] ), .Z(n17) );
  BUF_X1 U89 ( .A(B[2]), .Z(n9) );
  BUF_X1 U90 ( .A(B[2]), .Z(n10) );
  BUF_X1 U91 ( .A(A[1]), .Z(n11) );
  CLKBUF_X1 U92 ( .A(\PTMP[12][59] ), .Z(n12) );
  CLKBUF_X1 U93 ( .A(\PTMP[10][55] ), .Z(n19) );
  INV_X1 U94 ( .A(n17), .ZN(n20) );
  INV_X1 U95 ( .A(n20), .ZN(n21) );
  CLKBUF_X1 U96 ( .A(\PTMP[11][57] ), .Z(n22) );
endmodule

