
module BOOTHENC_NBIT64_i0 ( A, A_n, A_ns, A_s, B, O, A_so, A_nso );
  input [63:0] A;
  input [63:0] A_n;
  input [63:0] A_ns;
  input [63:0] A_s;
  input [63:0] B;
  output [63:0] O;
  output [63:0] A_so;
  output [63:0] A_nso;
  wire   \A_s[62] , \A_s[61] , \A_s[60] , \A_s[59] , \A_s[58] , \A_s[57] ,
         \A_s[56] , \A_s[55] , \A_s[54] , \A_s[53] , \A_s[52] , \A_s[51] ,
         \A_s[50] , \A_s[49] , \A_s[48] , \A_s[47] , \A_s[46] , \A_s[45] ,
         \A_s[44] , \A_s[43] , \A_s[42] , \A_s[41] , \A_s[40] , \A_s[39] ,
         \A_s[38] , \A_s[37] , \A_s[36] , \A_s[35] , \A_s[34] , \A_s[33] ,
         \A_s[32] , \A_s[31] , \A_s[30] , \A_s[29] , \A_s[28] , \A_s[27] ,
         \A_s[26] , \A_s[25] , \A_s[24] , \A_s[23] , \A_s[22] , \A_s[21] ,
         \A_s[20] , \A_s[19] , \A_s[18] , \A_s[17] , \A_s[16] , \A_s[15] ,
         \A_s[14] , \A_s[13] , \A_s[12] , \A_s[11] , \A_s[10] , \A_s[9] ,
         \A_s[8] , \A_s[7] , \A_s[6] , \A_s[5] , \A_s[4] , \A_s[3] , \A_s[2] ,
         \A_s[1] , \A_s[0] , n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399;
  assign A_nso[0] = 1'b0;
  assign A_so[0] = 1'b0;
  assign A_nso[63] = \A_s[62] ;
  assign A_so[63] = \A_s[62] ;
  assign \A_s[62]  = A_s[62];
  assign A_nso[62] = \A_s[61] ;
  assign A_so[62] = \A_s[61] ;
  assign \A_s[61]  = A_s[61];
  assign A_nso[61] = \A_s[60] ;
  assign A_so[61] = \A_s[60] ;
  assign \A_s[60]  = A_s[60];
  assign A_nso[60] = \A_s[59] ;
  assign A_so[60] = \A_s[59] ;
  assign \A_s[59]  = A_s[59];
  assign A_nso[59] = \A_s[58] ;
  assign A_so[59] = \A_s[58] ;
  assign \A_s[58]  = A_s[58];
  assign A_nso[58] = \A_s[57] ;
  assign A_so[58] = \A_s[57] ;
  assign \A_s[57]  = A_s[57];
  assign A_nso[57] = \A_s[56] ;
  assign A_so[57] = \A_s[56] ;
  assign \A_s[56]  = A_s[56];
  assign A_nso[56] = \A_s[55] ;
  assign A_so[56] = \A_s[55] ;
  assign \A_s[55]  = A_s[55];
  assign A_nso[55] = \A_s[54] ;
  assign A_so[55] = \A_s[54] ;
  assign \A_s[54]  = A_s[54];
  assign A_nso[54] = \A_s[53] ;
  assign A_so[54] = \A_s[53] ;
  assign \A_s[53]  = A_s[53];
  assign A_nso[53] = \A_s[52] ;
  assign A_so[53] = \A_s[52] ;
  assign \A_s[52]  = A_s[52];
  assign A_nso[52] = \A_s[51] ;
  assign A_so[52] = \A_s[51] ;
  assign \A_s[51]  = A_s[51];
  assign A_nso[51] = \A_s[50] ;
  assign A_so[51] = \A_s[50] ;
  assign \A_s[50]  = A_s[50];
  assign A_nso[50] = \A_s[49] ;
  assign A_so[50] = \A_s[49] ;
  assign \A_s[49]  = A_s[49];
  assign A_nso[49] = \A_s[48] ;
  assign A_so[49] = \A_s[48] ;
  assign \A_s[48]  = A_s[48];
  assign A_nso[48] = \A_s[47] ;
  assign A_so[48] = \A_s[47] ;
  assign \A_s[47]  = A_s[47];
  assign A_nso[47] = \A_s[46] ;
  assign A_so[47] = \A_s[46] ;
  assign \A_s[46]  = A_s[46];
  assign A_nso[46] = \A_s[45] ;
  assign A_so[46] = \A_s[45] ;
  assign \A_s[45]  = A_s[45];
  assign A_nso[45] = \A_s[44] ;
  assign A_so[45] = \A_s[44] ;
  assign \A_s[44]  = A_s[44];
  assign A_nso[44] = \A_s[43] ;
  assign A_so[44] = \A_s[43] ;
  assign \A_s[43]  = A_s[43];
  assign A_nso[43] = \A_s[42] ;
  assign A_so[43] = \A_s[42] ;
  assign \A_s[42]  = A_s[42];
  assign A_nso[42] = \A_s[41] ;
  assign A_so[42] = \A_s[41] ;
  assign \A_s[41]  = A_s[41];
  assign A_nso[41] = \A_s[40] ;
  assign A_so[41] = \A_s[40] ;
  assign \A_s[40]  = A_s[40];
  assign A_nso[40] = \A_s[39] ;
  assign A_so[40] = \A_s[39] ;
  assign \A_s[39]  = A_s[39];
  assign A_nso[39] = \A_s[38] ;
  assign A_so[39] = \A_s[38] ;
  assign \A_s[38]  = A_s[38];
  assign A_nso[38] = \A_s[37] ;
  assign A_so[38] = \A_s[37] ;
  assign \A_s[37]  = A_s[37];
  assign A_nso[37] = \A_s[36] ;
  assign A_so[37] = \A_s[36] ;
  assign \A_s[36]  = A_s[36];
  assign A_nso[36] = \A_s[35] ;
  assign A_so[36] = \A_s[35] ;
  assign \A_s[35]  = A_s[35];
  assign A_nso[35] = \A_s[34] ;
  assign A_so[35] = \A_s[34] ;
  assign \A_s[34]  = A_s[34];
  assign A_nso[34] = \A_s[33] ;
  assign A_so[34] = \A_s[33] ;
  assign \A_s[33]  = A_s[33];
  assign A_nso[33] = \A_s[32] ;
  assign A_so[33] = \A_s[32] ;
  assign \A_s[32]  = A_s[32];
  assign A_nso[32] = \A_s[31] ;
  assign A_so[32] = \A_s[31] ;
  assign \A_s[31]  = A_s[31];
  assign A_nso[31] = \A_s[30] ;
  assign A_so[31] = \A_s[30] ;
  assign \A_s[30]  = A_s[30];
  assign A_nso[30] = \A_s[29] ;
  assign A_so[30] = \A_s[29] ;
  assign \A_s[29]  = A_s[29];
  assign A_nso[29] = \A_s[28] ;
  assign A_so[29] = \A_s[28] ;
  assign \A_s[28]  = A_s[28];
  assign A_nso[28] = \A_s[27] ;
  assign A_so[28] = \A_s[27] ;
  assign \A_s[27]  = A_s[27];
  assign A_nso[27] = \A_s[26] ;
  assign A_so[27] = \A_s[26] ;
  assign \A_s[26]  = A_s[26];
  assign A_nso[26] = \A_s[25] ;
  assign A_so[26] = \A_s[25] ;
  assign \A_s[25]  = A_s[25];
  assign A_nso[25] = \A_s[24] ;
  assign A_so[25] = \A_s[24] ;
  assign \A_s[24]  = A_s[24];
  assign A_nso[24] = \A_s[23] ;
  assign A_so[24] = \A_s[23] ;
  assign \A_s[23]  = A_s[23];
  assign A_nso[23] = \A_s[22] ;
  assign A_so[23] = \A_s[22] ;
  assign \A_s[22]  = A_s[22];
  assign A_nso[22] = \A_s[21] ;
  assign A_so[22] = \A_s[21] ;
  assign \A_s[21]  = A_s[21];
  assign A_nso[21] = \A_s[20] ;
  assign A_so[21] = \A_s[20] ;
  assign \A_s[20]  = A_s[20];
  assign A_nso[20] = \A_s[19] ;
  assign A_so[20] = \A_s[19] ;
  assign \A_s[19]  = A_s[19];
  assign A_nso[19] = \A_s[18] ;
  assign A_so[19] = \A_s[18] ;
  assign \A_s[18]  = A_s[18];
  assign A_nso[18] = \A_s[17] ;
  assign A_so[18] = \A_s[17] ;
  assign \A_s[17]  = A_s[17];
  assign A_nso[17] = \A_s[16] ;
  assign A_so[17] = \A_s[16] ;
  assign \A_s[16]  = A_s[16];
  assign A_nso[16] = \A_s[15] ;
  assign A_so[16] = \A_s[15] ;
  assign \A_s[15]  = A_s[15];
  assign A_nso[15] = \A_s[14] ;
  assign A_so[15] = \A_s[14] ;
  assign \A_s[14]  = A_s[14];
  assign A_nso[14] = \A_s[13] ;
  assign A_so[14] = \A_s[13] ;
  assign \A_s[13]  = A_s[13];
  assign A_nso[13] = \A_s[12] ;
  assign A_so[13] = \A_s[12] ;
  assign \A_s[12]  = A_s[12];
  assign A_nso[12] = \A_s[11] ;
  assign A_so[12] = \A_s[11] ;
  assign \A_s[11]  = A_s[11];
  assign A_nso[11] = \A_s[10] ;
  assign A_so[11] = \A_s[10] ;
  assign \A_s[10]  = A_s[10];
  assign A_nso[10] = \A_s[9] ;
  assign A_so[10] = \A_s[9] ;
  assign \A_s[9]  = A_s[9];
  assign A_nso[9] = \A_s[8] ;
  assign A_so[9] = \A_s[8] ;
  assign \A_s[8]  = A_s[8];
  assign A_nso[8] = \A_s[7] ;
  assign A_so[8] = \A_s[7] ;
  assign \A_s[7]  = A_s[7];
  assign A_nso[7] = \A_s[6] ;
  assign A_so[7] = \A_s[6] ;
  assign \A_s[6]  = A_s[6];
  assign A_nso[6] = \A_s[5] ;
  assign A_so[6] = \A_s[5] ;
  assign \A_s[5]  = A_s[5];
  assign A_nso[5] = \A_s[4] ;
  assign A_so[5] = \A_s[4] ;
  assign \A_s[4]  = A_s[4];
  assign A_nso[4] = \A_s[3] ;
  assign A_so[4] = \A_s[3] ;
  assign \A_s[3]  = A_s[3];
  assign A_nso[3] = \A_s[2] ;
  assign A_so[3] = \A_s[2] ;
  assign \A_s[2]  = A_s[2];
  assign A_nso[2] = \A_s[1] ;
  assign A_so[2] = \A_s[1] ;
  assign \A_s[1]  = A_s[1];
  assign A_nso[1] = \A_s[0] ;
  assign A_so[1] = \A_s[0] ;
  assign \A_s[0]  = A_s[0];

  INV_X4 U3 ( .A(n280), .ZN(n272) );
  OR2_X4 U4 ( .A1(n398), .A2(B[0]), .ZN(n267) );
  NAND2_X4 U5 ( .A1(B[0]), .A2(n280), .ZN(n269) );
  OAI221_X1 U6 ( .B1(n267), .B2(n268), .C1(n269), .C2(n270), .A(n271), .ZN(
        O[9]) );
  NAND2_X1 U7 ( .A1(\A_s[9] ), .A2(n272), .ZN(n271) );
  OAI221_X1 U8 ( .B1(n267), .B2(n273), .C1(n268), .C2(n269), .A(n274), .ZN(
        O[8]) );
  NAND2_X1 U9 ( .A1(\A_s[8] ), .A2(n272), .ZN(n274) );
  INV_X1 U10 ( .A(A_ns[8]), .ZN(n268) );
  OAI221_X1 U11 ( .B1(n267), .B2(n275), .C1(n269), .C2(n273), .A(n276), .ZN(
        O[7]) );
  NAND2_X1 U12 ( .A1(\A_s[7] ), .A2(n272), .ZN(n276) );
  INV_X1 U13 ( .A(A_ns[7]), .ZN(n273) );
  OAI221_X1 U14 ( .B1(n267), .B2(n277), .C1(n269), .C2(n275), .A(n278), .ZN(
        O[6]) );
  NAND2_X1 U15 ( .A1(\A_s[6] ), .A2(n272), .ZN(n278) );
  INV_X1 U16 ( .A(A_ns[6]), .ZN(n275) );
  OAI222_X1 U17 ( .A1(n279), .A2(n280), .B1(n281), .B2(n267), .C1(n282), .C2(
        n269), .ZN(O[63]) );
  INV_X1 U18 ( .A(A_ns[63]), .ZN(n282) );
  INV_X1 U19 ( .A(A_s[63]), .ZN(n279) );
  OAI221_X1 U20 ( .B1(n267), .B2(n283), .C1(n269), .C2(n281), .A(n284), .ZN(
        O[62]) );
  NAND2_X1 U21 ( .A1(\A_s[62] ), .A2(n272), .ZN(n284) );
  INV_X1 U22 ( .A(A_ns[62]), .ZN(n281) );
  OAI221_X1 U23 ( .B1(n267), .B2(n285), .C1(n269), .C2(n283), .A(n286), .ZN(
        O[61]) );
  NAND2_X1 U24 ( .A1(\A_s[61] ), .A2(n272), .ZN(n286) );
  INV_X1 U25 ( .A(A_ns[61]), .ZN(n283) );
  OAI221_X1 U26 ( .B1(n267), .B2(n287), .C1(n269), .C2(n285), .A(n288), .ZN(
        O[60]) );
  NAND2_X1 U27 ( .A1(\A_s[60] ), .A2(n272), .ZN(n288) );
  INV_X1 U28 ( .A(A_ns[60]), .ZN(n285) );
  OAI221_X1 U29 ( .B1(n267), .B2(n289), .C1(n269), .C2(n277), .A(n290), .ZN(
        O[5]) );
  NAND2_X1 U30 ( .A1(\A_s[5] ), .A2(n272), .ZN(n290) );
  INV_X1 U31 ( .A(A_ns[5]), .ZN(n277) );
  OAI221_X1 U32 ( .B1(n267), .B2(n291), .C1(n269), .C2(n287), .A(n292), .ZN(
        O[59]) );
  NAND2_X1 U33 ( .A1(\A_s[59] ), .A2(n272), .ZN(n292) );
  INV_X1 U34 ( .A(A_ns[59]), .ZN(n287) );
  OAI221_X1 U35 ( .B1(n267), .B2(n293), .C1(n269), .C2(n291), .A(n294), .ZN(
        O[58]) );
  NAND2_X1 U36 ( .A1(\A_s[58] ), .A2(n272), .ZN(n294) );
  INV_X1 U37 ( .A(A_ns[58]), .ZN(n291) );
  OAI221_X1 U38 ( .B1(n267), .B2(n295), .C1(n269), .C2(n293), .A(n296), .ZN(
        O[57]) );
  NAND2_X1 U39 ( .A1(\A_s[57] ), .A2(n272), .ZN(n296) );
  INV_X1 U40 ( .A(A_ns[57]), .ZN(n293) );
  OAI221_X1 U41 ( .B1(n267), .B2(n297), .C1(n269), .C2(n295), .A(n298), .ZN(
        O[56]) );
  NAND2_X1 U42 ( .A1(\A_s[56] ), .A2(n272), .ZN(n298) );
  INV_X1 U43 ( .A(A_ns[56]), .ZN(n295) );
  OAI221_X1 U44 ( .B1(n267), .B2(n299), .C1(n269), .C2(n297), .A(n300), .ZN(
        O[55]) );
  NAND2_X1 U45 ( .A1(\A_s[55] ), .A2(n272), .ZN(n300) );
  INV_X1 U46 ( .A(A_ns[55]), .ZN(n297) );
  OAI221_X1 U47 ( .B1(n267), .B2(n301), .C1(n269), .C2(n299), .A(n302), .ZN(
        O[54]) );
  NAND2_X1 U48 ( .A1(\A_s[54] ), .A2(n272), .ZN(n302) );
  INV_X1 U49 ( .A(A_ns[54]), .ZN(n299) );
  OAI221_X1 U50 ( .B1(n267), .B2(n303), .C1(n269), .C2(n301), .A(n304), .ZN(
        O[53]) );
  NAND2_X1 U51 ( .A1(\A_s[53] ), .A2(n272), .ZN(n304) );
  INV_X1 U52 ( .A(A_ns[53]), .ZN(n301) );
  OAI221_X1 U53 ( .B1(n267), .B2(n305), .C1(n269), .C2(n303), .A(n306), .ZN(
        O[52]) );
  NAND2_X1 U54 ( .A1(\A_s[52] ), .A2(n272), .ZN(n306) );
  INV_X1 U55 ( .A(A_ns[52]), .ZN(n303) );
  OAI221_X1 U56 ( .B1(n267), .B2(n307), .C1(n269), .C2(n305), .A(n308), .ZN(
        O[51]) );
  NAND2_X1 U57 ( .A1(\A_s[51] ), .A2(n272), .ZN(n308) );
  INV_X1 U58 ( .A(A_ns[51]), .ZN(n305) );
  OAI221_X1 U59 ( .B1(n267), .B2(n309), .C1(n269), .C2(n307), .A(n310), .ZN(
        O[50]) );
  NAND2_X1 U60 ( .A1(\A_s[50] ), .A2(n272), .ZN(n310) );
  INV_X1 U61 ( .A(A_ns[50]), .ZN(n307) );
  OAI221_X1 U62 ( .B1(n267), .B2(n311), .C1(n269), .C2(n289), .A(n312), .ZN(
        O[4]) );
  NAND2_X1 U63 ( .A1(\A_s[4] ), .A2(n272), .ZN(n312) );
  INV_X1 U64 ( .A(A_ns[4]), .ZN(n289) );
  OAI221_X1 U65 ( .B1(n267), .B2(n313), .C1(n269), .C2(n309), .A(n314), .ZN(
        O[49]) );
  NAND2_X1 U66 ( .A1(\A_s[49] ), .A2(n272), .ZN(n314) );
  INV_X1 U67 ( .A(A_ns[49]), .ZN(n309) );
  OAI221_X1 U68 ( .B1(n267), .B2(n315), .C1(n269), .C2(n313), .A(n316), .ZN(
        O[48]) );
  NAND2_X1 U69 ( .A1(\A_s[48] ), .A2(n272), .ZN(n316) );
  INV_X1 U70 ( .A(A_ns[48]), .ZN(n313) );
  OAI221_X1 U71 ( .B1(n267), .B2(n317), .C1(n269), .C2(n315), .A(n318), .ZN(
        O[47]) );
  NAND2_X1 U72 ( .A1(\A_s[47] ), .A2(n272), .ZN(n318) );
  INV_X1 U73 ( .A(A_ns[47]), .ZN(n315) );
  OAI221_X1 U74 ( .B1(n267), .B2(n319), .C1(n269), .C2(n317), .A(n320), .ZN(
        O[46]) );
  NAND2_X1 U75 ( .A1(\A_s[46] ), .A2(n272), .ZN(n320) );
  INV_X1 U76 ( .A(A_ns[46]), .ZN(n317) );
  OAI221_X1 U77 ( .B1(n267), .B2(n321), .C1(n269), .C2(n319), .A(n322), .ZN(
        O[45]) );
  NAND2_X1 U78 ( .A1(\A_s[45] ), .A2(n272), .ZN(n322) );
  INV_X1 U79 ( .A(A_ns[45]), .ZN(n319) );
  OAI221_X1 U80 ( .B1(n267), .B2(n323), .C1(n269), .C2(n321), .A(n324), .ZN(
        O[44]) );
  NAND2_X1 U81 ( .A1(\A_s[44] ), .A2(n272), .ZN(n324) );
  INV_X1 U82 ( .A(A_ns[44]), .ZN(n321) );
  OAI221_X1 U83 ( .B1(n267), .B2(n325), .C1(n269), .C2(n323), .A(n326), .ZN(
        O[43]) );
  NAND2_X1 U84 ( .A1(\A_s[43] ), .A2(n272), .ZN(n326) );
  INV_X1 U85 ( .A(A_ns[43]), .ZN(n323) );
  OAI221_X1 U86 ( .B1(n267), .B2(n327), .C1(n269), .C2(n325), .A(n328), .ZN(
        O[42]) );
  NAND2_X1 U87 ( .A1(\A_s[42] ), .A2(n272), .ZN(n328) );
  INV_X1 U88 ( .A(A_ns[42]), .ZN(n325) );
  OAI221_X1 U89 ( .B1(n267), .B2(n329), .C1(n269), .C2(n327), .A(n330), .ZN(
        O[41]) );
  NAND2_X1 U90 ( .A1(\A_s[41] ), .A2(n272), .ZN(n330) );
  INV_X1 U91 ( .A(A_ns[41]), .ZN(n327) );
  OAI221_X1 U92 ( .B1(n267), .B2(n331), .C1(n269), .C2(n329), .A(n332), .ZN(
        O[40]) );
  NAND2_X1 U93 ( .A1(\A_s[40] ), .A2(n272), .ZN(n332) );
  INV_X1 U94 ( .A(A_ns[40]), .ZN(n329) );
  OAI221_X1 U95 ( .B1(n267), .B2(n333), .C1(n269), .C2(n311), .A(n334), .ZN(
        O[3]) );
  NAND2_X1 U96 ( .A1(\A_s[3] ), .A2(n272), .ZN(n334) );
  INV_X1 U97 ( .A(A_ns[3]), .ZN(n311) );
  OAI221_X1 U98 ( .B1(n267), .B2(n335), .C1(n269), .C2(n331), .A(n336), .ZN(
        O[39]) );
  NAND2_X1 U99 ( .A1(\A_s[39] ), .A2(n272), .ZN(n336) );
  INV_X1 U100 ( .A(A_ns[39]), .ZN(n331) );
  OAI221_X1 U101 ( .B1(n267), .B2(n337), .C1(n269), .C2(n335), .A(n338), .ZN(
        O[38]) );
  NAND2_X1 U102 ( .A1(\A_s[38] ), .A2(n272), .ZN(n338) );
  INV_X1 U103 ( .A(A_ns[38]), .ZN(n335) );
  OAI221_X1 U104 ( .B1(n267), .B2(n339), .C1(n269), .C2(n337), .A(n340), .ZN(
        O[37]) );
  NAND2_X1 U105 ( .A1(\A_s[37] ), .A2(n272), .ZN(n340) );
  INV_X1 U106 ( .A(A_ns[37]), .ZN(n337) );
  OAI221_X1 U107 ( .B1(n267), .B2(n341), .C1(n269), .C2(n339), .A(n342), .ZN(
        O[36]) );
  NAND2_X1 U108 ( .A1(\A_s[36] ), .A2(n272), .ZN(n342) );
  INV_X1 U109 ( .A(A_ns[36]), .ZN(n339) );
  OAI221_X1 U110 ( .B1(n267), .B2(n343), .C1(n269), .C2(n341), .A(n344), .ZN(
        O[35]) );
  NAND2_X1 U111 ( .A1(\A_s[35] ), .A2(n272), .ZN(n344) );
  INV_X1 U112 ( .A(A_ns[35]), .ZN(n341) );
  OAI221_X1 U113 ( .B1(n267), .B2(n345), .C1(n269), .C2(n343), .A(n346), .ZN(
        O[34]) );
  NAND2_X1 U114 ( .A1(\A_s[34] ), .A2(n272), .ZN(n346) );
  INV_X1 U115 ( .A(A_ns[34]), .ZN(n343) );
  OAI221_X1 U116 ( .B1(n267), .B2(n347), .C1(n269), .C2(n345), .A(n348), .ZN(
        O[33]) );
  NAND2_X1 U117 ( .A1(\A_s[33] ), .A2(n272), .ZN(n348) );
  INV_X1 U118 ( .A(A_ns[33]), .ZN(n345) );
  OAI221_X1 U119 ( .B1(n267), .B2(n349), .C1(n269), .C2(n347), .A(n350), .ZN(
        O[32]) );
  NAND2_X1 U120 ( .A1(\A_s[32] ), .A2(n272), .ZN(n350) );
  INV_X1 U121 ( .A(A_ns[32]), .ZN(n347) );
  OAI221_X1 U122 ( .B1(n267), .B2(n351), .C1(n269), .C2(n349), .A(n352), .ZN(
        O[31]) );
  NAND2_X1 U123 ( .A1(\A_s[31] ), .A2(n272), .ZN(n352) );
  INV_X1 U124 ( .A(A_ns[31]), .ZN(n349) );
  OAI221_X1 U125 ( .B1(n267), .B2(n353), .C1(n269), .C2(n351), .A(n354), .ZN(
        O[30]) );
  NAND2_X1 U126 ( .A1(\A_s[30] ), .A2(n272), .ZN(n354) );
  INV_X1 U127 ( .A(A_ns[30]), .ZN(n351) );
  OAI221_X1 U128 ( .B1(n267), .B2(n355), .C1(n269), .C2(n333), .A(n356), .ZN(
        O[2]) );
  NAND2_X1 U129 ( .A1(\A_s[2] ), .A2(n272), .ZN(n356) );
  INV_X1 U130 ( .A(A_ns[2]), .ZN(n333) );
  OAI221_X1 U131 ( .B1(n267), .B2(n357), .C1(n269), .C2(n353), .A(n358), .ZN(
        O[29]) );
  NAND2_X1 U132 ( .A1(\A_s[29] ), .A2(n272), .ZN(n358) );
  INV_X1 U133 ( .A(A_ns[29]), .ZN(n353) );
  OAI221_X1 U134 ( .B1(n267), .B2(n359), .C1(n269), .C2(n357), .A(n360), .ZN(
        O[28]) );
  NAND2_X1 U135 ( .A1(\A_s[28] ), .A2(n272), .ZN(n360) );
  INV_X1 U136 ( .A(A_ns[28]), .ZN(n357) );
  OAI221_X1 U137 ( .B1(n267), .B2(n361), .C1(n269), .C2(n359), .A(n362), .ZN(
        O[27]) );
  NAND2_X1 U138 ( .A1(\A_s[27] ), .A2(n272), .ZN(n362) );
  INV_X1 U139 ( .A(A_ns[27]), .ZN(n359) );
  OAI221_X1 U140 ( .B1(n267), .B2(n363), .C1(n269), .C2(n361), .A(n364), .ZN(
        O[26]) );
  NAND2_X1 U141 ( .A1(\A_s[26] ), .A2(n272), .ZN(n364) );
  INV_X1 U142 ( .A(A_ns[26]), .ZN(n361) );
  OAI221_X1 U143 ( .B1(n267), .B2(n365), .C1(n269), .C2(n363), .A(n366), .ZN(
        O[25]) );
  NAND2_X1 U144 ( .A1(\A_s[25] ), .A2(n272), .ZN(n366) );
  INV_X1 U145 ( .A(A_ns[25]), .ZN(n363) );
  OAI221_X1 U146 ( .B1(n267), .B2(n367), .C1(n269), .C2(n365), .A(n368), .ZN(
        O[24]) );
  NAND2_X1 U147 ( .A1(\A_s[24] ), .A2(n272), .ZN(n368) );
  INV_X1 U148 ( .A(A_ns[24]), .ZN(n365) );
  OAI221_X1 U149 ( .B1(n267), .B2(n369), .C1(n269), .C2(n367), .A(n370), .ZN(
        O[23]) );
  NAND2_X1 U150 ( .A1(\A_s[23] ), .A2(n272), .ZN(n370) );
  INV_X1 U151 ( .A(A_ns[23]), .ZN(n367) );
  OAI221_X1 U152 ( .B1(n267), .B2(n371), .C1(n269), .C2(n369), .A(n372), .ZN(
        O[22]) );
  NAND2_X1 U153 ( .A1(\A_s[22] ), .A2(n272), .ZN(n372) );
  INV_X1 U154 ( .A(A_ns[22]), .ZN(n369) );
  OAI221_X1 U155 ( .B1(n267), .B2(n373), .C1(n269), .C2(n371), .A(n374), .ZN(
        O[21]) );
  NAND2_X1 U156 ( .A1(\A_s[21] ), .A2(n272), .ZN(n374) );
  INV_X1 U157 ( .A(A_ns[21]), .ZN(n371) );
  OAI221_X1 U158 ( .B1(n267), .B2(n375), .C1(n269), .C2(n373), .A(n376), .ZN(
        O[20]) );
  NAND2_X1 U159 ( .A1(\A_s[20] ), .A2(n272), .ZN(n376) );
  INV_X1 U160 ( .A(A_ns[20]), .ZN(n373) );
  OAI221_X1 U161 ( .B1(n267), .B2(n377), .C1(n269), .C2(n355), .A(n378), .ZN(
        O[1]) );
  NAND2_X1 U162 ( .A1(\A_s[1] ), .A2(n272), .ZN(n378) );
  INV_X1 U163 ( .A(A_ns[1]), .ZN(n355) );
  OAI221_X1 U164 ( .B1(n267), .B2(n379), .C1(n269), .C2(n375), .A(n380), .ZN(
        O[19]) );
  NAND2_X1 U165 ( .A1(\A_s[19] ), .A2(n272), .ZN(n380) );
  INV_X1 U166 ( .A(A_ns[19]), .ZN(n375) );
  OAI221_X1 U167 ( .B1(n267), .B2(n381), .C1(n269), .C2(n379), .A(n382), .ZN(
        O[18]) );
  NAND2_X1 U168 ( .A1(\A_s[18] ), .A2(n272), .ZN(n382) );
  INV_X1 U169 ( .A(A_ns[18]), .ZN(n379) );
  OAI221_X1 U170 ( .B1(n267), .B2(n383), .C1(n269), .C2(n381), .A(n384), .ZN(
        O[17]) );
  NAND2_X1 U171 ( .A1(\A_s[17] ), .A2(n272), .ZN(n384) );
  INV_X1 U172 ( .A(A_ns[17]), .ZN(n381) );
  OAI221_X1 U173 ( .B1(n267), .B2(n385), .C1(n269), .C2(n383), .A(n386), .ZN(
        O[16]) );
  NAND2_X1 U174 ( .A1(\A_s[16] ), .A2(n272), .ZN(n386) );
  INV_X1 U175 ( .A(A_ns[16]), .ZN(n383) );
  OAI221_X1 U176 ( .B1(n267), .B2(n387), .C1(n269), .C2(n385), .A(n388), .ZN(
        O[15]) );
  NAND2_X1 U177 ( .A1(\A_s[15] ), .A2(n272), .ZN(n388) );
  INV_X1 U178 ( .A(A_ns[15]), .ZN(n385) );
  OAI221_X1 U179 ( .B1(n267), .B2(n389), .C1(n269), .C2(n387), .A(n390), .ZN(
        O[14]) );
  NAND2_X1 U180 ( .A1(\A_s[14] ), .A2(n272), .ZN(n390) );
  INV_X1 U181 ( .A(A_ns[14]), .ZN(n387) );
  OAI221_X1 U182 ( .B1(n267), .B2(n391), .C1(n269), .C2(n389), .A(n392), .ZN(
        O[13]) );
  NAND2_X1 U183 ( .A1(\A_s[13] ), .A2(n272), .ZN(n392) );
  INV_X1 U184 ( .A(A_ns[13]), .ZN(n389) );
  OAI221_X1 U185 ( .B1(n267), .B2(n393), .C1(n269), .C2(n391), .A(n394), .ZN(
        O[12]) );
  NAND2_X1 U186 ( .A1(\A_s[12] ), .A2(n272), .ZN(n394) );
  INV_X1 U187 ( .A(A_ns[12]), .ZN(n391) );
  OAI221_X1 U188 ( .B1(n267), .B2(n395), .C1(n269), .C2(n393), .A(n396), .ZN(
        O[11]) );
  NAND2_X1 U189 ( .A1(\A_s[11] ), .A2(n272), .ZN(n396) );
  INV_X1 U190 ( .A(A_ns[11]), .ZN(n393) );
  OAI221_X1 U191 ( .B1(n267), .B2(n270), .C1(n269), .C2(n395), .A(n397), .ZN(
        O[10]) );
  NAND2_X1 U192 ( .A1(\A_s[10] ), .A2(n272), .ZN(n397) );
  INV_X1 U193 ( .A(A_ns[10]), .ZN(n395) );
  INV_X1 U194 ( .A(A_ns[9]), .ZN(n270) );
  OAI22_X1 U195 ( .A1(n280), .A2(n399), .B1(n269), .B2(n377), .ZN(O[0]) );
  INV_X1 U196 ( .A(A_ns[0]), .ZN(n377) );
  INV_X1 U197 ( .A(\A_s[0] ), .ZN(n399) );
  NAND2_X1 U198 ( .A1(B[0]), .A2(n398), .ZN(n280) );
  INV_X1 U199 ( .A(B[1]), .ZN(n398) );
endmodule


module BOOTHENC_NBIT64_i2 ( A, A_n, A_ns, A_s, B, O, A_so, A_nso );
  input [63:0] A;
  input [63:0] A_n;
  input [63:0] A_ns;
  input [63:0] A_s;
  input [63:0] B;
  output [63:0] O;
  output [63:0] A_so;
  output [63:0] A_nso;
  wire   \A_s[61] , \A_s[60] , \A_s[59] , \A_s[58] , \A_s[57] , \A_s[56] ,
         \A_s[55] , \A_s[54] , \A_s[53] , \A_s[52] , \A_s[51] , \A_s[50] ,
         \A_s[49] , \A_s[48] , \A_s[47] , \A_s[46] , \A_s[45] , \A_s[44] ,
         \A_s[43] , \A_s[42] , \A_s[41] , \A_s[40] , \A_s[39] , \A_s[38] ,
         \A_s[37] , \A_s[36] , \A_s[35] , \A_s[34] , \A_s[33] , \A_s[32] ,
         \A_s[31] , \A_s[30] , \A_s[29] , \A_s[28] , \A_s[27] , \A_s[26] ,
         \A_s[25] , \A_s[24] , \A_s[23] , \A_s[22] , \A_s[21] , \A_s[20] ,
         \A_s[19] , \A_s[18] , \A_s[17] , \A_s[16] , \A_s[15] , \A_s[14] ,
         \A_s[13] , \A_s[12] , \A_s[11] , \A_s[10] , \A_s[9] , \A_s[8] ,
         \A_s[7] , \A_s[6] , \A_s[5] , \A_s[4] , \A_s[3] , \A_s[2] , \A_s[1] ,
         \A_s[0] , n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585;
  assign A_nso[0] = 1'b0;
  assign A_nso[1] = 1'b0;
  assign A_so[0] = 1'b0;
  assign A_so[1] = 1'b0;
  assign O[0] = 1'b0;
  assign A_nso[63] = \A_s[61] ;
  assign A_so[63] = \A_s[61] ;
  assign \A_s[61]  = A_s[61];
  assign A_nso[62] = \A_s[60] ;
  assign A_so[62] = \A_s[60] ;
  assign \A_s[60]  = A_s[60];
  assign A_nso[61] = \A_s[59] ;
  assign A_so[61] = \A_s[59] ;
  assign \A_s[59]  = A_s[59];
  assign A_nso[60] = \A_s[58] ;
  assign A_so[60] = \A_s[58] ;
  assign \A_s[58]  = A_s[58];
  assign A_nso[59] = \A_s[57] ;
  assign A_so[59] = \A_s[57] ;
  assign \A_s[57]  = A_s[57];
  assign A_nso[58] = \A_s[56] ;
  assign A_so[58] = \A_s[56] ;
  assign \A_s[56]  = A_s[56];
  assign A_nso[57] = \A_s[55] ;
  assign A_so[57] = \A_s[55] ;
  assign \A_s[55]  = A_s[55];
  assign A_nso[56] = \A_s[54] ;
  assign A_so[56] = \A_s[54] ;
  assign \A_s[54]  = A_s[54];
  assign A_nso[55] = \A_s[53] ;
  assign A_so[55] = \A_s[53] ;
  assign \A_s[53]  = A_s[53];
  assign A_nso[54] = \A_s[52] ;
  assign A_so[54] = \A_s[52] ;
  assign \A_s[52]  = A_s[52];
  assign A_nso[53] = \A_s[51] ;
  assign A_so[53] = \A_s[51] ;
  assign \A_s[51]  = A_s[51];
  assign A_nso[52] = \A_s[50] ;
  assign A_so[52] = \A_s[50] ;
  assign \A_s[50]  = A_s[50];
  assign A_nso[51] = \A_s[49] ;
  assign A_so[51] = \A_s[49] ;
  assign \A_s[49]  = A_s[49];
  assign A_nso[50] = \A_s[48] ;
  assign A_so[50] = \A_s[48] ;
  assign \A_s[48]  = A_s[48];
  assign A_nso[49] = \A_s[47] ;
  assign A_so[49] = \A_s[47] ;
  assign \A_s[47]  = A_s[47];
  assign A_nso[48] = \A_s[46] ;
  assign A_so[48] = \A_s[46] ;
  assign \A_s[46]  = A_s[46];
  assign A_nso[47] = \A_s[45] ;
  assign A_so[47] = \A_s[45] ;
  assign \A_s[45]  = A_s[45];
  assign A_nso[46] = \A_s[44] ;
  assign A_so[46] = \A_s[44] ;
  assign \A_s[44]  = A_s[44];
  assign A_nso[45] = \A_s[43] ;
  assign A_so[45] = \A_s[43] ;
  assign \A_s[43]  = A_s[43];
  assign A_nso[44] = \A_s[42] ;
  assign A_so[44] = \A_s[42] ;
  assign \A_s[42]  = A_s[42];
  assign A_nso[43] = \A_s[41] ;
  assign A_so[43] = \A_s[41] ;
  assign \A_s[41]  = A_s[41];
  assign A_nso[42] = \A_s[40] ;
  assign A_so[42] = \A_s[40] ;
  assign \A_s[40]  = A_s[40];
  assign A_nso[41] = \A_s[39] ;
  assign A_so[41] = \A_s[39] ;
  assign \A_s[39]  = A_s[39];
  assign A_nso[40] = \A_s[38] ;
  assign A_so[40] = \A_s[38] ;
  assign \A_s[38]  = A_s[38];
  assign A_nso[39] = \A_s[37] ;
  assign A_so[39] = \A_s[37] ;
  assign \A_s[37]  = A_s[37];
  assign A_nso[38] = \A_s[36] ;
  assign A_so[38] = \A_s[36] ;
  assign \A_s[36]  = A_s[36];
  assign A_nso[37] = \A_s[35] ;
  assign A_so[37] = \A_s[35] ;
  assign \A_s[35]  = A_s[35];
  assign A_nso[36] = \A_s[34] ;
  assign A_so[36] = \A_s[34] ;
  assign \A_s[34]  = A_s[34];
  assign A_nso[35] = \A_s[33] ;
  assign A_so[35] = \A_s[33] ;
  assign \A_s[33]  = A_s[33];
  assign A_nso[34] = \A_s[32] ;
  assign A_so[34] = \A_s[32] ;
  assign \A_s[32]  = A_s[32];
  assign A_nso[33] = \A_s[31] ;
  assign A_so[33] = \A_s[31] ;
  assign \A_s[31]  = A_s[31];
  assign A_nso[32] = \A_s[30] ;
  assign A_so[32] = \A_s[30] ;
  assign \A_s[30]  = A_s[30];
  assign A_nso[31] = \A_s[29] ;
  assign A_so[31] = \A_s[29] ;
  assign \A_s[29]  = A_s[29];
  assign A_nso[30] = \A_s[28] ;
  assign A_so[30] = \A_s[28] ;
  assign \A_s[28]  = A_s[28];
  assign A_nso[29] = \A_s[27] ;
  assign A_so[29] = \A_s[27] ;
  assign \A_s[27]  = A_s[27];
  assign A_nso[28] = \A_s[26] ;
  assign A_so[28] = \A_s[26] ;
  assign \A_s[26]  = A_s[26];
  assign A_nso[27] = \A_s[25] ;
  assign A_so[27] = \A_s[25] ;
  assign \A_s[25]  = A_s[25];
  assign A_nso[26] = \A_s[24] ;
  assign A_so[26] = \A_s[24] ;
  assign \A_s[24]  = A_s[24];
  assign A_nso[25] = \A_s[23] ;
  assign A_so[25] = \A_s[23] ;
  assign \A_s[23]  = A_s[23];
  assign A_nso[24] = \A_s[22] ;
  assign A_so[24] = \A_s[22] ;
  assign \A_s[22]  = A_s[22];
  assign A_nso[23] = \A_s[21] ;
  assign A_so[23] = \A_s[21] ;
  assign \A_s[21]  = A_s[21];
  assign A_nso[22] = \A_s[20] ;
  assign A_so[22] = \A_s[20] ;
  assign \A_s[20]  = A_s[20];
  assign A_nso[21] = \A_s[19] ;
  assign A_so[21] = \A_s[19] ;
  assign \A_s[19]  = A_s[19];
  assign A_nso[20] = \A_s[18] ;
  assign A_so[20] = \A_s[18] ;
  assign \A_s[18]  = A_s[18];
  assign A_nso[19] = \A_s[17] ;
  assign A_so[19] = \A_s[17] ;
  assign \A_s[17]  = A_s[17];
  assign A_nso[18] = \A_s[16] ;
  assign A_so[18] = \A_s[16] ;
  assign \A_s[16]  = A_s[16];
  assign A_nso[17] = \A_s[15] ;
  assign A_so[17] = \A_s[15] ;
  assign \A_s[15]  = A_s[15];
  assign A_nso[16] = \A_s[14] ;
  assign A_so[16] = \A_s[14] ;
  assign \A_s[14]  = A_s[14];
  assign A_nso[15] = \A_s[13] ;
  assign A_so[15] = \A_s[13] ;
  assign \A_s[13]  = A_s[13];
  assign A_nso[14] = \A_s[12] ;
  assign A_so[14] = \A_s[12] ;
  assign \A_s[12]  = A_s[12];
  assign A_nso[13] = \A_s[11] ;
  assign A_so[13] = \A_s[11] ;
  assign \A_s[11]  = A_s[11];
  assign A_nso[12] = \A_s[10] ;
  assign A_so[12] = \A_s[10] ;
  assign \A_s[10]  = A_s[10];
  assign A_nso[11] = \A_s[9] ;
  assign A_so[11] = \A_s[9] ;
  assign \A_s[9]  = A_s[9];
  assign A_nso[10] = \A_s[8] ;
  assign A_so[10] = \A_s[8] ;
  assign \A_s[8]  = A_s[8];
  assign A_nso[9] = \A_s[7] ;
  assign A_so[9] = \A_s[7] ;
  assign \A_s[7]  = A_s[7];
  assign A_nso[8] = \A_s[6] ;
  assign A_so[8] = \A_s[6] ;
  assign \A_s[6]  = A_s[6];
  assign A_nso[7] = \A_s[5] ;
  assign A_so[7] = \A_s[5] ;
  assign \A_s[5]  = A_s[5];
  assign A_nso[6] = \A_s[4] ;
  assign A_so[6] = \A_s[4] ;
  assign \A_s[4]  = A_s[4];
  assign A_nso[5] = \A_s[3] ;
  assign A_so[5] = \A_s[3] ;
  assign \A_s[3]  = A_s[3];
  assign A_nso[4] = \A_s[2] ;
  assign A_so[4] = \A_s[2] ;
  assign \A_s[2]  = A_s[2];
  assign A_nso[3] = \A_s[1] ;
  assign A_so[3] = \A_s[1] ;
  assign \A_s[1]  = A_s[1];
  assign A_nso[2] = \A_s[0] ;
  assign A_so[2] = \A_s[0] ;
  assign \A_s[0]  = A_s[0];

  AND3_X1 U2 ( .A1(B[2]), .A2(n585), .A3(B[1]), .ZN(n391) );
  INV_X4 U3 ( .A(n391), .ZN(n392) );
  INV_X4 U4 ( .A(n552), .ZN(n398) );
  OR3_X4 U5 ( .A1(B[1]), .A2(B[2]), .A3(n585), .ZN(n393) );
  INV_X4 U6 ( .A(n553), .ZN(n397) );
  OAI221_X1 U7 ( .B1(n393), .B2(n394), .C1(n392), .C2(n395), .A(n396), .ZN(
        O[9]) );
  AOI22_X1 U8 ( .A1(A_ns[8]), .A2(n397), .B1(\A_s[8] ), .B2(n398), .ZN(n396)
         );
  INV_X1 U9 ( .A(\A_s[7] ), .ZN(n395) );
  INV_X1 U10 ( .A(A_ns[7]), .ZN(n394) );
  OAI221_X1 U11 ( .B1(n393), .B2(n399), .C1(n392), .C2(n400), .A(n401), .ZN(
        O[8]) );
  AOI22_X1 U12 ( .A1(A_ns[7]), .A2(n397), .B1(\A_s[7] ), .B2(n398), .ZN(n401)
         );
  INV_X1 U13 ( .A(\A_s[6] ), .ZN(n400) );
  INV_X1 U14 ( .A(A_ns[6]), .ZN(n399) );
  OAI221_X1 U15 ( .B1(n393), .B2(n402), .C1(n392), .C2(n403), .A(n404), .ZN(
        O[7]) );
  AOI22_X1 U16 ( .A1(A_ns[6]), .A2(n397), .B1(\A_s[6] ), .B2(n398), .ZN(n404)
         );
  INV_X1 U17 ( .A(\A_s[5] ), .ZN(n403) );
  INV_X1 U18 ( .A(A_ns[5]), .ZN(n402) );
  OAI221_X1 U19 ( .B1(n393), .B2(n405), .C1(n392), .C2(n406), .A(n407), .ZN(
        O[6]) );
  AOI22_X1 U20 ( .A1(A_ns[5]), .A2(n397), .B1(\A_s[5] ), .B2(n398), .ZN(n407)
         );
  INV_X1 U21 ( .A(\A_s[4] ), .ZN(n406) );
  INV_X1 U22 ( .A(A_ns[4]), .ZN(n405) );
  OAI221_X1 U23 ( .B1(n393), .B2(n408), .C1(n392), .C2(n409), .A(n410), .ZN(
        O[63]) );
  AOI22_X1 U24 ( .A1(A_ns[62]), .A2(n397), .B1(A_s[62]), .B2(n398), .ZN(n410)
         );
  INV_X1 U25 ( .A(\A_s[61] ), .ZN(n409) );
  INV_X1 U26 ( .A(A_ns[61]), .ZN(n408) );
  OAI221_X1 U27 ( .B1(n393), .B2(n411), .C1(n392), .C2(n412), .A(n413), .ZN(
        O[62]) );
  AOI22_X1 U28 ( .A1(A_ns[61]), .A2(n397), .B1(\A_s[61] ), .B2(n398), .ZN(n413) );
  INV_X1 U29 ( .A(\A_s[60] ), .ZN(n412) );
  INV_X1 U30 ( .A(A_ns[60]), .ZN(n411) );
  OAI221_X1 U31 ( .B1(n393), .B2(n414), .C1(n392), .C2(n415), .A(n416), .ZN(
        O[61]) );
  AOI22_X1 U32 ( .A1(A_ns[60]), .A2(n397), .B1(\A_s[60] ), .B2(n398), .ZN(n416) );
  INV_X1 U33 ( .A(\A_s[59] ), .ZN(n415) );
  INV_X1 U34 ( .A(A_ns[59]), .ZN(n414) );
  OAI221_X1 U35 ( .B1(n393), .B2(n417), .C1(n392), .C2(n418), .A(n419), .ZN(
        O[60]) );
  AOI22_X1 U36 ( .A1(A_ns[59]), .A2(n397), .B1(\A_s[59] ), .B2(n398), .ZN(n419) );
  INV_X1 U37 ( .A(\A_s[58] ), .ZN(n418) );
  INV_X1 U38 ( .A(A_ns[58]), .ZN(n417) );
  OAI221_X1 U39 ( .B1(n393), .B2(n420), .C1(n392), .C2(n421), .A(n422), .ZN(
        O[5]) );
  AOI22_X1 U40 ( .A1(A_ns[4]), .A2(n397), .B1(\A_s[4] ), .B2(n398), .ZN(n422)
         );
  INV_X1 U41 ( .A(\A_s[3] ), .ZN(n421) );
  INV_X1 U42 ( .A(A_ns[3]), .ZN(n420) );
  OAI221_X1 U43 ( .B1(n393), .B2(n423), .C1(n392), .C2(n424), .A(n425), .ZN(
        O[59]) );
  AOI22_X1 U44 ( .A1(A_ns[58]), .A2(n397), .B1(\A_s[58] ), .B2(n398), .ZN(n425) );
  INV_X1 U45 ( .A(\A_s[57] ), .ZN(n424) );
  INV_X1 U46 ( .A(A_ns[57]), .ZN(n423) );
  OAI221_X1 U47 ( .B1(n393), .B2(n426), .C1(n392), .C2(n427), .A(n428), .ZN(
        O[58]) );
  AOI22_X1 U48 ( .A1(A_ns[57]), .A2(n397), .B1(\A_s[57] ), .B2(n398), .ZN(n428) );
  INV_X1 U49 ( .A(\A_s[56] ), .ZN(n427) );
  INV_X1 U50 ( .A(A_ns[56]), .ZN(n426) );
  OAI221_X1 U51 ( .B1(n393), .B2(n429), .C1(n392), .C2(n430), .A(n431), .ZN(
        O[57]) );
  AOI22_X1 U52 ( .A1(A_ns[56]), .A2(n397), .B1(\A_s[56] ), .B2(n398), .ZN(n431) );
  INV_X1 U53 ( .A(\A_s[55] ), .ZN(n430) );
  INV_X1 U54 ( .A(A_ns[55]), .ZN(n429) );
  OAI221_X1 U55 ( .B1(n393), .B2(n432), .C1(n392), .C2(n433), .A(n434), .ZN(
        O[56]) );
  AOI22_X1 U56 ( .A1(A_ns[55]), .A2(n397), .B1(\A_s[55] ), .B2(n398), .ZN(n434) );
  INV_X1 U57 ( .A(\A_s[54] ), .ZN(n433) );
  INV_X1 U58 ( .A(A_ns[54]), .ZN(n432) );
  OAI221_X1 U59 ( .B1(n393), .B2(n435), .C1(n392), .C2(n436), .A(n437), .ZN(
        O[55]) );
  AOI22_X1 U60 ( .A1(A_ns[54]), .A2(n397), .B1(\A_s[54] ), .B2(n398), .ZN(n437) );
  INV_X1 U61 ( .A(\A_s[53] ), .ZN(n436) );
  INV_X1 U62 ( .A(A_ns[53]), .ZN(n435) );
  OAI221_X1 U63 ( .B1(n393), .B2(n438), .C1(n392), .C2(n439), .A(n440), .ZN(
        O[54]) );
  AOI22_X1 U64 ( .A1(A_ns[53]), .A2(n397), .B1(\A_s[53] ), .B2(n398), .ZN(n440) );
  INV_X1 U65 ( .A(\A_s[52] ), .ZN(n439) );
  INV_X1 U66 ( .A(A_ns[52]), .ZN(n438) );
  OAI221_X1 U67 ( .B1(n393), .B2(n441), .C1(n392), .C2(n442), .A(n443), .ZN(
        O[53]) );
  AOI22_X1 U68 ( .A1(A_ns[52]), .A2(n397), .B1(\A_s[52] ), .B2(n398), .ZN(n443) );
  INV_X1 U69 ( .A(\A_s[51] ), .ZN(n442) );
  INV_X1 U70 ( .A(A_ns[51]), .ZN(n441) );
  OAI221_X1 U71 ( .B1(n393), .B2(n444), .C1(n392), .C2(n445), .A(n446), .ZN(
        O[52]) );
  AOI22_X1 U72 ( .A1(A_ns[51]), .A2(n397), .B1(\A_s[51] ), .B2(n398), .ZN(n446) );
  INV_X1 U73 ( .A(\A_s[50] ), .ZN(n445) );
  INV_X1 U74 ( .A(A_ns[50]), .ZN(n444) );
  OAI221_X1 U75 ( .B1(n393), .B2(n447), .C1(n392), .C2(n448), .A(n449), .ZN(
        O[51]) );
  AOI22_X1 U76 ( .A1(A_ns[50]), .A2(n397), .B1(\A_s[50] ), .B2(n398), .ZN(n449) );
  INV_X1 U77 ( .A(\A_s[49] ), .ZN(n448) );
  INV_X1 U78 ( .A(A_ns[49]), .ZN(n447) );
  OAI221_X1 U79 ( .B1(n393), .B2(n450), .C1(n392), .C2(n451), .A(n452), .ZN(
        O[50]) );
  AOI22_X1 U80 ( .A1(A_ns[49]), .A2(n397), .B1(\A_s[49] ), .B2(n398), .ZN(n452) );
  INV_X1 U81 ( .A(\A_s[48] ), .ZN(n451) );
  INV_X1 U82 ( .A(A_ns[48]), .ZN(n450) );
  OAI221_X1 U83 ( .B1(n393), .B2(n453), .C1(n392), .C2(n454), .A(n455), .ZN(
        O[4]) );
  AOI22_X1 U84 ( .A1(A_ns[3]), .A2(n397), .B1(\A_s[3] ), .B2(n398), .ZN(n455)
         );
  INV_X1 U85 ( .A(\A_s[2] ), .ZN(n454) );
  INV_X1 U86 ( .A(A_ns[2]), .ZN(n453) );
  OAI221_X1 U87 ( .B1(n393), .B2(n456), .C1(n392), .C2(n457), .A(n458), .ZN(
        O[49]) );
  AOI22_X1 U88 ( .A1(A_ns[48]), .A2(n397), .B1(\A_s[48] ), .B2(n398), .ZN(n458) );
  INV_X1 U89 ( .A(\A_s[47] ), .ZN(n457) );
  INV_X1 U90 ( .A(A_ns[47]), .ZN(n456) );
  OAI221_X1 U91 ( .B1(n393), .B2(n459), .C1(n392), .C2(n460), .A(n461), .ZN(
        O[48]) );
  AOI22_X1 U92 ( .A1(A_ns[47]), .A2(n397), .B1(\A_s[47] ), .B2(n398), .ZN(n461) );
  INV_X1 U93 ( .A(\A_s[46] ), .ZN(n460) );
  INV_X1 U94 ( .A(A_ns[46]), .ZN(n459) );
  OAI221_X1 U95 ( .B1(n393), .B2(n462), .C1(n392), .C2(n463), .A(n464), .ZN(
        O[47]) );
  AOI22_X1 U96 ( .A1(A_ns[46]), .A2(n397), .B1(\A_s[46] ), .B2(n398), .ZN(n464) );
  INV_X1 U97 ( .A(\A_s[45] ), .ZN(n463) );
  INV_X1 U98 ( .A(A_ns[45]), .ZN(n462) );
  OAI221_X1 U99 ( .B1(n393), .B2(n465), .C1(n392), .C2(n466), .A(n467), .ZN(
        O[46]) );
  AOI22_X1 U100 ( .A1(A_ns[45]), .A2(n397), .B1(\A_s[45] ), .B2(n398), .ZN(
        n467) );
  INV_X1 U101 ( .A(\A_s[44] ), .ZN(n466) );
  INV_X1 U102 ( .A(A_ns[44]), .ZN(n465) );
  OAI221_X1 U103 ( .B1(n393), .B2(n468), .C1(n392), .C2(n469), .A(n470), .ZN(
        O[45]) );
  AOI22_X1 U104 ( .A1(A_ns[44]), .A2(n397), .B1(\A_s[44] ), .B2(n398), .ZN(
        n470) );
  INV_X1 U105 ( .A(\A_s[43] ), .ZN(n469) );
  INV_X1 U106 ( .A(A_ns[43]), .ZN(n468) );
  OAI221_X1 U107 ( .B1(n393), .B2(n471), .C1(n392), .C2(n472), .A(n473), .ZN(
        O[44]) );
  AOI22_X1 U108 ( .A1(A_ns[43]), .A2(n397), .B1(\A_s[43] ), .B2(n398), .ZN(
        n473) );
  INV_X1 U109 ( .A(\A_s[42] ), .ZN(n472) );
  INV_X1 U110 ( .A(A_ns[42]), .ZN(n471) );
  OAI221_X1 U111 ( .B1(n393), .B2(n474), .C1(n392), .C2(n475), .A(n476), .ZN(
        O[43]) );
  AOI22_X1 U112 ( .A1(A_ns[42]), .A2(n397), .B1(\A_s[42] ), .B2(n398), .ZN(
        n476) );
  INV_X1 U113 ( .A(\A_s[41] ), .ZN(n475) );
  INV_X1 U114 ( .A(A_ns[41]), .ZN(n474) );
  OAI221_X1 U115 ( .B1(n393), .B2(n477), .C1(n392), .C2(n478), .A(n479), .ZN(
        O[42]) );
  AOI22_X1 U116 ( .A1(A_ns[41]), .A2(n397), .B1(\A_s[41] ), .B2(n398), .ZN(
        n479) );
  INV_X1 U117 ( .A(\A_s[40] ), .ZN(n478) );
  INV_X1 U118 ( .A(A_ns[40]), .ZN(n477) );
  OAI221_X1 U119 ( .B1(n393), .B2(n480), .C1(n392), .C2(n481), .A(n482), .ZN(
        O[41]) );
  AOI22_X1 U120 ( .A1(A_ns[40]), .A2(n397), .B1(\A_s[40] ), .B2(n398), .ZN(
        n482) );
  INV_X1 U121 ( .A(\A_s[39] ), .ZN(n481) );
  INV_X1 U122 ( .A(A_ns[39]), .ZN(n480) );
  OAI221_X1 U123 ( .B1(n393), .B2(n483), .C1(n392), .C2(n484), .A(n485), .ZN(
        O[40]) );
  AOI22_X1 U124 ( .A1(A_ns[39]), .A2(n397), .B1(\A_s[39] ), .B2(n398), .ZN(
        n485) );
  INV_X1 U125 ( .A(\A_s[38] ), .ZN(n484) );
  INV_X1 U126 ( .A(A_ns[38]), .ZN(n483) );
  OAI221_X1 U127 ( .B1(n393), .B2(n486), .C1(n392), .C2(n487), .A(n488), .ZN(
        O[3]) );
  AOI22_X1 U128 ( .A1(A_ns[2]), .A2(n397), .B1(\A_s[2] ), .B2(n398), .ZN(n488)
         );
  INV_X1 U129 ( .A(\A_s[1] ), .ZN(n487) );
  INV_X1 U130 ( .A(A_ns[1]), .ZN(n486) );
  OAI221_X1 U131 ( .B1(n393), .B2(n489), .C1(n392), .C2(n490), .A(n491), .ZN(
        O[39]) );
  AOI22_X1 U132 ( .A1(A_ns[38]), .A2(n397), .B1(\A_s[38] ), .B2(n398), .ZN(
        n491) );
  INV_X1 U133 ( .A(\A_s[37] ), .ZN(n490) );
  INV_X1 U134 ( .A(A_ns[37]), .ZN(n489) );
  OAI221_X1 U135 ( .B1(n393), .B2(n492), .C1(n392), .C2(n493), .A(n494), .ZN(
        O[38]) );
  AOI22_X1 U136 ( .A1(A_ns[37]), .A2(n397), .B1(\A_s[37] ), .B2(n398), .ZN(
        n494) );
  INV_X1 U137 ( .A(\A_s[36] ), .ZN(n493) );
  INV_X1 U138 ( .A(A_ns[36]), .ZN(n492) );
  OAI221_X1 U139 ( .B1(n393), .B2(n495), .C1(n392), .C2(n496), .A(n497), .ZN(
        O[37]) );
  AOI22_X1 U140 ( .A1(A_ns[36]), .A2(n397), .B1(\A_s[36] ), .B2(n398), .ZN(
        n497) );
  INV_X1 U141 ( .A(\A_s[35] ), .ZN(n496) );
  INV_X1 U142 ( .A(A_ns[35]), .ZN(n495) );
  OAI221_X1 U143 ( .B1(n393), .B2(n498), .C1(n392), .C2(n499), .A(n500), .ZN(
        O[36]) );
  AOI22_X1 U144 ( .A1(A_ns[35]), .A2(n397), .B1(\A_s[35] ), .B2(n398), .ZN(
        n500) );
  INV_X1 U145 ( .A(\A_s[34] ), .ZN(n499) );
  INV_X1 U146 ( .A(A_ns[34]), .ZN(n498) );
  OAI221_X1 U147 ( .B1(n393), .B2(n501), .C1(n392), .C2(n502), .A(n503), .ZN(
        O[35]) );
  AOI22_X1 U148 ( .A1(A_ns[34]), .A2(n397), .B1(\A_s[34] ), .B2(n398), .ZN(
        n503) );
  INV_X1 U149 ( .A(\A_s[33] ), .ZN(n502) );
  INV_X1 U150 ( .A(A_ns[33]), .ZN(n501) );
  OAI221_X1 U151 ( .B1(n393), .B2(n504), .C1(n392), .C2(n505), .A(n506), .ZN(
        O[34]) );
  AOI22_X1 U152 ( .A1(A_ns[33]), .A2(n397), .B1(\A_s[33] ), .B2(n398), .ZN(
        n506) );
  INV_X1 U153 ( .A(\A_s[32] ), .ZN(n505) );
  INV_X1 U154 ( .A(A_ns[32]), .ZN(n504) );
  OAI221_X1 U155 ( .B1(n393), .B2(n507), .C1(n392), .C2(n508), .A(n509), .ZN(
        O[33]) );
  AOI22_X1 U156 ( .A1(A_ns[32]), .A2(n397), .B1(\A_s[32] ), .B2(n398), .ZN(
        n509) );
  INV_X1 U157 ( .A(\A_s[31] ), .ZN(n508) );
  INV_X1 U158 ( .A(A_ns[31]), .ZN(n507) );
  OAI221_X1 U159 ( .B1(n393), .B2(n510), .C1(n392), .C2(n511), .A(n512), .ZN(
        O[32]) );
  AOI22_X1 U160 ( .A1(A_ns[31]), .A2(n397), .B1(\A_s[31] ), .B2(n398), .ZN(
        n512) );
  INV_X1 U161 ( .A(\A_s[30] ), .ZN(n511) );
  INV_X1 U162 ( .A(A_ns[30]), .ZN(n510) );
  OAI221_X1 U163 ( .B1(n393), .B2(n513), .C1(n392), .C2(n514), .A(n515), .ZN(
        O[31]) );
  AOI22_X1 U164 ( .A1(A_ns[30]), .A2(n397), .B1(\A_s[30] ), .B2(n398), .ZN(
        n515) );
  INV_X1 U165 ( .A(\A_s[29] ), .ZN(n514) );
  INV_X1 U166 ( .A(A_ns[29]), .ZN(n513) );
  OAI221_X1 U167 ( .B1(n393), .B2(n516), .C1(n392), .C2(n517), .A(n518), .ZN(
        O[30]) );
  AOI22_X1 U168 ( .A1(A_ns[29]), .A2(n397), .B1(\A_s[29] ), .B2(n398), .ZN(
        n518) );
  INV_X1 U169 ( .A(\A_s[28] ), .ZN(n517) );
  INV_X1 U170 ( .A(A_ns[28]), .ZN(n516) );
  OAI221_X1 U171 ( .B1(n393), .B2(n519), .C1(n392), .C2(n520), .A(n521), .ZN(
        O[2]) );
  AOI22_X1 U172 ( .A1(A_ns[1]), .A2(n397), .B1(\A_s[1] ), .B2(n398), .ZN(n521)
         );
  OAI221_X1 U173 ( .B1(n393), .B2(n522), .C1(n392), .C2(n523), .A(n524), .ZN(
        O[29]) );
  AOI22_X1 U174 ( .A1(A_ns[28]), .A2(n397), .B1(\A_s[28] ), .B2(n398), .ZN(
        n524) );
  INV_X1 U175 ( .A(\A_s[27] ), .ZN(n523) );
  INV_X1 U176 ( .A(A_ns[27]), .ZN(n522) );
  OAI221_X1 U177 ( .B1(n393), .B2(n525), .C1(n392), .C2(n526), .A(n527), .ZN(
        O[28]) );
  AOI22_X1 U178 ( .A1(A_ns[27]), .A2(n397), .B1(\A_s[27] ), .B2(n398), .ZN(
        n527) );
  INV_X1 U179 ( .A(\A_s[26] ), .ZN(n526) );
  INV_X1 U180 ( .A(A_ns[26]), .ZN(n525) );
  OAI221_X1 U181 ( .B1(n393), .B2(n528), .C1(n392), .C2(n529), .A(n530), .ZN(
        O[27]) );
  AOI22_X1 U182 ( .A1(A_ns[26]), .A2(n397), .B1(\A_s[26] ), .B2(n398), .ZN(
        n530) );
  INV_X1 U183 ( .A(\A_s[25] ), .ZN(n529) );
  INV_X1 U184 ( .A(A_ns[25]), .ZN(n528) );
  OAI221_X1 U185 ( .B1(n393), .B2(n531), .C1(n392), .C2(n532), .A(n533), .ZN(
        O[26]) );
  AOI22_X1 U186 ( .A1(A_ns[25]), .A2(n397), .B1(\A_s[25] ), .B2(n398), .ZN(
        n533) );
  INV_X1 U187 ( .A(\A_s[24] ), .ZN(n532) );
  INV_X1 U188 ( .A(A_ns[24]), .ZN(n531) );
  OAI221_X1 U189 ( .B1(n393), .B2(n534), .C1(n392), .C2(n535), .A(n536), .ZN(
        O[25]) );
  AOI22_X1 U190 ( .A1(A_ns[24]), .A2(n397), .B1(\A_s[24] ), .B2(n398), .ZN(
        n536) );
  INV_X1 U191 ( .A(\A_s[23] ), .ZN(n535) );
  INV_X1 U192 ( .A(A_ns[23]), .ZN(n534) );
  OAI221_X1 U193 ( .B1(n393), .B2(n537), .C1(n392), .C2(n538), .A(n539), .ZN(
        O[24]) );
  AOI22_X1 U194 ( .A1(A_ns[23]), .A2(n397), .B1(\A_s[23] ), .B2(n398), .ZN(
        n539) );
  INV_X1 U195 ( .A(\A_s[22] ), .ZN(n538) );
  INV_X1 U196 ( .A(A_ns[22]), .ZN(n537) );
  OAI221_X1 U197 ( .B1(n393), .B2(n540), .C1(n392), .C2(n541), .A(n542), .ZN(
        O[23]) );
  AOI22_X1 U198 ( .A1(A_ns[22]), .A2(n397), .B1(\A_s[22] ), .B2(n398), .ZN(
        n542) );
  INV_X1 U199 ( .A(\A_s[21] ), .ZN(n541) );
  INV_X1 U200 ( .A(A_ns[21]), .ZN(n540) );
  OAI221_X1 U201 ( .B1(n393), .B2(n543), .C1(n392), .C2(n544), .A(n545), .ZN(
        O[22]) );
  AOI22_X1 U202 ( .A1(A_ns[21]), .A2(n397), .B1(\A_s[21] ), .B2(n398), .ZN(
        n545) );
  INV_X1 U203 ( .A(\A_s[20] ), .ZN(n544) );
  INV_X1 U204 ( .A(A_ns[20]), .ZN(n543) );
  OAI221_X1 U205 ( .B1(n393), .B2(n546), .C1(n392), .C2(n547), .A(n548), .ZN(
        O[21]) );
  AOI22_X1 U206 ( .A1(A_ns[20]), .A2(n397), .B1(\A_s[20] ), .B2(n398), .ZN(
        n548) );
  INV_X1 U207 ( .A(\A_s[19] ), .ZN(n547) );
  INV_X1 U208 ( .A(A_ns[19]), .ZN(n546) );
  OAI221_X1 U209 ( .B1(n393), .B2(n549), .C1(n392), .C2(n550), .A(n551), .ZN(
        O[20]) );
  AOI22_X1 U210 ( .A1(A_ns[19]), .A2(n397), .B1(\A_s[19] ), .B2(n398), .ZN(
        n551) );
  INV_X1 U211 ( .A(\A_s[18] ), .ZN(n550) );
  INV_X1 U212 ( .A(A_ns[18]), .ZN(n549) );
  OAI22_X1 U213 ( .A1(n552), .A2(n520), .B1(n553), .B2(n519), .ZN(O[1]) );
  INV_X1 U214 ( .A(A_ns[0]), .ZN(n519) );
  INV_X1 U215 ( .A(\A_s[0] ), .ZN(n520) );
  OAI221_X1 U216 ( .B1(n393), .B2(n554), .C1(n392), .C2(n555), .A(n556), .ZN(
        O[19]) );
  AOI22_X1 U217 ( .A1(A_ns[18]), .A2(n397), .B1(\A_s[18] ), .B2(n398), .ZN(
        n556) );
  INV_X1 U218 ( .A(\A_s[17] ), .ZN(n555) );
  INV_X1 U219 ( .A(A_ns[17]), .ZN(n554) );
  OAI221_X1 U220 ( .B1(n393), .B2(n557), .C1(n392), .C2(n558), .A(n559), .ZN(
        O[18]) );
  AOI22_X1 U221 ( .A1(A_ns[17]), .A2(n397), .B1(\A_s[17] ), .B2(n398), .ZN(
        n559) );
  INV_X1 U222 ( .A(\A_s[16] ), .ZN(n558) );
  INV_X1 U223 ( .A(A_ns[16]), .ZN(n557) );
  OAI221_X1 U224 ( .B1(n393), .B2(n560), .C1(n392), .C2(n561), .A(n562), .ZN(
        O[17]) );
  AOI22_X1 U225 ( .A1(A_ns[16]), .A2(n397), .B1(\A_s[16] ), .B2(n398), .ZN(
        n562) );
  INV_X1 U226 ( .A(\A_s[15] ), .ZN(n561) );
  INV_X1 U227 ( .A(A_ns[15]), .ZN(n560) );
  OAI221_X1 U228 ( .B1(n393), .B2(n563), .C1(n392), .C2(n564), .A(n565), .ZN(
        O[16]) );
  AOI22_X1 U229 ( .A1(A_ns[15]), .A2(n397), .B1(\A_s[15] ), .B2(n398), .ZN(
        n565) );
  INV_X1 U230 ( .A(\A_s[14] ), .ZN(n564) );
  INV_X1 U231 ( .A(A_ns[14]), .ZN(n563) );
  OAI221_X1 U232 ( .B1(n393), .B2(n566), .C1(n392), .C2(n567), .A(n568), .ZN(
        O[15]) );
  AOI22_X1 U233 ( .A1(A_ns[14]), .A2(n397), .B1(\A_s[14] ), .B2(n398), .ZN(
        n568) );
  INV_X1 U234 ( .A(\A_s[13] ), .ZN(n567) );
  INV_X1 U235 ( .A(A_ns[13]), .ZN(n566) );
  OAI221_X1 U236 ( .B1(n393), .B2(n569), .C1(n392), .C2(n570), .A(n571), .ZN(
        O[14]) );
  AOI22_X1 U237 ( .A1(A_ns[13]), .A2(n397), .B1(\A_s[13] ), .B2(n398), .ZN(
        n571) );
  INV_X1 U238 ( .A(\A_s[12] ), .ZN(n570) );
  INV_X1 U239 ( .A(A_ns[12]), .ZN(n569) );
  OAI221_X1 U240 ( .B1(n393), .B2(n572), .C1(n392), .C2(n573), .A(n574), .ZN(
        O[13]) );
  AOI22_X1 U241 ( .A1(A_ns[12]), .A2(n397), .B1(\A_s[12] ), .B2(n398), .ZN(
        n574) );
  INV_X1 U242 ( .A(\A_s[11] ), .ZN(n573) );
  INV_X1 U243 ( .A(A_ns[11]), .ZN(n572) );
  OAI221_X1 U244 ( .B1(n393), .B2(n575), .C1(n392), .C2(n576), .A(n577), .ZN(
        O[12]) );
  AOI22_X1 U245 ( .A1(A_ns[11]), .A2(n397), .B1(\A_s[11] ), .B2(n398), .ZN(
        n577) );
  INV_X1 U246 ( .A(\A_s[10] ), .ZN(n576) );
  INV_X1 U247 ( .A(A_ns[10]), .ZN(n575) );
  OAI221_X1 U248 ( .B1(n393), .B2(n578), .C1(n392), .C2(n579), .A(n580), .ZN(
        O[11]) );
  AOI22_X1 U249 ( .A1(A_ns[10]), .A2(n397), .B1(\A_s[10] ), .B2(n398), .ZN(
        n580) );
  INV_X1 U250 ( .A(\A_s[9] ), .ZN(n579) );
  INV_X1 U251 ( .A(A_ns[9]), .ZN(n578) );
  OAI221_X1 U252 ( .B1(n581), .B2(n393), .C1(n582), .C2(n392), .A(n583), .ZN(
        O[10]) );
  AOI22_X1 U253 ( .A1(A_ns[9]), .A2(n397), .B1(\A_s[9] ), .B2(n398), .ZN(n583)
         );
  NAND2_X1 U254 ( .A1(n584), .A2(n552), .ZN(n553) );
  NAND2_X1 U255 ( .A1(n584), .A2(n585), .ZN(n552) );
  XOR2_X1 U256 ( .A(B[1]), .B(B[2]), .Z(n584) );
  INV_X1 U257 ( .A(\A_s[8] ), .ZN(n582) );
  INV_X1 U258 ( .A(B[3]), .ZN(n585) );
  INV_X1 U259 ( .A(A_ns[8]), .ZN(n581) );
endmodule


module BOOTHENC_NBIT64_i4 ( A, A_n, A_ns, A_s, B, O, A_so, A_nso );
  input [63:0] A;
  input [63:0] A_n;
  input [63:0] A_ns;
  input [63:0] A_s;
  input [63:0] B;
  output [63:0] O;
  output [63:0] A_so;
  output [63:0] A_nso;
  wire   \A_s[61] , \A_s[60] , \A_s[59] , \A_s[58] , \A_s[57] , \A_s[56] ,
         \A_s[55] , \A_s[54] , \A_s[53] , \A_s[52] , \A_s[51] , \A_s[50] ,
         \A_s[49] , \A_s[48] , \A_s[47] , \A_s[46] , \A_s[45] , \A_s[44] ,
         \A_s[43] , \A_s[42] , \A_s[41] , \A_s[40] , \A_s[39] , \A_s[38] ,
         \A_s[37] , \A_s[36] , \A_s[35] , \A_s[34] , \A_s[33] , \A_s[32] ,
         \A_s[31] , \A_s[30] , \A_s[29] , \A_s[28] , \A_s[27] , \A_s[26] ,
         \A_s[25] , \A_s[24] , \A_s[23] , \A_s[22] , \A_s[21] , \A_s[20] ,
         \A_s[19] , \A_s[18] , \A_s[17] , \A_s[16] , \A_s[15] , \A_s[14] ,
         \A_s[13] , \A_s[12] , \A_s[11] , \A_s[10] , \A_s[9] , \A_s[8] ,
         \A_s[7] , \A_s[6] , \A_s[5] , \A_s[4] , \A_s[3] , \A_s[2] , \A_s[1] ,
         \A_s[0] , n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585;
  assign A_nso[0] = 1'b0;
  assign A_nso[1] = 1'b0;
  assign A_so[0] = 1'b0;
  assign A_so[1] = 1'b0;
  assign O[0] = 1'b0;
  assign A_nso[63] = \A_s[61] ;
  assign A_so[63] = \A_s[61] ;
  assign \A_s[61]  = A_s[61];
  assign A_nso[62] = \A_s[60] ;
  assign A_so[62] = \A_s[60] ;
  assign \A_s[60]  = A_s[60];
  assign A_nso[61] = \A_s[59] ;
  assign A_so[61] = \A_s[59] ;
  assign \A_s[59]  = A_s[59];
  assign A_nso[60] = \A_s[58] ;
  assign A_so[60] = \A_s[58] ;
  assign \A_s[58]  = A_s[58];
  assign A_nso[59] = \A_s[57] ;
  assign A_so[59] = \A_s[57] ;
  assign \A_s[57]  = A_s[57];
  assign A_nso[58] = \A_s[56] ;
  assign A_so[58] = \A_s[56] ;
  assign \A_s[56]  = A_s[56];
  assign A_nso[57] = \A_s[55] ;
  assign A_so[57] = \A_s[55] ;
  assign \A_s[55]  = A_s[55];
  assign A_nso[56] = \A_s[54] ;
  assign A_so[56] = \A_s[54] ;
  assign \A_s[54]  = A_s[54];
  assign A_nso[55] = \A_s[53] ;
  assign A_so[55] = \A_s[53] ;
  assign \A_s[53]  = A_s[53];
  assign A_nso[54] = \A_s[52] ;
  assign A_so[54] = \A_s[52] ;
  assign \A_s[52]  = A_s[52];
  assign A_nso[53] = \A_s[51] ;
  assign A_so[53] = \A_s[51] ;
  assign \A_s[51]  = A_s[51];
  assign A_nso[52] = \A_s[50] ;
  assign A_so[52] = \A_s[50] ;
  assign \A_s[50]  = A_s[50];
  assign A_nso[51] = \A_s[49] ;
  assign A_so[51] = \A_s[49] ;
  assign \A_s[49]  = A_s[49];
  assign A_nso[50] = \A_s[48] ;
  assign A_so[50] = \A_s[48] ;
  assign \A_s[48]  = A_s[48];
  assign A_nso[49] = \A_s[47] ;
  assign A_so[49] = \A_s[47] ;
  assign \A_s[47]  = A_s[47];
  assign A_nso[48] = \A_s[46] ;
  assign A_so[48] = \A_s[46] ;
  assign \A_s[46]  = A_s[46];
  assign A_nso[47] = \A_s[45] ;
  assign A_so[47] = \A_s[45] ;
  assign \A_s[45]  = A_s[45];
  assign A_nso[46] = \A_s[44] ;
  assign A_so[46] = \A_s[44] ;
  assign \A_s[44]  = A_s[44];
  assign A_nso[45] = \A_s[43] ;
  assign A_so[45] = \A_s[43] ;
  assign \A_s[43]  = A_s[43];
  assign A_nso[44] = \A_s[42] ;
  assign A_so[44] = \A_s[42] ;
  assign \A_s[42]  = A_s[42];
  assign A_nso[43] = \A_s[41] ;
  assign A_so[43] = \A_s[41] ;
  assign \A_s[41]  = A_s[41];
  assign A_nso[42] = \A_s[40] ;
  assign A_so[42] = \A_s[40] ;
  assign \A_s[40]  = A_s[40];
  assign A_nso[41] = \A_s[39] ;
  assign A_so[41] = \A_s[39] ;
  assign \A_s[39]  = A_s[39];
  assign A_nso[40] = \A_s[38] ;
  assign A_so[40] = \A_s[38] ;
  assign \A_s[38]  = A_s[38];
  assign A_nso[39] = \A_s[37] ;
  assign A_so[39] = \A_s[37] ;
  assign \A_s[37]  = A_s[37];
  assign A_nso[38] = \A_s[36] ;
  assign A_so[38] = \A_s[36] ;
  assign \A_s[36]  = A_s[36];
  assign A_nso[37] = \A_s[35] ;
  assign A_so[37] = \A_s[35] ;
  assign \A_s[35]  = A_s[35];
  assign A_nso[36] = \A_s[34] ;
  assign A_so[36] = \A_s[34] ;
  assign \A_s[34]  = A_s[34];
  assign A_nso[35] = \A_s[33] ;
  assign A_so[35] = \A_s[33] ;
  assign \A_s[33]  = A_s[33];
  assign A_nso[34] = \A_s[32] ;
  assign A_so[34] = \A_s[32] ;
  assign \A_s[32]  = A_s[32];
  assign A_nso[33] = \A_s[31] ;
  assign A_so[33] = \A_s[31] ;
  assign \A_s[31]  = A_s[31];
  assign A_nso[32] = \A_s[30] ;
  assign A_so[32] = \A_s[30] ;
  assign \A_s[30]  = A_s[30];
  assign A_nso[31] = \A_s[29] ;
  assign A_so[31] = \A_s[29] ;
  assign \A_s[29]  = A_s[29];
  assign A_nso[30] = \A_s[28] ;
  assign A_so[30] = \A_s[28] ;
  assign \A_s[28]  = A_s[28];
  assign A_nso[29] = \A_s[27] ;
  assign A_so[29] = \A_s[27] ;
  assign \A_s[27]  = A_s[27];
  assign A_nso[28] = \A_s[26] ;
  assign A_so[28] = \A_s[26] ;
  assign \A_s[26]  = A_s[26];
  assign A_nso[27] = \A_s[25] ;
  assign A_so[27] = \A_s[25] ;
  assign \A_s[25]  = A_s[25];
  assign A_nso[26] = \A_s[24] ;
  assign A_so[26] = \A_s[24] ;
  assign \A_s[24]  = A_s[24];
  assign A_nso[25] = \A_s[23] ;
  assign A_so[25] = \A_s[23] ;
  assign \A_s[23]  = A_s[23];
  assign A_nso[24] = \A_s[22] ;
  assign A_so[24] = \A_s[22] ;
  assign \A_s[22]  = A_s[22];
  assign A_nso[23] = \A_s[21] ;
  assign A_so[23] = \A_s[21] ;
  assign \A_s[21]  = A_s[21];
  assign A_nso[22] = \A_s[20] ;
  assign A_so[22] = \A_s[20] ;
  assign \A_s[20]  = A_s[20];
  assign A_nso[21] = \A_s[19] ;
  assign A_so[21] = \A_s[19] ;
  assign \A_s[19]  = A_s[19];
  assign A_nso[20] = \A_s[18] ;
  assign A_so[20] = \A_s[18] ;
  assign \A_s[18]  = A_s[18];
  assign A_nso[19] = \A_s[17] ;
  assign A_so[19] = \A_s[17] ;
  assign \A_s[17]  = A_s[17];
  assign A_nso[18] = \A_s[16] ;
  assign A_so[18] = \A_s[16] ;
  assign \A_s[16]  = A_s[16];
  assign A_nso[17] = \A_s[15] ;
  assign A_so[17] = \A_s[15] ;
  assign \A_s[15]  = A_s[15];
  assign A_nso[16] = \A_s[14] ;
  assign A_so[16] = \A_s[14] ;
  assign \A_s[14]  = A_s[14];
  assign A_nso[15] = \A_s[13] ;
  assign A_so[15] = \A_s[13] ;
  assign \A_s[13]  = A_s[13];
  assign A_nso[14] = \A_s[12] ;
  assign A_so[14] = \A_s[12] ;
  assign \A_s[12]  = A_s[12];
  assign A_nso[13] = \A_s[11] ;
  assign A_so[13] = \A_s[11] ;
  assign \A_s[11]  = A_s[11];
  assign A_nso[12] = \A_s[10] ;
  assign A_so[12] = \A_s[10] ;
  assign \A_s[10]  = A_s[10];
  assign A_nso[11] = \A_s[9] ;
  assign A_so[11] = \A_s[9] ;
  assign \A_s[9]  = A_s[9];
  assign A_nso[10] = \A_s[8] ;
  assign A_so[10] = \A_s[8] ;
  assign \A_s[8]  = A_s[8];
  assign A_nso[9] = \A_s[7] ;
  assign A_so[9] = \A_s[7] ;
  assign \A_s[7]  = A_s[7];
  assign A_nso[8] = \A_s[6] ;
  assign A_so[8] = \A_s[6] ;
  assign \A_s[6]  = A_s[6];
  assign A_nso[7] = \A_s[5] ;
  assign A_so[7] = \A_s[5] ;
  assign \A_s[5]  = A_s[5];
  assign A_nso[6] = \A_s[4] ;
  assign A_so[6] = \A_s[4] ;
  assign \A_s[4]  = A_s[4];
  assign A_nso[5] = \A_s[3] ;
  assign A_so[5] = \A_s[3] ;
  assign \A_s[3]  = A_s[3];
  assign A_nso[4] = \A_s[2] ;
  assign A_so[4] = \A_s[2] ;
  assign \A_s[2]  = A_s[2];
  assign A_nso[3] = \A_s[1] ;
  assign A_so[3] = \A_s[1] ;
  assign \A_s[1]  = A_s[1];
  assign A_nso[2] = \A_s[0] ;
  assign A_so[2] = \A_s[0] ;
  assign \A_s[0]  = A_s[0];

  AND3_X1 U2 ( .A1(B[4]), .A2(n585), .A3(B[3]), .ZN(n391) );
  INV_X4 U3 ( .A(n391), .ZN(n392) );
  INV_X4 U4 ( .A(n552), .ZN(n398) );
  OR3_X4 U5 ( .A1(B[3]), .A2(B[4]), .A3(n585), .ZN(n393) );
  INV_X4 U6 ( .A(n553), .ZN(n397) );
  OAI221_X1 U7 ( .B1(n393), .B2(n394), .C1(n392), .C2(n395), .A(n396), .ZN(
        O[9]) );
  AOI22_X1 U8 ( .A1(A_ns[8]), .A2(n397), .B1(\A_s[8] ), .B2(n398), .ZN(n396)
         );
  INV_X1 U9 ( .A(\A_s[7] ), .ZN(n395) );
  INV_X1 U10 ( .A(A_ns[7]), .ZN(n394) );
  OAI221_X1 U11 ( .B1(n393), .B2(n399), .C1(n392), .C2(n400), .A(n401), .ZN(
        O[8]) );
  AOI22_X1 U12 ( .A1(A_ns[7]), .A2(n397), .B1(\A_s[7] ), .B2(n398), .ZN(n401)
         );
  INV_X1 U13 ( .A(\A_s[6] ), .ZN(n400) );
  INV_X1 U14 ( .A(A_ns[6]), .ZN(n399) );
  OAI221_X1 U15 ( .B1(n393), .B2(n402), .C1(n392), .C2(n403), .A(n404), .ZN(
        O[7]) );
  AOI22_X1 U16 ( .A1(A_ns[6]), .A2(n397), .B1(\A_s[6] ), .B2(n398), .ZN(n404)
         );
  INV_X1 U17 ( .A(\A_s[5] ), .ZN(n403) );
  INV_X1 U18 ( .A(A_ns[5]), .ZN(n402) );
  OAI221_X1 U19 ( .B1(n393), .B2(n405), .C1(n392), .C2(n406), .A(n407), .ZN(
        O[6]) );
  AOI22_X1 U20 ( .A1(A_ns[5]), .A2(n397), .B1(\A_s[5] ), .B2(n398), .ZN(n407)
         );
  INV_X1 U21 ( .A(\A_s[4] ), .ZN(n406) );
  INV_X1 U22 ( .A(A_ns[4]), .ZN(n405) );
  OAI221_X1 U23 ( .B1(n393), .B2(n408), .C1(n392), .C2(n409), .A(n410), .ZN(
        O[63]) );
  AOI22_X1 U24 ( .A1(A_ns[62]), .A2(n397), .B1(A_s[62]), .B2(n398), .ZN(n410)
         );
  INV_X1 U25 ( .A(\A_s[61] ), .ZN(n409) );
  INV_X1 U26 ( .A(A_ns[61]), .ZN(n408) );
  OAI221_X1 U27 ( .B1(n393), .B2(n411), .C1(n392), .C2(n412), .A(n413), .ZN(
        O[62]) );
  AOI22_X1 U28 ( .A1(A_ns[61]), .A2(n397), .B1(\A_s[61] ), .B2(n398), .ZN(n413) );
  INV_X1 U29 ( .A(\A_s[60] ), .ZN(n412) );
  INV_X1 U30 ( .A(A_ns[60]), .ZN(n411) );
  OAI221_X1 U31 ( .B1(n393), .B2(n414), .C1(n392), .C2(n415), .A(n416), .ZN(
        O[61]) );
  AOI22_X1 U32 ( .A1(A_ns[60]), .A2(n397), .B1(\A_s[60] ), .B2(n398), .ZN(n416) );
  INV_X1 U33 ( .A(\A_s[59] ), .ZN(n415) );
  INV_X1 U34 ( .A(A_ns[59]), .ZN(n414) );
  OAI221_X1 U35 ( .B1(n393), .B2(n417), .C1(n392), .C2(n418), .A(n419), .ZN(
        O[60]) );
  AOI22_X1 U36 ( .A1(A_ns[59]), .A2(n397), .B1(\A_s[59] ), .B2(n398), .ZN(n419) );
  INV_X1 U37 ( .A(\A_s[58] ), .ZN(n418) );
  INV_X1 U38 ( .A(A_ns[58]), .ZN(n417) );
  OAI221_X1 U39 ( .B1(n393), .B2(n420), .C1(n392), .C2(n421), .A(n422), .ZN(
        O[5]) );
  AOI22_X1 U40 ( .A1(A_ns[4]), .A2(n397), .B1(\A_s[4] ), .B2(n398), .ZN(n422)
         );
  INV_X1 U41 ( .A(\A_s[3] ), .ZN(n421) );
  INV_X1 U42 ( .A(A_ns[3]), .ZN(n420) );
  OAI221_X1 U43 ( .B1(n393), .B2(n423), .C1(n392), .C2(n424), .A(n425), .ZN(
        O[59]) );
  AOI22_X1 U44 ( .A1(A_ns[58]), .A2(n397), .B1(\A_s[58] ), .B2(n398), .ZN(n425) );
  INV_X1 U45 ( .A(\A_s[57] ), .ZN(n424) );
  INV_X1 U46 ( .A(A_ns[57]), .ZN(n423) );
  OAI221_X1 U47 ( .B1(n393), .B2(n426), .C1(n392), .C2(n427), .A(n428), .ZN(
        O[58]) );
  AOI22_X1 U48 ( .A1(A_ns[57]), .A2(n397), .B1(\A_s[57] ), .B2(n398), .ZN(n428) );
  INV_X1 U49 ( .A(\A_s[56] ), .ZN(n427) );
  INV_X1 U50 ( .A(A_ns[56]), .ZN(n426) );
  OAI221_X1 U51 ( .B1(n393), .B2(n429), .C1(n392), .C2(n430), .A(n431), .ZN(
        O[57]) );
  AOI22_X1 U52 ( .A1(A_ns[56]), .A2(n397), .B1(\A_s[56] ), .B2(n398), .ZN(n431) );
  INV_X1 U53 ( .A(\A_s[55] ), .ZN(n430) );
  INV_X1 U54 ( .A(A_ns[55]), .ZN(n429) );
  OAI221_X1 U55 ( .B1(n393), .B2(n432), .C1(n392), .C2(n433), .A(n434), .ZN(
        O[56]) );
  AOI22_X1 U56 ( .A1(A_ns[55]), .A2(n397), .B1(\A_s[55] ), .B2(n398), .ZN(n434) );
  INV_X1 U57 ( .A(\A_s[54] ), .ZN(n433) );
  INV_X1 U58 ( .A(A_ns[54]), .ZN(n432) );
  OAI221_X1 U59 ( .B1(n393), .B2(n435), .C1(n392), .C2(n436), .A(n437), .ZN(
        O[55]) );
  AOI22_X1 U60 ( .A1(A_ns[54]), .A2(n397), .B1(\A_s[54] ), .B2(n398), .ZN(n437) );
  INV_X1 U61 ( .A(\A_s[53] ), .ZN(n436) );
  INV_X1 U62 ( .A(A_ns[53]), .ZN(n435) );
  OAI221_X1 U63 ( .B1(n393), .B2(n438), .C1(n392), .C2(n439), .A(n440), .ZN(
        O[54]) );
  AOI22_X1 U64 ( .A1(A_ns[53]), .A2(n397), .B1(\A_s[53] ), .B2(n398), .ZN(n440) );
  INV_X1 U65 ( .A(\A_s[52] ), .ZN(n439) );
  INV_X1 U66 ( .A(A_ns[52]), .ZN(n438) );
  OAI221_X1 U67 ( .B1(n393), .B2(n441), .C1(n392), .C2(n442), .A(n443), .ZN(
        O[53]) );
  AOI22_X1 U68 ( .A1(A_ns[52]), .A2(n397), .B1(\A_s[52] ), .B2(n398), .ZN(n443) );
  INV_X1 U69 ( .A(\A_s[51] ), .ZN(n442) );
  INV_X1 U70 ( .A(A_ns[51]), .ZN(n441) );
  OAI221_X1 U71 ( .B1(n393), .B2(n444), .C1(n392), .C2(n445), .A(n446), .ZN(
        O[52]) );
  AOI22_X1 U72 ( .A1(A_ns[51]), .A2(n397), .B1(\A_s[51] ), .B2(n398), .ZN(n446) );
  INV_X1 U73 ( .A(\A_s[50] ), .ZN(n445) );
  INV_X1 U74 ( .A(A_ns[50]), .ZN(n444) );
  OAI221_X1 U75 ( .B1(n393), .B2(n447), .C1(n392), .C2(n448), .A(n449), .ZN(
        O[51]) );
  AOI22_X1 U76 ( .A1(A_ns[50]), .A2(n397), .B1(\A_s[50] ), .B2(n398), .ZN(n449) );
  INV_X1 U77 ( .A(\A_s[49] ), .ZN(n448) );
  INV_X1 U78 ( .A(A_ns[49]), .ZN(n447) );
  OAI221_X1 U79 ( .B1(n393), .B2(n450), .C1(n392), .C2(n451), .A(n452), .ZN(
        O[50]) );
  AOI22_X1 U80 ( .A1(A_ns[49]), .A2(n397), .B1(\A_s[49] ), .B2(n398), .ZN(n452) );
  INV_X1 U81 ( .A(\A_s[48] ), .ZN(n451) );
  INV_X1 U82 ( .A(A_ns[48]), .ZN(n450) );
  OAI221_X1 U83 ( .B1(n393), .B2(n453), .C1(n392), .C2(n454), .A(n455), .ZN(
        O[4]) );
  AOI22_X1 U84 ( .A1(A_ns[3]), .A2(n397), .B1(\A_s[3] ), .B2(n398), .ZN(n455)
         );
  INV_X1 U85 ( .A(\A_s[2] ), .ZN(n454) );
  INV_X1 U86 ( .A(A_ns[2]), .ZN(n453) );
  OAI221_X1 U87 ( .B1(n393), .B2(n456), .C1(n392), .C2(n457), .A(n458), .ZN(
        O[49]) );
  AOI22_X1 U88 ( .A1(A_ns[48]), .A2(n397), .B1(\A_s[48] ), .B2(n398), .ZN(n458) );
  INV_X1 U89 ( .A(\A_s[47] ), .ZN(n457) );
  INV_X1 U90 ( .A(A_ns[47]), .ZN(n456) );
  OAI221_X1 U91 ( .B1(n393), .B2(n459), .C1(n392), .C2(n460), .A(n461), .ZN(
        O[48]) );
  AOI22_X1 U92 ( .A1(A_ns[47]), .A2(n397), .B1(\A_s[47] ), .B2(n398), .ZN(n461) );
  INV_X1 U93 ( .A(\A_s[46] ), .ZN(n460) );
  INV_X1 U94 ( .A(A_ns[46]), .ZN(n459) );
  OAI221_X1 U95 ( .B1(n393), .B2(n462), .C1(n392), .C2(n463), .A(n464), .ZN(
        O[47]) );
  AOI22_X1 U96 ( .A1(A_ns[46]), .A2(n397), .B1(\A_s[46] ), .B2(n398), .ZN(n464) );
  INV_X1 U97 ( .A(\A_s[45] ), .ZN(n463) );
  INV_X1 U98 ( .A(A_ns[45]), .ZN(n462) );
  OAI221_X1 U99 ( .B1(n393), .B2(n465), .C1(n392), .C2(n466), .A(n467), .ZN(
        O[46]) );
  AOI22_X1 U100 ( .A1(A_ns[45]), .A2(n397), .B1(\A_s[45] ), .B2(n398), .ZN(
        n467) );
  INV_X1 U101 ( .A(\A_s[44] ), .ZN(n466) );
  INV_X1 U102 ( .A(A_ns[44]), .ZN(n465) );
  OAI221_X1 U103 ( .B1(n393), .B2(n468), .C1(n392), .C2(n469), .A(n470), .ZN(
        O[45]) );
  AOI22_X1 U104 ( .A1(A_ns[44]), .A2(n397), .B1(\A_s[44] ), .B2(n398), .ZN(
        n470) );
  INV_X1 U105 ( .A(\A_s[43] ), .ZN(n469) );
  INV_X1 U106 ( .A(A_ns[43]), .ZN(n468) );
  OAI221_X1 U107 ( .B1(n393), .B2(n471), .C1(n392), .C2(n472), .A(n473), .ZN(
        O[44]) );
  AOI22_X1 U108 ( .A1(A_ns[43]), .A2(n397), .B1(\A_s[43] ), .B2(n398), .ZN(
        n473) );
  INV_X1 U109 ( .A(\A_s[42] ), .ZN(n472) );
  INV_X1 U110 ( .A(A_ns[42]), .ZN(n471) );
  OAI221_X1 U111 ( .B1(n393), .B2(n474), .C1(n392), .C2(n475), .A(n476), .ZN(
        O[43]) );
  AOI22_X1 U112 ( .A1(A_ns[42]), .A2(n397), .B1(\A_s[42] ), .B2(n398), .ZN(
        n476) );
  INV_X1 U113 ( .A(\A_s[41] ), .ZN(n475) );
  INV_X1 U114 ( .A(A_ns[41]), .ZN(n474) );
  OAI221_X1 U115 ( .B1(n393), .B2(n477), .C1(n392), .C2(n478), .A(n479), .ZN(
        O[42]) );
  AOI22_X1 U116 ( .A1(A_ns[41]), .A2(n397), .B1(\A_s[41] ), .B2(n398), .ZN(
        n479) );
  INV_X1 U117 ( .A(\A_s[40] ), .ZN(n478) );
  INV_X1 U118 ( .A(A_ns[40]), .ZN(n477) );
  OAI221_X1 U119 ( .B1(n393), .B2(n480), .C1(n392), .C2(n481), .A(n482), .ZN(
        O[41]) );
  AOI22_X1 U120 ( .A1(A_ns[40]), .A2(n397), .B1(\A_s[40] ), .B2(n398), .ZN(
        n482) );
  INV_X1 U121 ( .A(\A_s[39] ), .ZN(n481) );
  INV_X1 U122 ( .A(A_ns[39]), .ZN(n480) );
  OAI221_X1 U123 ( .B1(n393), .B2(n483), .C1(n392), .C2(n484), .A(n485), .ZN(
        O[40]) );
  AOI22_X1 U124 ( .A1(A_ns[39]), .A2(n397), .B1(\A_s[39] ), .B2(n398), .ZN(
        n485) );
  INV_X1 U125 ( .A(\A_s[38] ), .ZN(n484) );
  INV_X1 U126 ( .A(A_ns[38]), .ZN(n483) );
  OAI221_X1 U127 ( .B1(n393), .B2(n486), .C1(n392), .C2(n487), .A(n488), .ZN(
        O[3]) );
  AOI22_X1 U128 ( .A1(A_ns[2]), .A2(n397), .B1(\A_s[2] ), .B2(n398), .ZN(n488)
         );
  INV_X1 U129 ( .A(\A_s[1] ), .ZN(n487) );
  INV_X1 U130 ( .A(A_ns[1]), .ZN(n486) );
  OAI221_X1 U131 ( .B1(n393), .B2(n489), .C1(n392), .C2(n490), .A(n491), .ZN(
        O[39]) );
  AOI22_X1 U132 ( .A1(A_ns[38]), .A2(n397), .B1(\A_s[38] ), .B2(n398), .ZN(
        n491) );
  INV_X1 U133 ( .A(\A_s[37] ), .ZN(n490) );
  INV_X1 U134 ( .A(A_ns[37]), .ZN(n489) );
  OAI221_X1 U135 ( .B1(n393), .B2(n492), .C1(n392), .C2(n493), .A(n494), .ZN(
        O[38]) );
  AOI22_X1 U136 ( .A1(A_ns[37]), .A2(n397), .B1(\A_s[37] ), .B2(n398), .ZN(
        n494) );
  INV_X1 U137 ( .A(\A_s[36] ), .ZN(n493) );
  INV_X1 U138 ( .A(A_ns[36]), .ZN(n492) );
  OAI221_X1 U139 ( .B1(n393), .B2(n495), .C1(n392), .C2(n496), .A(n497), .ZN(
        O[37]) );
  AOI22_X1 U140 ( .A1(A_ns[36]), .A2(n397), .B1(\A_s[36] ), .B2(n398), .ZN(
        n497) );
  INV_X1 U141 ( .A(\A_s[35] ), .ZN(n496) );
  INV_X1 U142 ( .A(A_ns[35]), .ZN(n495) );
  OAI221_X1 U143 ( .B1(n393), .B2(n498), .C1(n392), .C2(n499), .A(n500), .ZN(
        O[36]) );
  AOI22_X1 U144 ( .A1(A_ns[35]), .A2(n397), .B1(\A_s[35] ), .B2(n398), .ZN(
        n500) );
  INV_X1 U145 ( .A(\A_s[34] ), .ZN(n499) );
  INV_X1 U146 ( .A(A_ns[34]), .ZN(n498) );
  OAI221_X1 U147 ( .B1(n393), .B2(n501), .C1(n392), .C2(n502), .A(n503), .ZN(
        O[35]) );
  AOI22_X1 U148 ( .A1(A_ns[34]), .A2(n397), .B1(\A_s[34] ), .B2(n398), .ZN(
        n503) );
  INV_X1 U149 ( .A(\A_s[33] ), .ZN(n502) );
  INV_X1 U150 ( .A(A_ns[33]), .ZN(n501) );
  OAI221_X1 U151 ( .B1(n393), .B2(n504), .C1(n392), .C2(n505), .A(n506), .ZN(
        O[34]) );
  AOI22_X1 U152 ( .A1(A_ns[33]), .A2(n397), .B1(\A_s[33] ), .B2(n398), .ZN(
        n506) );
  INV_X1 U153 ( .A(\A_s[32] ), .ZN(n505) );
  INV_X1 U154 ( .A(A_ns[32]), .ZN(n504) );
  OAI221_X1 U155 ( .B1(n393), .B2(n507), .C1(n392), .C2(n508), .A(n509), .ZN(
        O[33]) );
  AOI22_X1 U156 ( .A1(A_ns[32]), .A2(n397), .B1(\A_s[32] ), .B2(n398), .ZN(
        n509) );
  INV_X1 U157 ( .A(\A_s[31] ), .ZN(n508) );
  INV_X1 U158 ( .A(A_ns[31]), .ZN(n507) );
  OAI221_X1 U159 ( .B1(n393), .B2(n510), .C1(n392), .C2(n511), .A(n512), .ZN(
        O[32]) );
  AOI22_X1 U160 ( .A1(A_ns[31]), .A2(n397), .B1(\A_s[31] ), .B2(n398), .ZN(
        n512) );
  INV_X1 U161 ( .A(\A_s[30] ), .ZN(n511) );
  INV_X1 U162 ( .A(A_ns[30]), .ZN(n510) );
  OAI221_X1 U163 ( .B1(n393), .B2(n513), .C1(n392), .C2(n514), .A(n515), .ZN(
        O[31]) );
  AOI22_X1 U164 ( .A1(A_ns[30]), .A2(n397), .B1(\A_s[30] ), .B2(n398), .ZN(
        n515) );
  INV_X1 U165 ( .A(\A_s[29] ), .ZN(n514) );
  INV_X1 U166 ( .A(A_ns[29]), .ZN(n513) );
  OAI221_X1 U167 ( .B1(n393), .B2(n516), .C1(n392), .C2(n517), .A(n518), .ZN(
        O[30]) );
  AOI22_X1 U168 ( .A1(A_ns[29]), .A2(n397), .B1(\A_s[29] ), .B2(n398), .ZN(
        n518) );
  INV_X1 U169 ( .A(\A_s[28] ), .ZN(n517) );
  INV_X1 U170 ( .A(A_ns[28]), .ZN(n516) );
  OAI221_X1 U171 ( .B1(n393), .B2(n519), .C1(n392), .C2(n520), .A(n521), .ZN(
        O[2]) );
  AOI22_X1 U172 ( .A1(A_ns[1]), .A2(n397), .B1(\A_s[1] ), .B2(n398), .ZN(n521)
         );
  OAI221_X1 U173 ( .B1(n393), .B2(n522), .C1(n392), .C2(n523), .A(n524), .ZN(
        O[29]) );
  AOI22_X1 U174 ( .A1(A_ns[28]), .A2(n397), .B1(\A_s[28] ), .B2(n398), .ZN(
        n524) );
  INV_X1 U175 ( .A(\A_s[27] ), .ZN(n523) );
  INV_X1 U176 ( .A(A_ns[27]), .ZN(n522) );
  OAI221_X1 U177 ( .B1(n393), .B2(n525), .C1(n392), .C2(n526), .A(n527), .ZN(
        O[28]) );
  AOI22_X1 U178 ( .A1(A_ns[27]), .A2(n397), .B1(\A_s[27] ), .B2(n398), .ZN(
        n527) );
  INV_X1 U179 ( .A(\A_s[26] ), .ZN(n526) );
  INV_X1 U180 ( .A(A_ns[26]), .ZN(n525) );
  OAI221_X1 U181 ( .B1(n393), .B2(n528), .C1(n392), .C2(n529), .A(n530), .ZN(
        O[27]) );
  AOI22_X1 U182 ( .A1(A_ns[26]), .A2(n397), .B1(\A_s[26] ), .B2(n398), .ZN(
        n530) );
  INV_X1 U183 ( .A(\A_s[25] ), .ZN(n529) );
  INV_X1 U184 ( .A(A_ns[25]), .ZN(n528) );
  OAI221_X1 U185 ( .B1(n393), .B2(n531), .C1(n392), .C2(n532), .A(n533), .ZN(
        O[26]) );
  AOI22_X1 U186 ( .A1(A_ns[25]), .A2(n397), .B1(\A_s[25] ), .B2(n398), .ZN(
        n533) );
  INV_X1 U187 ( .A(\A_s[24] ), .ZN(n532) );
  INV_X1 U188 ( .A(A_ns[24]), .ZN(n531) );
  OAI221_X1 U189 ( .B1(n393), .B2(n534), .C1(n392), .C2(n535), .A(n536), .ZN(
        O[25]) );
  AOI22_X1 U190 ( .A1(A_ns[24]), .A2(n397), .B1(\A_s[24] ), .B2(n398), .ZN(
        n536) );
  INV_X1 U191 ( .A(\A_s[23] ), .ZN(n535) );
  INV_X1 U192 ( .A(A_ns[23]), .ZN(n534) );
  OAI221_X1 U193 ( .B1(n393), .B2(n537), .C1(n392), .C2(n538), .A(n539), .ZN(
        O[24]) );
  AOI22_X1 U194 ( .A1(A_ns[23]), .A2(n397), .B1(\A_s[23] ), .B2(n398), .ZN(
        n539) );
  INV_X1 U195 ( .A(\A_s[22] ), .ZN(n538) );
  INV_X1 U196 ( .A(A_ns[22]), .ZN(n537) );
  OAI221_X1 U197 ( .B1(n393), .B2(n540), .C1(n392), .C2(n541), .A(n542), .ZN(
        O[23]) );
  AOI22_X1 U198 ( .A1(A_ns[22]), .A2(n397), .B1(\A_s[22] ), .B2(n398), .ZN(
        n542) );
  INV_X1 U199 ( .A(\A_s[21] ), .ZN(n541) );
  INV_X1 U200 ( .A(A_ns[21]), .ZN(n540) );
  OAI221_X1 U201 ( .B1(n393), .B2(n543), .C1(n392), .C2(n544), .A(n545), .ZN(
        O[22]) );
  AOI22_X1 U202 ( .A1(A_ns[21]), .A2(n397), .B1(\A_s[21] ), .B2(n398), .ZN(
        n545) );
  INV_X1 U203 ( .A(\A_s[20] ), .ZN(n544) );
  INV_X1 U204 ( .A(A_ns[20]), .ZN(n543) );
  OAI221_X1 U205 ( .B1(n393), .B2(n546), .C1(n392), .C2(n547), .A(n548), .ZN(
        O[21]) );
  AOI22_X1 U206 ( .A1(A_ns[20]), .A2(n397), .B1(\A_s[20] ), .B2(n398), .ZN(
        n548) );
  INV_X1 U207 ( .A(\A_s[19] ), .ZN(n547) );
  INV_X1 U208 ( .A(A_ns[19]), .ZN(n546) );
  OAI221_X1 U209 ( .B1(n393), .B2(n549), .C1(n392), .C2(n550), .A(n551), .ZN(
        O[20]) );
  AOI22_X1 U210 ( .A1(A_ns[19]), .A2(n397), .B1(\A_s[19] ), .B2(n398), .ZN(
        n551) );
  INV_X1 U211 ( .A(\A_s[18] ), .ZN(n550) );
  INV_X1 U212 ( .A(A_ns[18]), .ZN(n549) );
  OAI22_X1 U213 ( .A1(n552), .A2(n520), .B1(n553), .B2(n519), .ZN(O[1]) );
  INV_X1 U214 ( .A(A_ns[0]), .ZN(n519) );
  INV_X1 U215 ( .A(\A_s[0] ), .ZN(n520) );
  OAI221_X1 U216 ( .B1(n393), .B2(n554), .C1(n392), .C2(n555), .A(n556), .ZN(
        O[19]) );
  AOI22_X1 U217 ( .A1(A_ns[18]), .A2(n397), .B1(\A_s[18] ), .B2(n398), .ZN(
        n556) );
  INV_X1 U218 ( .A(\A_s[17] ), .ZN(n555) );
  INV_X1 U219 ( .A(A_ns[17]), .ZN(n554) );
  OAI221_X1 U220 ( .B1(n393), .B2(n557), .C1(n392), .C2(n558), .A(n559), .ZN(
        O[18]) );
  AOI22_X1 U221 ( .A1(A_ns[17]), .A2(n397), .B1(\A_s[17] ), .B2(n398), .ZN(
        n559) );
  INV_X1 U222 ( .A(\A_s[16] ), .ZN(n558) );
  INV_X1 U223 ( .A(A_ns[16]), .ZN(n557) );
  OAI221_X1 U224 ( .B1(n393), .B2(n560), .C1(n392), .C2(n561), .A(n562), .ZN(
        O[17]) );
  AOI22_X1 U225 ( .A1(A_ns[16]), .A2(n397), .B1(\A_s[16] ), .B2(n398), .ZN(
        n562) );
  INV_X1 U226 ( .A(\A_s[15] ), .ZN(n561) );
  INV_X1 U227 ( .A(A_ns[15]), .ZN(n560) );
  OAI221_X1 U228 ( .B1(n393), .B2(n563), .C1(n392), .C2(n564), .A(n565), .ZN(
        O[16]) );
  AOI22_X1 U229 ( .A1(A_ns[15]), .A2(n397), .B1(\A_s[15] ), .B2(n398), .ZN(
        n565) );
  INV_X1 U230 ( .A(\A_s[14] ), .ZN(n564) );
  INV_X1 U231 ( .A(A_ns[14]), .ZN(n563) );
  OAI221_X1 U232 ( .B1(n393), .B2(n566), .C1(n392), .C2(n567), .A(n568), .ZN(
        O[15]) );
  AOI22_X1 U233 ( .A1(A_ns[14]), .A2(n397), .B1(\A_s[14] ), .B2(n398), .ZN(
        n568) );
  INV_X1 U234 ( .A(\A_s[13] ), .ZN(n567) );
  INV_X1 U235 ( .A(A_ns[13]), .ZN(n566) );
  OAI221_X1 U236 ( .B1(n393), .B2(n569), .C1(n392), .C2(n570), .A(n571), .ZN(
        O[14]) );
  AOI22_X1 U237 ( .A1(A_ns[13]), .A2(n397), .B1(\A_s[13] ), .B2(n398), .ZN(
        n571) );
  INV_X1 U238 ( .A(\A_s[12] ), .ZN(n570) );
  INV_X1 U239 ( .A(A_ns[12]), .ZN(n569) );
  OAI221_X1 U240 ( .B1(n393), .B2(n572), .C1(n392), .C2(n573), .A(n574), .ZN(
        O[13]) );
  AOI22_X1 U241 ( .A1(A_ns[12]), .A2(n397), .B1(\A_s[12] ), .B2(n398), .ZN(
        n574) );
  INV_X1 U242 ( .A(\A_s[11] ), .ZN(n573) );
  INV_X1 U243 ( .A(A_ns[11]), .ZN(n572) );
  OAI221_X1 U244 ( .B1(n393), .B2(n575), .C1(n392), .C2(n576), .A(n577), .ZN(
        O[12]) );
  AOI22_X1 U245 ( .A1(A_ns[11]), .A2(n397), .B1(\A_s[11] ), .B2(n398), .ZN(
        n577) );
  INV_X1 U246 ( .A(\A_s[10] ), .ZN(n576) );
  INV_X1 U247 ( .A(A_ns[10]), .ZN(n575) );
  OAI221_X1 U248 ( .B1(n393), .B2(n578), .C1(n392), .C2(n579), .A(n580), .ZN(
        O[11]) );
  AOI22_X1 U249 ( .A1(A_ns[10]), .A2(n397), .B1(\A_s[10] ), .B2(n398), .ZN(
        n580) );
  INV_X1 U250 ( .A(\A_s[9] ), .ZN(n579) );
  INV_X1 U251 ( .A(A_ns[9]), .ZN(n578) );
  OAI221_X1 U252 ( .B1(n581), .B2(n393), .C1(n582), .C2(n392), .A(n583), .ZN(
        O[10]) );
  AOI22_X1 U253 ( .A1(A_ns[9]), .A2(n397), .B1(\A_s[9] ), .B2(n398), .ZN(n583)
         );
  NAND2_X1 U254 ( .A1(n584), .A2(n552), .ZN(n553) );
  NAND2_X1 U255 ( .A1(n584), .A2(n585), .ZN(n552) );
  XOR2_X1 U256 ( .A(B[3]), .B(B[4]), .Z(n584) );
  INV_X1 U257 ( .A(\A_s[8] ), .ZN(n582) );
  INV_X1 U258 ( .A(B[5]), .ZN(n585) );
  INV_X1 U259 ( .A(A_ns[8]), .ZN(n581) );
endmodule


module BOOTHENC_NBIT64_i6 ( A, A_n, A_ns, A_s, B, O, A_so, A_nso );
  input [63:0] A;
  input [63:0] A_n;
  input [63:0] A_ns;
  input [63:0] A_s;
  input [63:0] B;
  output [63:0] O;
  output [63:0] A_so;
  output [63:0] A_nso;
  wire   \A_s[61] , \A_s[60] , \A_s[59] , \A_s[58] , \A_s[57] , \A_s[56] ,
         \A_s[55] , \A_s[54] , \A_s[53] , \A_s[52] , \A_s[51] , \A_s[50] ,
         \A_s[49] , \A_s[48] , \A_s[47] , \A_s[46] , \A_s[45] , \A_s[44] ,
         \A_s[43] , \A_s[42] , \A_s[41] , \A_s[40] , \A_s[39] , \A_s[38] ,
         \A_s[37] , \A_s[36] , \A_s[35] , \A_s[34] , \A_s[33] , \A_s[32] ,
         \A_s[31] , \A_s[30] , \A_s[29] , \A_s[28] , \A_s[27] , \A_s[26] ,
         \A_s[25] , \A_s[24] , \A_s[23] , \A_s[22] , \A_s[21] , \A_s[20] ,
         \A_s[19] , \A_s[18] , \A_s[17] , \A_s[16] , \A_s[15] , \A_s[14] ,
         \A_s[13] , \A_s[12] , \A_s[11] , \A_s[10] , \A_s[9] , \A_s[8] ,
         \A_s[7] , \A_s[6] , \A_s[5] , \A_s[4] , \A_s[3] , \A_s[2] , \A_s[1] ,
         \A_s[0] , n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585;
  assign A_nso[0] = 1'b0;
  assign A_nso[1] = 1'b0;
  assign A_so[0] = 1'b0;
  assign A_so[1] = 1'b0;
  assign O[0] = 1'b0;
  assign A_nso[63] = \A_s[61] ;
  assign A_so[63] = \A_s[61] ;
  assign \A_s[61]  = A_s[61];
  assign A_nso[62] = \A_s[60] ;
  assign A_so[62] = \A_s[60] ;
  assign \A_s[60]  = A_s[60];
  assign A_nso[61] = \A_s[59] ;
  assign A_so[61] = \A_s[59] ;
  assign \A_s[59]  = A_s[59];
  assign A_nso[60] = \A_s[58] ;
  assign A_so[60] = \A_s[58] ;
  assign \A_s[58]  = A_s[58];
  assign A_nso[59] = \A_s[57] ;
  assign A_so[59] = \A_s[57] ;
  assign \A_s[57]  = A_s[57];
  assign A_nso[58] = \A_s[56] ;
  assign A_so[58] = \A_s[56] ;
  assign \A_s[56]  = A_s[56];
  assign A_nso[57] = \A_s[55] ;
  assign A_so[57] = \A_s[55] ;
  assign \A_s[55]  = A_s[55];
  assign A_nso[56] = \A_s[54] ;
  assign A_so[56] = \A_s[54] ;
  assign \A_s[54]  = A_s[54];
  assign A_nso[55] = \A_s[53] ;
  assign A_so[55] = \A_s[53] ;
  assign \A_s[53]  = A_s[53];
  assign A_nso[54] = \A_s[52] ;
  assign A_so[54] = \A_s[52] ;
  assign \A_s[52]  = A_s[52];
  assign A_nso[53] = \A_s[51] ;
  assign A_so[53] = \A_s[51] ;
  assign \A_s[51]  = A_s[51];
  assign A_nso[52] = \A_s[50] ;
  assign A_so[52] = \A_s[50] ;
  assign \A_s[50]  = A_s[50];
  assign A_nso[51] = \A_s[49] ;
  assign A_so[51] = \A_s[49] ;
  assign \A_s[49]  = A_s[49];
  assign A_nso[50] = \A_s[48] ;
  assign A_so[50] = \A_s[48] ;
  assign \A_s[48]  = A_s[48];
  assign A_nso[49] = \A_s[47] ;
  assign A_so[49] = \A_s[47] ;
  assign \A_s[47]  = A_s[47];
  assign A_nso[48] = \A_s[46] ;
  assign A_so[48] = \A_s[46] ;
  assign \A_s[46]  = A_s[46];
  assign A_nso[47] = \A_s[45] ;
  assign A_so[47] = \A_s[45] ;
  assign \A_s[45]  = A_s[45];
  assign A_nso[46] = \A_s[44] ;
  assign A_so[46] = \A_s[44] ;
  assign \A_s[44]  = A_s[44];
  assign A_nso[45] = \A_s[43] ;
  assign A_so[45] = \A_s[43] ;
  assign \A_s[43]  = A_s[43];
  assign A_nso[44] = \A_s[42] ;
  assign A_so[44] = \A_s[42] ;
  assign \A_s[42]  = A_s[42];
  assign A_nso[43] = \A_s[41] ;
  assign A_so[43] = \A_s[41] ;
  assign \A_s[41]  = A_s[41];
  assign A_nso[42] = \A_s[40] ;
  assign A_so[42] = \A_s[40] ;
  assign \A_s[40]  = A_s[40];
  assign A_nso[41] = \A_s[39] ;
  assign A_so[41] = \A_s[39] ;
  assign \A_s[39]  = A_s[39];
  assign A_nso[40] = \A_s[38] ;
  assign A_so[40] = \A_s[38] ;
  assign \A_s[38]  = A_s[38];
  assign A_nso[39] = \A_s[37] ;
  assign A_so[39] = \A_s[37] ;
  assign \A_s[37]  = A_s[37];
  assign A_nso[38] = \A_s[36] ;
  assign A_so[38] = \A_s[36] ;
  assign \A_s[36]  = A_s[36];
  assign A_nso[37] = \A_s[35] ;
  assign A_so[37] = \A_s[35] ;
  assign \A_s[35]  = A_s[35];
  assign A_nso[36] = \A_s[34] ;
  assign A_so[36] = \A_s[34] ;
  assign \A_s[34]  = A_s[34];
  assign A_nso[35] = \A_s[33] ;
  assign A_so[35] = \A_s[33] ;
  assign \A_s[33]  = A_s[33];
  assign A_nso[34] = \A_s[32] ;
  assign A_so[34] = \A_s[32] ;
  assign \A_s[32]  = A_s[32];
  assign A_nso[33] = \A_s[31] ;
  assign A_so[33] = \A_s[31] ;
  assign \A_s[31]  = A_s[31];
  assign A_nso[32] = \A_s[30] ;
  assign A_so[32] = \A_s[30] ;
  assign \A_s[30]  = A_s[30];
  assign A_nso[31] = \A_s[29] ;
  assign A_so[31] = \A_s[29] ;
  assign \A_s[29]  = A_s[29];
  assign A_nso[30] = \A_s[28] ;
  assign A_so[30] = \A_s[28] ;
  assign \A_s[28]  = A_s[28];
  assign A_nso[29] = \A_s[27] ;
  assign A_so[29] = \A_s[27] ;
  assign \A_s[27]  = A_s[27];
  assign A_nso[28] = \A_s[26] ;
  assign A_so[28] = \A_s[26] ;
  assign \A_s[26]  = A_s[26];
  assign A_nso[27] = \A_s[25] ;
  assign A_so[27] = \A_s[25] ;
  assign \A_s[25]  = A_s[25];
  assign A_nso[26] = \A_s[24] ;
  assign A_so[26] = \A_s[24] ;
  assign \A_s[24]  = A_s[24];
  assign A_nso[25] = \A_s[23] ;
  assign A_so[25] = \A_s[23] ;
  assign \A_s[23]  = A_s[23];
  assign A_nso[24] = \A_s[22] ;
  assign A_so[24] = \A_s[22] ;
  assign \A_s[22]  = A_s[22];
  assign A_nso[23] = \A_s[21] ;
  assign A_so[23] = \A_s[21] ;
  assign \A_s[21]  = A_s[21];
  assign A_nso[22] = \A_s[20] ;
  assign A_so[22] = \A_s[20] ;
  assign \A_s[20]  = A_s[20];
  assign A_nso[21] = \A_s[19] ;
  assign A_so[21] = \A_s[19] ;
  assign \A_s[19]  = A_s[19];
  assign A_nso[20] = \A_s[18] ;
  assign A_so[20] = \A_s[18] ;
  assign \A_s[18]  = A_s[18];
  assign A_nso[19] = \A_s[17] ;
  assign A_so[19] = \A_s[17] ;
  assign \A_s[17]  = A_s[17];
  assign A_nso[18] = \A_s[16] ;
  assign A_so[18] = \A_s[16] ;
  assign \A_s[16]  = A_s[16];
  assign A_nso[17] = \A_s[15] ;
  assign A_so[17] = \A_s[15] ;
  assign \A_s[15]  = A_s[15];
  assign A_nso[16] = \A_s[14] ;
  assign A_so[16] = \A_s[14] ;
  assign \A_s[14]  = A_s[14];
  assign A_nso[15] = \A_s[13] ;
  assign A_so[15] = \A_s[13] ;
  assign \A_s[13]  = A_s[13];
  assign A_nso[14] = \A_s[12] ;
  assign A_so[14] = \A_s[12] ;
  assign \A_s[12]  = A_s[12];
  assign A_nso[13] = \A_s[11] ;
  assign A_so[13] = \A_s[11] ;
  assign \A_s[11]  = A_s[11];
  assign A_nso[12] = \A_s[10] ;
  assign A_so[12] = \A_s[10] ;
  assign \A_s[10]  = A_s[10];
  assign A_nso[11] = \A_s[9] ;
  assign A_so[11] = \A_s[9] ;
  assign \A_s[9]  = A_s[9];
  assign A_nso[10] = \A_s[8] ;
  assign A_so[10] = \A_s[8] ;
  assign \A_s[8]  = A_s[8];
  assign A_nso[9] = \A_s[7] ;
  assign A_so[9] = \A_s[7] ;
  assign \A_s[7]  = A_s[7];
  assign A_nso[8] = \A_s[6] ;
  assign A_so[8] = \A_s[6] ;
  assign \A_s[6]  = A_s[6];
  assign A_nso[7] = \A_s[5] ;
  assign A_so[7] = \A_s[5] ;
  assign \A_s[5]  = A_s[5];
  assign A_nso[6] = \A_s[4] ;
  assign A_so[6] = \A_s[4] ;
  assign \A_s[4]  = A_s[4];
  assign A_nso[5] = \A_s[3] ;
  assign A_so[5] = \A_s[3] ;
  assign \A_s[3]  = A_s[3];
  assign A_nso[4] = \A_s[2] ;
  assign A_so[4] = \A_s[2] ;
  assign \A_s[2]  = A_s[2];
  assign A_nso[3] = \A_s[1] ;
  assign A_so[3] = \A_s[1] ;
  assign \A_s[1]  = A_s[1];
  assign A_nso[2] = \A_s[0] ;
  assign A_so[2] = \A_s[0] ;
  assign \A_s[0]  = A_s[0];

  AND3_X1 U2 ( .A1(B[6]), .A2(n585), .A3(B[5]), .ZN(n391) );
  INV_X4 U3 ( .A(n391), .ZN(n392) );
  INV_X4 U4 ( .A(n552), .ZN(n398) );
  OR3_X4 U5 ( .A1(B[5]), .A2(B[6]), .A3(n585), .ZN(n393) );
  INV_X4 U6 ( .A(n553), .ZN(n397) );
  OAI221_X1 U7 ( .B1(n393), .B2(n394), .C1(n392), .C2(n395), .A(n396), .ZN(
        O[9]) );
  AOI22_X1 U8 ( .A1(A_ns[8]), .A2(n397), .B1(\A_s[8] ), .B2(n398), .ZN(n396)
         );
  INV_X1 U9 ( .A(\A_s[7] ), .ZN(n395) );
  INV_X1 U10 ( .A(A_ns[7]), .ZN(n394) );
  OAI221_X1 U11 ( .B1(n393), .B2(n399), .C1(n392), .C2(n400), .A(n401), .ZN(
        O[8]) );
  AOI22_X1 U12 ( .A1(A_ns[7]), .A2(n397), .B1(\A_s[7] ), .B2(n398), .ZN(n401)
         );
  INV_X1 U13 ( .A(\A_s[6] ), .ZN(n400) );
  INV_X1 U14 ( .A(A_ns[6]), .ZN(n399) );
  OAI221_X1 U15 ( .B1(n393), .B2(n402), .C1(n392), .C2(n403), .A(n404), .ZN(
        O[7]) );
  AOI22_X1 U16 ( .A1(A_ns[6]), .A2(n397), .B1(\A_s[6] ), .B2(n398), .ZN(n404)
         );
  INV_X1 U17 ( .A(\A_s[5] ), .ZN(n403) );
  INV_X1 U18 ( .A(A_ns[5]), .ZN(n402) );
  OAI221_X1 U19 ( .B1(n393), .B2(n405), .C1(n392), .C2(n406), .A(n407), .ZN(
        O[6]) );
  AOI22_X1 U20 ( .A1(A_ns[5]), .A2(n397), .B1(\A_s[5] ), .B2(n398), .ZN(n407)
         );
  INV_X1 U21 ( .A(\A_s[4] ), .ZN(n406) );
  INV_X1 U22 ( .A(A_ns[4]), .ZN(n405) );
  OAI221_X1 U23 ( .B1(n393), .B2(n408), .C1(n392), .C2(n409), .A(n410), .ZN(
        O[63]) );
  AOI22_X1 U24 ( .A1(A_ns[62]), .A2(n397), .B1(A_s[62]), .B2(n398), .ZN(n410)
         );
  INV_X1 U25 ( .A(\A_s[61] ), .ZN(n409) );
  INV_X1 U26 ( .A(A_ns[61]), .ZN(n408) );
  OAI221_X1 U27 ( .B1(n393), .B2(n411), .C1(n392), .C2(n412), .A(n413), .ZN(
        O[62]) );
  AOI22_X1 U28 ( .A1(A_ns[61]), .A2(n397), .B1(\A_s[61] ), .B2(n398), .ZN(n413) );
  INV_X1 U29 ( .A(\A_s[60] ), .ZN(n412) );
  INV_X1 U30 ( .A(A_ns[60]), .ZN(n411) );
  OAI221_X1 U31 ( .B1(n393), .B2(n414), .C1(n392), .C2(n415), .A(n416), .ZN(
        O[61]) );
  AOI22_X1 U32 ( .A1(A_ns[60]), .A2(n397), .B1(\A_s[60] ), .B2(n398), .ZN(n416) );
  INV_X1 U33 ( .A(\A_s[59] ), .ZN(n415) );
  INV_X1 U34 ( .A(A_ns[59]), .ZN(n414) );
  OAI221_X1 U35 ( .B1(n393), .B2(n417), .C1(n392), .C2(n418), .A(n419), .ZN(
        O[60]) );
  AOI22_X1 U36 ( .A1(A_ns[59]), .A2(n397), .B1(\A_s[59] ), .B2(n398), .ZN(n419) );
  INV_X1 U37 ( .A(\A_s[58] ), .ZN(n418) );
  INV_X1 U38 ( .A(A_ns[58]), .ZN(n417) );
  OAI221_X1 U39 ( .B1(n393), .B2(n420), .C1(n392), .C2(n421), .A(n422), .ZN(
        O[5]) );
  AOI22_X1 U40 ( .A1(A_ns[4]), .A2(n397), .B1(\A_s[4] ), .B2(n398), .ZN(n422)
         );
  INV_X1 U41 ( .A(\A_s[3] ), .ZN(n421) );
  INV_X1 U42 ( .A(A_ns[3]), .ZN(n420) );
  OAI221_X1 U43 ( .B1(n393), .B2(n423), .C1(n392), .C2(n424), .A(n425), .ZN(
        O[59]) );
  AOI22_X1 U44 ( .A1(A_ns[58]), .A2(n397), .B1(\A_s[58] ), .B2(n398), .ZN(n425) );
  INV_X1 U45 ( .A(\A_s[57] ), .ZN(n424) );
  INV_X1 U46 ( .A(A_ns[57]), .ZN(n423) );
  OAI221_X1 U47 ( .B1(n393), .B2(n426), .C1(n392), .C2(n427), .A(n428), .ZN(
        O[58]) );
  AOI22_X1 U48 ( .A1(A_ns[57]), .A2(n397), .B1(\A_s[57] ), .B2(n398), .ZN(n428) );
  INV_X1 U49 ( .A(\A_s[56] ), .ZN(n427) );
  INV_X1 U50 ( .A(A_ns[56]), .ZN(n426) );
  OAI221_X1 U51 ( .B1(n393), .B2(n429), .C1(n392), .C2(n430), .A(n431), .ZN(
        O[57]) );
  AOI22_X1 U52 ( .A1(A_ns[56]), .A2(n397), .B1(\A_s[56] ), .B2(n398), .ZN(n431) );
  INV_X1 U53 ( .A(\A_s[55] ), .ZN(n430) );
  INV_X1 U54 ( .A(A_ns[55]), .ZN(n429) );
  OAI221_X1 U55 ( .B1(n393), .B2(n432), .C1(n392), .C2(n433), .A(n434), .ZN(
        O[56]) );
  AOI22_X1 U56 ( .A1(A_ns[55]), .A2(n397), .B1(\A_s[55] ), .B2(n398), .ZN(n434) );
  INV_X1 U57 ( .A(\A_s[54] ), .ZN(n433) );
  INV_X1 U58 ( .A(A_ns[54]), .ZN(n432) );
  OAI221_X1 U59 ( .B1(n393), .B2(n435), .C1(n392), .C2(n436), .A(n437), .ZN(
        O[55]) );
  AOI22_X1 U60 ( .A1(A_ns[54]), .A2(n397), .B1(\A_s[54] ), .B2(n398), .ZN(n437) );
  INV_X1 U61 ( .A(\A_s[53] ), .ZN(n436) );
  INV_X1 U62 ( .A(A_ns[53]), .ZN(n435) );
  OAI221_X1 U63 ( .B1(n393), .B2(n438), .C1(n392), .C2(n439), .A(n440), .ZN(
        O[54]) );
  AOI22_X1 U64 ( .A1(A_ns[53]), .A2(n397), .B1(\A_s[53] ), .B2(n398), .ZN(n440) );
  INV_X1 U65 ( .A(\A_s[52] ), .ZN(n439) );
  INV_X1 U66 ( .A(A_ns[52]), .ZN(n438) );
  OAI221_X1 U67 ( .B1(n393), .B2(n441), .C1(n392), .C2(n442), .A(n443), .ZN(
        O[53]) );
  AOI22_X1 U68 ( .A1(A_ns[52]), .A2(n397), .B1(\A_s[52] ), .B2(n398), .ZN(n443) );
  INV_X1 U69 ( .A(\A_s[51] ), .ZN(n442) );
  INV_X1 U70 ( .A(A_ns[51]), .ZN(n441) );
  OAI221_X1 U71 ( .B1(n393), .B2(n444), .C1(n392), .C2(n445), .A(n446), .ZN(
        O[52]) );
  AOI22_X1 U72 ( .A1(A_ns[51]), .A2(n397), .B1(\A_s[51] ), .B2(n398), .ZN(n446) );
  INV_X1 U73 ( .A(\A_s[50] ), .ZN(n445) );
  INV_X1 U74 ( .A(A_ns[50]), .ZN(n444) );
  OAI221_X1 U75 ( .B1(n393), .B2(n447), .C1(n392), .C2(n448), .A(n449), .ZN(
        O[51]) );
  AOI22_X1 U76 ( .A1(A_ns[50]), .A2(n397), .B1(\A_s[50] ), .B2(n398), .ZN(n449) );
  INV_X1 U77 ( .A(\A_s[49] ), .ZN(n448) );
  INV_X1 U78 ( .A(A_ns[49]), .ZN(n447) );
  OAI221_X1 U79 ( .B1(n393), .B2(n450), .C1(n392), .C2(n451), .A(n452), .ZN(
        O[50]) );
  AOI22_X1 U80 ( .A1(A_ns[49]), .A2(n397), .B1(\A_s[49] ), .B2(n398), .ZN(n452) );
  INV_X1 U81 ( .A(\A_s[48] ), .ZN(n451) );
  INV_X1 U82 ( .A(A_ns[48]), .ZN(n450) );
  OAI221_X1 U83 ( .B1(n393), .B2(n453), .C1(n392), .C2(n454), .A(n455), .ZN(
        O[4]) );
  AOI22_X1 U84 ( .A1(A_ns[3]), .A2(n397), .B1(\A_s[3] ), .B2(n398), .ZN(n455)
         );
  INV_X1 U85 ( .A(\A_s[2] ), .ZN(n454) );
  INV_X1 U86 ( .A(A_ns[2]), .ZN(n453) );
  OAI221_X1 U87 ( .B1(n393), .B2(n456), .C1(n392), .C2(n457), .A(n458), .ZN(
        O[49]) );
  AOI22_X1 U88 ( .A1(A_ns[48]), .A2(n397), .B1(\A_s[48] ), .B2(n398), .ZN(n458) );
  INV_X1 U89 ( .A(\A_s[47] ), .ZN(n457) );
  INV_X1 U90 ( .A(A_ns[47]), .ZN(n456) );
  OAI221_X1 U91 ( .B1(n393), .B2(n459), .C1(n392), .C2(n460), .A(n461), .ZN(
        O[48]) );
  AOI22_X1 U92 ( .A1(A_ns[47]), .A2(n397), .B1(\A_s[47] ), .B2(n398), .ZN(n461) );
  INV_X1 U93 ( .A(\A_s[46] ), .ZN(n460) );
  INV_X1 U94 ( .A(A_ns[46]), .ZN(n459) );
  OAI221_X1 U95 ( .B1(n393), .B2(n462), .C1(n392), .C2(n463), .A(n464), .ZN(
        O[47]) );
  AOI22_X1 U96 ( .A1(A_ns[46]), .A2(n397), .B1(\A_s[46] ), .B2(n398), .ZN(n464) );
  INV_X1 U97 ( .A(\A_s[45] ), .ZN(n463) );
  INV_X1 U98 ( .A(A_ns[45]), .ZN(n462) );
  OAI221_X1 U99 ( .B1(n393), .B2(n465), .C1(n392), .C2(n466), .A(n467), .ZN(
        O[46]) );
  AOI22_X1 U100 ( .A1(A_ns[45]), .A2(n397), .B1(\A_s[45] ), .B2(n398), .ZN(
        n467) );
  INV_X1 U101 ( .A(\A_s[44] ), .ZN(n466) );
  INV_X1 U102 ( .A(A_ns[44]), .ZN(n465) );
  OAI221_X1 U103 ( .B1(n393), .B2(n468), .C1(n392), .C2(n469), .A(n470), .ZN(
        O[45]) );
  AOI22_X1 U104 ( .A1(A_ns[44]), .A2(n397), .B1(\A_s[44] ), .B2(n398), .ZN(
        n470) );
  INV_X1 U105 ( .A(\A_s[43] ), .ZN(n469) );
  INV_X1 U106 ( .A(A_ns[43]), .ZN(n468) );
  OAI221_X1 U107 ( .B1(n393), .B2(n471), .C1(n392), .C2(n472), .A(n473), .ZN(
        O[44]) );
  AOI22_X1 U108 ( .A1(A_ns[43]), .A2(n397), .B1(\A_s[43] ), .B2(n398), .ZN(
        n473) );
  INV_X1 U109 ( .A(\A_s[42] ), .ZN(n472) );
  INV_X1 U110 ( .A(A_ns[42]), .ZN(n471) );
  OAI221_X1 U111 ( .B1(n393), .B2(n474), .C1(n392), .C2(n475), .A(n476), .ZN(
        O[43]) );
  AOI22_X1 U112 ( .A1(A_ns[42]), .A2(n397), .B1(\A_s[42] ), .B2(n398), .ZN(
        n476) );
  INV_X1 U113 ( .A(\A_s[41] ), .ZN(n475) );
  INV_X1 U114 ( .A(A_ns[41]), .ZN(n474) );
  OAI221_X1 U115 ( .B1(n393), .B2(n477), .C1(n392), .C2(n478), .A(n479), .ZN(
        O[42]) );
  AOI22_X1 U116 ( .A1(A_ns[41]), .A2(n397), .B1(\A_s[41] ), .B2(n398), .ZN(
        n479) );
  INV_X1 U117 ( .A(\A_s[40] ), .ZN(n478) );
  INV_X1 U118 ( .A(A_ns[40]), .ZN(n477) );
  OAI221_X1 U119 ( .B1(n393), .B2(n480), .C1(n392), .C2(n481), .A(n482), .ZN(
        O[41]) );
  AOI22_X1 U120 ( .A1(A_ns[40]), .A2(n397), .B1(\A_s[40] ), .B2(n398), .ZN(
        n482) );
  INV_X1 U121 ( .A(\A_s[39] ), .ZN(n481) );
  INV_X1 U122 ( .A(A_ns[39]), .ZN(n480) );
  OAI221_X1 U123 ( .B1(n393), .B2(n483), .C1(n392), .C2(n484), .A(n485), .ZN(
        O[40]) );
  AOI22_X1 U124 ( .A1(A_ns[39]), .A2(n397), .B1(\A_s[39] ), .B2(n398), .ZN(
        n485) );
  INV_X1 U125 ( .A(\A_s[38] ), .ZN(n484) );
  INV_X1 U126 ( .A(A_ns[38]), .ZN(n483) );
  OAI221_X1 U127 ( .B1(n393), .B2(n486), .C1(n392), .C2(n487), .A(n488), .ZN(
        O[3]) );
  AOI22_X1 U128 ( .A1(A_ns[2]), .A2(n397), .B1(\A_s[2] ), .B2(n398), .ZN(n488)
         );
  INV_X1 U129 ( .A(\A_s[1] ), .ZN(n487) );
  INV_X1 U130 ( .A(A_ns[1]), .ZN(n486) );
  OAI221_X1 U131 ( .B1(n393), .B2(n489), .C1(n392), .C2(n490), .A(n491), .ZN(
        O[39]) );
  AOI22_X1 U132 ( .A1(A_ns[38]), .A2(n397), .B1(\A_s[38] ), .B2(n398), .ZN(
        n491) );
  INV_X1 U133 ( .A(\A_s[37] ), .ZN(n490) );
  INV_X1 U134 ( .A(A_ns[37]), .ZN(n489) );
  OAI221_X1 U135 ( .B1(n393), .B2(n492), .C1(n392), .C2(n493), .A(n494), .ZN(
        O[38]) );
  AOI22_X1 U136 ( .A1(A_ns[37]), .A2(n397), .B1(\A_s[37] ), .B2(n398), .ZN(
        n494) );
  INV_X1 U137 ( .A(\A_s[36] ), .ZN(n493) );
  INV_X1 U138 ( .A(A_ns[36]), .ZN(n492) );
  OAI221_X1 U139 ( .B1(n393), .B2(n495), .C1(n392), .C2(n496), .A(n497), .ZN(
        O[37]) );
  AOI22_X1 U140 ( .A1(A_ns[36]), .A2(n397), .B1(\A_s[36] ), .B2(n398), .ZN(
        n497) );
  INV_X1 U141 ( .A(\A_s[35] ), .ZN(n496) );
  INV_X1 U142 ( .A(A_ns[35]), .ZN(n495) );
  OAI221_X1 U143 ( .B1(n393), .B2(n498), .C1(n392), .C2(n499), .A(n500), .ZN(
        O[36]) );
  AOI22_X1 U144 ( .A1(A_ns[35]), .A2(n397), .B1(\A_s[35] ), .B2(n398), .ZN(
        n500) );
  INV_X1 U145 ( .A(\A_s[34] ), .ZN(n499) );
  INV_X1 U146 ( .A(A_ns[34]), .ZN(n498) );
  OAI221_X1 U147 ( .B1(n393), .B2(n501), .C1(n392), .C2(n502), .A(n503), .ZN(
        O[35]) );
  AOI22_X1 U148 ( .A1(A_ns[34]), .A2(n397), .B1(\A_s[34] ), .B2(n398), .ZN(
        n503) );
  INV_X1 U149 ( .A(\A_s[33] ), .ZN(n502) );
  INV_X1 U150 ( .A(A_ns[33]), .ZN(n501) );
  OAI221_X1 U151 ( .B1(n393), .B2(n504), .C1(n392), .C2(n505), .A(n506), .ZN(
        O[34]) );
  AOI22_X1 U152 ( .A1(A_ns[33]), .A2(n397), .B1(\A_s[33] ), .B2(n398), .ZN(
        n506) );
  INV_X1 U153 ( .A(\A_s[32] ), .ZN(n505) );
  INV_X1 U154 ( .A(A_ns[32]), .ZN(n504) );
  OAI221_X1 U155 ( .B1(n393), .B2(n507), .C1(n392), .C2(n508), .A(n509), .ZN(
        O[33]) );
  AOI22_X1 U156 ( .A1(A_ns[32]), .A2(n397), .B1(\A_s[32] ), .B2(n398), .ZN(
        n509) );
  INV_X1 U157 ( .A(\A_s[31] ), .ZN(n508) );
  INV_X1 U158 ( .A(A_ns[31]), .ZN(n507) );
  OAI221_X1 U159 ( .B1(n393), .B2(n510), .C1(n392), .C2(n511), .A(n512), .ZN(
        O[32]) );
  AOI22_X1 U160 ( .A1(A_ns[31]), .A2(n397), .B1(\A_s[31] ), .B2(n398), .ZN(
        n512) );
  INV_X1 U161 ( .A(\A_s[30] ), .ZN(n511) );
  INV_X1 U162 ( .A(A_ns[30]), .ZN(n510) );
  OAI221_X1 U163 ( .B1(n393), .B2(n513), .C1(n392), .C2(n514), .A(n515), .ZN(
        O[31]) );
  AOI22_X1 U164 ( .A1(A_ns[30]), .A2(n397), .B1(\A_s[30] ), .B2(n398), .ZN(
        n515) );
  INV_X1 U165 ( .A(\A_s[29] ), .ZN(n514) );
  INV_X1 U166 ( .A(A_ns[29]), .ZN(n513) );
  OAI221_X1 U167 ( .B1(n393), .B2(n516), .C1(n392), .C2(n517), .A(n518), .ZN(
        O[30]) );
  AOI22_X1 U168 ( .A1(A_ns[29]), .A2(n397), .B1(\A_s[29] ), .B2(n398), .ZN(
        n518) );
  INV_X1 U169 ( .A(\A_s[28] ), .ZN(n517) );
  INV_X1 U170 ( .A(A_ns[28]), .ZN(n516) );
  OAI221_X1 U171 ( .B1(n393), .B2(n519), .C1(n392), .C2(n520), .A(n521), .ZN(
        O[2]) );
  AOI22_X1 U172 ( .A1(A_ns[1]), .A2(n397), .B1(\A_s[1] ), .B2(n398), .ZN(n521)
         );
  OAI221_X1 U173 ( .B1(n393), .B2(n522), .C1(n392), .C2(n523), .A(n524), .ZN(
        O[29]) );
  AOI22_X1 U174 ( .A1(A_ns[28]), .A2(n397), .B1(\A_s[28] ), .B2(n398), .ZN(
        n524) );
  INV_X1 U175 ( .A(\A_s[27] ), .ZN(n523) );
  INV_X1 U176 ( .A(A_ns[27]), .ZN(n522) );
  OAI221_X1 U177 ( .B1(n393), .B2(n525), .C1(n392), .C2(n526), .A(n527), .ZN(
        O[28]) );
  AOI22_X1 U178 ( .A1(A_ns[27]), .A2(n397), .B1(\A_s[27] ), .B2(n398), .ZN(
        n527) );
  INV_X1 U179 ( .A(\A_s[26] ), .ZN(n526) );
  INV_X1 U180 ( .A(A_ns[26]), .ZN(n525) );
  OAI221_X1 U181 ( .B1(n393), .B2(n528), .C1(n392), .C2(n529), .A(n530), .ZN(
        O[27]) );
  AOI22_X1 U182 ( .A1(A_ns[26]), .A2(n397), .B1(\A_s[26] ), .B2(n398), .ZN(
        n530) );
  INV_X1 U183 ( .A(\A_s[25] ), .ZN(n529) );
  INV_X1 U184 ( .A(A_ns[25]), .ZN(n528) );
  OAI221_X1 U185 ( .B1(n393), .B2(n531), .C1(n392), .C2(n532), .A(n533), .ZN(
        O[26]) );
  AOI22_X1 U186 ( .A1(A_ns[25]), .A2(n397), .B1(\A_s[25] ), .B2(n398), .ZN(
        n533) );
  INV_X1 U187 ( .A(\A_s[24] ), .ZN(n532) );
  INV_X1 U188 ( .A(A_ns[24]), .ZN(n531) );
  OAI221_X1 U189 ( .B1(n393), .B2(n534), .C1(n392), .C2(n535), .A(n536), .ZN(
        O[25]) );
  AOI22_X1 U190 ( .A1(A_ns[24]), .A2(n397), .B1(\A_s[24] ), .B2(n398), .ZN(
        n536) );
  INV_X1 U191 ( .A(\A_s[23] ), .ZN(n535) );
  INV_X1 U192 ( .A(A_ns[23]), .ZN(n534) );
  OAI221_X1 U193 ( .B1(n393), .B2(n537), .C1(n392), .C2(n538), .A(n539), .ZN(
        O[24]) );
  AOI22_X1 U194 ( .A1(A_ns[23]), .A2(n397), .B1(\A_s[23] ), .B2(n398), .ZN(
        n539) );
  INV_X1 U195 ( .A(\A_s[22] ), .ZN(n538) );
  INV_X1 U196 ( .A(A_ns[22]), .ZN(n537) );
  OAI221_X1 U197 ( .B1(n393), .B2(n540), .C1(n392), .C2(n541), .A(n542), .ZN(
        O[23]) );
  AOI22_X1 U198 ( .A1(A_ns[22]), .A2(n397), .B1(\A_s[22] ), .B2(n398), .ZN(
        n542) );
  INV_X1 U199 ( .A(\A_s[21] ), .ZN(n541) );
  INV_X1 U200 ( .A(A_ns[21]), .ZN(n540) );
  OAI221_X1 U201 ( .B1(n393), .B2(n543), .C1(n392), .C2(n544), .A(n545), .ZN(
        O[22]) );
  AOI22_X1 U202 ( .A1(A_ns[21]), .A2(n397), .B1(\A_s[21] ), .B2(n398), .ZN(
        n545) );
  INV_X1 U203 ( .A(\A_s[20] ), .ZN(n544) );
  INV_X1 U204 ( .A(A_ns[20]), .ZN(n543) );
  OAI221_X1 U205 ( .B1(n393), .B2(n546), .C1(n392), .C2(n547), .A(n548), .ZN(
        O[21]) );
  AOI22_X1 U206 ( .A1(A_ns[20]), .A2(n397), .B1(\A_s[20] ), .B2(n398), .ZN(
        n548) );
  INV_X1 U207 ( .A(\A_s[19] ), .ZN(n547) );
  INV_X1 U208 ( .A(A_ns[19]), .ZN(n546) );
  OAI221_X1 U209 ( .B1(n393), .B2(n549), .C1(n392), .C2(n550), .A(n551), .ZN(
        O[20]) );
  AOI22_X1 U210 ( .A1(A_ns[19]), .A2(n397), .B1(\A_s[19] ), .B2(n398), .ZN(
        n551) );
  INV_X1 U211 ( .A(\A_s[18] ), .ZN(n550) );
  INV_X1 U212 ( .A(A_ns[18]), .ZN(n549) );
  OAI22_X1 U213 ( .A1(n552), .A2(n520), .B1(n553), .B2(n519), .ZN(O[1]) );
  INV_X1 U214 ( .A(A_ns[0]), .ZN(n519) );
  INV_X1 U215 ( .A(\A_s[0] ), .ZN(n520) );
  OAI221_X1 U216 ( .B1(n393), .B2(n554), .C1(n392), .C2(n555), .A(n556), .ZN(
        O[19]) );
  AOI22_X1 U217 ( .A1(A_ns[18]), .A2(n397), .B1(\A_s[18] ), .B2(n398), .ZN(
        n556) );
  INV_X1 U218 ( .A(\A_s[17] ), .ZN(n555) );
  INV_X1 U219 ( .A(A_ns[17]), .ZN(n554) );
  OAI221_X1 U220 ( .B1(n393), .B2(n557), .C1(n392), .C2(n558), .A(n559), .ZN(
        O[18]) );
  AOI22_X1 U221 ( .A1(A_ns[17]), .A2(n397), .B1(\A_s[17] ), .B2(n398), .ZN(
        n559) );
  INV_X1 U222 ( .A(\A_s[16] ), .ZN(n558) );
  INV_X1 U223 ( .A(A_ns[16]), .ZN(n557) );
  OAI221_X1 U224 ( .B1(n393), .B2(n560), .C1(n392), .C2(n561), .A(n562), .ZN(
        O[17]) );
  AOI22_X1 U225 ( .A1(A_ns[16]), .A2(n397), .B1(\A_s[16] ), .B2(n398), .ZN(
        n562) );
  INV_X1 U226 ( .A(\A_s[15] ), .ZN(n561) );
  INV_X1 U227 ( .A(A_ns[15]), .ZN(n560) );
  OAI221_X1 U228 ( .B1(n393), .B2(n563), .C1(n392), .C2(n564), .A(n565), .ZN(
        O[16]) );
  AOI22_X1 U229 ( .A1(A_ns[15]), .A2(n397), .B1(\A_s[15] ), .B2(n398), .ZN(
        n565) );
  INV_X1 U230 ( .A(\A_s[14] ), .ZN(n564) );
  INV_X1 U231 ( .A(A_ns[14]), .ZN(n563) );
  OAI221_X1 U232 ( .B1(n393), .B2(n566), .C1(n392), .C2(n567), .A(n568), .ZN(
        O[15]) );
  AOI22_X1 U233 ( .A1(A_ns[14]), .A2(n397), .B1(\A_s[14] ), .B2(n398), .ZN(
        n568) );
  INV_X1 U234 ( .A(\A_s[13] ), .ZN(n567) );
  INV_X1 U235 ( .A(A_ns[13]), .ZN(n566) );
  OAI221_X1 U236 ( .B1(n393), .B2(n569), .C1(n392), .C2(n570), .A(n571), .ZN(
        O[14]) );
  AOI22_X1 U237 ( .A1(A_ns[13]), .A2(n397), .B1(\A_s[13] ), .B2(n398), .ZN(
        n571) );
  INV_X1 U238 ( .A(\A_s[12] ), .ZN(n570) );
  INV_X1 U239 ( .A(A_ns[12]), .ZN(n569) );
  OAI221_X1 U240 ( .B1(n393), .B2(n572), .C1(n392), .C2(n573), .A(n574), .ZN(
        O[13]) );
  AOI22_X1 U241 ( .A1(A_ns[12]), .A2(n397), .B1(\A_s[12] ), .B2(n398), .ZN(
        n574) );
  INV_X1 U242 ( .A(\A_s[11] ), .ZN(n573) );
  INV_X1 U243 ( .A(A_ns[11]), .ZN(n572) );
  OAI221_X1 U244 ( .B1(n393), .B2(n575), .C1(n392), .C2(n576), .A(n577), .ZN(
        O[12]) );
  AOI22_X1 U245 ( .A1(A_ns[11]), .A2(n397), .B1(\A_s[11] ), .B2(n398), .ZN(
        n577) );
  INV_X1 U246 ( .A(\A_s[10] ), .ZN(n576) );
  INV_X1 U247 ( .A(A_ns[10]), .ZN(n575) );
  OAI221_X1 U248 ( .B1(n393), .B2(n578), .C1(n392), .C2(n579), .A(n580), .ZN(
        O[11]) );
  AOI22_X1 U249 ( .A1(A_ns[10]), .A2(n397), .B1(\A_s[10] ), .B2(n398), .ZN(
        n580) );
  INV_X1 U250 ( .A(\A_s[9] ), .ZN(n579) );
  INV_X1 U251 ( .A(A_ns[9]), .ZN(n578) );
  OAI221_X1 U252 ( .B1(n581), .B2(n393), .C1(n582), .C2(n392), .A(n583), .ZN(
        O[10]) );
  AOI22_X1 U253 ( .A1(A_ns[9]), .A2(n397), .B1(\A_s[9] ), .B2(n398), .ZN(n583)
         );
  NAND2_X1 U254 ( .A1(n584), .A2(n552), .ZN(n553) );
  NAND2_X1 U255 ( .A1(n584), .A2(n585), .ZN(n552) );
  XOR2_X1 U256 ( .A(B[5]), .B(B[6]), .Z(n584) );
  INV_X1 U257 ( .A(\A_s[8] ), .ZN(n582) );
  INV_X1 U258 ( .A(B[7]), .ZN(n585) );
  INV_X1 U259 ( .A(A_ns[8]), .ZN(n581) );
endmodule


module BOOTHENC_NBIT64_i8 ( A, A_n, A_ns, A_s, B, O, A_so, A_nso );
  input [63:0] A;
  input [63:0] A_n;
  input [63:0] A_ns;
  input [63:0] A_s;
  input [63:0] B;
  output [63:0] O;
  output [63:0] A_so;
  output [63:0] A_nso;
  wire   \A_s[61] , \A_s[60] , \A_s[59] , \A_s[58] , \A_s[57] , \A_s[56] ,
         \A_s[55] , \A_s[54] , \A_s[53] , \A_s[52] , \A_s[51] , \A_s[50] ,
         \A_s[49] , \A_s[48] , \A_s[47] , \A_s[46] , \A_s[45] , \A_s[44] ,
         \A_s[43] , \A_s[42] , \A_s[41] , \A_s[40] , \A_s[39] , \A_s[38] ,
         \A_s[37] , \A_s[36] , \A_s[35] , \A_s[34] , \A_s[33] , \A_s[32] ,
         \A_s[31] , \A_s[30] , \A_s[29] , \A_s[28] , \A_s[27] , \A_s[26] ,
         \A_s[25] , \A_s[24] , \A_s[23] , \A_s[22] , \A_s[21] , \A_s[20] ,
         \A_s[19] , \A_s[18] , \A_s[17] , \A_s[16] , \A_s[15] , \A_s[14] ,
         \A_s[13] , \A_s[12] , \A_s[11] , \A_s[10] , \A_s[9] , \A_s[8] ,
         \A_s[7] , \A_s[6] , \A_s[5] , \A_s[4] , \A_s[3] , \A_s[2] , \A_s[1] ,
         \A_s[0] , n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585;
  assign A_nso[0] = 1'b0;
  assign A_nso[1] = 1'b0;
  assign A_so[0] = 1'b0;
  assign A_so[1] = 1'b0;
  assign O[0] = 1'b0;
  assign A_nso[63] = \A_s[61] ;
  assign A_so[63] = \A_s[61] ;
  assign \A_s[61]  = A_s[61];
  assign A_nso[62] = \A_s[60] ;
  assign A_so[62] = \A_s[60] ;
  assign \A_s[60]  = A_s[60];
  assign A_nso[61] = \A_s[59] ;
  assign A_so[61] = \A_s[59] ;
  assign \A_s[59]  = A_s[59];
  assign A_nso[60] = \A_s[58] ;
  assign A_so[60] = \A_s[58] ;
  assign \A_s[58]  = A_s[58];
  assign A_nso[59] = \A_s[57] ;
  assign A_so[59] = \A_s[57] ;
  assign \A_s[57]  = A_s[57];
  assign A_nso[58] = \A_s[56] ;
  assign A_so[58] = \A_s[56] ;
  assign \A_s[56]  = A_s[56];
  assign A_nso[57] = \A_s[55] ;
  assign A_so[57] = \A_s[55] ;
  assign \A_s[55]  = A_s[55];
  assign A_nso[56] = \A_s[54] ;
  assign A_so[56] = \A_s[54] ;
  assign \A_s[54]  = A_s[54];
  assign A_nso[55] = \A_s[53] ;
  assign A_so[55] = \A_s[53] ;
  assign \A_s[53]  = A_s[53];
  assign A_nso[54] = \A_s[52] ;
  assign A_so[54] = \A_s[52] ;
  assign \A_s[52]  = A_s[52];
  assign A_nso[53] = \A_s[51] ;
  assign A_so[53] = \A_s[51] ;
  assign \A_s[51]  = A_s[51];
  assign A_nso[52] = \A_s[50] ;
  assign A_so[52] = \A_s[50] ;
  assign \A_s[50]  = A_s[50];
  assign A_nso[51] = \A_s[49] ;
  assign A_so[51] = \A_s[49] ;
  assign \A_s[49]  = A_s[49];
  assign A_nso[50] = \A_s[48] ;
  assign A_so[50] = \A_s[48] ;
  assign \A_s[48]  = A_s[48];
  assign A_nso[49] = \A_s[47] ;
  assign A_so[49] = \A_s[47] ;
  assign \A_s[47]  = A_s[47];
  assign A_nso[48] = \A_s[46] ;
  assign A_so[48] = \A_s[46] ;
  assign \A_s[46]  = A_s[46];
  assign A_nso[47] = \A_s[45] ;
  assign A_so[47] = \A_s[45] ;
  assign \A_s[45]  = A_s[45];
  assign A_nso[46] = \A_s[44] ;
  assign A_so[46] = \A_s[44] ;
  assign \A_s[44]  = A_s[44];
  assign A_nso[45] = \A_s[43] ;
  assign A_so[45] = \A_s[43] ;
  assign \A_s[43]  = A_s[43];
  assign A_nso[44] = \A_s[42] ;
  assign A_so[44] = \A_s[42] ;
  assign \A_s[42]  = A_s[42];
  assign A_nso[43] = \A_s[41] ;
  assign A_so[43] = \A_s[41] ;
  assign \A_s[41]  = A_s[41];
  assign A_nso[42] = \A_s[40] ;
  assign A_so[42] = \A_s[40] ;
  assign \A_s[40]  = A_s[40];
  assign A_nso[41] = \A_s[39] ;
  assign A_so[41] = \A_s[39] ;
  assign \A_s[39]  = A_s[39];
  assign A_nso[40] = \A_s[38] ;
  assign A_so[40] = \A_s[38] ;
  assign \A_s[38]  = A_s[38];
  assign A_nso[39] = \A_s[37] ;
  assign A_so[39] = \A_s[37] ;
  assign \A_s[37]  = A_s[37];
  assign A_nso[38] = \A_s[36] ;
  assign A_so[38] = \A_s[36] ;
  assign \A_s[36]  = A_s[36];
  assign A_nso[37] = \A_s[35] ;
  assign A_so[37] = \A_s[35] ;
  assign \A_s[35]  = A_s[35];
  assign A_nso[36] = \A_s[34] ;
  assign A_so[36] = \A_s[34] ;
  assign \A_s[34]  = A_s[34];
  assign A_nso[35] = \A_s[33] ;
  assign A_so[35] = \A_s[33] ;
  assign \A_s[33]  = A_s[33];
  assign A_nso[34] = \A_s[32] ;
  assign A_so[34] = \A_s[32] ;
  assign \A_s[32]  = A_s[32];
  assign A_nso[33] = \A_s[31] ;
  assign A_so[33] = \A_s[31] ;
  assign \A_s[31]  = A_s[31];
  assign A_nso[32] = \A_s[30] ;
  assign A_so[32] = \A_s[30] ;
  assign \A_s[30]  = A_s[30];
  assign A_nso[31] = \A_s[29] ;
  assign A_so[31] = \A_s[29] ;
  assign \A_s[29]  = A_s[29];
  assign A_nso[30] = \A_s[28] ;
  assign A_so[30] = \A_s[28] ;
  assign \A_s[28]  = A_s[28];
  assign A_nso[29] = \A_s[27] ;
  assign A_so[29] = \A_s[27] ;
  assign \A_s[27]  = A_s[27];
  assign A_nso[28] = \A_s[26] ;
  assign A_so[28] = \A_s[26] ;
  assign \A_s[26]  = A_s[26];
  assign A_nso[27] = \A_s[25] ;
  assign A_so[27] = \A_s[25] ;
  assign \A_s[25]  = A_s[25];
  assign A_nso[26] = \A_s[24] ;
  assign A_so[26] = \A_s[24] ;
  assign \A_s[24]  = A_s[24];
  assign A_nso[25] = \A_s[23] ;
  assign A_so[25] = \A_s[23] ;
  assign \A_s[23]  = A_s[23];
  assign A_nso[24] = \A_s[22] ;
  assign A_so[24] = \A_s[22] ;
  assign \A_s[22]  = A_s[22];
  assign A_nso[23] = \A_s[21] ;
  assign A_so[23] = \A_s[21] ;
  assign \A_s[21]  = A_s[21];
  assign A_nso[22] = \A_s[20] ;
  assign A_so[22] = \A_s[20] ;
  assign \A_s[20]  = A_s[20];
  assign A_nso[21] = \A_s[19] ;
  assign A_so[21] = \A_s[19] ;
  assign \A_s[19]  = A_s[19];
  assign A_nso[20] = \A_s[18] ;
  assign A_so[20] = \A_s[18] ;
  assign \A_s[18]  = A_s[18];
  assign A_nso[19] = \A_s[17] ;
  assign A_so[19] = \A_s[17] ;
  assign \A_s[17]  = A_s[17];
  assign A_nso[18] = \A_s[16] ;
  assign A_so[18] = \A_s[16] ;
  assign \A_s[16]  = A_s[16];
  assign A_nso[17] = \A_s[15] ;
  assign A_so[17] = \A_s[15] ;
  assign \A_s[15]  = A_s[15];
  assign A_nso[16] = \A_s[14] ;
  assign A_so[16] = \A_s[14] ;
  assign \A_s[14]  = A_s[14];
  assign A_nso[15] = \A_s[13] ;
  assign A_so[15] = \A_s[13] ;
  assign \A_s[13]  = A_s[13];
  assign A_nso[14] = \A_s[12] ;
  assign A_so[14] = \A_s[12] ;
  assign \A_s[12]  = A_s[12];
  assign A_nso[13] = \A_s[11] ;
  assign A_so[13] = \A_s[11] ;
  assign \A_s[11]  = A_s[11];
  assign A_nso[12] = \A_s[10] ;
  assign A_so[12] = \A_s[10] ;
  assign \A_s[10]  = A_s[10];
  assign A_nso[11] = \A_s[9] ;
  assign A_so[11] = \A_s[9] ;
  assign \A_s[9]  = A_s[9];
  assign A_nso[10] = \A_s[8] ;
  assign A_so[10] = \A_s[8] ;
  assign \A_s[8]  = A_s[8];
  assign A_nso[9] = \A_s[7] ;
  assign A_so[9] = \A_s[7] ;
  assign \A_s[7]  = A_s[7];
  assign A_nso[8] = \A_s[6] ;
  assign A_so[8] = \A_s[6] ;
  assign \A_s[6]  = A_s[6];
  assign A_nso[7] = \A_s[5] ;
  assign A_so[7] = \A_s[5] ;
  assign \A_s[5]  = A_s[5];
  assign A_nso[6] = \A_s[4] ;
  assign A_so[6] = \A_s[4] ;
  assign \A_s[4]  = A_s[4];
  assign A_nso[5] = \A_s[3] ;
  assign A_so[5] = \A_s[3] ;
  assign \A_s[3]  = A_s[3];
  assign A_nso[4] = \A_s[2] ;
  assign A_so[4] = \A_s[2] ;
  assign \A_s[2]  = A_s[2];
  assign A_nso[3] = \A_s[1] ;
  assign A_so[3] = \A_s[1] ;
  assign \A_s[1]  = A_s[1];
  assign A_nso[2] = \A_s[0] ;
  assign A_so[2] = \A_s[0] ;
  assign \A_s[0]  = A_s[0];

  AND3_X1 U2 ( .A1(B[8]), .A2(n585), .A3(B[7]), .ZN(n391) );
  INV_X4 U3 ( .A(n391), .ZN(n392) );
  INV_X4 U4 ( .A(n552), .ZN(n398) );
  OR3_X4 U5 ( .A1(B[7]), .A2(B[8]), .A3(n585), .ZN(n393) );
  INV_X4 U6 ( .A(n553), .ZN(n397) );
  OAI221_X1 U7 ( .B1(n393), .B2(n394), .C1(n392), .C2(n395), .A(n396), .ZN(
        O[9]) );
  AOI22_X1 U8 ( .A1(A_ns[8]), .A2(n397), .B1(\A_s[8] ), .B2(n398), .ZN(n396)
         );
  INV_X1 U9 ( .A(\A_s[7] ), .ZN(n395) );
  INV_X1 U10 ( .A(A_ns[7]), .ZN(n394) );
  OAI221_X1 U11 ( .B1(n393), .B2(n399), .C1(n392), .C2(n400), .A(n401), .ZN(
        O[8]) );
  AOI22_X1 U12 ( .A1(A_ns[7]), .A2(n397), .B1(\A_s[7] ), .B2(n398), .ZN(n401)
         );
  INV_X1 U13 ( .A(\A_s[6] ), .ZN(n400) );
  INV_X1 U14 ( .A(A_ns[6]), .ZN(n399) );
  OAI221_X1 U15 ( .B1(n393), .B2(n402), .C1(n392), .C2(n403), .A(n404), .ZN(
        O[7]) );
  AOI22_X1 U16 ( .A1(A_ns[6]), .A2(n397), .B1(\A_s[6] ), .B2(n398), .ZN(n404)
         );
  INV_X1 U17 ( .A(\A_s[5] ), .ZN(n403) );
  INV_X1 U18 ( .A(A_ns[5]), .ZN(n402) );
  OAI221_X1 U19 ( .B1(n393), .B2(n405), .C1(n392), .C2(n406), .A(n407), .ZN(
        O[6]) );
  AOI22_X1 U20 ( .A1(A_ns[5]), .A2(n397), .B1(\A_s[5] ), .B2(n398), .ZN(n407)
         );
  INV_X1 U21 ( .A(\A_s[4] ), .ZN(n406) );
  INV_X1 U22 ( .A(A_ns[4]), .ZN(n405) );
  OAI221_X1 U23 ( .B1(n393), .B2(n408), .C1(n392), .C2(n409), .A(n410), .ZN(
        O[63]) );
  AOI22_X1 U24 ( .A1(A_ns[62]), .A2(n397), .B1(A_s[62]), .B2(n398), .ZN(n410)
         );
  INV_X1 U25 ( .A(\A_s[61] ), .ZN(n409) );
  INV_X1 U26 ( .A(A_ns[61]), .ZN(n408) );
  OAI221_X1 U27 ( .B1(n393), .B2(n411), .C1(n392), .C2(n412), .A(n413), .ZN(
        O[62]) );
  AOI22_X1 U28 ( .A1(A_ns[61]), .A2(n397), .B1(\A_s[61] ), .B2(n398), .ZN(n413) );
  INV_X1 U29 ( .A(\A_s[60] ), .ZN(n412) );
  INV_X1 U30 ( .A(A_ns[60]), .ZN(n411) );
  OAI221_X1 U31 ( .B1(n393), .B2(n414), .C1(n392), .C2(n415), .A(n416), .ZN(
        O[61]) );
  AOI22_X1 U32 ( .A1(A_ns[60]), .A2(n397), .B1(\A_s[60] ), .B2(n398), .ZN(n416) );
  INV_X1 U33 ( .A(\A_s[59] ), .ZN(n415) );
  INV_X1 U34 ( .A(A_ns[59]), .ZN(n414) );
  OAI221_X1 U35 ( .B1(n393), .B2(n417), .C1(n392), .C2(n418), .A(n419), .ZN(
        O[60]) );
  AOI22_X1 U36 ( .A1(A_ns[59]), .A2(n397), .B1(\A_s[59] ), .B2(n398), .ZN(n419) );
  INV_X1 U37 ( .A(\A_s[58] ), .ZN(n418) );
  INV_X1 U38 ( .A(A_ns[58]), .ZN(n417) );
  OAI221_X1 U39 ( .B1(n393), .B2(n420), .C1(n392), .C2(n421), .A(n422), .ZN(
        O[5]) );
  AOI22_X1 U40 ( .A1(A_ns[4]), .A2(n397), .B1(\A_s[4] ), .B2(n398), .ZN(n422)
         );
  INV_X1 U41 ( .A(\A_s[3] ), .ZN(n421) );
  INV_X1 U42 ( .A(A_ns[3]), .ZN(n420) );
  OAI221_X1 U43 ( .B1(n393), .B2(n423), .C1(n392), .C2(n424), .A(n425), .ZN(
        O[59]) );
  AOI22_X1 U44 ( .A1(A_ns[58]), .A2(n397), .B1(\A_s[58] ), .B2(n398), .ZN(n425) );
  INV_X1 U45 ( .A(\A_s[57] ), .ZN(n424) );
  INV_X1 U46 ( .A(A_ns[57]), .ZN(n423) );
  OAI221_X1 U47 ( .B1(n393), .B2(n426), .C1(n392), .C2(n427), .A(n428), .ZN(
        O[58]) );
  AOI22_X1 U48 ( .A1(A_ns[57]), .A2(n397), .B1(\A_s[57] ), .B2(n398), .ZN(n428) );
  INV_X1 U49 ( .A(\A_s[56] ), .ZN(n427) );
  INV_X1 U50 ( .A(A_ns[56]), .ZN(n426) );
  OAI221_X1 U51 ( .B1(n393), .B2(n429), .C1(n392), .C2(n430), .A(n431), .ZN(
        O[57]) );
  AOI22_X1 U52 ( .A1(A_ns[56]), .A2(n397), .B1(\A_s[56] ), .B2(n398), .ZN(n431) );
  INV_X1 U53 ( .A(\A_s[55] ), .ZN(n430) );
  INV_X1 U54 ( .A(A_ns[55]), .ZN(n429) );
  OAI221_X1 U55 ( .B1(n393), .B2(n432), .C1(n392), .C2(n433), .A(n434), .ZN(
        O[56]) );
  AOI22_X1 U56 ( .A1(A_ns[55]), .A2(n397), .B1(\A_s[55] ), .B2(n398), .ZN(n434) );
  INV_X1 U57 ( .A(\A_s[54] ), .ZN(n433) );
  INV_X1 U58 ( .A(A_ns[54]), .ZN(n432) );
  OAI221_X1 U59 ( .B1(n393), .B2(n435), .C1(n392), .C2(n436), .A(n437), .ZN(
        O[55]) );
  AOI22_X1 U60 ( .A1(A_ns[54]), .A2(n397), .B1(\A_s[54] ), .B2(n398), .ZN(n437) );
  INV_X1 U61 ( .A(\A_s[53] ), .ZN(n436) );
  INV_X1 U62 ( .A(A_ns[53]), .ZN(n435) );
  OAI221_X1 U63 ( .B1(n393), .B2(n438), .C1(n392), .C2(n439), .A(n440), .ZN(
        O[54]) );
  AOI22_X1 U64 ( .A1(A_ns[53]), .A2(n397), .B1(\A_s[53] ), .B2(n398), .ZN(n440) );
  INV_X1 U65 ( .A(\A_s[52] ), .ZN(n439) );
  INV_X1 U66 ( .A(A_ns[52]), .ZN(n438) );
  OAI221_X1 U67 ( .B1(n393), .B2(n441), .C1(n392), .C2(n442), .A(n443), .ZN(
        O[53]) );
  AOI22_X1 U68 ( .A1(A_ns[52]), .A2(n397), .B1(\A_s[52] ), .B2(n398), .ZN(n443) );
  INV_X1 U69 ( .A(\A_s[51] ), .ZN(n442) );
  INV_X1 U70 ( .A(A_ns[51]), .ZN(n441) );
  OAI221_X1 U71 ( .B1(n393), .B2(n444), .C1(n392), .C2(n445), .A(n446), .ZN(
        O[52]) );
  AOI22_X1 U72 ( .A1(A_ns[51]), .A2(n397), .B1(\A_s[51] ), .B2(n398), .ZN(n446) );
  INV_X1 U73 ( .A(\A_s[50] ), .ZN(n445) );
  INV_X1 U74 ( .A(A_ns[50]), .ZN(n444) );
  OAI221_X1 U75 ( .B1(n393), .B2(n447), .C1(n392), .C2(n448), .A(n449), .ZN(
        O[51]) );
  AOI22_X1 U76 ( .A1(A_ns[50]), .A2(n397), .B1(\A_s[50] ), .B2(n398), .ZN(n449) );
  INV_X1 U77 ( .A(\A_s[49] ), .ZN(n448) );
  INV_X1 U78 ( .A(A_ns[49]), .ZN(n447) );
  OAI221_X1 U79 ( .B1(n393), .B2(n450), .C1(n392), .C2(n451), .A(n452), .ZN(
        O[50]) );
  AOI22_X1 U80 ( .A1(A_ns[49]), .A2(n397), .B1(\A_s[49] ), .B2(n398), .ZN(n452) );
  INV_X1 U81 ( .A(\A_s[48] ), .ZN(n451) );
  INV_X1 U82 ( .A(A_ns[48]), .ZN(n450) );
  OAI221_X1 U83 ( .B1(n393), .B2(n453), .C1(n392), .C2(n454), .A(n455), .ZN(
        O[4]) );
  AOI22_X1 U84 ( .A1(A_ns[3]), .A2(n397), .B1(\A_s[3] ), .B2(n398), .ZN(n455)
         );
  INV_X1 U85 ( .A(\A_s[2] ), .ZN(n454) );
  INV_X1 U86 ( .A(A_ns[2]), .ZN(n453) );
  OAI221_X1 U87 ( .B1(n393), .B2(n456), .C1(n392), .C2(n457), .A(n458), .ZN(
        O[49]) );
  AOI22_X1 U88 ( .A1(A_ns[48]), .A2(n397), .B1(\A_s[48] ), .B2(n398), .ZN(n458) );
  INV_X1 U89 ( .A(\A_s[47] ), .ZN(n457) );
  INV_X1 U90 ( .A(A_ns[47]), .ZN(n456) );
  OAI221_X1 U91 ( .B1(n393), .B2(n459), .C1(n392), .C2(n460), .A(n461), .ZN(
        O[48]) );
  AOI22_X1 U92 ( .A1(A_ns[47]), .A2(n397), .B1(\A_s[47] ), .B2(n398), .ZN(n461) );
  INV_X1 U93 ( .A(\A_s[46] ), .ZN(n460) );
  INV_X1 U94 ( .A(A_ns[46]), .ZN(n459) );
  OAI221_X1 U95 ( .B1(n393), .B2(n462), .C1(n392), .C2(n463), .A(n464), .ZN(
        O[47]) );
  AOI22_X1 U96 ( .A1(A_ns[46]), .A2(n397), .B1(\A_s[46] ), .B2(n398), .ZN(n464) );
  INV_X1 U97 ( .A(\A_s[45] ), .ZN(n463) );
  INV_X1 U98 ( .A(A_ns[45]), .ZN(n462) );
  OAI221_X1 U99 ( .B1(n393), .B2(n465), .C1(n392), .C2(n466), .A(n467), .ZN(
        O[46]) );
  AOI22_X1 U100 ( .A1(A_ns[45]), .A2(n397), .B1(\A_s[45] ), .B2(n398), .ZN(
        n467) );
  INV_X1 U101 ( .A(\A_s[44] ), .ZN(n466) );
  INV_X1 U102 ( .A(A_ns[44]), .ZN(n465) );
  OAI221_X1 U103 ( .B1(n393), .B2(n468), .C1(n392), .C2(n469), .A(n470), .ZN(
        O[45]) );
  AOI22_X1 U104 ( .A1(A_ns[44]), .A2(n397), .B1(\A_s[44] ), .B2(n398), .ZN(
        n470) );
  INV_X1 U105 ( .A(\A_s[43] ), .ZN(n469) );
  INV_X1 U106 ( .A(A_ns[43]), .ZN(n468) );
  OAI221_X1 U107 ( .B1(n393), .B2(n471), .C1(n392), .C2(n472), .A(n473), .ZN(
        O[44]) );
  AOI22_X1 U108 ( .A1(A_ns[43]), .A2(n397), .B1(\A_s[43] ), .B2(n398), .ZN(
        n473) );
  INV_X1 U109 ( .A(\A_s[42] ), .ZN(n472) );
  INV_X1 U110 ( .A(A_ns[42]), .ZN(n471) );
  OAI221_X1 U111 ( .B1(n393), .B2(n474), .C1(n392), .C2(n475), .A(n476), .ZN(
        O[43]) );
  AOI22_X1 U112 ( .A1(A_ns[42]), .A2(n397), .B1(\A_s[42] ), .B2(n398), .ZN(
        n476) );
  INV_X1 U113 ( .A(\A_s[41] ), .ZN(n475) );
  INV_X1 U114 ( .A(A_ns[41]), .ZN(n474) );
  OAI221_X1 U115 ( .B1(n393), .B2(n477), .C1(n392), .C2(n478), .A(n479), .ZN(
        O[42]) );
  AOI22_X1 U116 ( .A1(A_ns[41]), .A2(n397), .B1(\A_s[41] ), .B2(n398), .ZN(
        n479) );
  INV_X1 U117 ( .A(\A_s[40] ), .ZN(n478) );
  INV_X1 U118 ( .A(A_ns[40]), .ZN(n477) );
  OAI221_X1 U119 ( .B1(n393), .B2(n480), .C1(n392), .C2(n481), .A(n482), .ZN(
        O[41]) );
  AOI22_X1 U120 ( .A1(A_ns[40]), .A2(n397), .B1(\A_s[40] ), .B2(n398), .ZN(
        n482) );
  INV_X1 U121 ( .A(\A_s[39] ), .ZN(n481) );
  INV_X1 U122 ( .A(A_ns[39]), .ZN(n480) );
  OAI221_X1 U123 ( .B1(n393), .B2(n483), .C1(n392), .C2(n484), .A(n485), .ZN(
        O[40]) );
  AOI22_X1 U124 ( .A1(A_ns[39]), .A2(n397), .B1(\A_s[39] ), .B2(n398), .ZN(
        n485) );
  INV_X1 U125 ( .A(\A_s[38] ), .ZN(n484) );
  INV_X1 U126 ( .A(A_ns[38]), .ZN(n483) );
  OAI221_X1 U127 ( .B1(n393), .B2(n486), .C1(n392), .C2(n487), .A(n488), .ZN(
        O[3]) );
  AOI22_X1 U128 ( .A1(A_ns[2]), .A2(n397), .B1(\A_s[2] ), .B2(n398), .ZN(n488)
         );
  INV_X1 U129 ( .A(\A_s[1] ), .ZN(n487) );
  INV_X1 U130 ( .A(A_ns[1]), .ZN(n486) );
  OAI221_X1 U131 ( .B1(n393), .B2(n489), .C1(n392), .C2(n490), .A(n491), .ZN(
        O[39]) );
  AOI22_X1 U132 ( .A1(A_ns[38]), .A2(n397), .B1(\A_s[38] ), .B2(n398), .ZN(
        n491) );
  INV_X1 U133 ( .A(\A_s[37] ), .ZN(n490) );
  INV_X1 U134 ( .A(A_ns[37]), .ZN(n489) );
  OAI221_X1 U135 ( .B1(n393), .B2(n492), .C1(n392), .C2(n493), .A(n494), .ZN(
        O[38]) );
  AOI22_X1 U136 ( .A1(A_ns[37]), .A2(n397), .B1(\A_s[37] ), .B2(n398), .ZN(
        n494) );
  INV_X1 U137 ( .A(\A_s[36] ), .ZN(n493) );
  INV_X1 U138 ( .A(A_ns[36]), .ZN(n492) );
  OAI221_X1 U139 ( .B1(n393), .B2(n495), .C1(n392), .C2(n496), .A(n497), .ZN(
        O[37]) );
  AOI22_X1 U140 ( .A1(A_ns[36]), .A2(n397), .B1(\A_s[36] ), .B2(n398), .ZN(
        n497) );
  INV_X1 U141 ( .A(\A_s[35] ), .ZN(n496) );
  INV_X1 U142 ( .A(A_ns[35]), .ZN(n495) );
  OAI221_X1 U143 ( .B1(n393), .B2(n498), .C1(n392), .C2(n499), .A(n500), .ZN(
        O[36]) );
  AOI22_X1 U144 ( .A1(A_ns[35]), .A2(n397), .B1(\A_s[35] ), .B2(n398), .ZN(
        n500) );
  INV_X1 U145 ( .A(\A_s[34] ), .ZN(n499) );
  INV_X1 U146 ( .A(A_ns[34]), .ZN(n498) );
  OAI221_X1 U147 ( .B1(n393), .B2(n501), .C1(n392), .C2(n502), .A(n503), .ZN(
        O[35]) );
  AOI22_X1 U148 ( .A1(A_ns[34]), .A2(n397), .B1(\A_s[34] ), .B2(n398), .ZN(
        n503) );
  INV_X1 U149 ( .A(\A_s[33] ), .ZN(n502) );
  INV_X1 U150 ( .A(A_ns[33]), .ZN(n501) );
  OAI221_X1 U151 ( .B1(n393), .B2(n504), .C1(n392), .C2(n505), .A(n506), .ZN(
        O[34]) );
  AOI22_X1 U152 ( .A1(A_ns[33]), .A2(n397), .B1(\A_s[33] ), .B2(n398), .ZN(
        n506) );
  INV_X1 U153 ( .A(\A_s[32] ), .ZN(n505) );
  INV_X1 U154 ( .A(A_ns[32]), .ZN(n504) );
  OAI221_X1 U155 ( .B1(n393), .B2(n507), .C1(n392), .C2(n508), .A(n509), .ZN(
        O[33]) );
  AOI22_X1 U156 ( .A1(A_ns[32]), .A2(n397), .B1(\A_s[32] ), .B2(n398), .ZN(
        n509) );
  INV_X1 U157 ( .A(\A_s[31] ), .ZN(n508) );
  INV_X1 U158 ( .A(A_ns[31]), .ZN(n507) );
  OAI221_X1 U159 ( .B1(n393), .B2(n510), .C1(n392), .C2(n511), .A(n512), .ZN(
        O[32]) );
  AOI22_X1 U160 ( .A1(A_ns[31]), .A2(n397), .B1(\A_s[31] ), .B2(n398), .ZN(
        n512) );
  INV_X1 U161 ( .A(\A_s[30] ), .ZN(n511) );
  INV_X1 U162 ( .A(A_ns[30]), .ZN(n510) );
  OAI221_X1 U163 ( .B1(n393), .B2(n513), .C1(n392), .C2(n514), .A(n515), .ZN(
        O[31]) );
  AOI22_X1 U164 ( .A1(A_ns[30]), .A2(n397), .B1(\A_s[30] ), .B2(n398), .ZN(
        n515) );
  INV_X1 U165 ( .A(\A_s[29] ), .ZN(n514) );
  INV_X1 U166 ( .A(A_ns[29]), .ZN(n513) );
  OAI221_X1 U167 ( .B1(n393), .B2(n516), .C1(n392), .C2(n517), .A(n518), .ZN(
        O[30]) );
  AOI22_X1 U168 ( .A1(A_ns[29]), .A2(n397), .B1(\A_s[29] ), .B2(n398), .ZN(
        n518) );
  INV_X1 U169 ( .A(\A_s[28] ), .ZN(n517) );
  INV_X1 U170 ( .A(A_ns[28]), .ZN(n516) );
  OAI221_X1 U171 ( .B1(n393), .B2(n519), .C1(n392), .C2(n520), .A(n521), .ZN(
        O[2]) );
  AOI22_X1 U172 ( .A1(A_ns[1]), .A2(n397), .B1(\A_s[1] ), .B2(n398), .ZN(n521)
         );
  OAI221_X1 U173 ( .B1(n393), .B2(n522), .C1(n392), .C2(n523), .A(n524), .ZN(
        O[29]) );
  AOI22_X1 U174 ( .A1(A_ns[28]), .A2(n397), .B1(\A_s[28] ), .B2(n398), .ZN(
        n524) );
  INV_X1 U175 ( .A(\A_s[27] ), .ZN(n523) );
  INV_X1 U176 ( .A(A_ns[27]), .ZN(n522) );
  OAI221_X1 U177 ( .B1(n393), .B2(n525), .C1(n392), .C2(n526), .A(n527), .ZN(
        O[28]) );
  AOI22_X1 U178 ( .A1(A_ns[27]), .A2(n397), .B1(\A_s[27] ), .B2(n398), .ZN(
        n527) );
  INV_X1 U179 ( .A(\A_s[26] ), .ZN(n526) );
  INV_X1 U180 ( .A(A_ns[26]), .ZN(n525) );
  OAI221_X1 U181 ( .B1(n393), .B2(n528), .C1(n392), .C2(n529), .A(n530), .ZN(
        O[27]) );
  AOI22_X1 U182 ( .A1(A_ns[26]), .A2(n397), .B1(\A_s[26] ), .B2(n398), .ZN(
        n530) );
  INV_X1 U183 ( .A(\A_s[25] ), .ZN(n529) );
  INV_X1 U184 ( .A(A_ns[25]), .ZN(n528) );
  OAI221_X1 U185 ( .B1(n393), .B2(n531), .C1(n392), .C2(n532), .A(n533), .ZN(
        O[26]) );
  AOI22_X1 U186 ( .A1(A_ns[25]), .A2(n397), .B1(\A_s[25] ), .B2(n398), .ZN(
        n533) );
  INV_X1 U187 ( .A(\A_s[24] ), .ZN(n532) );
  INV_X1 U188 ( .A(A_ns[24]), .ZN(n531) );
  OAI221_X1 U189 ( .B1(n393), .B2(n534), .C1(n392), .C2(n535), .A(n536), .ZN(
        O[25]) );
  AOI22_X1 U190 ( .A1(A_ns[24]), .A2(n397), .B1(\A_s[24] ), .B2(n398), .ZN(
        n536) );
  INV_X1 U191 ( .A(\A_s[23] ), .ZN(n535) );
  INV_X1 U192 ( .A(A_ns[23]), .ZN(n534) );
  OAI221_X1 U193 ( .B1(n393), .B2(n537), .C1(n392), .C2(n538), .A(n539), .ZN(
        O[24]) );
  AOI22_X1 U194 ( .A1(A_ns[23]), .A2(n397), .B1(\A_s[23] ), .B2(n398), .ZN(
        n539) );
  INV_X1 U195 ( .A(\A_s[22] ), .ZN(n538) );
  INV_X1 U196 ( .A(A_ns[22]), .ZN(n537) );
  OAI221_X1 U197 ( .B1(n393), .B2(n540), .C1(n392), .C2(n541), .A(n542), .ZN(
        O[23]) );
  AOI22_X1 U198 ( .A1(A_ns[22]), .A2(n397), .B1(\A_s[22] ), .B2(n398), .ZN(
        n542) );
  INV_X1 U199 ( .A(\A_s[21] ), .ZN(n541) );
  INV_X1 U200 ( .A(A_ns[21]), .ZN(n540) );
  OAI221_X1 U201 ( .B1(n393), .B2(n543), .C1(n392), .C2(n544), .A(n545), .ZN(
        O[22]) );
  AOI22_X1 U202 ( .A1(A_ns[21]), .A2(n397), .B1(\A_s[21] ), .B2(n398), .ZN(
        n545) );
  INV_X1 U203 ( .A(\A_s[20] ), .ZN(n544) );
  INV_X1 U204 ( .A(A_ns[20]), .ZN(n543) );
  OAI221_X1 U205 ( .B1(n393), .B2(n546), .C1(n392), .C2(n547), .A(n548), .ZN(
        O[21]) );
  AOI22_X1 U206 ( .A1(A_ns[20]), .A2(n397), .B1(\A_s[20] ), .B2(n398), .ZN(
        n548) );
  INV_X1 U207 ( .A(\A_s[19] ), .ZN(n547) );
  INV_X1 U208 ( .A(A_ns[19]), .ZN(n546) );
  OAI221_X1 U209 ( .B1(n393), .B2(n549), .C1(n392), .C2(n550), .A(n551), .ZN(
        O[20]) );
  AOI22_X1 U210 ( .A1(A_ns[19]), .A2(n397), .B1(\A_s[19] ), .B2(n398), .ZN(
        n551) );
  INV_X1 U211 ( .A(\A_s[18] ), .ZN(n550) );
  INV_X1 U212 ( .A(A_ns[18]), .ZN(n549) );
  OAI22_X1 U213 ( .A1(n552), .A2(n520), .B1(n553), .B2(n519), .ZN(O[1]) );
  INV_X1 U214 ( .A(A_ns[0]), .ZN(n519) );
  INV_X1 U215 ( .A(\A_s[0] ), .ZN(n520) );
  OAI221_X1 U216 ( .B1(n393), .B2(n554), .C1(n392), .C2(n555), .A(n556), .ZN(
        O[19]) );
  AOI22_X1 U217 ( .A1(A_ns[18]), .A2(n397), .B1(\A_s[18] ), .B2(n398), .ZN(
        n556) );
  INV_X1 U218 ( .A(\A_s[17] ), .ZN(n555) );
  INV_X1 U219 ( .A(A_ns[17]), .ZN(n554) );
  OAI221_X1 U220 ( .B1(n393), .B2(n557), .C1(n392), .C2(n558), .A(n559), .ZN(
        O[18]) );
  AOI22_X1 U221 ( .A1(A_ns[17]), .A2(n397), .B1(\A_s[17] ), .B2(n398), .ZN(
        n559) );
  INV_X1 U222 ( .A(\A_s[16] ), .ZN(n558) );
  INV_X1 U223 ( .A(A_ns[16]), .ZN(n557) );
  OAI221_X1 U224 ( .B1(n393), .B2(n560), .C1(n392), .C2(n561), .A(n562), .ZN(
        O[17]) );
  AOI22_X1 U225 ( .A1(A_ns[16]), .A2(n397), .B1(\A_s[16] ), .B2(n398), .ZN(
        n562) );
  INV_X1 U226 ( .A(\A_s[15] ), .ZN(n561) );
  INV_X1 U227 ( .A(A_ns[15]), .ZN(n560) );
  OAI221_X1 U228 ( .B1(n393), .B2(n563), .C1(n392), .C2(n564), .A(n565), .ZN(
        O[16]) );
  AOI22_X1 U229 ( .A1(A_ns[15]), .A2(n397), .B1(\A_s[15] ), .B2(n398), .ZN(
        n565) );
  INV_X1 U230 ( .A(\A_s[14] ), .ZN(n564) );
  INV_X1 U231 ( .A(A_ns[14]), .ZN(n563) );
  OAI221_X1 U232 ( .B1(n393), .B2(n566), .C1(n392), .C2(n567), .A(n568), .ZN(
        O[15]) );
  AOI22_X1 U233 ( .A1(A_ns[14]), .A2(n397), .B1(\A_s[14] ), .B2(n398), .ZN(
        n568) );
  INV_X1 U234 ( .A(\A_s[13] ), .ZN(n567) );
  INV_X1 U235 ( .A(A_ns[13]), .ZN(n566) );
  OAI221_X1 U236 ( .B1(n393), .B2(n569), .C1(n392), .C2(n570), .A(n571), .ZN(
        O[14]) );
  AOI22_X1 U237 ( .A1(A_ns[13]), .A2(n397), .B1(\A_s[13] ), .B2(n398), .ZN(
        n571) );
  INV_X1 U238 ( .A(\A_s[12] ), .ZN(n570) );
  INV_X1 U239 ( .A(A_ns[12]), .ZN(n569) );
  OAI221_X1 U240 ( .B1(n393), .B2(n572), .C1(n392), .C2(n573), .A(n574), .ZN(
        O[13]) );
  AOI22_X1 U241 ( .A1(A_ns[12]), .A2(n397), .B1(\A_s[12] ), .B2(n398), .ZN(
        n574) );
  INV_X1 U242 ( .A(\A_s[11] ), .ZN(n573) );
  INV_X1 U243 ( .A(A_ns[11]), .ZN(n572) );
  OAI221_X1 U244 ( .B1(n393), .B2(n575), .C1(n392), .C2(n576), .A(n577), .ZN(
        O[12]) );
  AOI22_X1 U245 ( .A1(A_ns[11]), .A2(n397), .B1(\A_s[11] ), .B2(n398), .ZN(
        n577) );
  INV_X1 U246 ( .A(\A_s[10] ), .ZN(n576) );
  INV_X1 U247 ( .A(A_ns[10]), .ZN(n575) );
  OAI221_X1 U248 ( .B1(n393), .B2(n578), .C1(n392), .C2(n579), .A(n580), .ZN(
        O[11]) );
  AOI22_X1 U249 ( .A1(A_ns[10]), .A2(n397), .B1(\A_s[10] ), .B2(n398), .ZN(
        n580) );
  INV_X1 U250 ( .A(\A_s[9] ), .ZN(n579) );
  INV_X1 U251 ( .A(A_ns[9]), .ZN(n578) );
  OAI221_X1 U252 ( .B1(n581), .B2(n393), .C1(n582), .C2(n392), .A(n583), .ZN(
        O[10]) );
  AOI22_X1 U253 ( .A1(A_ns[9]), .A2(n397), .B1(\A_s[9] ), .B2(n398), .ZN(n583)
         );
  NAND2_X1 U254 ( .A1(n584), .A2(n552), .ZN(n553) );
  NAND2_X1 U255 ( .A1(n584), .A2(n585), .ZN(n552) );
  XOR2_X1 U256 ( .A(B[7]), .B(B[8]), .Z(n584) );
  INV_X1 U257 ( .A(\A_s[8] ), .ZN(n582) );
  INV_X1 U258 ( .A(B[9]), .ZN(n585) );
  INV_X1 U259 ( .A(A_ns[8]), .ZN(n581) );
endmodule


module BOOTHENC_NBIT64_i10 ( A, A_n, A_ns, A_s, B, O, A_so, A_nso );
  input [63:0] A;
  input [63:0] A_n;
  input [63:0] A_ns;
  input [63:0] A_s;
  input [63:0] B;
  output [63:0] O;
  output [63:0] A_so;
  output [63:0] A_nso;
  wire   \A_s[61] , \A_s[60] , \A_s[59] , \A_s[58] , \A_s[57] , \A_s[56] ,
         \A_s[55] , \A_s[54] , \A_s[53] , \A_s[52] , \A_s[51] , \A_s[50] ,
         \A_s[49] , \A_s[48] , \A_s[47] , \A_s[46] , \A_s[45] , \A_s[44] ,
         \A_s[43] , \A_s[42] , \A_s[41] , \A_s[40] , \A_s[39] , \A_s[38] ,
         \A_s[37] , \A_s[36] , \A_s[35] , \A_s[34] , \A_s[33] , \A_s[32] ,
         \A_s[31] , \A_s[30] , \A_s[29] , \A_s[28] , \A_s[27] , \A_s[26] ,
         \A_s[25] , \A_s[24] , \A_s[23] , \A_s[22] , \A_s[21] , \A_s[20] ,
         \A_s[19] , \A_s[18] , \A_s[17] , \A_s[16] , \A_s[15] , \A_s[14] ,
         \A_s[13] , \A_s[12] , \A_s[11] , \A_s[10] , \A_s[9] , \A_s[8] ,
         \A_s[7] , \A_s[6] , \A_s[5] , \A_s[4] , \A_s[3] , \A_s[2] , \A_s[1] ,
         \A_s[0] , n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585;
  assign A_nso[0] = 1'b0;
  assign A_nso[1] = 1'b0;
  assign A_so[0] = 1'b0;
  assign A_so[1] = 1'b0;
  assign O[0] = 1'b0;
  assign A_nso[63] = \A_s[61] ;
  assign A_so[63] = \A_s[61] ;
  assign \A_s[61]  = A_s[61];
  assign A_nso[62] = \A_s[60] ;
  assign A_so[62] = \A_s[60] ;
  assign \A_s[60]  = A_s[60];
  assign A_nso[61] = \A_s[59] ;
  assign A_so[61] = \A_s[59] ;
  assign \A_s[59]  = A_s[59];
  assign A_nso[60] = \A_s[58] ;
  assign A_so[60] = \A_s[58] ;
  assign \A_s[58]  = A_s[58];
  assign A_nso[59] = \A_s[57] ;
  assign A_so[59] = \A_s[57] ;
  assign \A_s[57]  = A_s[57];
  assign A_nso[58] = \A_s[56] ;
  assign A_so[58] = \A_s[56] ;
  assign \A_s[56]  = A_s[56];
  assign A_nso[57] = \A_s[55] ;
  assign A_so[57] = \A_s[55] ;
  assign \A_s[55]  = A_s[55];
  assign A_nso[56] = \A_s[54] ;
  assign A_so[56] = \A_s[54] ;
  assign \A_s[54]  = A_s[54];
  assign A_nso[55] = \A_s[53] ;
  assign A_so[55] = \A_s[53] ;
  assign \A_s[53]  = A_s[53];
  assign A_nso[54] = \A_s[52] ;
  assign A_so[54] = \A_s[52] ;
  assign \A_s[52]  = A_s[52];
  assign A_nso[53] = \A_s[51] ;
  assign A_so[53] = \A_s[51] ;
  assign \A_s[51]  = A_s[51];
  assign A_nso[52] = \A_s[50] ;
  assign A_so[52] = \A_s[50] ;
  assign \A_s[50]  = A_s[50];
  assign A_nso[51] = \A_s[49] ;
  assign A_so[51] = \A_s[49] ;
  assign \A_s[49]  = A_s[49];
  assign A_nso[50] = \A_s[48] ;
  assign A_so[50] = \A_s[48] ;
  assign \A_s[48]  = A_s[48];
  assign A_nso[49] = \A_s[47] ;
  assign A_so[49] = \A_s[47] ;
  assign \A_s[47]  = A_s[47];
  assign A_nso[48] = \A_s[46] ;
  assign A_so[48] = \A_s[46] ;
  assign \A_s[46]  = A_s[46];
  assign A_nso[47] = \A_s[45] ;
  assign A_so[47] = \A_s[45] ;
  assign \A_s[45]  = A_s[45];
  assign A_nso[46] = \A_s[44] ;
  assign A_so[46] = \A_s[44] ;
  assign \A_s[44]  = A_s[44];
  assign A_nso[45] = \A_s[43] ;
  assign A_so[45] = \A_s[43] ;
  assign \A_s[43]  = A_s[43];
  assign A_nso[44] = \A_s[42] ;
  assign A_so[44] = \A_s[42] ;
  assign \A_s[42]  = A_s[42];
  assign A_nso[43] = \A_s[41] ;
  assign A_so[43] = \A_s[41] ;
  assign \A_s[41]  = A_s[41];
  assign A_nso[42] = \A_s[40] ;
  assign A_so[42] = \A_s[40] ;
  assign \A_s[40]  = A_s[40];
  assign A_nso[41] = \A_s[39] ;
  assign A_so[41] = \A_s[39] ;
  assign \A_s[39]  = A_s[39];
  assign A_nso[40] = \A_s[38] ;
  assign A_so[40] = \A_s[38] ;
  assign \A_s[38]  = A_s[38];
  assign A_nso[39] = \A_s[37] ;
  assign A_so[39] = \A_s[37] ;
  assign \A_s[37]  = A_s[37];
  assign A_nso[38] = \A_s[36] ;
  assign A_so[38] = \A_s[36] ;
  assign \A_s[36]  = A_s[36];
  assign A_nso[37] = \A_s[35] ;
  assign A_so[37] = \A_s[35] ;
  assign \A_s[35]  = A_s[35];
  assign A_nso[36] = \A_s[34] ;
  assign A_so[36] = \A_s[34] ;
  assign \A_s[34]  = A_s[34];
  assign A_nso[35] = \A_s[33] ;
  assign A_so[35] = \A_s[33] ;
  assign \A_s[33]  = A_s[33];
  assign A_nso[34] = \A_s[32] ;
  assign A_so[34] = \A_s[32] ;
  assign \A_s[32]  = A_s[32];
  assign A_nso[33] = \A_s[31] ;
  assign A_so[33] = \A_s[31] ;
  assign \A_s[31]  = A_s[31];
  assign A_nso[32] = \A_s[30] ;
  assign A_so[32] = \A_s[30] ;
  assign \A_s[30]  = A_s[30];
  assign A_nso[31] = \A_s[29] ;
  assign A_so[31] = \A_s[29] ;
  assign \A_s[29]  = A_s[29];
  assign A_nso[30] = \A_s[28] ;
  assign A_so[30] = \A_s[28] ;
  assign \A_s[28]  = A_s[28];
  assign A_nso[29] = \A_s[27] ;
  assign A_so[29] = \A_s[27] ;
  assign \A_s[27]  = A_s[27];
  assign A_nso[28] = \A_s[26] ;
  assign A_so[28] = \A_s[26] ;
  assign \A_s[26]  = A_s[26];
  assign A_nso[27] = \A_s[25] ;
  assign A_so[27] = \A_s[25] ;
  assign \A_s[25]  = A_s[25];
  assign A_nso[26] = \A_s[24] ;
  assign A_so[26] = \A_s[24] ;
  assign \A_s[24]  = A_s[24];
  assign A_nso[25] = \A_s[23] ;
  assign A_so[25] = \A_s[23] ;
  assign \A_s[23]  = A_s[23];
  assign A_nso[24] = \A_s[22] ;
  assign A_so[24] = \A_s[22] ;
  assign \A_s[22]  = A_s[22];
  assign A_nso[23] = \A_s[21] ;
  assign A_so[23] = \A_s[21] ;
  assign \A_s[21]  = A_s[21];
  assign A_nso[22] = \A_s[20] ;
  assign A_so[22] = \A_s[20] ;
  assign \A_s[20]  = A_s[20];
  assign A_nso[21] = \A_s[19] ;
  assign A_so[21] = \A_s[19] ;
  assign \A_s[19]  = A_s[19];
  assign A_nso[20] = \A_s[18] ;
  assign A_so[20] = \A_s[18] ;
  assign \A_s[18]  = A_s[18];
  assign A_nso[19] = \A_s[17] ;
  assign A_so[19] = \A_s[17] ;
  assign \A_s[17]  = A_s[17];
  assign A_nso[18] = \A_s[16] ;
  assign A_so[18] = \A_s[16] ;
  assign \A_s[16]  = A_s[16];
  assign A_nso[17] = \A_s[15] ;
  assign A_so[17] = \A_s[15] ;
  assign \A_s[15]  = A_s[15];
  assign A_nso[16] = \A_s[14] ;
  assign A_so[16] = \A_s[14] ;
  assign \A_s[14]  = A_s[14];
  assign A_nso[15] = \A_s[13] ;
  assign A_so[15] = \A_s[13] ;
  assign \A_s[13]  = A_s[13];
  assign A_nso[14] = \A_s[12] ;
  assign A_so[14] = \A_s[12] ;
  assign \A_s[12]  = A_s[12];
  assign A_nso[13] = \A_s[11] ;
  assign A_so[13] = \A_s[11] ;
  assign \A_s[11]  = A_s[11];
  assign A_nso[12] = \A_s[10] ;
  assign A_so[12] = \A_s[10] ;
  assign \A_s[10]  = A_s[10];
  assign A_nso[11] = \A_s[9] ;
  assign A_so[11] = \A_s[9] ;
  assign \A_s[9]  = A_s[9];
  assign A_nso[10] = \A_s[8] ;
  assign A_so[10] = \A_s[8] ;
  assign \A_s[8]  = A_s[8];
  assign A_nso[9] = \A_s[7] ;
  assign A_so[9] = \A_s[7] ;
  assign \A_s[7]  = A_s[7];
  assign A_nso[8] = \A_s[6] ;
  assign A_so[8] = \A_s[6] ;
  assign \A_s[6]  = A_s[6];
  assign A_nso[7] = \A_s[5] ;
  assign A_so[7] = \A_s[5] ;
  assign \A_s[5]  = A_s[5];
  assign A_nso[6] = \A_s[4] ;
  assign A_so[6] = \A_s[4] ;
  assign \A_s[4]  = A_s[4];
  assign A_nso[5] = \A_s[3] ;
  assign A_so[5] = \A_s[3] ;
  assign \A_s[3]  = A_s[3];
  assign A_nso[4] = \A_s[2] ;
  assign A_so[4] = \A_s[2] ;
  assign \A_s[2]  = A_s[2];
  assign A_nso[3] = \A_s[1] ;
  assign A_so[3] = \A_s[1] ;
  assign \A_s[1]  = A_s[1];
  assign A_nso[2] = \A_s[0] ;
  assign A_so[2] = \A_s[0] ;
  assign \A_s[0]  = A_s[0];

  AND3_X1 U2 ( .A1(B[9]), .A2(n585), .A3(B[10]), .ZN(n391) );
  INV_X4 U3 ( .A(n391), .ZN(n392) );
  INV_X4 U4 ( .A(n552), .ZN(n398) );
  OR3_X4 U5 ( .A1(B[10]), .A2(B[9]), .A3(n585), .ZN(n393) );
  INV_X4 U6 ( .A(n553), .ZN(n397) );
  OAI221_X1 U7 ( .B1(n393), .B2(n394), .C1(n392), .C2(n395), .A(n396), .ZN(
        O[9]) );
  AOI22_X1 U8 ( .A1(A_ns[8]), .A2(n397), .B1(\A_s[8] ), .B2(n398), .ZN(n396)
         );
  INV_X1 U9 ( .A(\A_s[7] ), .ZN(n395) );
  INV_X1 U10 ( .A(A_ns[7]), .ZN(n394) );
  OAI221_X1 U11 ( .B1(n393), .B2(n399), .C1(n392), .C2(n400), .A(n401), .ZN(
        O[8]) );
  AOI22_X1 U12 ( .A1(A_ns[7]), .A2(n397), .B1(\A_s[7] ), .B2(n398), .ZN(n401)
         );
  INV_X1 U13 ( .A(\A_s[6] ), .ZN(n400) );
  INV_X1 U14 ( .A(A_ns[6]), .ZN(n399) );
  OAI221_X1 U15 ( .B1(n393), .B2(n402), .C1(n392), .C2(n403), .A(n404), .ZN(
        O[7]) );
  AOI22_X1 U16 ( .A1(A_ns[6]), .A2(n397), .B1(\A_s[6] ), .B2(n398), .ZN(n404)
         );
  INV_X1 U17 ( .A(\A_s[5] ), .ZN(n403) );
  INV_X1 U18 ( .A(A_ns[5]), .ZN(n402) );
  OAI221_X1 U19 ( .B1(n393), .B2(n405), .C1(n392), .C2(n406), .A(n407), .ZN(
        O[6]) );
  AOI22_X1 U20 ( .A1(A_ns[5]), .A2(n397), .B1(\A_s[5] ), .B2(n398), .ZN(n407)
         );
  INV_X1 U21 ( .A(\A_s[4] ), .ZN(n406) );
  INV_X1 U22 ( .A(A_ns[4]), .ZN(n405) );
  OAI221_X1 U23 ( .B1(n393), .B2(n408), .C1(n392), .C2(n409), .A(n410), .ZN(
        O[63]) );
  AOI22_X1 U24 ( .A1(A_ns[62]), .A2(n397), .B1(A_s[62]), .B2(n398), .ZN(n410)
         );
  INV_X1 U25 ( .A(\A_s[61] ), .ZN(n409) );
  INV_X1 U26 ( .A(A_ns[61]), .ZN(n408) );
  OAI221_X1 U27 ( .B1(n393), .B2(n411), .C1(n392), .C2(n412), .A(n413), .ZN(
        O[62]) );
  AOI22_X1 U28 ( .A1(A_ns[61]), .A2(n397), .B1(\A_s[61] ), .B2(n398), .ZN(n413) );
  INV_X1 U29 ( .A(\A_s[60] ), .ZN(n412) );
  INV_X1 U30 ( .A(A_ns[60]), .ZN(n411) );
  OAI221_X1 U31 ( .B1(n393), .B2(n414), .C1(n392), .C2(n415), .A(n416), .ZN(
        O[61]) );
  AOI22_X1 U32 ( .A1(A_ns[60]), .A2(n397), .B1(\A_s[60] ), .B2(n398), .ZN(n416) );
  INV_X1 U33 ( .A(\A_s[59] ), .ZN(n415) );
  INV_X1 U34 ( .A(A_ns[59]), .ZN(n414) );
  OAI221_X1 U35 ( .B1(n393), .B2(n417), .C1(n392), .C2(n418), .A(n419), .ZN(
        O[60]) );
  AOI22_X1 U36 ( .A1(A_ns[59]), .A2(n397), .B1(\A_s[59] ), .B2(n398), .ZN(n419) );
  INV_X1 U37 ( .A(\A_s[58] ), .ZN(n418) );
  INV_X1 U38 ( .A(A_ns[58]), .ZN(n417) );
  OAI221_X1 U39 ( .B1(n393), .B2(n420), .C1(n392), .C2(n421), .A(n422), .ZN(
        O[5]) );
  AOI22_X1 U40 ( .A1(A_ns[4]), .A2(n397), .B1(\A_s[4] ), .B2(n398), .ZN(n422)
         );
  INV_X1 U41 ( .A(\A_s[3] ), .ZN(n421) );
  INV_X1 U42 ( .A(A_ns[3]), .ZN(n420) );
  OAI221_X1 U43 ( .B1(n393), .B2(n423), .C1(n392), .C2(n424), .A(n425), .ZN(
        O[59]) );
  AOI22_X1 U44 ( .A1(A_ns[58]), .A2(n397), .B1(\A_s[58] ), .B2(n398), .ZN(n425) );
  INV_X1 U45 ( .A(\A_s[57] ), .ZN(n424) );
  INV_X1 U46 ( .A(A_ns[57]), .ZN(n423) );
  OAI221_X1 U47 ( .B1(n393), .B2(n426), .C1(n392), .C2(n427), .A(n428), .ZN(
        O[58]) );
  AOI22_X1 U48 ( .A1(A_ns[57]), .A2(n397), .B1(\A_s[57] ), .B2(n398), .ZN(n428) );
  INV_X1 U49 ( .A(\A_s[56] ), .ZN(n427) );
  INV_X1 U50 ( .A(A_ns[56]), .ZN(n426) );
  OAI221_X1 U51 ( .B1(n393), .B2(n429), .C1(n392), .C2(n430), .A(n431), .ZN(
        O[57]) );
  AOI22_X1 U52 ( .A1(A_ns[56]), .A2(n397), .B1(\A_s[56] ), .B2(n398), .ZN(n431) );
  INV_X1 U53 ( .A(\A_s[55] ), .ZN(n430) );
  INV_X1 U54 ( .A(A_ns[55]), .ZN(n429) );
  OAI221_X1 U55 ( .B1(n393), .B2(n432), .C1(n392), .C2(n433), .A(n434), .ZN(
        O[56]) );
  AOI22_X1 U56 ( .A1(A_ns[55]), .A2(n397), .B1(\A_s[55] ), .B2(n398), .ZN(n434) );
  INV_X1 U57 ( .A(\A_s[54] ), .ZN(n433) );
  INV_X1 U58 ( .A(A_ns[54]), .ZN(n432) );
  OAI221_X1 U59 ( .B1(n393), .B2(n435), .C1(n392), .C2(n436), .A(n437), .ZN(
        O[55]) );
  AOI22_X1 U60 ( .A1(A_ns[54]), .A2(n397), .B1(\A_s[54] ), .B2(n398), .ZN(n437) );
  INV_X1 U61 ( .A(\A_s[53] ), .ZN(n436) );
  INV_X1 U62 ( .A(A_ns[53]), .ZN(n435) );
  OAI221_X1 U63 ( .B1(n393), .B2(n438), .C1(n392), .C2(n439), .A(n440), .ZN(
        O[54]) );
  AOI22_X1 U64 ( .A1(A_ns[53]), .A2(n397), .B1(\A_s[53] ), .B2(n398), .ZN(n440) );
  INV_X1 U65 ( .A(\A_s[52] ), .ZN(n439) );
  INV_X1 U66 ( .A(A_ns[52]), .ZN(n438) );
  OAI221_X1 U67 ( .B1(n393), .B2(n441), .C1(n392), .C2(n442), .A(n443), .ZN(
        O[53]) );
  AOI22_X1 U68 ( .A1(A_ns[52]), .A2(n397), .B1(\A_s[52] ), .B2(n398), .ZN(n443) );
  INV_X1 U69 ( .A(\A_s[51] ), .ZN(n442) );
  INV_X1 U70 ( .A(A_ns[51]), .ZN(n441) );
  OAI221_X1 U71 ( .B1(n393), .B2(n444), .C1(n392), .C2(n445), .A(n446), .ZN(
        O[52]) );
  AOI22_X1 U72 ( .A1(A_ns[51]), .A2(n397), .B1(\A_s[51] ), .B2(n398), .ZN(n446) );
  INV_X1 U73 ( .A(\A_s[50] ), .ZN(n445) );
  INV_X1 U74 ( .A(A_ns[50]), .ZN(n444) );
  OAI221_X1 U75 ( .B1(n393), .B2(n447), .C1(n392), .C2(n448), .A(n449), .ZN(
        O[51]) );
  AOI22_X1 U76 ( .A1(A_ns[50]), .A2(n397), .B1(\A_s[50] ), .B2(n398), .ZN(n449) );
  INV_X1 U77 ( .A(\A_s[49] ), .ZN(n448) );
  INV_X1 U78 ( .A(A_ns[49]), .ZN(n447) );
  OAI221_X1 U79 ( .B1(n393), .B2(n450), .C1(n392), .C2(n451), .A(n452), .ZN(
        O[50]) );
  AOI22_X1 U80 ( .A1(A_ns[49]), .A2(n397), .B1(\A_s[49] ), .B2(n398), .ZN(n452) );
  INV_X1 U81 ( .A(\A_s[48] ), .ZN(n451) );
  INV_X1 U82 ( .A(A_ns[48]), .ZN(n450) );
  OAI221_X1 U83 ( .B1(n393), .B2(n453), .C1(n392), .C2(n454), .A(n455), .ZN(
        O[4]) );
  AOI22_X1 U84 ( .A1(A_ns[3]), .A2(n397), .B1(\A_s[3] ), .B2(n398), .ZN(n455)
         );
  INV_X1 U85 ( .A(\A_s[2] ), .ZN(n454) );
  INV_X1 U86 ( .A(A_ns[2]), .ZN(n453) );
  OAI221_X1 U87 ( .B1(n393), .B2(n456), .C1(n392), .C2(n457), .A(n458), .ZN(
        O[49]) );
  AOI22_X1 U88 ( .A1(A_ns[48]), .A2(n397), .B1(\A_s[48] ), .B2(n398), .ZN(n458) );
  INV_X1 U89 ( .A(\A_s[47] ), .ZN(n457) );
  INV_X1 U90 ( .A(A_ns[47]), .ZN(n456) );
  OAI221_X1 U91 ( .B1(n393), .B2(n459), .C1(n392), .C2(n460), .A(n461), .ZN(
        O[48]) );
  AOI22_X1 U92 ( .A1(A_ns[47]), .A2(n397), .B1(\A_s[47] ), .B2(n398), .ZN(n461) );
  INV_X1 U93 ( .A(\A_s[46] ), .ZN(n460) );
  INV_X1 U94 ( .A(A_ns[46]), .ZN(n459) );
  OAI221_X1 U95 ( .B1(n393), .B2(n462), .C1(n392), .C2(n463), .A(n464), .ZN(
        O[47]) );
  AOI22_X1 U96 ( .A1(A_ns[46]), .A2(n397), .B1(\A_s[46] ), .B2(n398), .ZN(n464) );
  INV_X1 U97 ( .A(\A_s[45] ), .ZN(n463) );
  INV_X1 U98 ( .A(A_ns[45]), .ZN(n462) );
  OAI221_X1 U99 ( .B1(n393), .B2(n465), .C1(n392), .C2(n466), .A(n467), .ZN(
        O[46]) );
  AOI22_X1 U100 ( .A1(A_ns[45]), .A2(n397), .B1(\A_s[45] ), .B2(n398), .ZN(
        n467) );
  INV_X1 U101 ( .A(\A_s[44] ), .ZN(n466) );
  INV_X1 U102 ( .A(A_ns[44]), .ZN(n465) );
  OAI221_X1 U103 ( .B1(n393), .B2(n468), .C1(n392), .C2(n469), .A(n470), .ZN(
        O[45]) );
  AOI22_X1 U104 ( .A1(A_ns[44]), .A2(n397), .B1(\A_s[44] ), .B2(n398), .ZN(
        n470) );
  INV_X1 U105 ( .A(\A_s[43] ), .ZN(n469) );
  INV_X1 U106 ( .A(A_ns[43]), .ZN(n468) );
  OAI221_X1 U107 ( .B1(n393), .B2(n471), .C1(n392), .C2(n472), .A(n473), .ZN(
        O[44]) );
  AOI22_X1 U108 ( .A1(A_ns[43]), .A2(n397), .B1(\A_s[43] ), .B2(n398), .ZN(
        n473) );
  INV_X1 U109 ( .A(\A_s[42] ), .ZN(n472) );
  INV_X1 U110 ( .A(A_ns[42]), .ZN(n471) );
  OAI221_X1 U111 ( .B1(n393), .B2(n474), .C1(n392), .C2(n475), .A(n476), .ZN(
        O[43]) );
  AOI22_X1 U112 ( .A1(A_ns[42]), .A2(n397), .B1(\A_s[42] ), .B2(n398), .ZN(
        n476) );
  INV_X1 U113 ( .A(\A_s[41] ), .ZN(n475) );
  INV_X1 U114 ( .A(A_ns[41]), .ZN(n474) );
  OAI221_X1 U115 ( .B1(n393), .B2(n477), .C1(n392), .C2(n478), .A(n479), .ZN(
        O[42]) );
  AOI22_X1 U116 ( .A1(A_ns[41]), .A2(n397), .B1(\A_s[41] ), .B2(n398), .ZN(
        n479) );
  INV_X1 U117 ( .A(\A_s[40] ), .ZN(n478) );
  INV_X1 U118 ( .A(A_ns[40]), .ZN(n477) );
  OAI221_X1 U119 ( .B1(n393), .B2(n480), .C1(n392), .C2(n481), .A(n482), .ZN(
        O[41]) );
  AOI22_X1 U120 ( .A1(A_ns[40]), .A2(n397), .B1(\A_s[40] ), .B2(n398), .ZN(
        n482) );
  INV_X1 U121 ( .A(\A_s[39] ), .ZN(n481) );
  INV_X1 U122 ( .A(A_ns[39]), .ZN(n480) );
  OAI221_X1 U123 ( .B1(n393), .B2(n483), .C1(n392), .C2(n484), .A(n485), .ZN(
        O[40]) );
  AOI22_X1 U124 ( .A1(A_ns[39]), .A2(n397), .B1(\A_s[39] ), .B2(n398), .ZN(
        n485) );
  INV_X1 U125 ( .A(\A_s[38] ), .ZN(n484) );
  INV_X1 U126 ( .A(A_ns[38]), .ZN(n483) );
  OAI221_X1 U127 ( .B1(n393), .B2(n486), .C1(n392), .C2(n487), .A(n488), .ZN(
        O[3]) );
  AOI22_X1 U128 ( .A1(A_ns[2]), .A2(n397), .B1(\A_s[2] ), .B2(n398), .ZN(n488)
         );
  INV_X1 U129 ( .A(\A_s[1] ), .ZN(n487) );
  INV_X1 U130 ( .A(A_ns[1]), .ZN(n486) );
  OAI221_X1 U131 ( .B1(n393), .B2(n489), .C1(n392), .C2(n490), .A(n491), .ZN(
        O[39]) );
  AOI22_X1 U132 ( .A1(A_ns[38]), .A2(n397), .B1(\A_s[38] ), .B2(n398), .ZN(
        n491) );
  INV_X1 U133 ( .A(\A_s[37] ), .ZN(n490) );
  INV_X1 U134 ( .A(A_ns[37]), .ZN(n489) );
  OAI221_X1 U135 ( .B1(n393), .B2(n492), .C1(n392), .C2(n493), .A(n494), .ZN(
        O[38]) );
  AOI22_X1 U136 ( .A1(A_ns[37]), .A2(n397), .B1(\A_s[37] ), .B2(n398), .ZN(
        n494) );
  INV_X1 U137 ( .A(\A_s[36] ), .ZN(n493) );
  INV_X1 U138 ( .A(A_ns[36]), .ZN(n492) );
  OAI221_X1 U139 ( .B1(n393), .B2(n495), .C1(n392), .C2(n496), .A(n497), .ZN(
        O[37]) );
  AOI22_X1 U140 ( .A1(A_ns[36]), .A2(n397), .B1(\A_s[36] ), .B2(n398), .ZN(
        n497) );
  INV_X1 U141 ( .A(\A_s[35] ), .ZN(n496) );
  INV_X1 U142 ( .A(A_ns[35]), .ZN(n495) );
  OAI221_X1 U143 ( .B1(n393), .B2(n498), .C1(n392), .C2(n499), .A(n500), .ZN(
        O[36]) );
  AOI22_X1 U144 ( .A1(A_ns[35]), .A2(n397), .B1(\A_s[35] ), .B2(n398), .ZN(
        n500) );
  INV_X1 U145 ( .A(\A_s[34] ), .ZN(n499) );
  INV_X1 U146 ( .A(A_ns[34]), .ZN(n498) );
  OAI221_X1 U147 ( .B1(n393), .B2(n501), .C1(n392), .C2(n502), .A(n503), .ZN(
        O[35]) );
  AOI22_X1 U148 ( .A1(A_ns[34]), .A2(n397), .B1(\A_s[34] ), .B2(n398), .ZN(
        n503) );
  INV_X1 U149 ( .A(\A_s[33] ), .ZN(n502) );
  INV_X1 U150 ( .A(A_ns[33]), .ZN(n501) );
  OAI221_X1 U151 ( .B1(n393), .B2(n504), .C1(n392), .C2(n505), .A(n506), .ZN(
        O[34]) );
  AOI22_X1 U152 ( .A1(A_ns[33]), .A2(n397), .B1(\A_s[33] ), .B2(n398), .ZN(
        n506) );
  INV_X1 U153 ( .A(\A_s[32] ), .ZN(n505) );
  INV_X1 U154 ( .A(A_ns[32]), .ZN(n504) );
  OAI221_X1 U155 ( .B1(n393), .B2(n507), .C1(n392), .C2(n508), .A(n509), .ZN(
        O[33]) );
  AOI22_X1 U156 ( .A1(A_ns[32]), .A2(n397), .B1(\A_s[32] ), .B2(n398), .ZN(
        n509) );
  INV_X1 U157 ( .A(\A_s[31] ), .ZN(n508) );
  INV_X1 U158 ( .A(A_ns[31]), .ZN(n507) );
  OAI221_X1 U159 ( .B1(n393), .B2(n510), .C1(n392), .C2(n511), .A(n512), .ZN(
        O[32]) );
  AOI22_X1 U160 ( .A1(A_ns[31]), .A2(n397), .B1(\A_s[31] ), .B2(n398), .ZN(
        n512) );
  INV_X1 U161 ( .A(\A_s[30] ), .ZN(n511) );
  INV_X1 U162 ( .A(A_ns[30]), .ZN(n510) );
  OAI221_X1 U163 ( .B1(n393), .B2(n513), .C1(n392), .C2(n514), .A(n515), .ZN(
        O[31]) );
  AOI22_X1 U164 ( .A1(A_ns[30]), .A2(n397), .B1(\A_s[30] ), .B2(n398), .ZN(
        n515) );
  INV_X1 U165 ( .A(\A_s[29] ), .ZN(n514) );
  INV_X1 U166 ( .A(A_ns[29]), .ZN(n513) );
  OAI221_X1 U167 ( .B1(n393), .B2(n516), .C1(n392), .C2(n517), .A(n518), .ZN(
        O[30]) );
  AOI22_X1 U168 ( .A1(A_ns[29]), .A2(n397), .B1(\A_s[29] ), .B2(n398), .ZN(
        n518) );
  INV_X1 U169 ( .A(\A_s[28] ), .ZN(n517) );
  INV_X1 U170 ( .A(A_ns[28]), .ZN(n516) );
  OAI221_X1 U171 ( .B1(n393), .B2(n519), .C1(n392), .C2(n520), .A(n521), .ZN(
        O[2]) );
  AOI22_X1 U172 ( .A1(A_ns[1]), .A2(n397), .B1(\A_s[1] ), .B2(n398), .ZN(n521)
         );
  OAI221_X1 U173 ( .B1(n393), .B2(n522), .C1(n392), .C2(n523), .A(n524), .ZN(
        O[29]) );
  AOI22_X1 U174 ( .A1(A_ns[28]), .A2(n397), .B1(\A_s[28] ), .B2(n398), .ZN(
        n524) );
  INV_X1 U175 ( .A(\A_s[27] ), .ZN(n523) );
  INV_X1 U176 ( .A(A_ns[27]), .ZN(n522) );
  OAI221_X1 U177 ( .B1(n393), .B2(n525), .C1(n392), .C2(n526), .A(n527), .ZN(
        O[28]) );
  AOI22_X1 U178 ( .A1(A_ns[27]), .A2(n397), .B1(\A_s[27] ), .B2(n398), .ZN(
        n527) );
  INV_X1 U179 ( .A(\A_s[26] ), .ZN(n526) );
  INV_X1 U180 ( .A(A_ns[26]), .ZN(n525) );
  OAI221_X1 U181 ( .B1(n393), .B2(n528), .C1(n392), .C2(n529), .A(n530), .ZN(
        O[27]) );
  AOI22_X1 U182 ( .A1(A_ns[26]), .A2(n397), .B1(\A_s[26] ), .B2(n398), .ZN(
        n530) );
  INV_X1 U183 ( .A(\A_s[25] ), .ZN(n529) );
  INV_X1 U184 ( .A(A_ns[25]), .ZN(n528) );
  OAI221_X1 U185 ( .B1(n393), .B2(n531), .C1(n392), .C2(n532), .A(n533), .ZN(
        O[26]) );
  AOI22_X1 U186 ( .A1(A_ns[25]), .A2(n397), .B1(\A_s[25] ), .B2(n398), .ZN(
        n533) );
  INV_X1 U187 ( .A(\A_s[24] ), .ZN(n532) );
  INV_X1 U188 ( .A(A_ns[24]), .ZN(n531) );
  OAI221_X1 U189 ( .B1(n393), .B2(n534), .C1(n392), .C2(n535), .A(n536), .ZN(
        O[25]) );
  AOI22_X1 U190 ( .A1(A_ns[24]), .A2(n397), .B1(\A_s[24] ), .B2(n398), .ZN(
        n536) );
  INV_X1 U191 ( .A(\A_s[23] ), .ZN(n535) );
  INV_X1 U192 ( .A(A_ns[23]), .ZN(n534) );
  OAI221_X1 U193 ( .B1(n393), .B2(n537), .C1(n392), .C2(n538), .A(n539), .ZN(
        O[24]) );
  AOI22_X1 U194 ( .A1(A_ns[23]), .A2(n397), .B1(\A_s[23] ), .B2(n398), .ZN(
        n539) );
  INV_X1 U195 ( .A(\A_s[22] ), .ZN(n538) );
  INV_X1 U196 ( .A(A_ns[22]), .ZN(n537) );
  OAI221_X1 U197 ( .B1(n393), .B2(n540), .C1(n392), .C2(n541), .A(n542), .ZN(
        O[23]) );
  AOI22_X1 U198 ( .A1(A_ns[22]), .A2(n397), .B1(\A_s[22] ), .B2(n398), .ZN(
        n542) );
  INV_X1 U199 ( .A(\A_s[21] ), .ZN(n541) );
  INV_X1 U200 ( .A(A_ns[21]), .ZN(n540) );
  OAI221_X1 U201 ( .B1(n393), .B2(n543), .C1(n392), .C2(n544), .A(n545), .ZN(
        O[22]) );
  AOI22_X1 U202 ( .A1(A_ns[21]), .A2(n397), .B1(\A_s[21] ), .B2(n398), .ZN(
        n545) );
  INV_X1 U203 ( .A(\A_s[20] ), .ZN(n544) );
  INV_X1 U204 ( .A(A_ns[20]), .ZN(n543) );
  OAI221_X1 U205 ( .B1(n393), .B2(n546), .C1(n392), .C2(n547), .A(n548), .ZN(
        O[21]) );
  AOI22_X1 U206 ( .A1(A_ns[20]), .A2(n397), .B1(\A_s[20] ), .B2(n398), .ZN(
        n548) );
  INV_X1 U207 ( .A(\A_s[19] ), .ZN(n547) );
  INV_X1 U208 ( .A(A_ns[19]), .ZN(n546) );
  OAI221_X1 U209 ( .B1(n393), .B2(n549), .C1(n392), .C2(n550), .A(n551), .ZN(
        O[20]) );
  AOI22_X1 U210 ( .A1(A_ns[19]), .A2(n397), .B1(\A_s[19] ), .B2(n398), .ZN(
        n551) );
  INV_X1 U211 ( .A(\A_s[18] ), .ZN(n550) );
  INV_X1 U212 ( .A(A_ns[18]), .ZN(n549) );
  OAI22_X1 U213 ( .A1(n552), .A2(n520), .B1(n553), .B2(n519), .ZN(O[1]) );
  INV_X1 U214 ( .A(A_ns[0]), .ZN(n519) );
  INV_X1 U215 ( .A(\A_s[0] ), .ZN(n520) );
  OAI221_X1 U216 ( .B1(n393), .B2(n554), .C1(n392), .C2(n555), .A(n556), .ZN(
        O[19]) );
  AOI22_X1 U217 ( .A1(A_ns[18]), .A2(n397), .B1(\A_s[18] ), .B2(n398), .ZN(
        n556) );
  INV_X1 U218 ( .A(\A_s[17] ), .ZN(n555) );
  INV_X1 U219 ( .A(A_ns[17]), .ZN(n554) );
  OAI221_X1 U220 ( .B1(n393), .B2(n557), .C1(n392), .C2(n558), .A(n559), .ZN(
        O[18]) );
  AOI22_X1 U221 ( .A1(A_ns[17]), .A2(n397), .B1(\A_s[17] ), .B2(n398), .ZN(
        n559) );
  INV_X1 U222 ( .A(\A_s[16] ), .ZN(n558) );
  INV_X1 U223 ( .A(A_ns[16]), .ZN(n557) );
  OAI221_X1 U224 ( .B1(n393), .B2(n560), .C1(n392), .C2(n561), .A(n562), .ZN(
        O[17]) );
  AOI22_X1 U225 ( .A1(A_ns[16]), .A2(n397), .B1(\A_s[16] ), .B2(n398), .ZN(
        n562) );
  INV_X1 U226 ( .A(\A_s[15] ), .ZN(n561) );
  INV_X1 U227 ( .A(A_ns[15]), .ZN(n560) );
  OAI221_X1 U228 ( .B1(n393), .B2(n563), .C1(n392), .C2(n564), .A(n565), .ZN(
        O[16]) );
  AOI22_X1 U229 ( .A1(A_ns[15]), .A2(n397), .B1(\A_s[15] ), .B2(n398), .ZN(
        n565) );
  INV_X1 U230 ( .A(\A_s[14] ), .ZN(n564) );
  INV_X1 U231 ( .A(A_ns[14]), .ZN(n563) );
  OAI221_X1 U232 ( .B1(n393), .B2(n566), .C1(n392), .C2(n567), .A(n568), .ZN(
        O[15]) );
  AOI22_X1 U233 ( .A1(A_ns[14]), .A2(n397), .B1(\A_s[14] ), .B2(n398), .ZN(
        n568) );
  INV_X1 U234 ( .A(\A_s[13] ), .ZN(n567) );
  INV_X1 U235 ( .A(A_ns[13]), .ZN(n566) );
  OAI221_X1 U236 ( .B1(n393), .B2(n569), .C1(n392), .C2(n570), .A(n571), .ZN(
        O[14]) );
  AOI22_X1 U237 ( .A1(A_ns[13]), .A2(n397), .B1(\A_s[13] ), .B2(n398), .ZN(
        n571) );
  INV_X1 U238 ( .A(\A_s[12] ), .ZN(n570) );
  INV_X1 U239 ( .A(A_ns[12]), .ZN(n569) );
  OAI221_X1 U240 ( .B1(n393), .B2(n572), .C1(n392), .C2(n573), .A(n574), .ZN(
        O[13]) );
  AOI22_X1 U241 ( .A1(A_ns[12]), .A2(n397), .B1(\A_s[12] ), .B2(n398), .ZN(
        n574) );
  INV_X1 U242 ( .A(\A_s[11] ), .ZN(n573) );
  INV_X1 U243 ( .A(A_ns[11]), .ZN(n572) );
  OAI221_X1 U244 ( .B1(n393), .B2(n575), .C1(n392), .C2(n576), .A(n577), .ZN(
        O[12]) );
  AOI22_X1 U245 ( .A1(A_ns[11]), .A2(n397), .B1(\A_s[11] ), .B2(n398), .ZN(
        n577) );
  INV_X1 U246 ( .A(\A_s[10] ), .ZN(n576) );
  INV_X1 U247 ( .A(A_ns[10]), .ZN(n575) );
  OAI221_X1 U248 ( .B1(n393), .B2(n578), .C1(n392), .C2(n579), .A(n580), .ZN(
        O[11]) );
  AOI22_X1 U249 ( .A1(A_ns[10]), .A2(n397), .B1(\A_s[10] ), .B2(n398), .ZN(
        n580) );
  INV_X1 U250 ( .A(\A_s[9] ), .ZN(n579) );
  INV_X1 U251 ( .A(A_ns[9]), .ZN(n578) );
  OAI221_X1 U252 ( .B1(n581), .B2(n393), .C1(n582), .C2(n392), .A(n583), .ZN(
        O[10]) );
  AOI22_X1 U253 ( .A1(A_ns[9]), .A2(n397), .B1(\A_s[9] ), .B2(n398), .ZN(n583)
         );
  NAND2_X1 U254 ( .A1(n584), .A2(n552), .ZN(n553) );
  NAND2_X1 U255 ( .A1(n584), .A2(n585), .ZN(n552) );
  XOR2_X1 U256 ( .A(B[10]), .B(B[9]), .Z(n584) );
  INV_X1 U257 ( .A(\A_s[8] ), .ZN(n582) );
  INV_X1 U258 ( .A(B[11]), .ZN(n585) );
  INV_X1 U259 ( .A(A_ns[8]), .ZN(n581) );
endmodule


module BOOTHENC_NBIT64_i12 ( A, A_n, A_ns, A_s, B, O, A_so, A_nso );
  input [63:0] A;
  input [63:0] A_n;
  input [63:0] A_ns;
  input [63:0] A_s;
  input [63:0] B;
  output [63:0] O;
  output [63:0] A_so;
  output [63:0] A_nso;
  wire   \A_s[61] , \A_s[60] , \A_s[59] , \A_s[58] , \A_s[57] , \A_s[56] ,
         \A_s[55] , \A_s[54] , \A_s[53] , \A_s[52] , \A_s[51] , \A_s[50] ,
         \A_s[49] , \A_s[48] , \A_s[47] , \A_s[46] , \A_s[45] , \A_s[44] ,
         \A_s[43] , \A_s[42] , \A_s[41] , \A_s[40] , \A_s[39] , \A_s[38] ,
         \A_s[37] , \A_s[36] , \A_s[35] , \A_s[34] , \A_s[33] , \A_s[32] ,
         \A_s[31] , \A_s[30] , \A_s[29] , \A_s[28] , \A_s[27] , \A_s[26] ,
         \A_s[25] , \A_s[24] , \A_s[23] , \A_s[22] , \A_s[21] , \A_s[20] ,
         \A_s[19] , \A_s[18] , \A_s[17] , \A_s[16] , \A_s[15] , \A_s[14] ,
         \A_s[13] , \A_s[12] , \A_s[11] , \A_s[10] , \A_s[9] , \A_s[8] ,
         \A_s[7] , \A_s[6] , \A_s[5] , \A_s[4] , \A_s[3] , \A_s[2] , \A_s[1] ,
         \A_s[0] , n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585;
  assign A_nso[0] = 1'b0;
  assign A_nso[1] = 1'b0;
  assign A_so[0] = 1'b0;
  assign A_so[1] = 1'b0;
  assign O[0] = 1'b0;
  assign A_nso[63] = \A_s[61] ;
  assign A_so[63] = \A_s[61] ;
  assign \A_s[61]  = A_s[61];
  assign A_nso[62] = \A_s[60] ;
  assign A_so[62] = \A_s[60] ;
  assign \A_s[60]  = A_s[60];
  assign A_nso[61] = \A_s[59] ;
  assign A_so[61] = \A_s[59] ;
  assign \A_s[59]  = A_s[59];
  assign A_nso[60] = \A_s[58] ;
  assign A_so[60] = \A_s[58] ;
  assign \A_s[58]  = A_s[58];
  assign A_nso[59] = \A_s[57] ;
  assign A_so[59] = \A_s[57] ;
  assign \A_s[57]  = A_s[57];
  assign A_nso[58] = \A_s[56] ;
  assign A_so[58] = \A_s[56] ;
  assign \A_s[56]  = A_s[56];
  assign A_nso[57] = \A_s[55] ;
  assign A_so[57] = \A_s[55] ;
  assign \A_s[55]  = A_s[55];
  assign A_nso[56] = \A_s[54] ;
  assign A_so[56] = \A_s[54] ;
  assign \A_s[54]  = A_s[54];
  assign A_nso[55] = \A_s[53] ;
  assign A_so[55] = \A_s[53] ;
  assign \A_s[53]  = A_s[53];
  assign A_nso[54] = \A_s[52] ;
  assign A_so[54] = \A_s[52] ;
  assign \A_s[52]  = A_s[52];
  assign A_nso[53] = \A_s[51] ;
  assign A_so[53] = \A_s[51] ;
  assign \A_s[51]  = A_s[51];
  assign A_nso[52] = \A_s[50] ;
  assign A_so[52] = \A_s[50] ;
  assign \A_s[50]  = A_s[50];
  assign A_nso[51] = \A_s[49] ;
  assign A_so[51] = \A_s[49] ;
  assign \A_s[49]  = A_s[49];
  assign A_nso[50] = \A_s[48] ;
  assign A_so[50] = \A_s[48] ;
  assign \A_s[48]  = A_s[48];
  assign A_nso[49] = \A_s[47] ;
  assign A_so[49] = \A_s[47] ;
  assign \A_s[47]  = A_s[47];
  assign A_nso[48] = \A_s[46] ;
  assign A_so[48] = \A_s[46] ;
  assign \A_s[46]  = A_s[46];
  assign A_nso[47] = \A_s[45] ;
  assign A_so[47] = \A_s[45] ;
  assign \A_s[45]  = A_s[45];
  assign A_nso[46] = \A_s[44] ;
  assign A_so[46] = \A_s[44] ;
  assign \A_s[44]  = A_s[44];
  assign A_nso[45] = \A_s[43] ;
  assign A_so[45] = \A_s[43] ;
  assign \A_s[43]  = A_s[43];
  assign A_nso[44] = \A_s[42] ;
  assign A_so[44] = \A_s[42] ;
  assign \A_s[42]  = A_s[42];
  assign A_nso[43] = \A_s[41] ;
  assign A_so[43] = \A_s[41] ;
  assign \A_s[41]  = A_s[41];
  assign A_nso[42] = \A_s[40] ;
  assign A_so[42] = \A_s[40] ;
  assign \A_s[40]  = A_s[40];
  assign A_nso[41] = \A_s[39] ;
  assign A_so[41] = \A_s[39] ;
  assign \A_s[39]  = A_s[39];
  assign A_nso[40] = \A_s[38] ;
  assign A_so[40] = \A_s[38] ;
  assign \A_s[38]  = A_s[38];
  assign A_nso[39] = \A_s[37] ;
  assign A_so[39] = \A_s[37] ;
  assign \A_s[37]  = A_s[37];
  assign A_nso[38] = \A_s[36] ;
  assign A_so[38] = \A_s[36] ;
  assign \A_s[36]  = A_s[36];
  assign A_nso[37] = \A_s[35] ;
  assign A_so[37] = \A_s[35] ;
  assign \A_s[35]  = A_s[35];
  assign A_nso[36] = \A_s[34] ;
  assign A_so[36] = \A_s[34] ;
  assign \A_s[34]  = A_s[34];
  assign A_nso[35] = \A_s[33] ;
  assign A_so[35] = \A_s[33] ;
  assign \A_s[33]  = A_s[33];
  assign A_nso[34] = \A_s[32] ;
  assign A_so[34] = \A_s[32] ;
  assign \A_s[32]  = A_s[32];
  assign A_nso[33] = \A_s[31] ;
  assign A_so[33] = \A_s[31] ;
  assign \A_s[31]  = A_s[31];
  assign A_nso[32] = \A_s[30] ;
  assign A_so[32] = \A_s[30] ;
  assign \A_s[30]  = A_s[30];
  assign A_nso[31] = \A_s[29] ;
  assign A_so[31] = \A_s[29] ;
  assign \A_s[29]  = A_s[29];
  assign A_nso[30] = \A_s[28] ;
  assign A_so[30] = \A_s[28] ;
  assign \A_s[28]  = A_s[28];
  assign A_nso[29] = \A_s[27] ;
  assign A_so[29] = \A_s[27] ;
  assign \A_s[27]  = A_s[27];
  assign A_nso[28] = \A_s[26] ;
  assign A_so[28] = \A_s[26] ;
  assign \A_s[26]  = A_s[26];
  assign A_nso[27] = \A_s[25] ;
  assign A_so[27] = \A_s[25] ;
  assign \A_s[25]  = A_s[25];
  assign A_nso[26] = \A_s[24] ;
  assign A_so[26] = \A_s[24] ;
  assign \A_s[24]  = A_s[24];
  assign A_nso[25] = \A_s[23] ;
  assign A_so[25] = \A_s[23] ;
  assign \A_s[23]  = A_s[23];
  assign A_nso[24] = \A_s[22] ;
  assign A_so[24] = \A_s[22] ;
  assign \A_s[22]  = A_s[22];
  assign A_nso[23] = \A_s[21] ;
  assign A_so[23] = \A_s[21] ;
  assign \A_s[21]  = A_s[21];
  assign A_nso[22] = \A_s[20] ;
  assign A_so[22] = \A_s[20] ;
  assign \A_s[20]  = A_s[20];
  assign A_nso[21] = \A_s[19] ;
  assign A_so[21] = \A_s[19] ;
  assign \A_s[19]  = A_s[19];
  assign A_nso[20] = \A_s[18] ;
  assign A_so[20] = \A_s[18] ;
  assign \A_s[18]  = A_s[18];
  assign A_nso[19] = \A_s[17] ;
  assign A_so[19] = \A_s[17] ;
  assign \A_s[17]  = A_s[17];
  assign A_nso[18] = \A_s[16] ;
  assign A_so[18] = \A_s[16] ;
  assign \A_s[16]  = A_s[16];
  assign A_nso[17] = \A_s[15] ;
  assign A_so[17] = \A_s[15] ;
  assign \A_s[15]  = A_s[15];
  assign A_nso[16] = \A_s[14] ;
  assign A_so[16] = \A_s[14] ;
  assign \A_s[14]  = A_s[14];
  assign A_nso[15] = \A_s[13] ;
  assign A_so[15] = \A_s[13] ;
  assign \A_s[13]  = A_s[13];
  assign A_nso[14] = \A_s[12] ;
  assign A_so[14] = \A_s[12] ;
  assign \A_s[12]  = A_s[12];
  assign A_nso[13] = \A_s[11] ;
  assign A_so[13] = \A_s[11] ;
  assign \A_s[11]  = A_s[11];
  assign A_nso[12] = \A_s[10] ;
  assign A_so[12] = \A_s[10] ;
  assign \A_s[10]  = A_s[10];
  assign A_nso[11] = \A_s[9] ;
  assign A_so[11] = \A_s[9] ;
  assign \A_s[9]  = A_s[9];
  assign A_nso[10] = \A_s[8] ;
  assign A_so[10] = \A_s[8] ;
  assign \A_s[8]  = A_s[8];
  assign A_nso[9] = \A_s[7] ;
  assign A_so[9] = \A_s[7] ;
  assign \A_s[7]  = A_s[7];
  assign A_nso[8] = \A_s[6] ;
  assign A_so[8] = \A_s[6] ;
  assign \A_s[6]  = A_s[6];
  assign A_nso[7] = \A_s[5] ;
  assign A_so[7] = \A_s[5] ;
  assign \A_s[5]  = A_s[5];
  assign A_nso[6] = \A_s[4] ;
  assign A_so[6] = \A_s[4] ;
  assign \A_s[4]  = A_s[4];
  assign A_nso[5] = \A_s[3] ;
  assign A_so[5] = \A_s[3] ;
  assign \A_s[3]  = A_s[3];
  assign A_nso[4] = \A_s[2] ;
  assign A_so[4] = \A_s[2] ;
  assign \A_s[2]  = A_s[2];
  assign A_nso[3] = \A_s[1] ;
  assign A_so[3] = \A_s[1] ;
  assign \A_s[1]  = A_s[1];
  assign A_nso[2] = \A_s[0] ;
  assign A_so[2] = \A_s[0] ;
  assign \A_s[0]  = A_s[0];

  AND3_X1 U2 ( .A1(B[12]), .A2(n585), .A3(B[11]), .ZN(n391) );
  INV_X4 U3 ( .A(n391), .ZN(n392) );
  INV_X4 U4 ( .A(n552), .ZN(n398) );
  OR3_X4 U5 ( .A1(B[11]), .A2(B[12]), .A3(n585), .ZN(n393) );
  INV_X4 U6 ( .A(n553), .ZN(n397) );
  OAI221_X1 U7 ( .B1(n393), .B2(n394), .C1(n392), .C2(n395), .A(n396), .ZN(
        O[9]) );
  AOI22_X1 U8 ( .A1(A_ns[8]), .A2(n397), .B1(\A_s[8] ), .B2(n398), .ZN(n396)
         );
  INV_X1 U9 ( .A(\A_s[7] ), .ZN(n395) );
  INV_X1 U10 ( .A(A_ns[7]), .ZN(n394) );
  OAI221_X1 U11 ( .B1(n393), .B2(n399), .C1(n392), .C2(n400), .A(n401), .ZN(
        O[8]) );
  AOI22_X1 U12 ( .A1(A_ns[7]), .A2(n397), .B1(\A_s[7] ), .B2(n398), .ZN(n401)
         );
  INV_X1 U13 ( .A(\A_s[6] ), .ZN(n400) );
  INV_X1 U14 ( .A(A_ns[6]), .ZN(n399) );
  OAI221_X1 U15 ( .B1(n393), .B2(n402), .C1(n392), .C2(n403), .A(n404), .ZN(
        O[7]) );
  AOI22_X1 U16 ( .A1(A_ns[6]), .A2(n397), .B1(\A_s[6] ), .B2(n398), .ZN(n404)
         );
  INV_X1 U17 ( .A(\A_s[5] ), .ZN(n403) );
  INV_X1 U18 ( .A(A_ns[5]), .ZN(n402) );
  OAI221_X1 U19 ( .B1(n393), .B2(n405), .C1(n392), .C2(n406), .A(n407), .ZN(
        O[6]) );
  AOI22_X1 U20 ( .A1(A_ns[5]), .A2(n397), .B1(\A_s[5] ), .B2(n398), .ZN(n407)
         );
  INV_X1 U21 ( .A(\A_s[4] ), .ZN(n406) );
  INV_X1 U22 ( .A(A_ns[4]), .ZN(n405) );
  OAI221_X1 U23 ( .B1(n393), .B2(n408), .C1(n392), .C2(n409), .A(n410), .ZN(
        O[63]) );
  AOI22_X1 U24 ( .A1(A_ns[62]), .A2(n397), .B1(A_s[62]), .B2(n398), .ZN(n410)
         );
  INV_X1 U25 ( .A(\A_s[61] ), .ZN(n409) );
  INV_X1 U26 ( .A(A_ns[61]), .ZN(n408) );
  OAI221_X1 U27 ( .B1(n393), .B2(n411), .C1(n392), .C2(n412), .A(n413), .ZN(
        O[62]) );
  AOI22_X1 U28 ( .A1(A_ns[61]), .A2(n397), .B1(\A_s[61] ), .B2(n398), .ZN(n413) );
  INV_X1 U29 ( .A(\A_s[60] ), .ZN(n412) );
  INV_X1 U30 ( .A(A_ns[60]), .ZN(n411) );
  OAI221_X1 U31 ( .B1(n393), .B2(n414), .C1(n392), .C2(n415), .A(n416), .ZN(
        O[61]) );
  AOI22_X1 U32 ( .A1(A_ns[60]), .A2(n397), .B1(\A_s[60] ), .B2(n398), .ZN(n416) );
  INV_X1 U33 ( .A(\A_s[59] ), .ZN(n415) );
  INV_X1 U34 ( .A(A_ns[59]), .ZN(n414) );
  OAI221_X1 U35 ( .B1(n393), .B2(n417), .C1(n392), .C2(n418), .A(n419), .ZN(
        O[60]) );
  AOI22_X1 U36 ( .A1(A_ns[59]), .A2(n397), .B1(\A_s[59] ), .B2(n398), .ZN(n419) );
  INV_X1 U37 ( .A(\A_s[58] ), .ZN(n418) );
  INV_X1 U38 ( .A(A_ns[58]), .ZN(n417) );
  OAI221_X1 U39 ( .B1(n393), .B2(n420), .C1(n392), .C2(n421), .A(n422), .ZN(
        O[5]) );
  AOI22_X1 U40 ( .A1(A_ns[4]), .A2(n397), .B1(\A_s[4] ), .B2(n398), .ZN(n422)
         );
  INV_X1 U41 ( .A(\A_s[3] ), .ZN(n421) );
  INV_X1 U42 ( .A(A_ns[3]), .ZN(n420) );
  OAI221_X1 U43 ( .B1(n393), .B2(n423), .C1(n392), .C2(n424), .A(n425), .ZN(
        O[59]) );
  AOI22_X1 U44 ( .A1(A_ns[58]), .A2(n397), .B1(\A_s[58] ), .B2(n398), .ZN(n425) );
  INV_X1 U45 ( .A(\A_s[57] ), .ZN(n424) );
  INV_X1 U46 ( .A(A_ns[57]), .ZN(n423) );
  OAI221_X1 U47 ( .B1(n393), .B2(n426), .C1(n392), .C2(n427), .A(n428), .ZN(
        O[58]) );
  AOI22_X1 U48 ( .A1(A_ns[57]), .A2(n397), .B1(\A_s[57] ), .B2(n398), .ZN(n428) );
  INV_X1 U49 ( .A(\A_s[56] ), .ZN(n427) );
  INV_X1 U50 ( .A(A_ns[56]), .ZN(n426) );
  OAI221_X1 U51 ( .B1(n393), .B2(n429), .C1(n392), .C2(n430), .A(n431), .ZN(
        O[57]) );
  AOI22_X1 U52 ( .A1(A_ns[56]), .A2(n397), .B1(\A_s[56] ), .B2(n398), .ZN(n431) );
  INV_X1 U53 ( .A(\A_s[55] ), .ZN(n430) );
  INV_X1 U54 ( .A(A_ns[55]), .ZN(n429) );
  OAI221_X1 U55 ( .B1(n393), .B2(n432), .C1(n392), .C2(n433), .A(n434), .ZN(
        O[56]) );
  AOI22_X1 U56 ( .A1(A_ns[55]), .A2(n397), .B1(\A_s[55] ), .B2(n398), .ZN(n434) );
  INV_X1 U57 ( .A(\A_s[54] ), .ZN(n433) );
  INV_X1 U58 ( .A(A_ns[54]), .ZN(n432) );
  OAI221_X1 U59 ( .B1(n393), .B2(n435), .C1(n392), .C2(n436), .A(n437), .ZN(
        O[55]) );
  AOI22_X1 U60 ( .A1(A_ns[54]), .A2(n397), .B1(\A_s[54] ), .B2(n398), .ZN(n437) );
  INV_X1 U61 ( .A(\A_s[53] ), .ZN(n436) );
  INV_X1 U62 ( .A(A_ns[53]), .ZN(n435) );
  OAI221_X1 U63 ( .B1(n393), .B2(n438), .C1(n392), .C2(n439), .A(n440), .ZN(
        O[54]) );
  AOI22_X1 U64 ( .A1(A_ns[53]), .A2(n397), .B1(\A_s[53] ), .B2(n398), .ZN(n440) );
  INV_X1 U65 ( .A(\A_s[52] ), .ZN(n439) );
  INV_X1 U66 ( .A(A_ns[52]), .ZN(n438) );
  OAI221_X1 U67 ( .B1(n393), .B2(n441), .C1(n392), .C2(n442), .A(n443), .ZN(
        O[53]) );
  AOI22_X1 U68 ( .A1(A_ns[52]), .A2(n397), .B1(\A_s[52] ), .B2(n398), .ZN(n443) );
  INV_X1 U69 ( .A(\A_s[51] ), .ZN(n442) );
  INV_X1 U70 ( .A(A_ns[51]), .ZN(n441) );
  OAI221_X1 U71 ( .B1(n393), .B2(n444), .C1(n392), .C2(n445), .A(n446), .ZN(
        O[52]) );
  AOI22_X1 U72 ( .A1(A_ns[51]), .A2(n397), .B1(\A_s[51] ), .B2(n398), .ZN(n446) );
  INV_X1 U73 ( .A(\A_s[50] ), .ZN(n445) );
  INV_X1 U74 ( .A(A_ns[50]), .ZN(n444) );
  OAI221_X1 U75 ( .B1(n393), .B2(n447), .C1(n392), .C2(n448), .A(n449), .ZN(
        O[51]) );
  AOI22_X1 U76 ( .A1(A_ns[50]), .A2(n397), .B1(\A_s[50] ), .B2(n398), .ZN(n449) );
  INV_X1 U77 ( .A(\A_s[49] ), .ZN(n448) );
  INV_X1 U78 ( .A(A_ns[49]), .ZN(n447) );
  OAI221_X1 U79 ( .B1(n393), .B2(n450), .C1(n392), .C2(n451), .A(n452), .ZN(
        O[50]) );
  AOI22_X1 U80 ( .A1(A_ns[49]), .A2(n397), .B1(\A_s[49] ), .B2(n398), .ZN(n452) );
  INV_X1 U81 ( .A(\A_s[48] ), .ZN(n451) );
  INV_X1 U82 ( .A(A_ns[48]), .ZN(n450) );
  OAI221_X1 U83 ( .B1(n393), .B2(n453), .C1(n392), .C2(n454), .A(n455), .ZN(
        O[4]) );
  AOI22_X1 U84 ( .A1(A_ns[3]), .A2(n397), .B1(\A_s[3] ), .B2(n398), .ZN(n455)
         );
  INV_X1 U85 ( .A(\A_s[2] ), .ZN(n454) );
  INV_X1 U86 ( .A(A_ns[2]), .ZN(n453) );
  OAI221_X1 U87 ( .B1(n393), .B2(n456), .C1(n392), .C2(n457), .A(n458), .ZN(
        O[49]) );
  AOI22_X1 U88 ( .A1(A_ns[48]), .A2(n397), .B1(\A_s[48] ), .B2(n398), .ZN(n458) );
  INV_X1 U89 ( .A(\A_s[47] ), .ZN(n457) );
  INV_X1 U90 ( .A(A_ns[47]), .ZN(n456) );
  OAI221_X1 U91 ( .B1(n393), .B2(n459), .C1(n392), .C2(n460), .A(n461), .ZN(
        O[48]) );
  AOI22_X1 U92 ( .A1(A_ns[47]), .A2(n397), .B1(\A_s[47] ), .B2(n398), .ZN(n461) );
  INV_X1 U93 ( .A(\A_s[46] ), .ZN(n460) );
  INV_X1 U94 ( .A(A_ns[46]), .ZN(n459) );
  OAI221_X1 U95 ( .B1(n393), .B2(n462), .C1(n392), .C2(n463), .A(n464), .ZN(
        O[47]) );
  AOI22_X1 U96 ( .A1(A_ns[46]), .A2(n397), .B1(\A_s[46] ), .B2(n398), .ZN(n464) );
  INV_X1 U97 ( .A(\A_s[45] ), .ZN(n463) );
  INV_X1 U98 ( .A(A_ns[45]), .ZN(n462) );
  OAI221_X1 U99 ( .B1(n393), .B2(n465), .C1(n392), .C2(n466), .A(n467), .ZN(
        O[46]) );
  AOI22_X1 U100 ( .A1(A_ns[45]), .A2(n397), .B1(\A_s[45] ), .B2(n398), .ZN(
        n467) );
  INV_X1 U101 ( .A(\A_s[44] ), .ZN(n466) );
  INV_X1 U102 ( .A(A_ns[44]), .ZN(n465) );
  OAI221_X1 U103 ( .B1(n393), .B2(n468), .C1(n392), .C2(n469), .A(n470), .ZN(
        O[45]) );
  AOI22_X1 U104 ( .A1(A_ns[44]), .A2(n397), .B1(\A_s[44] ), .B2(n398), .ZN(
        n470) );
  INV_X1 U105 ( .A(\A_s[43] ), .ZN(n469) );
  INV_X1 U106 ( .A(A_ns[43]), .ZN(n468) );
  OAI221_X1 U107 ( .B1(n393), .B2(n471), .C1(n392), .C2(n472), .A(n473), .ZN(
        O[44]) );
  AOI22_X1 U108 ( .A1(A_ns[43]), .A2(n397), .B1(\A_s[43] ), .B2(n398), .ZN(
        n473) );
  INV_X1 U109 ( .A(\A_s[42] ), .ZN(n472) );
  INV_X1 U110 ( .A(A_ns[42]), .ZN(n471) );
  OAI221_X1 U111 ( .B1(n393), .B2(n474), .C1(n392), .C2(n475), .A(n476), .ZN(
        O[43]) );
  AOI22_X1 U112 ( .A1(A_ns[42]), .A2(n397), .B1(\A_s[42] ), .B2(n398), .ZN(
        n476) );
  INV_X1 U113 ( .A(\A_s[41] ), .ZN(n475) );
  INV_X1 U114 ( .A(A_ns[41]), .ZN(n474) );
  OAI221_X1 U115 ( .B1(n393), .B2(n477), .C1(n392), .C2(n478), .A(n479), .ZN(
        O[42]) );
  AOI22_X1 U116 ( .A1(A_ns[41]), .A2(n397), .B1(\A_s[41] ), .B2(n398), .ZN(
        n479) );
  INV_X1 U117 ( .A(\A_s[40] ), .ZN(n478) );
  INV_X1 U118 ( .A(A_ns[40]), .ZN(n477) );
  OAI221_X1 U119 ( .B1(n393), .B2(n480), .C1(n392), .C2(n481), .A(n482), .ZN(
        O[41]) );
  AOI22_X1 U120 ( .A1(A_ns[40]), .A2(n397), .B1(\A_s[40] ), .B2(n398), .ZN(
        n482) );
  INV_X1 U121 ( .A(\A_s[39] ), .ZN(n481) );
  INV_X1 U122 ( .A(A_ns[39]), .ZN(n480) );
  OAI221_X1 U123 ( .B1(n393), .B2(n483), .C1(n392), .C2(n484), .A(n485), .ZN(
        O[40]) );
  AOI22_X1 U124 ( .A1(A_ns[39]), .A2(n397), .B1(\A_s[39] ), .B2(n398), .ZN(
        n485) );
  INV_X1 U125 ( .A(\A_s[38] ), .ZN(n484) );
  INV_X1 U126 ( .A(A_ns[38]), .ZN(n483) );
  OAI221_X1 U127 ( .B1(n393), .B2(n486), .C1(n392), .C2(n487), .A(n488), .ZN(
        O[3]) );
  AOI22_X1 U128 ( .A1(A_ns[2]), .A2(n397), .B1(\A_s[2] ), .B2(n398), .ZN(n488)
         );
  INV_X1 U129 ( .A(\A_s[1] ), .ZN(n487) );
  INV_X1 U130 ( .A(A_ns[1]), .ZN(n486) );
  OAI221_X1 U131 ( .B1(n393), .B2(n489), .C1(n392), .C2(n490), .A(n491), .ZN(
        O[39]) );
  AOI22_X1 U132 ( .A1(A_ns[38]), .A2(n397), .B1(\A_s[38] ), .B2(n398), .ZN(
        n491) );
  INV_X1 U133 ( .A(\A_s[37] ), .ZN(n490) );
  INV_X1 U134 ( .A(A_ns[37]), .ZN(n489) );
  OAI221_X1 U135 ( .B1(n393), .B2(n492), .C1(n392), .C2(n493), .A(n494), .ZN(
        O[38]) );
  AOI22_X1 U136 ( .A1(A_ns[37]), .A2(n397), .B1(\A_s[37] ), .B2(n398), .ZN(
        n494) );
  INV_X1 U137 ( .A(\A_s[36] ), .ZN(n493) );
  INV_X1 U138 ( .A(A_ns[36]), .ZN(n492) );
  OAI221_X1 U139 ( .B1(n393), .B2(n495), .C1(n392), .C2(n496), .A(n497), .ZN(
        O[37]) );
  AOI22_X1 U140 ( .A1(A_ns[36]), .A2(n397), .B1(\A_s[36] ), .B2(n398), .ZN(
        n497) );
  INV_X1 U141 ( .A(\A_s[35] ), .ZN(n496) );
  INV_X1 U142 ( .A(A_ns[35]), .ZN(n495) );
  OAI221_X1 U143 ( .B1(n393), .B2(n498), .C1(n392), .C2(n499), .A(n500), .ZN(
        O[36]) );
  AOI22_X1 U144 ( .A1(A_ns[35]), .A2(n397), .B1(\A_s[35] ), .B2(n398), .ZN(
        n500) );
  INV_X1 U145 ( .A(\A_s[34] ), .ZN(n499) );
  INV_X1 U146 ( .A(A_ns[34]), .ZN(n498) );
  OAI221_X1 U147 ( .B1(n393), .B2(n501), .C1(n392), .C2(n502), .A(n503), .ZN(
        O[35]) );
  AOI22_X1 U148 ( .A1(A_ns[34]), .A2(n397), .B1(\A_s[34] ), .B2(n398), .ZN(
        n503) );
  INV_X1 U149 ( .A(\A_s[33] ), .ZN(n502) );
  INV_X1 U150 ( .A(A_ns[33]), .ZN(n501) );
  OAI221_X1 U151 ( .B1(n393), .B2(n504), .C1(n392), .C2(n505), .A(n506), .ZN(
        O[34]) );
  AOI22_X1 U152 ( .A1(A_ns[33]), .A2(n397), .B1(\A_s[33] ), .B2(n398), .ZN(
        n506) );
  INV_X1 U153 ( .A(\A_s[32] ), .ZN(n505) );
  INV_X1 U154 ( .A(A_ns[32]), .ZN(n504) );
  OAI221_X1 U155 ( .B1(n393), .B2(n507), .C1(n392), .C2(n508), .A(n509), .ZN(
        O[33]) );
  AOI22_X1 U156 ( .A1(A_ns[32]), .A2(n397), .B1(\A_s[32] ), .B2(n398), .ZN(
        n509) );
  INV_X1 U157 ( .A(\A_s[31] ), .ZN(n508) );
  INV_X1 U158 ( .A(A_ns[31]), .ZN(n507) );
  OAI221_X1 U159 ( .B1(n393), .B2(n510), .C1(n392), .C2(n511), .A(n512), .ZN(
        O[32]) );
  AOI22_X1 U160 ( .A1(A_ns[31]), .A2(n397), .B1(\A_s[31] ), .B2(n398), .ZN(
        n512) );
  INV_X1 U161 ( .A(\A_s[30] ), .ZN(n511) );
  INV_X1 U162 ( .A(A_ns[30]), .ZN(n510) );
  OAI221_X1 U163 ( .B1(n393), .B2(n513), .C1(n392), .C2(n514), .A(n515), .ZN(
        O[31]) );
  AOI22_X1 U164 ( .A1(A_ns[30]), .A2(n397), .B1(\A_s[30] ), .B2(n398), .ZN(
        n515) );
  INV_X1 U165 ( .A(\A_s[29] ), .ZN(n514) );
  INV_X1 U166 ( .A(A_ns[29]), .ZN(n513) );
  OAI221_X1 U167 ( .B1(n393), .B2(n516), .C1(n392), .C2(n517), .A(n518), .ZN(
        O[30]) );
  AOI22_X1 U168 ( .A1(A_ns[29]), .A2(n397), .B1(\A_s[29] ), .B2(n398), .ZN(
        n518) );
  INV_X1 U169 ( .A(\A_s[28] ), .ZN(n517) );
  INV_X1 U170 ( .A(A_ns[28]), .ZN(n516) );
  OAI221_X1 U171 ( .B1(n393), .B2(n519), .C1(n392), .C2(n520), .A(n521), .ZN(
        O[2]) );
  AOI22_X1 U172 ( .A1(A_ns[1]), .A2(n397), .B1(\A_s[1] ), .B2(n398), .ZN(n521)
         );
  OAI221_X1 U173 ( .B1(n393), .B2(n522), .C1(n392), .C2(n523), .A(n524), .ZN(
        O[29]) );
  AOI22_X1 U174 ( .A1(A_ns[28]), .A2(n397), .B1(\A_s[28] ), .B2(n398), .ZN(
        n524) );
  INV_X1 U175 ( .A(\A_s[27] ), .ZN(n523) );
  INV_X1 U176 ( .A(A_ns[27]), .ZN(n522) );
  OAI221_X1 U177 ( .B1(n393), .B2(n525), .C1(n392), .C2(n526), .A(n527), .ZN(
        O[28]) );
  AOI22_X1 U178 ( .A1(A_ns[27]), .A2(n397), .B1(\A_s[27] ), .B2(n398), .ZN(
        n527) );
  INV_X1 U179 ( .A(\A_s[26] ), .ZN(n526) );
  INV_X1 U180 ( .A(A_ns[26]), .ZN(n525) );
  OAI221_X1 U181 ( .B1(n393), .B2(n528), .C1(n392), .C2(n529), .A(n530), .ZN(
        O[27]) );
  AOI22_X1 U182 ( .A1(A_ns[26]), .A2(n397), .B1(\A_s[26] ), .B2(n398), .ZN(
        n530) );
  INV_X1 U183 ( .A(\A_s[25] ), .ZN(n529) );
  INV_X1 U184 ( .A(A_ns[25]), .ZN(n528) );
  OAI221_X1 U185 ( .B1(n393), .B2(n531), .C1(n392), .C2(n532), .A(n533), .ZN(
        O[26]) );
  AOI22_X1 U186 ( .A1(A_ns[25]), .A2(n397), .B1(\A_s[25] ), .B2(n398), .ZN(
        n533) );
  INV_X1 U187 ( .A(\A_s[24] ), .ZN(n532) );
  INV_X1 U188 ( .A(A_ns[24]), .ZN(n531) );
  OAI221_X1 U189 ( .B1(n393), .B2(n534), .C1(n392), .C2(n535), .A(n536), .ZN(
        O[25]) );
  AOI22_X1 U190 ( .A1(A_ns[24]), .A2(n397), .B1(\A_s[24] ), .B2(n398), .ZN(
        n536) );
  INV_X1 U191 ( .A(\A_s[23] ), .ZN(n535) );
  INV_X1 U192 ( .A(A_ns[23]), .ZN(n534) );
  OAI221_X1 U193 ( .B1(n393), .B2(n537), .C1(n392), .C2(n538), .A(n539), .ZN(
        O[24]) );
  AOI22_X1 U194 ( .A1(A_ns[23]), .A2(n397), .B1(\A_s[23] ), .B2(n398), .ZN(
        n539) );
  INV_X1 U195 ( .A(\A_s[22] ), .ZN(n538) );
  INV_X1 U196 ( .A(A_ns[22]), .ZN(n537) );
  OAI221_X1 U197 ( .B1(n393), .B2(n540), .C1(n392), .C2(n541), .A(n542), .ZN(
        O[23]) );
  AOI22_X1 U198 ( .A1(A_ns[22]), .A2(n397), .B1(\A_s[22] ), .B2(n398), .ZN(
        n542) );
  INV_X1 U199 ( .A(\A_s[21] ), .ZN(n541) );
  INV_X1 U200 ( .A(A_ns[21]), .ZN(n540) );
  OAI221_X1 U201 ( .B1(n393), .B2(n543), .C1(n392), .C2(n544), .A(n545), .ZN(
        O[22]) );
  AOI22_X1 U202 ( .A1(A_ns[21]), .A2(n397), .B1(\A_s[21] ), .B2(n398), .ZN(
        n545) );
  INV_X1 U203 ( .A(\A_s[20] ), .ZN(n544) );
  INV_X1 U204 ( .A(A_ns[20]), .ZN(n543) );
  OAI221_X1 U205 ( .B1(n393), .B2(n546), .C1(n392), .C2(n547), .A(n548), .ZN(
        O[21]) );
  AOI22_X1 U206 ( .A1(A_ns[20]), .A2(n397), .B1(\A_s[20] ), .B2(n398), .ZN(
        n548) );
  INV_X1 U207 ( .A(\A_s[19] ), .ZN(n547) );
  INV_X1 U208 ( .A(A_ns[19]), .ZN(n546) );
  OAI221_X1 U209 ( .B1(n393), .B2(n549), .C1(n392), .C2(n550), .A(n551), .ZN(
        O[20]) );
  AOI22_X1 U210 ( .A1(A_ns[19]), .A2(n397), .B1(\A_s[19] ), .B2(n398), .ZN(
        n551) );
  INV_X1 U211 ( .A(\A_s[18] ), .ZN(n550) );
  INV_X1 U212 ( .A(A_ns[18]), .ZN(n549) );
  OAI22_X1 U213 ( .A1(n552), .A2(n520), .B1(n553), .B2(n519), .ZN(O[1]) );
  INV_X1 U214 ( .A(A_ns[0]), .ZN(n519) );
  INV_X1 U215 ( .A(\A_s[0] ), .ZN(n520) );
  OAI221_X1 U216 ( .B1(n393), .B2(n554), .C1(n392), .C2(n555), .A(n556), .ZN(
        O[19]) );
  AOI22_X1 U217 ( .A1(A_ns[18]), .A2(n397), .B1(\A_s[18] ), .B2(n398), .ZN(
        n556) );
  INV_X1 U218 ( .A(\A_s[17] ), .ZN(n555) );
  INV_X1 U219 ( .A(A_ns[17]), .ZN(n554) );
  OAI221_X1 U220 ( .B1(n393), .B2(n557), .C1(n392), .C2(n558), .A(n559), .ZN(
        O[18]) );
  AOI22_X1 U221 ( .A1(A_ns[17]), .A2(n397), .B1(\A_s[17] ), .B2(n398), .ZN(
        n559) );
  INV_X1 U222 ( .A(\A_s[16] ), .ZN(n558) );
  INV_X1 U223 ( .A(A_ns[16]), .ZN(n557) );
  OAI221_X1 U224 ( .B1(n393), .B2(n560), .C1(n392), .C2(n561), .A(n562), .ZN(
        O[17]) );
  AOI22_X1 U225 ( .A1(A_ns[16]), .A2(n397), .B1(\A_s[16] ), .B2(n398), .ZN(
        n562) );
  INV_X1 U226 ( .A(\A_s[15] ), .ZN(n561) );
  INV_X1 U227 ( .A(A_ns[15]), .ZN(n560) );
  OAI221_X1 U228 ( .B1(n393), .B2(n563), .C1(n392), .C2(n564), .A(n565), .ZN(
        O[16]) );
  AOI22_X1 U229 ( .A1(A_ns[15]), .A2(n397), .B1(\A_s[15] ), .B2(n398), .ZN(
        n565) );
  INV_X1 U230 ( .A(\A_s[14] ), .ZN(n564) );
  INV_X1 U231 ( .A(A_ns[14]), .ZN(n563) );
  OAI221_X1 U232 ( .B1(n393), .B2(n566), .C1(n392), .C2(n567), .A(n568), .ZN(
        O[15]) );
  AOI22_X1 U233 ( .A1(A_ns[14]), .A2(n397), .B1(\A_s[14] ), .B2(n398), .ZN(
        n568) );
  INV_X1 U234 ( .A(\A_s[13] ), .ZN(n567) );
  INV_X1 U235 ( .A(A_ns[13]), .ZN(n566) );
  OAI221_X1 U236 ( .B1(n393), .B2(n569), .C1(n392), .C2(n570), .A(n571), .ZN(
        O[14]) );
  AOI22_X1 U237 ( .A1(A_ns[13]), .A2(n397), .B1(\A_s[13] ), .B2(n398), .ZN(
        n571) );
  INV_X1 U238 ( .A(\A_s[12] ), .ZN(n570) );
  INV_X1 U239 ( .A(A_ns[12]), .ZN(n569) );
  OAI221_X1 U240 ( .B1(n393), .B2(n572), .C1(n392), .C2(n573), .A(n574), .ZN(
        O[13]) );
  AOI22_X1 U241 ( .A1(A_ns[12]), .A2(n397), .B1(\A_s[12] ), .B2(n398), .ZN(
        n574) );
  INV_X1 U242 ( .A(\A_s[11] ), .ZN(n573) );
  INV_X1 U243 ( .A(A_ns[11]), .ZN(n572) );
  OAI221_X1 U244 ( .B1(n393), .B2(n575), .C1(n392), .C2(n576), .A(n577), .ZN(
        O[12]) );
  AOI22_X1 U245 ( .A1(A_ns[11]), .A2(n397), .B1(\A_s[11] ), .B2(n398), .ZN(
        n577) );
  INV_X1 U246 ( .A(\A_s[10] ), .ZN(n576) );
  INV_X1 U247 ( .A(A_ns[10]), .ZN(n575) );
  OAI221_X1 U248 ( .B1(n393), .B2(n578), .C1(n392), .C2(n579), .A(n580), .ZN(
        O[11]) );
  AOI22_X1 U249 ( .A1(A_ns[10]), .A2(n397), .B1(\A_s[10] ), .B2(n398), .ZN(
        n580) );
  INV_X1 U250 ( .A(\A_s[9] ), .ZN(n579) );
  INV_X1 U251 ( .A(A_ns[9]), .ZN(n578) );
  OAI221_X1 U252 ( .B1(n581), .B2(n393), .C1(n582), .C2(n392), .A(n583), .ZN(
        O[10]) );
  AOI22_X1 U253 ( .A1(A_ns[9]), .A2(n397), .B1(\A_s[9] ), .B2(n398), .ZN(n583)
         );
  NAND2_X1 U254 ( .A1(n584), .A2(n552), .ZN(n553) );
  NAND2_X1 U255 ( .A1(n584), .A2(n585), .ZN(n552) );
  XOR2_X1 U256 ( .A(B[11]), .B(B[12]), .Z(n584) );
  INV_X1 U257 ( .A(\A_s[8] ), .ZN(n582) );
  INV_X1 U258 ( .A(B[13]), .ZN(n585) );
  INV_X1 U259 ( .A(A_ns[8]), .ZN(n581) );
endmodule


module BOOTHENC_NBIT64_i14 ( A, A_n, A_ns, A_s, B, O, A_so, A_nso );
  input [63:0] A;
  input [63:0] A_n;
  input [63:0] A_ns;
  input [63:0] A_s;
  input [63:0] B;
  output [63:0] O;
  output [63:0] A_so;
  output [63:0] A_nso;
  wire   \A_s[61] , \A_s[60] , \A_s[59] , \A_s[58] , \A_s[57] , \A_s[56] ,
         \A_s[55] , \A_s[54] , \A_s[53] , \A_s[52] , \A_s[51] , \A_s[50] ,
         \A_s[49] , \A_s[48] , \A_s[47] , \A_s[46] , \A_s[45] , \A_s[44] ,
         \A_s[43] , \A_s[42] , \A_s[41] , \A_s[40] , \A_s[39] , \A_s[38] ,
         \A_s[37] , \A_s[36] , \A_s[35] , \A_s[34] , \A_s[33] , \A_s[32] ,
         \A_s[31] , \A_s[30] , \A_s[29] , \A_s[28] , \A_s[27] , \A_s[26] ,
         \A_s[25] , \A_s[24] , \A_s[23] , \A_s[22] , \A_s[21] , \A_s[20] ,
         \A_s[19] , \A_s[18] , \A_s[17] , \A_s[16] , \A_s[15] , \A_s[14] ,
         \A_s[13] , \A_s[12] , \A_s[11] , \A_s[10] , \A_s[9] , \A_s[8] ,
         \A_s[7] , \A_s[6] , \A_s[5] , \A_s[4] , \A_s[3] , \A_s[2] , \A_s[1] ,
         \A_s[0] , n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585;
  assign A_nso[0] = 1'b0;
  assign A_nso[1] = 1'b0;
  assign A_so[0] = 1'b0;
  assign A_so[1] = 1'b0;
  assign O[0] = 1'b0;
  assign A_nso[63] = \A_s[61] ;
  assign A_so[63] = \A_s[61] ;
  assign \A_s[61]  = A_s[61];
  assign A_nso[62] = \A_s[60] ;
  assign A_so[62] = \A_s[60] ;
  assign \A_s[60]  = A_s[60];
  assign A_nso[61] = \A_s[59] ;
  assign A_so[61] = \A_s[59] ;
  assign \A_s[59]  = A_s[59];
  assign A_nso[60] = \A_s[58] ;
  assign A_so[60] = \A_s[58] ;
  assign \A_s[58]  = A_s[58];
  assign A_nso[59] = \A_s[57] ;
  assign A_so[59] = \A_s[57] ;
  assign \A_s[57]  = A_s[57];
  assign A_nso[58] = \A_s[56] ;
  assign A_so[58] = \A_s[56] ;
  assign \A_s[56]  = A_s[56];
  assign A_nso[57] = \A_s[55] ;
  assign A_so[57] = \A_s[55] ;
  assign \A_s[55]  = A_s[55];
  assign A_nso[56] = \A_s[54] ;
  assign A_so[56] = \A_s[54] ;
  assign \A_s[54]  = A_s[54];
  assign A_nso[55] = \A_s[53] ;
  assign A_so[55] = \A_s[53] ;
  assign \A_s[53]  = A_s[53];
  assign A_nso[54] = \A_s[52] ;
  assign A_so[54] = \A_s[52] ;
  assign \A_s[52]  = A_s[52];
  assign A_nso[53] = \A_s[51] ;
  assign A_so[53] = \A_s[51] ;
  assign \A_s[51]  = A_s[51];
  assign A_nso[52] = \A_s[50] ;
  assign A_so[52] = \A_s[50] ;
  assign \A_s[50]  = A_s[50];
  assign A_nso[51] = \A_s[49] ;
  assign A_so[51] = \A_s[49] ;
  assign \A_s[49]  = A_s[49];
  assign A_nso[50] = \A_s[48] ;
  assign A_so[50] = \A_s[48] ;
  assign \A_s[48]  = A_s[48];
  assign A_nso[49] = \A_s[47] ;
  assign A_so[49] = \A_s[47] ;
  assign \A_s[47]  = A_s[47];
  assign A_nso[48] = \A_s[46] ;
  assign A_so[48] = \A_s[46] ;
  assign \A_s[46]  = A_s[46];
  assign A_nso[47] = \A_s[45] ;
  assign A_so[47] = \A_s[45] ;
  assign \A_s[45]  = A_s[45];
  assign A_nso[46] = \A_s[44] ;
  assign A_so[46] = \A_s[44] ;
  assign \A_s[44]  = A_s[44];
  assign A_nso[45] = \A_s[43] ;
  assign A_so[45] = \A_s[43] ;
  assign \A_s[43]  = A_s[43];
  assign A_nso[44] = \A_s[42] ;
  assign A_so[44] = \A_s[42] ;
  assign \A_s[42]  = A_s[42];
  assign A_nso[43] = \A_s[41] ;
  assign A_so[43] = \A_s[41] ;
  assign \A_s[41]  = A_s[41];
  assign A_nso[42] = \A_s[40] ;
  assign A_so[42] = \A_s[40] ;
  assign \A_s[40]  = A_s[40];
  assign A_nso[41] = \A_s[39] ;
  assign A_so[41] = \A_s[39] ;
  assign \A_s[39]  = A_s[39];
  assign A_nso[40] = \A_s[38] ;
  assign A_so[40] = \A_s[38] ;
  assign \A_s[38]  = A_s[38];
  assign A_nso[39] = \A_s[37] ;
  assign A_so[39] = \A_s[37] ;
  assign \A_s[37]  = A_s[37];
  assign A_nso[38] = \A_s[36] ;
  assign A_so[38] = \A_s[36] ;
  assign \A_s[36]  = A_s[36];
  assign A_nso[37] = \A_s[35] ;
  assign A_so[37] = \A_s[35] ;
  assign \A_s[35]  = A_s[35];
  assign A_nso[36] = \A_s[34] ;
  assign A_so[36] = \A_s[34] ;
  assign \A_s[34]  = A_s[34];
  assign A_nso[35] = \A_s[33] ;
  assign A_so[35] = \A_s[33] ;
  assign \A_s[33]  = A_s[33];
  assign A_nso[34] = \A_s[32] ;
  assign A_so[34] = \A_s[32] ;
  assign \A_s[32]  = A_s[32];
  assign A_nso[33] = \A_s[31] ;
  assign A_so[33] = \A_s[31] ;
  assign \A_s[31]  = A_s[31];
  assign A_nso[32] = \A_s[30] ;
  assign A_so[32] = \A_s[30] ;
  assign \A_s[30]  = A_s[30];
  assign A_nso[31] = \A_s[29] ;
  assign A_so[31] = \A_s[29] ;
  assign \A_s[29]  = A_s[29];
  assign A_nso[30] = \A_s[28] ;
  assign A_so[30] = \A_s[28] ;
  assign \A_s[28]  = A_s[28];
  assign A_nso[29] = \A_s[27] ;
  assign A_so[29] = \A_s[27] ;
  assign \A_s[27]  = A_s[27];
  assign A_nso[28] = \A_s[26] ;
  assign A_so[28] = \A_s[26] ;
  assign \A_s[26]  = A_s[26];
  assign A_nso[27] = \A_s[25] ;
  assign A_so[27] = \A_s[25] ;
  assign \A_s[25]  = A_s[25];
  assign A_nso[26] = \A_s[24] ;
  assign A_so[26] = \A_s[24] ;
  assign \A_s[24]  = A_s[24];
  assign A_nso[25] = \A_s[23] ;
  assign A_so[25] = \A_s[23] ;
  assign \A_s[23]  = A_s[23];
  assign A_nso[24] = \A_s[22] ;
  assign A_so[24] = \A_s[22] ;
  assign \A_s[22]  = A_s[22];
  assign A_nso[23] = \A_s[21] ;
  assign A_so[23] = \A_s[21] ;
  assign \A_s[21]  = A_s[21];
  assign A_nso[22] = \A_s[20] ;
  assign A_so[22] = \A_s[20] ;
  assign \A_s[20]  = A_s[20];
  assign A_nso[21] = \A_s[19] ;
  assign A_so[21] = \A_s[19] ;
  assign \A_s[19]  = A_s[19];
  assign A_nso[20] = \A_s[18] ;
  assign A_so[20] = \A_s[18] ;
  assign \A_s[18]  = A_s[18];
  assign A_nso[19] = \A_s[17] ;
  assign A_so[19] = \A_s[17] ;
  assign \A_s[17]  = A_s[17];
  assign A_nso[18] = \A_s[16] ;
  assign A_so[18] = \A_s[16] ;
  assign \A_s[16]  = A_s[16];
  assign A_nso[17] = \A_s[15] ;
  assign A_so[17] = \A_s[15] ;
  assign \A_s[15]  = A_s[15];
  assign A_nso[16] = \A_s[14] ;
  assign A_so[16] = \A_s[14] ;
  assign \A_s[14]  = A_s[14];
  assign A_nso[15] = \A_s[13] ;
  assign A_so[15] = \A_s[13] ;
  assign \A_s[13]  = A_s[13];
  assign A_nso[14] = \A_s[12] ;
  assign A_so[14] = \A_s[12] ;
  assign \A_s[12]  = A_s[12];
  assign A_nso[13] = \A_s[11] ;
  assign A_so[13] = \A_s[11] ;
  assign \A_s[11]  = A_s[11];
  assign A_nso[12] = \A_s[10] ;
  assign A_so[12] = \A_s[10] ;
  assign \A_s[10]  = A_s[10];
  assign A_nso[11] = \A_s[9] ;
  assign A_so[11] = \A_s[9] ;
  assign \A_s[9]  = A_s[9];
  assign A_nso[10] = \A_s[8] ;
  assign A_so[10] = \A_s[8] ;
  assign \A_s[8]  = A_s[8];
  assign A_nso[9] = \A_s[7] ;
  assign A_so[9] = \A_s[7] ;
  assign \A_s[7]  = A_s[7];
  assign A_nso[8] = \A_s[6] ;
  assign A_so[8] = \A_s[6] ;
  assign \A_s[6]  = A_s[6];
  assign A_nso[7] = \A_s[5] ;
  assign A_so[7] = \A_s[5] ;
  assign \A_s[5]  = A_s[5];
  assign A_nso[6] = \A_s[4] ;
  assign A_so[6] = \A_s[4] ;
  assign \A_s[4]  = A_s[4];
  assign A_nso[5] = \A_s[3] ;
  assign A_so[5] = \A_s[3] ;
  assign \A_s[3]  = A_s[3];
  assign A_nso[4] = \A_s[2] ;
  assign A_so[4] = \A_s[2] ;
  assign \A_s[2]  = A_s[2];
  assign A_nso[3] = \A_s[1] ;
  assign A_so[3] = \A_s[1] ;
  assign \A_s[1]  = A_s[1];
  assign A_nso[2] = \A_s[0] ;
  assign A_so[2] = \A_s[0] ;
  assign \A_s[0]  = A_s[0];

  AND3_X1 U2 ( .A1(B[14]), .A2(n585), .A3(B[13]), .ZN(n391) );
  INV_X4 U3 ( .A(n391), .ZN(n392) );
  INV_X4 U4 ( .A(n552), .ZN(n398) );
  OR3_X4 U5 ( .A1(B[13]), .A2(B[14]), .A3(n585), .ZN(n393) );
  INV_X4 U6 ( .A(n553), .ZN(n397) );
  OAI221_X1 U7 ( .B1(n393), .B2(n394), .C1(n392), .C2(n395), .A(n396), .ZN(
        O[9]) );
  AOI22_X1 U8 ( .A1(A_ns[8]), .A2(n397), .B1(\A_s[8] ), .B2(n398), .ZN(n396)
         );
  INV_X1 U9 ( .A(\A_s[7] ), .ZN(n395) );
  INV_X1 U10 ( .A(A_ns[7]), .ZN(n394) );
  OAI221_X1 U11 ( .B1(n393), .B2(n399), .C1(n392), .C2(n400), .A(n401), .ZN(
        O[8]) );
  AOI22_X1 U12 ( .A1(A_ns[7]), .A2(n397), .B1(\A_s[7] ), .B2(n398), .ZN(n401)
         );
  INV_X1 U13 ( .A(\A_s[6] ), .ZN(n400) );
  INV_X1 U14 ( .A(A_ns[6]), .ZN(n399) );
  OAI221_X1 U15 ( .B1(n393), .B2(n402), .C1(n392), .C2(n403), .A(n404), .ZN(
        O[7]) );
  AOI22_X1 U16 ( .A1(A_ns[6]), .A2(n397), .B1(\A_s[6] ), .B2(n398), .ZN(n404)
         );
  INV_X1 U17 ( .A(\A_s[5] ), .ZN(n403) );
  INV_X1 U18 ( .A(A_ns[5]), .ZN(n402) );
  OAI221_X1 U19 ( .B1(n393), .B2(n405), .C1(n392), .C2(n406), .A(n407), .ZN(
        O[6]) );
  AOI22_X1 U20 ( .A1(A_ns[5]), .A2(n397), .B1(\A_s[5] ), .B2(n398), .ZN(n407)
         );
  INV_X1 U21 ( .A(\A_s[4] ), .ZN(n406) );
  INV_X1 U22 ( .A(A_ns[4]), .ZN(n405) );
  OAI221_X1 U23 ( .B1(n393), .B2(n408), .C1(n392), .C2(n409), .A(n410), .ZN(
        O[63]) );
  AOI22_X1 U24 ( .A1(A_ns[62]), .A2(n397), .B1(A_s[62]), .B2(n398), .ZN(n410)
         );
  INV_X1 U25 ( .A(\A_s[61] ), .ZN(n409) );
  INV_X1 U26 ( .A(A_ns[61]), .ZN(n408) );
  OAI221_X1 U27 ( .B1(n393), .B2(n411), .C1(n392), .C2(n412), .A(n413), .ZN(
        O[62]) );
  AOI22_X1 U28 ( .A1(A_ns[61]), .A2(n397), .B1(\A_s[61] ), .B2(n398), .ZN(n413) );
  INV_X1 U29 ( .A(\A_s[60] ), .ZN(n412) );
  INV_X1 U30 ( .A(A_ns[60]), .ZN(n411) );
  OAI221_X1 U31 ( .B1(n393), .B2(n414), .C1(n392), .C2(n415), .A(n416), .ZN(
        O[61]) );
  AOI22_X1 U32 ( .A1(A_ns[60]), .A2(n397), .B1(\A_s[60] ), .B2(n398), .ZN(n416) );
  INV_X1 U33 ( .A(\A_s[59] ), .ZN(n415) );
  INV_X1 U34 ( .A(A_ns[59]), .ZN(n414) );
  OAI221_X1 U35 ( .B1(n393), .B2(n417), .C1(n392), .C2(n418), .A(n419), .ZN(
        O[60]) );
  AOI22_X1 U36 ( .A1(A_ns[59]), .A2(n397), .B1(\A_s[59] ), .B2(n398), .ZN(n419) );
  INV_X1 U37 ( .A(\A_s[58] ), .ZN(n418) );
  INV_X1 U38 ( .A(A_ns[58]), .ZN(n417) );
  OAI221_X1 U39 ( .B1(n393), .B2(n420), .C1(n392), .C2(n421), .A(n422), .ZN(
        O[5]) );
  AOI22_X1 U40 ( .A1(A_ns[4]), .A2(n397), .B1(\A_s[4] ), .B2(n398), .ZN(n422)
         );
  INV_X1 U41 ( .A(\A_s[3] ), .ZN(n421) );
  INV_X1 U42 ( .A(A_ns[3]), .ZN(n420) );
  OAI221_X1 U43 ( .B1(n393), .B2(n423), .C1(n392), .C2(n424), .A(n425), .ZN(
        O[59]) );
  AOI22_X1 U44 ( .A1(A_ns[58]), .A2(n397), .B1(\A_s[58] ), .B2(n398), .ZN(n425) );
  INV_X1 U45 ( .A(\A_s[57] ), .ZN(n424) );
  INV_X1 U46 ( .A(A_ns[57]), .ZN(n423) );
  OAI221_X1 U47 ( .B1(n393), .B2(n426), .C1(n392), .C2(n427), .A(n428), .ZN(
        O[58]) );
  AOI22_X1 U48 ( .A1(A_ns[57]), .A2(n397), .B1(\A_s[57] ), .B2(n398), .ZN(n428) );
  INV_X1 U49 ( .A(\A_s[56] ), .ZN(n427) );
  INV_X1 U50 ( .A(A_ns[56]), .ZN(n426) );
  OAI221_X1 U51 ( .B1(n393), .B2(n429), .C1(n392), .C2(n430), .A(n431), .ZN(
        O[57]) );
  AOI22_X1 U52 ( .A1(A_ns[56]), .A2(n397), .B1(\A_s[56] ), .B2(n398), .ZN(n431) );
  INV_X1 U53 ( .A(\A_s[55] ), .ZN(n430) );
  INV_X1 U54 ( .A(A_ns[55]), .ZN(n429) );
  OAI221_X1 U55 ( .B1(n393), .B2(n432), .C1(n392), .C2(n433), .A(n434), .ZN(
        O[56]) );
  AOI22_X1 U56 ( .A1(A_ns[55]), .A2(n397), .B1(\A_s[55] ), .B2(n398), .ZN(n434) );
  INV_X1 U57 ( .A(\A_s[54] ), .ZN(n433) );
  INV_X1 U58 ( .A(A_ns[54]), .ZN(n432) );
  OAI221_X1 U59 ( .B1(n393), .B2(n435), .C1(n392), .C2(n436), .A(n437), .ZN(
        O[55]) );
  AOI22_X1 U60 ( .A1(A_ns[54]), .A2(n397), .B1(\A_s[54] ), .B2(n398), .ZN(n437) );
  INV_X1 U61 ( .A(\A_s[53] ), .ZN(n436) );
  INV_X1 U62 ( .A(A_ns[53]), .ZN(n435) );
  OAI221_X1 U63 ( .B1(n393), .B2(n438), .C1(n392), .C2(n439), .A(n440), .ZN(
        O[54]) );
  AOI22_X1 U64 ( .A1(A_ns[53]), .A2(n397), .B1(\A_s[53] ), .B2(n398), .ZN(n440) );
  INV_X1 U65 ( .A(\A_s[52] ), .ZN(n439) );
  INV_X1 U66 ( .A(A_ns[52]), .ZN(n438) );
  OAI221_X1 U67 ( .B1(n393), .B2(n441), .C1(n392), .C2(n442), .A(n443), .ZN(
        O[53]) );
  AOI22_X1 U68 ( .A1(A_ns[52]), .A2(n397), .B1(\A_s[52] ), .B2(n398), .ZN(n443) );
  INV_X1 U69 ( .A(\A_s[51] ), .ZN(n442) );
  INV_X1 U70 ( .A(A_ns[51]), .ZN(n441) );
  OAI221_X1 U71 ( .B1(n393), .B2(n444), .C1(n392), .C2(n445), .A(n446), .ZN(
        O[52]) );
  AOI22_X1 U72 ( .A1(A_ns[51]), .A2(n397), .B1(\A_s[51] ), .B2(n398), .ZN(n446) );
  INV_X1 U73 ( .A(\A_s[50] ), .ZN(n445) );
  INV_X1 U74 ( .A(A_ns[50]), .ZN(n444) );
  OAI221_X1 U75 ( .B1(n393), .B2(n447), .C1(n392), .C2(n448), .A(n449), .ZN(
        O[51]) );
  AOI22_X1 U76 ( .A1(A_ns[50]), .A2(n397), .B1(\A_s[50] ), .B2(n398), .ZN(n449) );
  INV_X1 U77 ( .A(\A_s[49] ), .ZN(n448) );
  INV_X1 U78 ( .A(A_ns[49]), .ZN(n447) );
  OAI221_X1 U79 ( .B1(n393), .B2(n450), .C1(n392), .C2(n451), .A(n452), .ZN(
        O[50]) );
  AOI22_X1 U80 ( .A1(A_ns[49]), .A2(n397), .B1(\A_s[49] ), .B2(n398), .ZN(n452) );
  INV_X1 U81 ( .A(\A_s[48] ), .ZN(n451) );
  INV_X1 U82 ( .A(A_ns[48]), .ZN(n450) );
  OAI221_X1 U83 ( .B1(n393), .B2(n453), .C1(n392), .C2(n454), .A(n455), .ZN(
        O[4]) );
  AOI22_X1 U84 ( .A1(A_ns[3]), .A2(n397), .B1(\A_s[3] ), .B2(n398), .ZN(n455)
         );
  INV_X1 U85 ( .A(\A_s[2] ), .ZN(n454) );
  INV_X1 U86 ( .A(A_ns[2]), .ZN(n453) );
  OAI221_X1 U87 ( .B1(n393), .B2(n456), .C1(n392), .C2(n457), .A(n458), .ZN(
        O[49]) );
  AOI22_X1 U88 ( .A1(A_ns[48]), .A2(n397), .B1(\A_s[48] ), .B2(n398), .ZN(n458) );
  INV_X1 U89 ( .A(\A_s[47] ), .ZN(n457) );
  INV_X1 U90 ( .A(A_ns[47]), .ZN(n456) );
  OAI221_X1 U91 ( .B1(n393), .B2(n459), .C1(n392), .C2(n460), .A(n461), .ZN(
        O[48]) );
  AOI22_X1 U92 ( .A1(A_ns[47]), .A2(n397), .B1(\A_s[47] ), .B2(n398), .ZN(n461) );
  INV_X1 U93 ( .A(\A_s[46] ), .ZN(n460) );
  INV_X1 U94 ( .A(A_ns[46]), .ZN(n459) );
  OAI221_X1 U95 ( .B1(n393), .B2(n462), .C1(n392), .C2(n463), .A(n464), .ZN(
        O[47]) );
  AOI22_X1 U96 ( .A1(A_ns[46]), .A2(n397), .B1(\A_s[46] ), .B2(n398), .ZN(n464) );
  INV_X1 U97 ( .A(\A_s[45] ), .ZN(n463) );
  INV_X1 U98 ( .A(A_ns[45]), .ZN(n462) );
  OAI221_X1 U99 ( .B1(n393), .B2(n465), .C1(n392), .C2(n466), .A(n467), .ZN(
        O[46]) );
  AOI22_X1 U100 ( .A1(A_ns[45]), .A2(n397), .B1(\A_s[45] ), .B2(n398), .ZN(
        n467) );
  INV_X1 U101 ( .A(\A_s[44] ), .ZN(n466) );
  INV_X1 U102 ( .A(A_ns[44]), .ZN(n465) );
  OAI221_X1 U103 ( .B1(n393), .B2(n468), .C1(n392), .C2(n469), .A(n470), .ZN(
        O[45]) );
  AOI22_X1 U104 ( .A1(A_ns[44]), .A2(n397), .B1(\A_s[44] ), .B2(n398), .ZN(
        n470) );
  INV_X1 U105 ( .A(\A_s[43] ), .ZN(n469) );
  INV_X1 U106 ( .A(A_ns[43]), .ZN(n468) );
  OAI221_X1 U107 ( .B1(n393), .B2(n471), .C1(n392), .C2(n472), .A(n473), .ZN(
        O[44]) );
  AOI22_X1 U108 ( .A1(A_ns[43]), .A2(n397), .B1(\A_s[43] ), .B2(n398), .ZN(
        n473) );
  INV_X1 U109 ( .A(\A_s[42] ), .ZN(n472) );
  INV_X1 U110 ( .A(A_ns[42]), .ZN(n471) );
  OAI221_X1 U111 ( .B1(n393), .B2(n474), .C1(n392), .C2(n475), .A(n476), .ZN(
        O[43]) );
  AOI22_X1 U112 ( .A1(A_ns[42]), .A2(n397), .B1(\A_s[42] ), .B2(n398), .ZN(
        n476) );
  INV_X1 U113 ( .A(\A_s[41] ), .ZN(n475) );
  INV_X1 U114 ( .A(A_ns[41]), .ZN(n474) );
  OAI221_X1 U115 ( .B1(n393), .B2(n477), .C1(n392), .C2(n478), .A(n479), .ZN(
        O[42]) );
  AOI22_X1 U116 ( .A1(A_ns[41]), .A2(n397), .B1(\A_s[41] ), .B2(n398), .ZN(
        n479) );
  INV_X1 U117 ( .A(\A_s[40] ), .ZN(n478) );
  INV_X1 U118 ( .A(A_ns[40]), .ZN(n477) );
  OAI221_X1 U119 ( .B1(n393), .B2(n480), .C1(n392), .C2(n481), .A(n482), .ZN(
        O[41]) );
  AOI22_X1 U120 ( .A1(A_ns[40]), .A2(n397), .B1(\A_s[40] ), .B2(n398), .ZN(
        n482) );
  INV_X1 U121 ( .A(\A_s[39] ), .ZN(n481) );
  INV_X1 U122 ( .A(A_ns[39]), .ZN(n480) );
  OAI221_X1 U123 ( .B1(n393), .B2(n483), .C1(n392), .C2(n484), .A(n485), .ZN(
        O[40]) );
  AOI22_X1 U124 ( .A1(A_ns[39]), .A2(n397), .B1(\A_s[39] ), .B2(n398), .ZN(
        n485) );
  INV_X1 U125 ( .A(\A_s[38] ), .ZN(n484) );
  INV_X1 U126 ( .A(A_ns[38]), .ZN(n483) );
  OAI221_X1 U127 ( .B1(n393), .B2(n486), .C1(n392), .C2(n487), .A(n488), .ZN(
        O[3]) );
  AOI22_X1 U128 ( .A1(A_ns[2]), .A2(n397), .B1(\A_s[2] ), .B2(n398), .ZN(n488)
         );
  INV_X1 U129 ( .A(\A_s[1] ), .ZN(n487) );
  INV_X1 U130 ( .A(A_ns[1]), .ZN(n486) );
  OAI221_X1 U131 ( .B1(n393), .B2(n489), .C1(n392), .C2(n490), .A(n491), .ZN(
        O[39]) );
  AOI22_X1 U132 ( .A1(A_ns[38]), .A2(n397), .B1(\A_s[38] ), .B2(n398), .ZN(
        n491) );
  INV_X1 U133 ( .A(\A_s[37] ), .ZN(n490) );
  INV_X1 U134 ( .A(A_ns[37]), .ZN(n489) );
  OAI221_X1 U135 ( .B1(n393), .B2(n492), .C1(n392), .C2(n493), .A(n494), .ZN(
        O[38]) );
  AOI22_X1 U136 ( .A1(A_ns[37]), .A2(n397), .B1(\A_s[37] ), .B2(n398), .ZN(
        n494) );
  INV_X1 U137 ( .A(\A_s[36] ), .ZN(n493) );
  INV_X1 U138 ( .A(A_ns[36]), .ZN(n492) );
  OAI221_X1 U139 ( .B1(n393), .B2(n495), .C1(n392), .C2(n496), .A(n497), .ZN(
        O[37]) );
  AOI22_X1 U140 ( .A1(A_ns[36]), .A2(n397), .B1(\A_s[36] ), .B2(n398), .ZN(
        n497) );
  INV_X1 U141 ( .A(\A_s[35] ), .ZN(n496) );
  INV_X1 U142 ( .A(A_ns[35]), .ZN(n495) );
  OAI221_X1 U143 ( .B1(n393), .B2(n498), .C1(n392), .C2(n499), .A(n500), .ZN(
        O[36]) );
  AOI22_X1 U144 ( .A1(A_ns[35]), .A2(n397), .B1(\A_s[35] ), .B2(n398), .ZN(
        n500) );
  INV_X1 U145 ( .A(\A_s[34] ), .ZN(n499) );
  INV_X1 U146 ( .A(A_ns[34]), .ZN(n498) );
  OAI221_X1 U147 ( .B1(n393), .B2(n501), .C1(n392), .C2(n502), .A(n503), .ZN(
        O[35]) );
  AOI22_X1 U148 ( .A1(A_ns[34]), .A2(n397), .B1(\A_s[34] ), .B2(n398), .ZN(
        n503) );
  INV_X1 U149 ( .A(\A_s[33] ), .ZN(n502) );
  INV_X1 U150 ( .A(A_ns[33]), .ZN(n501) );
  OAI221_X1 U151 ( .B1(n393), .B2(n504), .C1(n392), .C2(n505), .A(n506), .ZN(
        O[34]) );
  AOI22_X1 U152 ( .A1(A_ns[33]), .A2(n397), .B1(\A_s[33] ), .B2(n398), .ZN(
        n506) );
  INV_X1 U153 ( .A(\A_s[32] ), .ZN(n505) );
  INV_X1 U154 ( .A(A_ns[32]), .ZN(n504) );
  OAI221_X1 U155 ( .B1(n393), .B2(n507), .C1(n392), .C2(n508), .A(n509), .ZN(
        O[33]) );
  AOI22_X1 U156 ( .A1(A_ns[32]), .A2(n397), .B1(\A_s[32] ), .B2(n398), .ZN(
        n509) );
  INV_X1 U157 ( .A(\A_s[31] ), .ZN(n508) );
  INV_X1 U158 ( .A(A_ns[31]), .ZN(n507) );
  OAI221_X1 U159 ( .B1(n393), .B2(n510), .C1(n392), .C2(n511), .A(n512), .ZN(
        O[32]) );
  AOI22_X1 U160 ( .A1(A_ns[31]), .A2(n397), .B1(\A_s[31] ), .B2(n398), .ZN(
        n512) );
  INV_X1 U161 ( .A(\A_s[30] ), .ZN(n511) );
  INV_X1 U162 ( .A(A_ns[30]), .ZN(n510) );
  OAI221_X1 U163 ( .B1(n393), .B2(n513), .C1(n392), .C2(n514), .A(n515), .ZN(
        O[31]) );
  AOI22_X1 U164 ( .A1(A_ns[30]), .A2(n397), .B1(\A_s[30] ), .B2(n398), .ZN(
        n515) );
  INV_X1 U165 ( .A(\A_s[29] ), .ZN(n514) );
  INV_X1 U166 ( .A(A_ns[29]), .ZN(n513) );
  OAI221_X1 U167 ( .B1(n393), .B2(n516), .C1(n392), .C2(n517), .A(n518), .ZN(
        O[30]) );
  AOI22_X1 U168 ( .A1(A_ns[29]), .A2(n397), .B1(\A_s[29] ), .B2(n398), .ZN(
        n518) );
  INV_X1 U169 ( .A(\A_s[28] ), .ZN(n517) );
  INV_X1 U170 ( .A(A_ns[28]), .ZN(n516) );
  OAI221_X1 U171 ( .B1(n393), .B2(n519), .C1(n392), .C2(n520), .A(n521), .ZN(
        O[2]) );
  AOI22_X1 U172 ( .A1(A_ns[1]), .A2(n397), .B1(\A_s[1] ), .B2(n398), .ZN(n521)
         );
  OAI221_X1 U173 ( .B1(n393), .B2(n522), .C1(n392), .C2(n523), .A(n524), .ZN(
        O[29]) );
  AOI22_X1 U174 ( .A1(A_ns[28]), .A2(n397), .B1(\A_s[28] ), .B2(n398), .ZN(
        n524) );
  INV_X1 U175 ( .A(\A_s[27] ), .ZN(n523) );
  INV_X1 U176 ( .A(A_ns[27]), .ZN(n522) );
  OAI221_X1 U177 ( .B1(n393), .B2(n525), .C1(n392), .C2(n526), .A(n527), .ZN(
        O[28]) );
  AOI22_X1 U178 ( .A1(A_ns[27]), .A2(n397), .B1(\A_s[27] ), .B2(n398), .ZN(
        n527) );
  INV_X1 U179 ( .A(\A_s[26] ), .ZN(n526) );
  INV_X1 U180 ( .A(A_ns[26]), .ZN(n525) );
  OAI221_X1 U181 ( .B1(n393), .B2(n528), .C1(n392), .C2(n529), .A(n530), .ZN(
        O[27]) );
  AOI22_X1 U182 ( .A1(A_ns[26]), .A2(n397), .B1(\A_s[26] ), .B2(n398), .ZN(
        n530) );
  INV_X1 U183 ( .A(\A_s[25] ), .ZN(n529) );
  INV_X1 U184 ( .A(A_ns[25]), .ZN(n528) );
  OAI221_X1 U185 ( .B1(n393), .B2(n531), .C1(n392), .C2(n532), .A(n533), .ZN(
        O[26]) );
  AOI22_X1 U186 ( .A1(A_ns[25]), .A2(n397), .B1(\A_s[25] ), .B2(n398), .ZN(
        n533) );
  INV_X1 U187 ( .A(\A_s[24] ), .ZN(n532) );
  INV_X1 U188 ( .A(A_ns[24]), .ZN(n531) );
  OAI221_X1 U189 ( .B1(n393), .B2(n534), .C1(n392), .C2(n535), .A(n536), .ZN(
        O[25]) );
  AOI22_X1 U190 ( .A1(A_ns[24]), .A2(n397), .B1(\A_s[24] ), .B2(n398), .ZN(
        n536) );
  INV_X1 U191 ( .A(\A_s[23] ), .ZN(n535) );
  INV_X1 U192 ( .A(A_ns[23]), .ZN(n534) );
  OAI221_X1 U193 ( .B1(n393), .B2(n537), .C1(n392), .C2(n538), .A(n539), .ZN(
        O[24]) );
  AOI22_X1 U194 ( .A1(A_ns[23]), .A2(n397), .B1(\A_s[23] ), .B2(n398), .ZN(
        n539) );
  INV_X1 U195 ( .A(\A_s[22] ), .ZN(n538) );
  INV_X1 U196 ( .A(A_ns[22]), .ZN(n537) );
  OAI221_X1 U197 ( .B1(n393), .B2(n540), .C1(n392), .C2(n541), .A(n542), .ZN(
        O[23]) );
  AOI22_X1 U198 ( .A1(A_ns[22]), .A2(n397), .B1(\A_s[22] ), .B2(n398), .ZN(
        n542) );
  INV_X1 U199 ( .A(\A_s[21] ), .ZN(n541) );
  INV_X1 U200 ( .A(A_ns[21]), .ZN(n540) );
  OAI221_X1 U201 ( .B1(n393), .B2(n543), .C1(n392), .C2(n544), .A(n545), .ZN(
        O[22]) );
  AOI22_X1 U202 ( .A1(A_ns[21]), .A2(n397), .B1(\A_s[21] ), .B2(n398), .ZN(
        n545) );
  INV_X1 U203 ( .A(\A_s[20] ), .ZN(n544) );
  INV_X1 U204 ( .A(A_ns[20]), .ZN(n543) );
  OAI221_X1 U205 ( .B1(n393), .B2(n546), .C1(n392), .C2(n547), .A(n548), .ZN(
        O[21]) );
  AOI22_X1 U206 ( .A1(A_ns[20]), .A2(n397), .B1(\A_s[20] ), .B2(n398), .ZN(
        n548) );
  INV_X1 U207 ( .A(\A_s[19] ), .ZN(n547) );
  INV_X1 U208 ( .A(A_ns[19]), .ZN(n546) );
  OAI221_X1 U209 ( .B1(n393), .B2(n549), .C1(n392), .C2(n550), .A(n551), .ZN(
        O[20]) );
  AOI22_X1 U210 ( .A1(A_ns[19]), .A2(n397), .B1(\A_s[19] ), .B2(n398), .ZN(
        n551) );
  INV_X1 U211 ( .A(\A_s[18] ), .ZN(n550) );
  INV_X1 U212 ( .A(A_ns[18]), .ZN(n549) );
  OAI22_X1 U213 ( .A1(n552), .A2(n520), .B1(n553), .B2(n519), .ZN(O[1]) );
  INV_X1 U214 ( .A(A_ns[0]), .ZN(n519) );
  INV_X1 U215 ( .A(\A_s[0] ), .ZN(n520) );
  OAI221_X1 U216 ( .B1(n393), .B2(n554), .C1(n392), .C2(n555), .A(n556), .ZN(
        O[19]) );
  AOI22_X1 U217 ( .A1(A_ns[18]), .A2(n397), .B1(\A_s[18] ), .B2(n398), .ZN(
        n556) );
  INV_X1 U218 ( .A(\A_s[17] ), .ZN(n555) );
  INV_X1 U219 ( .A(A_ns[17]), .ZN(n554) );
  OAI221_X1 U220 ( .B1(n393), .B2(n557), .C1(n392), .C2(n558), .A(n559), .ZN(
        O[18]) );
  AOI22_X1 U221 ( .A1(A_ns[17]), .A2(n397), .B1(\A_s[17] ), .B2(n398), .ZN(
        n559) );
  INV_X1 U222 ( .A(\A_s[16] ), .ZN(n558) );
  INV_X1 U223 ( .A(A_ns[16]), .ZN(n557) );
  OAI221_X1 U224 ( .B1(n393), .B2(n560), .C1(n392), .C2(n561), .A(n562), .ZN(
        O[17]) );
  AOI22_X1 U225 ( .A1(A_ns[16]), .A2(n397), .B1(\A_s[16] ), .B2(n398), .ZN(
        n562) );
  INV_X1 U226 ( .A(\A_s[15] ), .ZN(n561) );
  INV_X1 U227 ( .A(A_ns[15]), .ZN(n560) );
  OAI221_X1 U228 ( .B1(n393), .B2(n563), .C1(n392), .C2(n564), .A(n565), .ZN(
        O[16]) );
  AOI22_X1 U229 ( .A1(A_ns[15]), .A2(n397), .B1(\A_s[15] ), .B2(n398), .ZN(
        n565) );
  INV_X1 U230 ( .A(\A_s[14] ), .ZN(n564) );
  INV_X1 U231 ( .A(A_ns[14]), .ZN(n563) );
  OAI221_X1 U232 ( .B1(n393), .B2(n566), .C1(n392), .C2(n567), .A(n568), .ZN(
        O[15]) );
  AOI22_X1 U233 ( .A1(A_ns[14]), .A2(n397), .B1(\A_s[14] ), .B2(n398), .ZN(
        n568) );
  INV_X1 U234 ( .A(\A_s[13] ), .ZN(n567) );
  INV_X1 U235 ( .A(A_ns[13]), .ZN(n566) );
  OAI221_X1 U236 ( .B1(n393), .B2(n569), .C1(n392), .C2(n570), .A(n571), .ZN(
        O[14]) );
  AOI22_X1 U237 ( .A1(A_ns[13]), .A2(n397), .B1(\A_s[13] ), .B2(n398), .ZN(
        n571) );
  INV_X1 U238 ( .A(\A_s[12] ), .ZN(n570) );
  INV_X1 U239 ( .A(A_ns[12]), .ZN(n569) );
  OAI221_X1 U240 ( .B1(n393), .B2(n572), .C1(n392), .C2(n573), .A(n574), .ZN(
        O[13]) );
  AOI22_X1 U241 ( .A1(A_ns[12]), .A2(n397), .B1(\A_s[12] ), .B2(n398), .ZN(
        n574) );
  INV_X1 U242 ( .A(\A_s[11] ), .ZN(n573) );
  INV_X1 U243 ( .A(A_ns[11]), .ZN(n572) );
  OAI221_X1 U244 ( .B1(n393), .B2(n575), .C1(n392), .C2(n576), .A(n577), .ZN(
        O[12]) );
  AOI22_X1 U245 ( .A1(A_ns[11]), .A2(n397), .B1(\A_s[11] ), .B2(n398), .ZN(
        n577) );
  INV_X1 U246 ( .A(\A_s[10] ), .ZN(n576) );
  INV_X1 U247 ( .A(A_ns[10]), .ZN(n575) );
  OAI221_X1 U248 ( .B1(n393), .B2(n578), .C1(n392), .C2(n579), .A(n580), .ZN(
        O[11]) );
  AOI22_X1 U249 ( .A1(A_ns[10]), .A2(n397), .B1(\A_s[10] ), .B2(n398), .ZN(
        n580) );
  INV_X1 U250 ( .A(\A_s[9] ), .ZN(n579) );
  INV_X1 U251 ( .A(A_ns[9]), .ZN(n578) );
  OAI221_X1 U252 ( .B1(n581), .B2(n393), .C1(n582), .C2(n392), .A(n583), .ZN(
        O[10]) );
  AOI22_X1 U253 ( .A1(A_ns[9]), .A2(n397), .B1(\A_s[9] ), .B2(n398), .ZN(n583)
         );
  NAND2_X1 U254 ( .A1(n584), .A2(n552), .ZN(n553) );
  NAND2_X1 U255 ( .A1(n584), .A2(n585), .ZN(n552) );
  XOR2_X1 U256 ( .A(B[13]), .B(B[14]), .Z(n584) );
  INV_X1 U257 ( .A(\A_s[8] ), .ZN(n582) );
  INV_X1 U258 ( .A(B[15]), .ZN(n585) );
  INV_X1 U259 ( .A(A_ns[8]), .ZN(n581) );
endmodule


module BOOTHENC_NBIT64_i16 ( A, A_n, A_ns, A_s, B, O, A_so, A_nso );
  input [63:0] A;
  input [63:0] A_n;
  input [63:0] A_ns;
  input [63:0] A_s;
  input [63:0] B;
  output [63:0] O;
  output [63:0] A_so;
  output [63:0] A_nso;
  wire   \A_s[61] , \A_s[60] , \A_s[59] , \A_s[58] , \A_s[57] , \A_s[56] ,
         \A_s[55] , \A_s[54] , \A_s[53] , \A_s[52] , \A_s[51] , \A_s[50] ,
         \A_s[49] , \A_s[48] , \A_s[47] , \A_s[46] , \A_s[45] , \A_s[44] ,
         \A_s[43] , \A_s[42] , \A_s[41] , \A_s[40] , \A_s[39] , \A_s[38] ,
         \A_s[37] , \A_s[36] , \A_s[35] , \A_s[34] , \A_s[33] , \A_s[32] ,
         \A_s[31] , \A_s[30] , \A_s[29] , \A_s[28] , \A_s[27] , \A_s[26] ,
         \A_s[25] , \A_s[24] , \A_s[23] , \A_s[22] , \A_s[21] , \A_s[20] ,
         \A_s[19] , \A_s[18] , \A_s[17] , \A_s[16] , \A_s[15] , \A_s[14] ,
         \A_s[13] , \A_s[12] , \A_s[11] , \A_s[10] , \A_s[9] , \A_s[8] ,
         \A_s[7] , \A_s[6] , \A_s[5] , \A_s[4] , \A_s[3] , \A_s[2] , \A_s[1] ,
         \A_s[0] , n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585;
  assign A_nso[0] = 1'b0;
  assign A_nso[1] = 1'b0;
  assign A_so[0] = 1'b0;
  assign A_so[1] = 1'b0;
  assign O[0] = 1'b0;
  assign A_nso[63] = \A_s[61] ;
  assign A_so[63] = \A_s[61] ;
  assign \A_s[61]  = A_s[61];
  assign A_nso[62] = \A_s[60] ;
  assign A_so[62] = \A_s[60] ;
  assign \A_s[60]  = A_s[60];
  assign A_nso[61] = \A_s[59] ;
  assign A_so[61] = \A_s[59] ;
  assign \A_s[59]  = A_s[59];
  assign A_nso[60] = \A_s[58] ;
  assign A_so[60] = \A_s[58] ;
  assign \A_s[58]  = A_s[58];
  assign A_nso[59] = \A_s[57] ;
  assign A_so[59] = \A_s[57] ;
  assign \A_s[57]  = A_s[57];
  assign A_nso[58] = \A_s[56] ;
  assign A_so[58] = \A_s[56] ;
  assign \A_s[56]  = A_s[56];
  assign A_nso[57] = \A_s[55] ;
  assign A_so[57] = \A_s[55] ;
  assign \A_s[55]  = A_s[55];
  assign A_nso[56] = \A_s[54] ;
  assign A_so[56] = \A_s[54] ;
  assign \A_s[54]  = A_s[54];
  assign A_nso[55] = \A_s[53] ;
  assign A_so[55] = \A_s[53] ;
  assign \A_s[53]  = A_s[53];
  assign A_nso[54] = \A_s[52] ;
  assign A_so[54] = \A_s[52] ;
  assign \A_s[52]  = A_s[52];
  assign A_nso[53] = \A_s[51] ;
  assign A_so[53] = \A_s[51] ;
  assign \A_s[51]  = A_s[51];
  assign A_nso[52] = \A_s[50] ;
  assign A_so[52] = \A_s[50] ;
  assign \A_s[50]  = A_s[50];
  assign A_nso[51] = \A_s[49] ;
  assign A_so[51] = \A_s[49] ;
  assign \A_s[49]  = A_s[49];
  assign A_nso[50] = \A_s[48] ;
  assign A_so[50] = \A_s[48] ;
  assign \A_s[48]  = A_s[48];
  assign A_nso[49] = \A_s[47] ;
  assign A_so[49] = \A_s[47] ;
  assign \A_s[47]  = A_s[47];
  assign A_nso[48] = \A_s[46] ;
  assign A_so[48] = \A_s[46] ;
  assign \A_s[46]  = A_s[46];
  assign A_nso[47] = \A_s[45] ;
  assign A_so[47] = \A_s[45] ;
  assign \A_s[45]  = A_s[45];
  assign A_nso[46] = \A_s[44] ;
  assign A_so[46] = \A_s[44] ;
  assign \A_s[44]  = A_s[44];
  assign A_nso[45] = \A_s[43] ;
  assign A_so[45] = \A_s[43] ;
  assign \A_s[43]  = A_s[43];
  assign A_nso[44] = \A_s[42] ;
  assign A_so[44] = \A_s[42] ;
  assign \A_s[42]  = A_s[42];
  assign A_nso[43] = \A_s[41] ;
  assign A_so[43] = \A_s[41] ;
  assign \A_s[41]  = A_s[41];
  assign A_nso[42] = \A_s[40] ;
  assign A_so[42] = \A_s[40] ;
  assign \A_s[40]  = A_s[40];
  assign A_nso[41] = \A_s[39] ;
  assign A_so[41] = \A_s[39] ;
  assign \A_s[39]  = A_s[39];
  assign A_nso[40] = \A_s[38] ;
  assign A_so[40] = \A_s[38] ;
  assign \A_s[38]  = A_s[38];
  assign A_nso[39] = \A_s[37] ;
  assign A_so[39] = \A_s[37] ;
  assign \A_s[37]  = A_s[37];
  assign A_nso[38] = \A_s[36] ;
  assign A_so[38] = \A_s[36] ;
  assign \A_s[36]  = A_s[36];
  assign A_nso[37] = \A_s[35] ;
  assign A_so[37] = \A_s[35] ;
  assign \A_s[35]  = A_s[35];
  assign A_nso[36] = \A_s[34] ;
  assign A_so[36] = \A_s[34] ;
  assign \A_s[34]  = A_s[34];
  assign A_nso[35] = \A_s[33] ;
  assign A_so[35] = \A_s[33] ;
  assign \A_s[33]  = A_s[33];
  assign A_nso[34] = \A_s[32] ;
  assign A_so[34] = \A_s[32] ;
  assign \A_s[32]  = A_s[32];
  assign A_nso[33] = \A_s[31] ;
  assign A_so[33] = \A_s[31] ;
  assign \A_s[31]  = A_s[31];
  assign A_nso[32] = \A_s[30] ;
  assign A_so[32] = \A_s[30] ;
  assign \A_s[30]  = A_s[30];
  assign A_nso[31] = \A_s[29] ;
  assign A_so[31] = \A_s[29] ;
  assign \A_s[29]  = A_s[29];
  assign A_nso[30] = \A_s[28] ;
  assign A_so[30] = \A_s[28] ;
  assign \A_s[28]  = A_s[28];
  assign A_nso[29] = \A_s[27] ;
  assign A_so[29] = \A_s[27] ;
  assign \A_s[27]  = A_s[27];
  assign A_nso[28] = \A_s[26] ;
  assign A_so[28] = \A_s[26] ;
  assign \A_s[26]  = A_s[26];
  assign A_nso[27] = \A_s[25] ;
  assign A_so[27] = \A_s[25] ;
  assign \A_s[25]  = A_s[25];
  assign A_nso[26] = \A_s[24] ;
  assign A_so[26] = \A_s[24] ;
  assign \A_s[24]  = A_s[24];
  assign A_nso[25] = \A_s[23] ;
  assign A_so[25] = \A_s[23] ;
  assign \A_s[23]  = A_s[23];
  assign A_nso[24] = \A_s[22] ;
  assign A_so[24] = \A_s[22] ;
  assign \A_s[22]  = A_s[22];
  assign A_nso[23] = \A_s[21] ;
  assign A_so[23] = \A_s[21] ;
  assign \A_s[21]  = A_s[21];
  assign A_nso[22] = \A_s[20] ;
  assign A_so[22] = \A_s[20] ;
  assign \A_s[20]  = A_s[20];
  assign A_nso[21] = \A_s[19] ;
  assign A_so[21] = \A_s[19] ;
  assign \A_s[19]  = A_s[19];
  assign A_nso[20] = \A_s[18] ;
  assign A_so[20] = \A_s[18] ;
  assign \A_s[18]  = A_s[18];
  assign A_nso[19] = \A_s[17] ;
  assign A_so[19] = \A_s[17] ;
  assign \A_s[17]  = A_s[17];
  assign A_nso[18] = \A_s[16] ;
  assign A_so[18] = \A_s[16] ;
  assign \A_s[16]  = A_s[16];
  assign A_nso[17] = \A_s[15] ;
  assign A_so[17] = \A_s[15] ;
  assign \A_s[15]  = A_s[15];
  assign A_nso[16] = \A_s[14] ;
  assign A_so[16] = \A_s[14] ;
  assign \A_s[14]  = A_s[14];
  assign A_nso[15] = \A_s[13] ;
  assign A_so[15] = \A_s[13] ;
  assign \A_s[13]  = A_s[13];
  assign A_nso[14] = \A_s[12] ;
  assign A_so[14] = \A_s[12] ;
  assign \A_s[12]  = A_s[12];
  assign A_nso[13] = \A_s[11] ;
  assign A_so[13] = \A_s[11] ;
  assign \A_s[11]  = A_s[11];
  assign A_nso[12] = \A_s[10] ;
  assign A_so[12] = \A_s[10] ;
  assign \A_s[10]  = A_s[10];
  assign A_nso[11] = \A_s[9] ;
  assign A_so[11] = \A_s[9] ;
  assign \A_s[9]  = A_s[9];
  assign A_nso[10] = \A_s[8] ;
  assign A_so[10] = \A_s[8] ;
  assign \A_s[8]  = A_s[8];
  assign A_nso[9] = \A_s[7] ;
  assign A_so[9] = \A_s[7] ;
  assign \A_s[7]  = A_s[7];
  assign A_nso[8] = \A_s[6] ;
  assign A_so[8] = \A_s[6] ;
  assign \A_s[6]  = A_s[6];
  assign A_nso[7] = \A_s[5] ;
  assign A_so[7] = \A_s[5] ;
  assign \A_s[5]  = A_s[5];
  assign A_nso[6] = \A_s[4] ;
  assign A_so[6] = \A_s[4] ;
  assign \A_s[4]  = A_s[4];
  assign A_nso[5] = \A_s[3] ;
  assign A_so[5] = \A_s[3] ;
  assign \A_s[3]  = A_s[3];
  assign A_nso[4] = \A_s[2] ;
  assign A_so[4] = \A_s[2] ;
  assign \A_s[2]  = A_s[2];
  assign A_nso[3] = \A_s[1] ;
  assign A_so[3] = \A_s[1] ;
  assign \A_s[1]  = A_s[1];
  assign A_nso[2] = \A_s[0] ;
  assign A_so[2] = \A_s[0] ;
  assign \A_s[0]  = A_s[0];

  AND3_X1 U2 ( .A1(B[16]), .A2(n585), .A3(B[15]), .ZN(n391) );
  INV_X4 U3 ( .A(n391), .ZN(n392) );
  INV_X4 U4 ( .A(n552), .ZN(n398) );
  OR3_X4 U5 ( .A1(B[15]), .A2(B[16]), .A3(n585), .ZN(n393) );
  INV_X4 U6 ( .A(n553), .ZN(n397) );
  OAI221_X1 U7 ( .B1(n393), .B2(n394), .C1(n392), .C2(n395), .A(n396), .ZN(
        O[9]) );
  AOI22_X1 U8 ( .A1(A_ns[8]), .A2(n397), .B1(\A_s[8] ), .B2(n398), .ZN(n396)
         );
  INV_X1 U9 ( .A(\A_s[7] ), .ZN(n395) );
  INV_X1 U10 ( .A(A_ns[7]), .ZN(n394) );
  OAI221_X1 U11 ( .B1(n393), .B2(n399), .C1(n392), .C2(n400), .A(n401), .ZN(
        O[8]) );
  AOI22_X1 U12 ( .A1(A_ns[7]), .A2(n397), .B1(\A_s[7] ), .B2(n398), .ZN(n401)
         );
  INV_X1 U13 ( .A(\A_s[6] ), .ZN(n400) );
  INV_X1 U14 ( .A(A_ns[6]), .ZN(n399) );
  OAI221_X1 U15 ( .B1(n393), .B2(n402), .C1(n392), .C2(n403), .A(n404), .ZN(
        O[7]) );
  AOI22_X1 U16 ( .A1(A_ns[6]), .A2(n397), .B1(\A_s[6] ), .B2(n398), .ZN(n404)
         );
  INV_X1 U17 ( .A(\A_s[5] ), .ZN(n403) );
  INV_X1 U18 ( .A(A_ns[5]), .ZN(n402) );
  OAI221_X1 U19 ( .B1(n393), .B2(n405), .C1(n392), .C2(n406), .A(n407), .ZN(
        O[6]) );
  AOI22_X1 U20 ( .A1(A_ns[5]), .A2(n397), .B1(\A_s[5] ), .B2(n398), .ZN(n407)
         );
  INV_X1 U21 ( .A(\A_s[4] ), .ZN(n406) );
  INV_X1 U22 ( .A(A_ns[4]), .ZN(n405) );
  OAI221_X1 U23 ( .B1(n393), .B2(n408), .C1(n392), .C2(n409), .A(n410), .ZN(
        O[63]) );
  AOI22_X1 U24 ( .A1(A_ns[62]), .A2(n397), .B1(A_s[62]), .B2(n398), .ZN(n410)
         );
  INV_X1 U25 ( .A(\A_s[61] ), .ZN(n409) );
  INV_X1 U26 ( .A(A_ns[61]), .ZN(n408) );
  OAI221_X1 U27 ( .B1(n393), .B2(n411), .C1(n392), .C2(n412), .A(n413), .ZN(
        O[62]) );
  AOI22_X1 U28 ( .A1(A_ns[61]), .A2(n397), .B1(\A_s[61] ), .B2(n398), .ZN(n413) );
  INV_X1 U29 ( .A(\A_s[60] ), .ZN(n412) );
  INV_X1 U30 ( .A(A_ns[60]), .ZN(n411) );
  OAI221_X1 U31 ( .B1(n393), .B2(n414), .C1(n392), .C2(n415), .A(n416), .ZN(
        O[61]) );
  AOI22_X1 U32 ( .A1(A_ns[60]), .A2(n397), .B1(\A_s[60] ), .B2(n398), .ZN(n416) );
  INV_X1 U33 ( .A(\A_s[59] ), .ZN(n415) );
  INV_X1 U34 ( .A(A_ns[59]), .ZN(n414) );
  OAI221_X1 U35 ( .B1(n393), .B2(n417), .C1(n392), .C2(n418), .A(n419), .ZN(
        O[60]) );
  AOI22_X1 U36 ( .A1(A_ns[59]), .A2(n397), .B1(\A_s[59] ), .B2(n398), .ZN(n419) );
  INV_X1 U37 ( .A(\A_s[58] ), .ZN(n418) );
  INV_X1 U38 ( .A(A_ns[58]), .ZN(n417) );
  OAI221_X1 U39 ( .B1(n393), .B2(n420), .C1(n392), .C2(n421), .A(n422), .ZN(
        O[5]) );
  AOI22_X1 U40 ( .A1(A_ns[4]), .A2(n397), .B1(\A_s[4] ), .B2(n398), .ZN(n422)
         );
  INV_X1 U41 ( .A(\A_s[3] ), .ZN(n421) );
  INV_X1 U42 ( .A(A_ns[3]), .ZN(n420) );
  OAI221_X1 U43 ( .B1(n393), .B2(n423), .C1(n392), .C2(n424), .A(n425), .ZN(
        O[59]) );
  AOI22_X1 U44 ( .A1(A_ns[58]), .A2(n397), .B1(\A_s[58] ), .B2(n398), .ZN(n425) );
  INV_X1 U45 ( .A(\A_s[57] ), .ZN(n424) );
  INV_X1 U46 ( .A(A_ns[57]), .ZN(n423) );
  OAI221_X1 U47 ( .B1(n393), .B2(n426), .C1(n392), .C2(n427), .A(n428), .ZN(
        O[58]) );
  AOI22_X1 U48 ( .A1(A_ns[57]), .A2(n397), .B1(\A_s[57] ), .B2(n398), .ZN(n428) );
  INV_X1 U49 ( .A(\A_s[56] ), .ZN(n427) );
  INV_X1 U50 ( .A(A_ns[56]), .ZN(n426) );
  OAI221_X1 U51 ( .B1(n393), .B2(n429), .C1(n392), .C2(n430), .A(n431), .ZN(
        O[57]) );
  AOI22_X1 U52 ( .A1(A_ns[56]), .A2(n397), .B1(\A_s[56] ), .B2(n398), .ZN(n431) );
  INV_X1 U53 ( .A(\A_s[55] ), .ZN(n430) );
  INV_X1 U54 ( .A(A_ns[55]), .ZN(n429) );
  OAI221_X1 U55 ( .B1(n393), .B2(n432), .C1(n392), .C2(n433), .A(n434), .ZN(
        O[56]) );
  AOI22_X1 U56 ( .A1(A_ns[55]), .A2(n397), .B1(\A_s[55] ), .B2(n398), .ZN(n434) );
  INV_X1 U57 ( .A(\A_s[54] ), .ZN(n433) );
  INV_X1 U58 ( .A(A_ns[54]), .ZN(n432) );
  OAI221_X1 U59 ( .B1(n393), .B2(n435), .C1(n392), .C2(n436), .A(n437), .ZN(
        O[55]) );
  AOI22_X1 U60 ( .A1(A_ns[54]), .A2(n397), .B1(\A_s[54] ), .B2(n398), .ZN(n437) );
  INV_X1 U61 ( .A(\A_s[53] ), .ZN(n436) );
  INV_X1 U62 ( .A(A_ns[53]), .ZN(n435) );
  OAI221_X1 U63 ( .B1(n393), .B2(n438), .C1(n392), .C2(n439), .A(n440), .ZN(
        O[54]) );
  AOI22_X1 U64 ( .A1(A_ns[53]), .A2(n397), .B1(\A_s[53] ), .B2(n398), .ZN(n440) );
  INV_X1 U65 ( .A(\A_s[52] ), .ZN(n439) );
  INV_X1 U66 ( .A(A_ns[52]), .ZN(n438) );
  OAI221_X1 U67 ( .B1(n393), .B2(n441), .C1(n392), .C2(n442), .A(n443), .ZN(
        O[53]) );
  AOI22_X1 U68 ( .A1(A_ns[52]), .A2(n397), .B1(\A_s[52] ), .B2(n398), .ZN(n443) );
  INV_X1 U69 ( .A(\A_s[51] ), .ZN(n442) );
  INV_X1 U70 ( .A(A_ns[51]), .ZN(n441) );
  OAI221_X1 U71 ( .B1(n393), .B2(n444), .C1(n392), .C2(n445), .A(n446), .ZN(
        O[52]) );
  AOI22_X1 U72 ( .A1(A_ns[51]), .A2(n397), .B1(\A_s[51] ), .B2(n398), .ZN(n446) );
  INV_X1 U73 ( .A(\A_s[50] ), .ZN(n445) );
  INV_X1 U74 ( .A(A_ns[50]), .ZN(n444) );
  OAI221_X1 U75 ( .B1(n393), .B2(n447), .C1(n392), .C2(n448), .A(n449), .ZN(
        O[51]) );
  AOI22_X1 U76 ( .A1(A_ns[50]), .A2(n397), .B1(\A_s[50] ), .B2(n398), .ZN(n449) );
  INV_X1 U77 ( .A(\A_s[49] ), .ZN(n448) );
  INV_X1 U78 ( .A(A_ns[49]), .ZN(n447) );
  OAI221_X1 U79 ( .B1(n393), .B2(n450), .C1(n392), .C2(n451), .A(n452), .ZN(
        O[50]) );
  AOI22_X1 U80 ( .A1(A_ns[49]), .A2(n397), .B1(\A_s[49] ), .B2(n398), .ZN(n452) );
  INV_X1 U81 ( .A(\A_s[48] ), .ZN(n451) );
  INV_X1 U82 ( .A(A_ns[48]), .ZN(n450) );
  OAI221_X1 U83 ( .B1(n393), .B2(n453), .C1(n392), .C2(n454), .A(n455), .ZN(
        O[4]) );
  AOI22_X1 U84 ( .A1(A_ns[3]), .A2(n397), .B1(\A_s[3] ), .B2(n398), .ZN(n455)
         );
  INV_X1 U85 ( .A(\A_s[2] ), .ZN(n454) );
  INV_X1 U86 ( .A(A_ns[2]), .ZN(n453) );
  OAI221_X1 U87 ( .B1(n393), .B2(n456), .C1(n392), .C2(n457), .A(n458), .ZN(
        O[49]) );
  AOI22_X1 U88 ( .A1(A_ns[48]), .A2(n397), .B1(\A_s[48] ), .B2(n398), .ZN(n458) );
  INV_X1 U89 ( .A(\A_s[47] ), .ZN(n457) );
  INV_X1 U90 ( .A(A_ns[47]), .ZN(n456) );
  OAI221_X1 U91 ( .B1(n393), .B2(n459), .C1(n392), .C2(n460), .A(n461), .ZN(
        O[48]) );
  AOI22_X1 U92 ( .A1(A_ns[47]), .A2(n397), .B1(\A_s[47] ), .B2(n398), .ZN(n461) );
  INV_X1 U93 ( .A(\A_s[46] ), .ZN(n460) );
  INV_X1 U94 ( .A(A_ns[46]), .ZN(n459) );
  OAI221_X1 U95 ( .B1(n393), .B2(n462), .C1(n392), .C2(n463), .A(n464), .ZN(
        O[47]) );
  AOI22_X1 U96 ( .A1(A_ns[46]), .A2(n397), .B1(\A_s[46] ), .B2(n398), .ZN(n464) );
  INV_X1 U97 ( .A(\A_s[45] ), .ZN(n463) );
  INV_X1 U98 ( .A(A_ns[45]), .ZN(n462) );
  OAI221_X1 U99 ( .B1(n393), .B2(n465), .C1(n392), .C2(n466), .A(n467), .ZN(
        O[46]) );
  AOI22_X1 U100 ( .A1(A_ns[45]), .A2(n397), .B1(\A_s[45] ), .B2(n398), .ZN(
        n467) );
  INV_X1 U101 ( .A(\A_s[44] ), .ZN(n466) );
  INV_X1 U102 ( .A(A_ns[44]), .ZN(n465) );
  OAI221_X1 U103 ( .B1(n393), .B2(n468), .C1(n392), .C2(n469), .A(n470), .ZN(
        O[45]) );
  AOI22_X1 U104 ( .A1(A_ns[44]), .A2(n397), .B1(\A_s[44] ), .B2(n398), .ZN(
        n470) );
  INV_X1 U105 ( .A(\A_s[43] ), .ZN(n469) );
  INV_X1 U106 ( .A(A_ns[43]), .ZN(n468) );
  OAI221_X1 U107 ( .B1(n393), .B2(n471), .C1(n392), .C2(n472), .A(n473), .ZN(
        O[44]) );
  AOI22_X1 U108 ( .A1(A_ns[43]), .A2(n397), .B1(\A_s[43] ), .B2(n398), .ZN(
        n473) );
  INV_X1 U109 ( .A(\A_s[42] ), .ZN(n472) );
  INV_X1 U110 ( .A(A_ns[42]), .ZN(n471) );
  OAI221_X1 U111 ( .B1(n393), .B2(n474), .C1(n392), .C2(n475), .A(n476), .ZN(
        O[43]) );
  AOI22_X1 U112 ( .A1(A_ns[42]), .A2(n397), .B1(\A_s[42] ), .B2(n398), .ZN(
        n476) );
  INV_X1 U113 ( .A(\A_s[41] ), .ZN(n475) );
  INV_X1 U114 ( .A(A_ns[41]), .ZN(n474) );
  OAI221_X1 U115 ( .B1(n393), .B2(n477), .C1(n392), .C2(n478), .A(n479), .ZN(
        O[42]) );
  AOI22_X1 U116 ( .A1(A_ns[41]), .A2(n397), .B1(\A_s[41] ), .B2(n398), .ZN(
        n479) );
  INV_X1 U117 ( .A(\A_s[40] ), .ZN(n478) );
  INV_X1 U118 ( .A(A_ns[40]), .ZN(n477) );
  OAI221_X1 U119 ( .B1(n393), .B2(n480), .C1(n392), .C2(n481), .A(n482), .ZN(
        O[41]) );
  AOI22_X1 U120 ( .A1(A_ns[40]), .A2(n397), .B1(\A_s[40] ), .B2(n398), .ZN(
        n482) );
  INV_X1 U121 ( .A(\A_s[39] ), .ZN(n481) );
  INV_X1 U122 ( .A(A_ns[39]), .ZN(n480) );
  OAI221_X1 U123 ( .B1(n393), .B2(n483), .C1(n392), .C2(n484), .A(n485), .ZN(
        O[40]) );
  AOI22_X1 U124 ( .A1(A_ns[39]), .A2(n397), .B1(\A_s[39] ), .B2(n398), .ZN(
        n485) );
  INV_X1 U125 ( .A(\A_s[38] ), .ZN(n484) );
  INV_X1 U126 ( .A(A_ns[38]), .ZN(n483) );
  OAI221_X1 U127 ( .B1(n393), .B2(n486), .C1(n392), .C2(n487), .A(n488), .ZN(
        O[3]) );
  AOI22_X1 U128 ( .A1(A_ns[2]), .A2(n397), .B1(\A_s[2] ), .B2(n398), .ZN(n488)
         );
  INV_X1 U129 ( .A(\A_s[1] ), .ZN(n487) );
  INV_X1 U130 ( .A(A_ns[1]), .ZN(n486) );
  OAI221_X1 U131 ( .B1(n393), .B2(n489), .C1(n392), .C2(n490), .A(n491), .ZN(
        O[39]) );
  AOI22_X1 U132 ( .A1(A_ns[38]), .A2(n397), .B1(\A_s[38] ), .B2(n398), .ZN(
        n491) );
  INV_X1 U133 ( .A(\A_s[37] ), .ZN(n490) );
  INV_X1 U134 ( .A(A_ns[37]), .ZN(n489) );
  OAI221_X1 U135 ( .B1(n393), .B2(n492), .C1(n392), .C2(n493), .A(n494), .ZN(
        O[38]) );
  AOI22_X1 U136 ( .A1(A_ns[37]), .A2(n397), .B1(\A_s[37] ), .B2(n398), .ZN(
        n494) );
  INV_X1 U137 ( .A(\A_s[36] ), .ZN(n493) );
  INV_X1 U138 ( .A(A_ns[36]), .ZN(n492) );
  OAI221_X1 U139 ( .B1(n393), .B2(n495), .C1(n392), .C2(n496), .A(n497), .ZN(
        O[37]) );
  AOI22_X1 U140 ( .A1(A_ns[36]), .A2(n397), .B1(\A_s[36] ), .B2(n398), .ZN(
        n497) );
  INV_X1 U141 ( .A(\A_s[35] ), .ZN(n496) );
  INV_X1 U142 ( .A(A_ns[35]), .ZN(n495) );
  OAI221_X1 U143 ( .B1(n393), .B2(n498), .C1(n392), .C2(n499), .A(n500), .ZN(
        O[36]) );
  AOI22_X1 U144 ( .A1(A_ns[35]), .A2(n397), .B1(\A_s[35] ), .B2(n398), .ZN(
        n500) );
  INV_X1 U145 ( .A(\A_s[34] ), .ZN(n499) );
  INV_X1 U146 ( .A(A_ns[34]), .ZN(n498) );
  OAI221_X1 U147 ( .B1(n393), .B2(n501), .C1(n392), .C2(n502), .A(n503), .ZN(
        O[35]) );
  AOI22_X1 U148 ( .A1(A_ns[34]), .A2(n397), .B1(\A_s[34] ), .B2(n398), .ZN(
        n503) );
  INV_X1 U149 ( .A(\A_s[33] ), .ZN(n502) );
  INV_X1 U150 ( .A(A_ns[33]), .ZN(n501) );
  OAI221_X1 U151 ( .B1(n393), .B2(n504), .C1(n392), .C2(n505), .A(n506), .ZN(
        O[34]) );
  AOI22_X1 U152 ( .A1(A_ns[33]), .A2(n397), .B1(\A_s[33] ), .B2(n398), .ZN(
        n506) );
  INV_X1 U153 ( .A(\A_s[32] ), .ZN(n505) );
  INV_X1 U154 ( .A(A_ns[32]), .ZN(n504) );
  OAI221_X1 U155 ( .B1(n393), .B2(n507), .C1(n392), .C2(n508), .A(n509), .ZN(
        O[33]) );
  AOI22_X1 U156 ( .A1(A_ns[32]), .A2(n397), .B1(\A_s[32] ), .B2(n398), .ZN(
        n509) );
  INV_X1 U157 ( .A(\A_s[31] ), .ZN(n508) );
  INV_X1 U158 ( .A(A_ns[31]), .ZN(n507) );
  OAI221_X1 U159 ( .B1(n393), .B2(n510), .C1(n392), .C2(n511), .A(n512), .ZN(
        O[32]) );
  AOI22_X1 U160 ( .A1(A_ns[31]), .A2(n397), .B1(\A_s[31] ), .B2(n398), .ZN(
        n512) );
  INV_X1 U161 ( .A(\A_s[30] ), .ZN(n511) );
  INV_X1 U162 ( .A(A_ns[30]), .ZN(n510) );
  OAI221_X1 U163 ( .B1(n393), .B2(n513), .C1(n392), .C2(n514), .A(n515), .ZN(
        O[31]) );
  AOI22_X1 U164 ( .A1(A_ns[30]), .A2(n397), .B1(\A_s[30] ), .B2(n398), .ZN(
        n515) );
  INV_X1 U165 ( .A(\A_s[29] ), .ZN(n514) );
  INV_X1 U166 ( .A(A_ns[29]), .ZN(n513) );
  OAI221_X1 U167 ( .B1(n393), .B2(n516), .C1(n392), .C2(n517), .A(n518), .ZN(
        O[30]) );
  AOI22_X1 U168 ( .A1(A_ns[29]), .A2(n397), .B1(\A_s[29] ), .B2(n398), .ZN(
        n518) );
  INV_X1 U169 ( .A(\A_s[28] ), .ZN(n517) );
  INV_X1 U170 ( .A(A_ns[28]), .ZN(n516) );
  OAI221_X1 U171 ( .B1(n393), .B2(n519), .C1(n392), .C2(n520), .A(n521), .ZN(
        O[2]) );
  AOI22_X1 U172 ( .A1(A_ns[1]), .A2(n397), .B1(\A_s[1] ), .B2(n398), .ZN(n521)
         );
  OAI221_X1 U173 ( .B1(n393), .B2(n522), .C1(n392), .C2(n523), .A(n524), .ZN(
        O[29]) );
  AOI22_X1 U174 ( .A1(A_ns[28]), .A2(n397), .B1(\A_s[28] ), .B2(n398), .ZN(
        n524) );
  INV_X1 U175 ( .A(\A_s[27] ), .ZN(n523) );
  INV_X1 U176 ( .A(A_ns[27]), .ZN(n522) );
  OAI221_X1 U177 ( .B1(n393), .B2(n525), .C1(n392), .C2(n526), .A(n527), .ZN(
        O[28]) );
  AOI22_X1 U178 ( .A1(A_ns[27]), .A2(n397), .B1(\A_s[27] ), .B2(n398), .ZN(
        n527) );
  INV_X1 U179 ( .A(\A_s[26] ), .ZN(n526) );
  INV_X1 U180 ( .A(A_ns[26]), .ZN(n525) );
  OAI221_X1 U181 ( .B1(n393), .B2(n528), .C1(n392), .C2(n529), .A(n530), .ZN(
        O[27]) );
  AOI22_X1 U182 ( .A1(A_ns[26]), .A2(n397), .B1(\A_s[26] ), .B2(n398), .ZN(
        n530) );
  INV_X1 U183 ( .A(\A_s[25] ), .ZN(n529) );
  INV_X1 U184 ( .A(A_ns[25]), .ZN(n528) );
  OAI221_X1 U185 ( .B1(n393), .B2(n531), .C1(n392), .C2(n532), .A(n533), .ZN(
        O[26]) );
  AOI22_X1 U186 ( .A1(A_ns[25]), .A2(n397), .B1(\A_s[25] ), .B2(n398), .ZN(
        n533) );
  INV_X1 U187 ( .A(\A_s[24] ), .ZN(n532) );
  INV_X1 U188 ( .A(A_ns[24]), .ZN(n531) );
  OAI221_X1 U189 ( .B1(n393), .B2(n534), .C1(n392), .C2(n535), .A(n536), .ZN(
        O[25]) );
  AOI22_X1 U190 ( .A1(A_ns[24]), .A2(n397), .B1(\A_s[24] ), .B2(n398), .ZN(
        n536) );
  INV_X1 U191 ( .A(\A_s[23] ), .ZN(n535) );
  INV_X1 U192 ( .A(A_ns[23]), .ZN(n534) );
  OAI221_X1 U193 ( .B1(n393), .B2(n537), .C1(n392), .C2(n538), .A(n539), .ZN(
        O[24]) );
  AOI22_X1 U194 ( .A1(A_ns[23]), .A2(n397), .B1(\A_s[23] ), .B2(n398), .ZN(
        n539) );
  INV_X1 U195 ( .A(\A_s[22] ), .ZN(n538) );
  INV_X1 U196 ( .A(A_ns[22]), .ZN(n537) );
  OAI221_X1 U197 ( .B1(n393), .B2(n540), .C1(n392), .C2(n541), .A(n542), .ZN(
        O[23]) );
  AOI22_X1 U198 ( .A1(A_ns[22]), .A2(n397), .B1(\A_s[22] ), .B2(n398), .ZN(
        n542) );
  INV_X1 U199 ( .A(\A_s[21] ), .ZN(n541) );
  INV_X1 U200 ( .A(A_ns[21]), .ZN(n540) );
  OAI221_X1 U201 ( .B1(n393), .B2(n543), .C1(n392), .C2(n544), .A(n545), .ZN(
        O[22]) );
  AOI22_X1 U202 ( .A1(A_ns[21]), .A2(n397), .B1(\A_s[21] ), .B2(n398), .ZN(
        n545) );
  INV_X1 U203 ( .A(\A_s[20] ), .ZN(n544) );
  INV_X1 U204 ( .A(A_ns[20]), .ZN(n543) );
  OAI221_X1 U205 ( .B1(n393), .B2(n546), .C1(n392), .C2(n547), .A(n548), .ZN(
        O[21]) );
  AOI22_X1 U206 ( .A1(A_ns[20]), .A2(n397), .B1(\A_s[20] ), .B2(n398), .ZN(
        n548) );
  INV_X1 U207 ( .A(\A_s[19] ), .ZN(n547) );
  INV_X1 U208 ( .A(A_ns[19]), .ZN(n546) );
  OAI221_X1 U209 ( .B1(n393), .B2(n549), .C1(n392), .C2(n550), .A(n551), .ZN(
        O[20]) );
  AOI22_X1 U210 ( .A1(A_ns[19]), .A2(n397), .B1(\A_s[19] ), .B2(n398), .ZN(
        n551) );
  INV_X1 U211 ( .A(\A_s[18] ), .ZN(n550) );
  INV_X1 U212 ( .A(A_ns[18]), .ZN(n549) );
  OAI22_X1 U213 ( .A1(n552), .A2(n520), .B1(n553), .B2(n519), .ZN(O[1]) );
  INV_X1 U214 ( .A(A_ns[0]), .ZN(n519) );
  INV_X1 U215 ( .A(\A_s[0] ), .ZN(n520) );
  OAI221_X1 U216 ( .B1(n393), .B2(n554), .C1(n392), .C2(n555), .A(n556), .ZN(
        O[19]) );
  AOI22_X1 U217 ( .A1(A_ns[18]), .A2(n397), .B1(\A_s[18] ), .B2(n398), .ZN(
        n556) );
  INV_X1 U218 ( .A(\A_s[17] ), .ZN(n555) );
  INV_X1 U219 ( .A(A_ns[17]), .ZN(n554) );
  OAI221_X1 U220 ( .B1(n393), .B2(n557), .C1(n392), .C2(n558), .A(n559), .ZN(
        O[18]) );
  AOI22_X1 U221 ( .A1(A_ns[17]), .A2(n397), .B1(\A_s[17] ), .B2(n398), .ZN(
        n559) );
  INV_X1 U222 ( .A(\A_s[16] ), .ZN(n558) );
  INV_X1 U223 ( .A(A_ns[16]), .ZN(n557) );
  OAI221_X1 U224 ( .B1(n393), .B2(n560), .C1(n392), .C2(n561), .A(n562), .ZN(
        O[17]) );
  AOI22_X1 U225 ( .A1(A_ns[16]), .A2(n397), .B1(\A_s[16] ), .B2(n398), .ZN(
        n562) );
  INV_X1 U226 ( .A(\A_s[15] ), .ZN(n561) );
  INV_X1 U227 ( .A(A_ns[15]), .ZN(n560) );
  OAI221_X1 U228 ( .B1(n393), .B2(n563), .C1(n392), .C2(n564), .A(n565), .ZN(
        O[16]) );
  AOI22_X1 U229 ( .A1(A_ns[15]), .A2(n397), .B1(\A_s[15] ), .B2(n398), .ZN(
        n565) );
  INV_X1 U230 ( .A(\A_s[14] ), .ZN(n564) );
  INV_X1 U231 ( .A(A_ns[14]), .ZN(n563) );
  OAI221_X1 U232 ( .B1(n393), .B2(n566), .C1(n392), .C2(n567), .A(n568), .ZN(
        O[15]) );
  AOI22_X1 U233 ( .A1(A_ns[14]), .A2(n397), .B1(\A_s[14] ), .B2(n398), .ZN(
        n568) );
  INV_X1 U234 ( .A(\A_s[13] ), .ZN(n567) );
  INV_X1 U235 ( .A(A_ns[13]), .ZN(n566) );
  OAI221_X1 U236 ( .B1(n393), .B2(n569), .C1(n392), .C2(n570), .A(n571), .ZN(
        O[14]) );
  AOI22_X1 U237 ( .A1(A_ns[13]), .A2(n397), .B1(\A_s[13] ), .B2(n398), .ZN(
        n571) );
  INV_X1 U238 ( .A(\A_s[12] ), .ZN(n570) );
  INV_X1 U239 ( .A(A_ns[12]), .ZN(n569) );
  OAI221_X1 U240 ( .B1(n393), .B2(n572), .C1(n392), .C2(n573), .A(n574), .ZN(
        O[13]) );
  AOI22_X1 U241 ( .A1(A_ns[12]), .A2(n397), .B1(\A_s[12] ), .B2(n398), .ZN(
        n574) );
  INV_X1 U242 ( .A(\A_s[11] ), .ZN(n573) );
  INV_X1 U243 ( .A(A_ns[11]), .ZN(n572) );
  OAI221_X1 U244 ( .B1(n393), .B2(n575), .C1(n392), .C2(n576), .A(n577), .ZN(
        O[12]) );
  AOI22_X1 U245 ( .A1(A_ns[11]), .A2(n397), .B1(\A_s[11] ), .B2(n398), .ZN(
        n577) );
  INV_X1 U246 ( .A(\A_s[10] ), .ZN(n576) );
  INV_X1 U247 ( .A(A_ns[10]), .ZN(n575) );
  OAI221_X1 U248 ( .B1(n393), .B2(n578), .C1(n392), .C2(n579), .A(n580), .ZN(
        O[11]) );
  AOI22_X1 U249 ( .A1(A_ns[10]), .A2(n397), .B1(\A_s[10] ), .B2(n398), .ZN(
        n580) );
  INV_X1 U250 ( .A(\A_s[9] ), .ZN(n579) );
  INV_X1 U251 ( .A(A_ns[9]), .ZN(n578) );
  OAI221_X1 U252 ( .B1(n581), .B2(n393), .C1(n582), .C2(n392), .A(n583), .ZN(
        O[10]) );
  AOI22_X1 U253 ( .A1(A_ns[9]), .A2(n397), .B1(\A_s[9] ), .B2(n398), .ZN(n583)
         );
  NAND2_X1 U254 ( .A1(n584), .A2(n552), .ZN(n553) );
  NAND2_X1 U255 ( .A1(n584), .A2(n585), .ZN(n552) );
  XOR2_X1 U256 ( .A(B[15]), .B(B[16]), .Z(n584) );
  INV_X1 U257 ( .A(\A_s[8] ), .ZN(n582) );
  INV_X1 U258 ( .A(B[17]), .ZN(n585) );
  INV_X1 U259 ( .A(A_ns[8]), .ZN(n581) );
endmodule


module BOOTHENC_NBIT64_i18 ( A, A_n, A_ns, A_s, B, O, A_so, A_nso );
  input [63:0] A;
  input [63:0] A_n;
  input [63:0] A_ns;
  input [63:0] A_s;
  input [63:0] B;
  output [63:0] O;
  output [63:0] A_so;
  output [63:0] A_nso;
  wire   \A_s[61] , \A_s[60] , \A_s[59] , \A_s[58] , \A_s[57] , \A_s[56] ,
         \A_s[55] , \A_s[54] , \A_s[53] , \A_s[52] , \A_s[51] , \A_s[50] ,
         \A_s[49] , \A_s[48] , \A_s[47] , \A_s[46] , \A_s[45] , \A_s[44] ,
         \A_s[43] , \A_s[42] , \A_s[41] , \A_s[40] , \A_s[39] , \A_s[38] ,
         \A_s[37] , \A_s[36] , \A_s[35] , \A_s[34] , \A_s[33] , \A_s[32] ,
         \A_s[31] , \A_s[30] , \A_s[29] , \A_s[28] , \A_s[27] , \A_s[26] ,
         \A_s[25] , \A_s[24] , \A_s[23] , \A_s[22] , \A_s[21] , \A_s[20] ,
         \A_s[19] , \A_s[18] , \A_s[17] , \A_s[16] , \A_s[15] , \A_s[14] ,
         \A_s[13] , \A_s[12] , \A_s[11] , \A_s[10] , \A_s[9] , \A_s[8] ,
         \A_s[7] , \A_s[6] , \A_s[5] , \A_s[4] , \A_s[3] , \A_s[2] , \A_s[1] ,
         \A_s[0] , n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585;
  assign A_nso[0] = 1'b0;
  assign A_nso[1] = 1'b0;
  assign A_so[0] = 1'b0;
  assign A_so[1] = 1'b0;
  assign O[0] = 1'b0;
  assign A_nso[63] = \A_s[61] ;
  assign A_so[63] = \A_s[61] ;
  assign \A_s[61]  = A_s[61];
  assign A_nso[62] = \A_s[60] ;
  assign A_so[62] = \A_s[60] ;
  assign \A_s[60]  = A_s[60];
  assign A_nso[61] = \A_s[59] ;
  assign A_so[61] = \A_s[59] ;
  assign \A_s[59]  = A_s[59];
  assign A_nso[60] = \A_s[58] ;
  assign A_so[60] = \A_s[58] ;
  assign \A_s[58]  = A_s[58];
  assign A_nso[59] = \A_s[57] ;
  assign A_so[59] = \A_s[57] ;
  assign \A_s[57]  = A_s[57];
  assign A_nso[58] = \A_s[56] ;
  assign A_so[58] = \A_s[56] ;
  assign \A_s[56]  = A_s[56];
  assign A_nso[57] = \A_s[55] ;
  assign A_so[57] = \A_s[55] ;
  assign \A_s[55]  = A_s[55];
  assign A_nso[56] = \A_s[54] ;
  assign A_so[56] = \A_s[54] ;
  assign \A_s[54]  = A_s[54];
  assign A_nso[55] = \A_s[53] ;
  assign A_so[55] = \A_s[53] ;
  assign \A_s[53]  = A_s[53];
  assign A_nso[54] = \A_s[52] ;
  assign A_so[54] = \A_s[52] ;
  assign \A_s[52]  = A_s[52];
  assign A_nso[53] = \A_s[51] ;
  assign A_so[53] = \A_s[51] ;
  assign \A_s[51]  = A_s[51];
  assign A_nso[52] = \A_s[50] ;
  assign A_so[52] = \A_s[50] ;
  assign \A_s[50]  = A_s[50];
  assign A_nso[51] = \A_s[49] ;
  assign A_so[51] = \A_s[49] ;
  assign \A_s[49]  = A_s[49];
  assign A_nso[50] = \A_s[48] ;
  assign A_so[50] = \A_s[48] ;
  assign \A_s[48]  = A_s[48];
  assign A_nso[49] = \A_s[47] ;
  assign A_so[49] = \A_s[47] ;
  assign \A_s[47]  = A_s[47];
  assign A_nso[48] = \A_s[46] ;
  assign A_so[48] = \A_s[46] ;
  assign \A_s[46]  = A_s[46];
  assign A_nso[47] = \A_s[45] ;
  assign A_so[47] = \A_s[45] ;
  assign \A_s[45]  = A_s[45];
  assign A_nso[46] = \A_s[44] ;
  assign A_so[46] = \A_s[44] ;
  assign \A_s[44]  = A_s[44];
  assign A_nso[45] = \A_s[43] ;
  assign A_so[45] = \A_s[43] ;
  assign \A_s[43]  = A_s[43];
  assign A_nso[44] = \A_s[42] ;
  assign A_so[44] = \A_s[42] ;
  assign \A_s[42]  = A_s[42];
  assign A_nso[43] = \A_s[41] ;
  assign A_so[43] = \A_s[41] ;
  assign \A_s[41]  = A_s[41];
  assign A_nso[42] = \A_s[40] ;
  assign A_so[42] = \A_s[40] ;
  assign \A_s[40]  = A_s[40];
  assign A_nso[41] = \A_s[39] ;
  assign A_so[41] = \A_s[39] ;
  assign \A_s[39]  = A_s[39];
  assign A_nso[40] = \A_s[38] ;
  assign A_so[40] = \A_s[38] ;
  assign \A_s[38]  = A_s[38];
  assign A_nso[39] = \A_s[37] ;
  assign A_so[39] = \A_s[37] ;
  assign \A_s[37]  = A_s[37];
  assign A_nso[38] = \A_s[36] ;
  assign A_so[38] = \A_s[36] ;
  assign \A_s[36]  = A_s[36];
  assign A_nso[37] = \A_s[35] ;
  assign A_so[37] = \A_s[35] ;
  assign \A_s[35]  = A_s[35];
  assign A_nso[36] = \A_s[34] ;
  assign A_so[36] = \A_s[34] ;
  assign \A_s[34]  = A_s[34];
  assign A_nso[35] = \A_s[33] ;
  assign A_so[35] = \A_s[33] ;
  assign \A_s[33]  = A_s[33];
  assign A_nso[34] = \A_s[32] ;
  assign A_so[34] = \A_s[32] ;
  assign \A_s[32]  = A_s[32];
  assign A_nso[33] = \A_s[31] ;
  assign A_so[33] = \A_s[31] ;
  assign \A_s[31]  = A_s[31];
  assign A_nso[32] = \A_s[30] ;
  assign A_so[32] = \A_s[30] ;
  assign \A_s[30]  = A_s[30];
  assign A_nso[31] = \A_s[29] ;
  assign A_so[31] = \A_s[29] ;
  assign \A_s[29]  = A_s[29];
  assign A_nso[30] = \A_s[28] ;
  assign A_so[30] = \A_s[28] ;
  assign \A_s[28]  = A_s[28];
  assign A_nso[29] = \A_s[27] ;
  assign A_so[29] = \A_s[27] ;
  assign \A_s[27]  = A_s[27];
  assign A_nso[28] = \A_s[26] ;
  assign A_so[28] = \A_s[26] ;
  assign \A_s[26]  = A_s[26];
  assign A_nso[27] = \A_s[25] ;
  assign A_so[27] = \A_s[25] ;
  assign \A_s[25]  = A_s[25];
  assign A_nso[26] = \A_s[24] ;
  assign A_so[26] = \A_s[24] ;
  assign \A_s[24]  = A_s[24];
  assign A_nso[25] = \A_s[23] ;
  assign A_so[25] = \A_s[23] ;
  assign \A_s[23]  = A_s[23];
  assign A_nso[24] = \A_s[22] ;
  assign A_so[24] = \A_s[22] ;
  assign \A_s[22]  = A_s[22];
  assign A_nso[23] = \A_s[21] ;
  assign A_so[23] = \A_s[21] ;
  assign \A_s[21]  = A_s[21];
  assign A_nso[22] = \A_s[20] ;
  assign A_so[22] = \A_s[20] ;
  assign \A_s[20]  = A_s[20];
  assign A_nso[21] = \A_s[19] ;
  assign A_so[21] = \A_s[19] ;
  assign \A_s[19]  = A_s[19];
  assign A_nso[20] = \A_s[18] ;
  assign A_so[20] = \A_s[18] ;
  assign \A_s[18]  = A_s[18];
  assign A_nso[19] = \A_s[17] ;
  assign A_so[19] = \A_s[17] ;
  assign \A_s[17]  = A_s[17];
  assign A_nso[18] = \A_s[16] ;
  assign A_so[18] = \A_s[16] ;
  assign \A_s[16]  = A_s[16];
  assign A_nso[17] = \A_s[15] ;
  assign A_so[17] = \A_s[15] ;
  assign \A_s[15]  = A_s[15];
  assign A_nso[16] = \A_s[14] ;
  assign A_so[16] = \A_s[14] ;
  assign \A_s[14]  = A_s[14];
  assign A_nso[15] = \A_s[13] ;
  assign A_so[15] = \A_s[13] ;
  assign \A_s[13]  = A_s[13];
  assign A_nso[14] = \A_s[12] ;
  assign A_so[14] = \A_s[12] ;
  assign \A_s[12]  = A_s[12];
  assign A_nso[13] = \A_s[11] ;
  assign A_so[13] = \A_s[11] ;
  assign \A_s[11]  = A_s[11];
  assign A_nso[12] = \A_s[10] ;
  assign A_so[12] = \A_s[10] ;
  assign \A_s[10]  = A_s[10];
  assign A_nso[11] = \A_s[9] ;
  assign A_so[11] = \A_s[9] ;
  assign \A_s[9]  = A_s[9];
  assign A_nso[10] = \A_s[8] ;
  assign A_so[10] = \A_s[8] ;
  assign \A_s[8]  = A_s[8];
  assign A_nso[9] = \A_s[7] ;
  assign A_so[9] = \A_s[7] ;
  assign \A_s[7]  = A_s[7];
  assign A_nso[8] = \A_s[6] ;
  assign A_so[8] = \A_s[6] ;
  assign \A_s[6]  = A_s[6];
  assign A_nso[7] = \A_s[5] ;
  assign A_so[7] = \A_s[5] ;
  assign \A_s[5]  = A_s[5];
  assign A_nso[6] = \A_s[4] ;
  assign A_so[6] = \A_s[4] ;
  assign \A_s[4]  = A_s[4];
  assign A_nso[5] = \A_s[3] ;
  assign A_so[5] = \A_s[3] ;
  assign \A_s[3]  = A_s[3];
  assign A_nso[4] = \A_s[2] ;
  assign A_so[4] = \A_s[2] ;
  assign \A_s[2]  = A_s[2];
  assign A_nso[3] = \A_s[1] ;
  assign A_so[3] = \A_s[1] ;
  assign \A_s[1]  = A_s[1];
  assign A_nso[2] = \A_s[0] ;
  assign A_so[2] = \A_s[0] ;
  assign \A_s[0]  = A_s[0];

  AND3_X1 U2 ( .A1(B[18]), .A2(n585), .A3(B[17]), .ZN(n391) );
  INV_X4 U3 ( .A(n391), .ZN(n392) );
  INV_X4 U4 ( .A(n552), .ZN(n398) );
  OR3_X4 U5 ( .A1(B[17]), .A2(B[18]), .A3(n585), .ZN(n393) );
  INV_X4 U6 ( .A(n553), .ZN(n397) );
  OAI221_X1 U7 ( .B1(n393), .B2(n394), .C1(n392), .C2(n395), .A(n396), .ZN(
        O[9]) );
  AOI22_X1 U8 ( .A1(A_ns[8]), .A2(n397), .B1(\A_s[8] ), .B2(n398), .ZN(n396)
         );
  INV_X1 U9 ( .A(\A_s[7] ), .ZN(n395) );
  INV_X1 U10 ( .A(A_ns[7]), .ZN(n394) );
  OAI221_X1 U11 ( .B1(n393), .B2(n399), .C1(n392), .C2(n400), .A(n401), .ZN(
        O[8]) );
  AOI22_X1 U12 ( .A1(A_ns[7]), .A2(n397), .B1(\A_s[7] ), .B2(n398), .ZN(n401)
         );
  INV_X1 U13 ( .A(\A_s[6] ), .ZN(n400) );
  INV_X1 U14 ( .A(A_ns[6]), .ZN(n399) );
  OAI221_X1 U15 ( .B1(n393), .B2(n402), .C1(n392), .C2(n403), .A(n404), .ZN(
        O[7]) );
  AOI22_X1 U16 ( .A1(A_ns[6]), .A2(n397), .B1(\A_s[6] ), .B2(n398), .ZN(n404)
         );
  INV_X1 U17 ( .A(\A_s[5] ), .ZN(n403) );
  INV_X1 U18 ( .A(A_ns[5]), .ZN(n402) );
  OAI221_X1 U19 ( .B1(n393), .B2(n405), .C1(n392), .C2(n406), .A(n407), .ZN(
        O[6]) );
  AOI22_X1 U20 ( .A1(A_ns[5]), .A2(n397), .B1(\A_s[5] ), .B2(n398), .ZN(n407)
         );
  INV_X1 U21 ( .A(\A_s[4] ), .ZN(n406) );
  INV_X1 U22 ( .A(A_ns[4]), .ZN(n405) );
  OAI221_X1 U23 ( .B1(n393), .B2(n408), .C1(n392), .C2(n409), .A(n410), .ZN(
        O[63]) );
  AOI22_X1 U24 ( .A1(A_ns[62]), .A2(n397), .B1(A_s[62]), .B2(n398), .ZN(n410)
         );
  INV_X1 U25 ( .A(\A_s[61] ), .ZN(n409) );
  INV_X1 U26 ( .A(A_ns[61]), .ZN(n408) );
  OAI221_X1 U27 ( .B1(n393), .B2(n411), .C1(n392), .C2(n412), .A(n413), .ZN(
        O[62]) );
  AOI22_X1 U28 ( .A1(A_ns[61]), .A2(n397), .B1(\A_s[61] ), .B2(n398), .ZN(n413) );
  INV_X1 U29 ( .A(\A_s[60] ), .ZN(n412) );
  INV_X1 U30 ( .A(A_ns[60]), .ZN(n411) );
  OAI221_X1 U31 ( .B1(n393), .B2(n414), .C1(n392), .C2(n415), .A(n416), .ZN(
        O[61]) );
  AOI22_X1 U32 ( .A1(A_ns[60]), .A2(n397), .B1(\A_s[60] ), .B2(n398), .ZN(n416) );
  INV_X1 U33 ( .A(\A_s[59] ), .ZN(n415) );
  INV_X1 U34 ( .A(A_ns[59]), .ZN(n414) );
  OAI221_X1 U35 ( .B1(n393), .B2(n417), .C1(n392), .C2(n418), .A(n419), .ZN(
        O[60]) );
  AOI22_X1 U36 ( .A1(A_ns[59]), .A2(n397), .B1(\A_s[59] ), .B2(n398), .ZN(n419) );
  INV_X1 U37 ( .A(\A_s[58] ), .ZN(n418) );
  INV_X1 U38 ( .A(A_ns[58]), .ZN(n417) );
  OAI221_X1 U39 ( .B1(n393), .B2(n420), .C1(n392), .C2(n421), .A(n422), .ZN(
        O[5]) );
  AOI22_X1 U40 ( .A1(A_ns[4]), .A2(n397), .B1(\A_s[4] ), .B2(n398), .ZN(n422)
         );
  INV_X1 U41 ( .A(\A_s[3] ), .ZN(n421) );
  INV_X1 U42 ( .A(A_ns[3]), .ZN(n420) );
  OAI221_X1 U43 ( .B1(n393), .B2(n423), .C1(n392), .C2(n424), .A(n425), .ZN(
        O[59]) );
  AOI22_X1 U44 ( .A1(A_ns[58]), .A2(n397), .B1(\A_s[58] ), .B2(n398), .ZN(n425) );
  INV_X1 U45 ( .A(\A_s[57] ), .ZN(n424) );
  INV_X1 U46 ( .A(A_ns[57]), .ZN(n423) );
  OAI221_X1 U47 ( .B1(n393), .B2(n426), .C1(n392), .C2(n427), .A(n428), .ZN(
        O[58]) );
  AOI22_X1 U48 ( .A1(A_ns[57]), .A2(n397), .B1(\A_s[57] ), .B2(n398), .ZN(n428) );
  INV_X1 U49 ( .A(\A_s[56] ), .ZN(n427) );
  INV_X1 U50 ( .A(A_ns[56]), .ZN(n426) );
  OAI221_X1 U51 ( .B1(n393), .B2(n429), .C1(n392), .C2(n430), .A(n431), .ZN(
        O[57]) );
  AOI22_X1 U52 ( .A1(A_ns[56]), .A2(n397), .B1(\A_s[56] ), .B2(n398), .ZN(n431) );
  INV_X1 U53 ( .A(\A_s[55] ), .ZN(n430) );
  INV_X1 U54 ( .A(A_ns[55]), .ZN(n429) );
  OAI221_X1 U55 ( .B1(n393), .B2(n432), .C1(n392), .C2(n433), .A(n434), .ZN(
        O[56]) );
  AOI22_X1 U56 ( .A1(A_ns[55]), .A2(n397), .B1(\A_s[55] ), .B2(n398), .ZN(n434) );
  INV_X1 U57 ( .A(\A_s[54] ), .ZN(n433) );
  INV_X1 U58 ( .A(A_ns[54]), .ZN(n432) );
  OAI221_X1 U59 ( .B1(n393), .B2(n435), .C1(n392), .C2(n436), .A(n437), .ZN(
        O[55]) );
  AOI22_X1 U60 ( .A1(A_ns[54]), .A2(n397), .B1(\A_s[54] ), .B2(n398), .ZN(n437) );
  INV_X1 U61 ( .A(\A_s[53] ), .ZN(n436) );
  INV_X1 U62 ( .A(A_ns[53]), .ZN(n435) );
  OAI221_X1 U63 ( .B1(n393), .B2(n438), .C1(n392), .C2(n439), .A(n440), .ZN(
        O[54]) );
  AOI22_X1 U64 ( .A1(A_ns[53]), .A2(n397), .B1(\A_s[53] ), .B2(n398), .ZN(n440) );
  INV_X1 U65 ( .A(\A_s[52] ), .ZN(n439) );
  INV_X1 U66 ( .A(A_ns[52]), .ZN(n438) );
  OAI221_X1 U67 ( .B1(n393), .B2(n441), .C1(n392), .C2(n442), .A(n443), .ZN(
        O[53]) );
  AOI22_X1 U68 ( .A1(A_ns[52]), .A2(n397), .B1(\A_s[52] ), .B2(n398), .ZN(n443) );
  INV_X1 U69 ( .A(\A_s[51] ), .ZN(n442) );
  INV_X1 U70 ( .A(A_ns[51]), .ZN(n441) );
  OAI221_X1 U71 ( .B1(n393), .B2(n444), .C1(n392), .C2(n445), .A(n446), .ZN(
        O[52]) );
  AOI22_X1 U72 ( .A1(A_ns[51]), .A2(n397), .B1(\A_s[51] ), .B2(n398), .ZN(n446) );
  INV_X1 U73 ( .A(\A_s[50] ), .ZN(n445) );
  INV_X1 U74 ( .A(A_ns[50]), .ZN(n444) );
  OAI221_X1 U75 ( .B1(n393), .B2(n447), .C1(n392), .C2(n448), .A(n449), .ZN(
        O[51]) );
  AOI22_X1 U76 ( .A1(A_ns[50]), .A2(n397), .B1(\A_s[50] ), .B2(n398), .ZN(n449) );
  INV_X1 U77 ( .A(\A_s[49] ), .ZN(n448) );
  INV_X1 U78 ( .A(A_ns[49]), .ZN(n447) );
  OAI221_X1 U79 ( .B1(n393), .B2(n450), .C1(n392), .C2(n451), .A(n452), .ZN(
        O[50]) );
  AOI22_X1 U80 ( .A1(A_ns[49]), .A2(n397), .B1(\A_s[49] ), .B2(n398), .ZN(n452) );
  INV_X1 U81 ( .A(\A_s[48] ), .ZN(n451) );
  INV_X1 U82 ( .A(A_ns[48]), .ZN(n450) );
  OAI221_X1 U83 ( .B1(n393), .B2(n453), .C1(n392), .C2(n454), .A(n455), .ZN(
        O[4]) );
  AOI22_X1 U84 ( .A1(A_ns[3]), .A2(n397), .B1(\A_s[3] ), .B2(n398), .ZN(n455)
         );
  INV_X1 U85 ( .A(\A_s[2] ), .ZN(n454) );
  INV_X1 U86 ( .A(A_ns[2]), .ZN(n453) );
  OAI221_X1 U87 ( .B1(n393), .B2(n456), .C1(n392), .C2(n457), .A(n458), .ZN(
        O[49]) );
  AOI22_X1 U88 ( .A1(A_ns[48]), .A2(n397), .B1(\A_s[48] ), .B2(n398), .ZN(n458) );
  INV_X1 U89 ( .A(\A_s[47] ), .ZN(n457) );
  INV_X1 U90 ( .A(A_ns[47]), .ZN(n456) );
  OAI221_X1 U91 ( .B1(n393), .B2(n459), .C1(n392), .C2(n460), .A(n461), .ZN(
        O[48]) );
  AOI22_X1 U92 ( .A1(A_ns[47]), .A2(n397), .B1(\A_s[47] ), .B2(n398), .ZN(n461) );
  INV_X1 U93 ( .A(\A_s[46] ), .ZN(n460) );
  INV_X1 U94 ( .A(A_ns[46]), .ZN(n459) );
  OAI221_X1 U95 ( .B1(n393), .B2(n462), .C1(n392), .C2(n463), .A(n464), .ZN(
        O[47]) );
  AOI22_X1 U96 ( .A1(A_ns[46]), .A2(n397), .B1(\A_s[46] ), .B2(n398), .ZN(n464) );
  INV_X1 U97 ( .A(\A_s[45] ), .ZN(n463) );
  INV_X1 U98 ( .A(A_ns[45]), .ZN(n462) );
  OAI221_X1 U99 ( .B1(n393), .B2(n465), .C1(n392), .C2(n466), .A(n467), .ZN(
        O[46]) );
  AOI22_X1 U100 ( .A1(A_ns[45]), .A2(n397), .B1(\A_s[45] ), .B2(n398), .ZN(
        n467) );
  INV_X1 U101 ( .A(\A_s[44] ), .ZN(n466) );
  INV_X1 U102 ( .A(A_ns[44]), .ZN(n465) );
  OAI221_X1 U103 ( .B1(n393), .B2(n468), .C1(n392), .C2(n469), .A(n470), .ZN(
        O[45]) );
  AOI22_X1 U104 ( .A1(A_ns[44]), .A2(n397), .B1(\A_s[44] ), .B2(n398), .ZN(
        n470) );
  INV_X1 U105 ( .A(\A_s[43] ), .ZN(n469) );
  INV_X1 U106 ( .A(A_ns[43]), .ZN(n468) );
  OAI221_X1 U107 ( .B1(n393), .B2(n471), .C1(n392), .C2(n472), .A(n473), .ZN(
        O[44]) );
  AOI22_X1 U108 ( .A1(A_ns[43]), .A2(n397), .B1(\A_s[43] ), .B2(n398), .ZN(
        n473) );
  INV_X1 U109 ( .A(\A_s[42] ), .ZN(n472) );
  INV_X1 U110 ( .A(A_ns[42]), .ZN(n471) );
  OAI221_X1 U111 ( .B1(n393), .B2(n474), .C1(n392), .C2(n475), .A(n476), .ZN(
        O[43]) );
  AOI22_X1 U112 ( .A1(A_ns[42]), .A2(n397), .B1(\A_s[42] ), .B2(n398), .ZN(
        n476) );
  INV_X1 U113 ( .A(\A_s[41] ), .ZN(n475) );
  INV_X1 U114 ( .A(A_ns[41]), .ZN(n474) );
  OAI221_X1 U115 ( .B1(n393), .B2(n477), .C1(n392), .C2(n478), .A(n479), .ZN(
        O[42]) );
  AOI22_X1 U116 ( .A1(A_ns[41]), .A2(n397), .B1(\A_s[41] ), .B2(n398), .ZN(
        n479) );
  INV_X1 U117 ( .A(\A_s[40] ), .ZN(n478) );
  INV_X1 U118 ( .A(A_ns[40]), .ZN(n477) );
  OAI221_X1 U119 ( .B1(n393), .B2(n480), .C1(n392), .C2(n481), .A(n482), .ZN(
        O[41]) );
  AOI22_X1 U120 ( .A1(A_ns[40]), .A2(n397), .B1(\A_s[40] ), .B2(n398), .ZN(
        n482) );
  INV_X1 U121 ( .A(\A_s[39] ), .ZN(n481) );
  INV_X1 U122 ( .A(A_ns[39]), .ZN(n480) );
  OAI221_X1 U123 ( .B1(n393), .B2(n483), .C1(n392), .C2(n484), .A(n485), .ZN(
        O[40]) );
  AOI22_X1 U124 ( .A1(A_ns[39]), .A2(n397), .B1(\A_s[39] ), .B2(n398), .ZN(
        n485) );
  INV_X1 U125 ( .A(\A_s[38] ), .ZN(n484) );
  INV_X1 U126 ( .A(A_ns[38]), .ZN(n483) );
  OAI221_X1 U127 ( .B1(n393), .B2(n486), .C1(n392), .C2(n487), .A(n488), .ZN(
        O[3]) );
  AOI22_X1 U128 ( .A1(A_ns[2]), .A2(n397), .B1(\A_s[2] ), .B2(n398), .ZN(n488)
         );
  INV_X1 U129 ( .A(\A_s[1] ), .ZN(n487) );
  INV_X1 U130 ( .A(A_ns[1]), .ZN(n486) );
  OAI221_X1 U131 ( .B1(n393), .B2(n489), .C1(n392), .C2(n490), .A(n491), .ZN(
        O[39]) );
  AOI22_X1 U132 ( .A1(A_ns[38]), .A2(n397), .B1(\A_s[38] ), .B2(n398), .ZN(
        n491) );
  INV_X1 U133 ( .A(\A_s[37] ), .ZN(n490) );
  INV_X1 U134 ( .A(A_ns[37]), .ZN(n489) );
  OAI221_X1 U135 ( .B1(n393), .B2(n492), .C1(n392), .C2(n493), .A(n494), .ZN(
        O[38]) );
  AOI22_X1 U136 ( .A1(A_ns[37]), .A2(n397), .B1(\A_s[37] ), .B2(n398), .ZN(
        n494) );
  INV_X1 U137 ( .A(\A_s[36] ), .ZN(n493) );
  INV_X1 U138 ( .A(A_ns[36]), .ZN(n492) );
  OAI221_X1 U139 ( .B1(n393), .B2(n495), .C1(n392), .C2(n496), .A(n497), .ZN(
        O[37]) );
  AOI22_X1 U140 ( .A1(A_ns[36]), .A2(n397), .B1(\A_s[36] ), .B2(n398), .ZN(
        n497) );
  INV_X1 U141 ( .A(\A_s[35] ), .ZN(n496) );
  INV_X1 U142 ( .A(A_ns[35]), .ZN(n495) );
  OAI221_X1 U143 ( .B1(n393), .B2(n498), .C1(n392), .C2(n499), .A(n500), .ZN(
        O[36]) );
  AOI22_X1 U144 ( .A1(A_ns[35]), .A2(n397), .B1(\A_s[35] ), .B2(n398), .ZN(
        n500) );
  INV_X1 U145 ( .A(\A_s[34] ), .ZN(n499) );
  INV_X1 U146 ( .A(A_ns[34]), .ZN(n498) );
  OAI221_X1 U147 ( .B1(n393), .B2(n501), .C1(n392), .C2(n502), .A(n503), .ZN(
        O[35]) );
  AOI22_X1 U148 ( .A1(A_ns[34]), .A2(n397), .B1(\A_s[34] ), .B2(n398), .ZN(
        n503) );
  INV_X1 U149 ( .A(\A_s[33] ), .ZN(n502) );
  INV_X1 U150 ( .A(A_ns[33]), .ZN(n501) );
  OAI221_X1 U151 ( .B1(n393), .B2(n504), .C1(n392), .C2(n505), .A(n506), .ZN(
        O[34]) );
  AOI22_X1 U152 ( .A1(A_ns[33]), .A2(n397), .B1(\A_s[33] ), .B2(n398), .ZN(
        n506) );
  INV_X1 U153 ( .A(\A_s[32] ), .ZN(n505) );
  INV_X1 U154 ( .A(A_ns[32]), .ZN(n504) );
  OAI221_X1 U155 ( .B1(n393), .B2(n507), .C1(n392), .C2(n508), .A(n509), .ZN(
        O[33]) );
  AOI22_X1 U156 ( .A1(A_ns[32]), .A2(n397), .B1(\A_s[32] ), .B2(n398), .ZN(
        n509) );
  INV_X1 U157 ( .A(\A_s[31] ), .ZN(n508) );
  INV_X1 U158 ( .A(A_ns[31]), .ZN(n507) );
  OAI221_X1 U159 ( .B1(n393), .B2(n510), .C1(n392), .C2(n511), .A(n512), .ZN(
        O[32]) );
  AOI22_X1 U160 ( .A1(A_ns[31]), .A2(n397), .B1(\A_s[31] ), .B2(n398), .ZN(
        n512) );
  INV_X1 U161 ( .A(\A_s[30] ), .ZN(n511) );
  INV_X1 U162 ( .A(A_ns[30]), .ZN(n510) );
  OAI221_X1 U163 ( .B1(n393), .B2(n513), .C1(n392), .C2(n514), .A(n515), .ZN(
        O[31]) );
  AOI22_X1 U164 ( .A1(A_ns[30]), .A2(n397), .B1(\A_s[30] ), .B2(n398), .ZN(
        n515) );
  INV_X1 U165 ( .A(\A_s[29] ), .ZN(n514) );
  INV_X1 U166 ( .A(A_ns[29]), .ZN(n513) );
  OAI221_X1 U167 ( .B1(n393), .B2(n516), .C1(n392), .C2(n517), .A(n518), .ZN(
        O[30]) );
  AOI22_X1 U168 ( .A1(A_ns[29]), .A2(n397), .B1(\A_s[29] ), .B2(n398), .ZN(
        n518) );
  INV_X1 U169 ( .A(\A_s[28] ), .ZN(n517) );
  INV_X1 U170 ( .A(A_ns[28]), .ZN(n516) );
  OAI221_X1 U171 ( .B1(n393), .B2(n519), .C1(n392), .C2(n520), .A(n521), .ZN(
        O[2]) );
  AOI22_X1 U172 ( .A1(A_ns[1]), .A2(n397), .B1(\A_s[1] ), .B2(n398), .ZN(n521)
         );
  OAI221_X1 U173 ( .B1(n393), .B2(n522), .C1(n392), .C2(n523), .A(n524), .ZN(
        O[29]) );
  AOI22_X1 U174 ( .A1(A_ns[28]), .A2(n397), .B1(\A_s[28] ), .B2(n398), .ZN(
        n524) );
  INV_X1 U175 ( .A(\A_s[27] ), .ZN(n523) );
  INV_X1 U176 ( .A(A_ns[27]), .ZN(n522) );
  OAI221_X1 U177 ( .B1(n393), .B2(n525), .C1(n392), .C2(n526), .A(n527), .ZN(
        O[28]) );
  AOI22_X1 U178 ( .A1(A_ns[27]), .A2(n397), .B1(\A_s[27] ), .B2(n398), .ZN(
        n527) );
  INV_X1 U179 ( .A(\A_s[26] ), .ZN(n526) );
  INV_X1 U180 ( .A(A_ns[26]), .ZN(n525) );
  OAI221_X1 U181 ( .B1(n393), .B2(n528), .C1(n392), .C2(n529), .A(n530), .ZN(
        O[27]) );
  AOI22_X1 U182 ( .A1(A_ns[26]), .A2(n397), .B1(\A_s[26] ), .B2(n398), .ZN(
        n530) );
  INV_X1 U183 ( .A(\A_s[25] ), .ZN(n529) );
  INV_X1 U184 ( .A(A_ns[25]), .ZN(n528) );
  OAI221_X1 U185 ( .B1(n393), .B2(n531), .C1(n392), .C2(n532), .A(n533), .ZN(
        O[26]) );
  AOI22_X1 U186 ( .A1(A_ns[25]), .A2(n397), .B1(\A_s[25] ), .B2(n398), .ZN(
        n533) );
  INV_X1 U187 ( .A(\A_s[24] ), .ZN(n532) );
  INV_X1 U188 ( .A(A_ns[24]), .ZN(n531) );
  OAI221_X1 U189 ( .B1(n393), .B2(n534), .C1(n392), .C2(n535), .A(n536), .ZN(
        O[25]) );
  AOI22_X1 U190 ( .A1(A_ns[24]), .A2(n397), .B1(\A_s[24] ), .B2(n398), .ZN(
        n536) );
  INV_X1 U191 ( .A(\A_s[23] ), .ZN(n535) );
  INV_X1 U192 ( .A(A_ns[23]), .ZN(n534) );
  OAI221_X1 U193 ( .B1(n393), .B2(n537), .C1(n392), .C2(n538), .A(n539), .ZN(
        O[24]) );
  AOI22_X1 U194 ( .A1(A_ns[23]), .A2(n397), .B1(\A_s[23] ), .B2(n398), .ZN(
        n539) );
  INV_X1 U195 ( .A(\A_s[22] ), .ZN(n538) );
  INV_X1 U196 ( .A(A_ns[22]), .ZN(n537) );
  OAI221_X1 U197 ( .B1(n393), .B2(n540), .C1(n392), .C2(n541), .A(n542), .ZN(
        O[23]) );
  AOI22_X1 U198 ( .A1(A_ns[22]), .A2(n397), .B1(\A_s[22] ), .B2(n398), .ZN(
        n542) );
  INV_X1 U199 ( .A(\A_s[21] ), .ZN(n541) );
  INV_X1 U200 ( .A(A_ns[21]), .ZN(n540) );
  OAI221_X1 U201 ( .B1(n393), .B2(n543), .C1(n392), .C2(n544), .A(n545), .ZN(
        O[22]) );
  AOI22_X1 U202 ( .A1(A_ns[21]), .A2(n397), .B1(\A_s[21] ), .B2(n398), .ZN(
        n545) );
  INV_X1 U203 ( .A(\A_s[20] ), .ZN(n544) );
  INV_X1 U204 ( .A(A_ns[20]), .ZN(n543) );
  OAI221_X1 U205 ( .B1(n393), .B2(n546), .C1(n392), .C2(n547), .A(n548), .ZN(
        O[21]) );
  AOI22_X1 U206 ( .A1(A_ns[20]), .A2(n397), .B1(\A_s[20] ), .B2(n398), .ZN(
        n548) );
  INV_X1 U207 ( .A(\A_s[19] ), .ZN(n547) );
  INV_X1 U208 ( .A(A_ns[19]), .ZN(n546) );
  OAI221_X1 U209 ( .B1(n393), .B2(n549), .C1(n392), .C2(n550), .A(n551), .ZN(
        O[20]) );
  AOI22_X1 U210 ( .A1(A_ns[19]), .A2(n397), .B1(\A_s[19] ), .B2(n398), .ZN(
        n551) );
  INV_X1 U211 ( .A(\A_s[18] ), .ZN(n550) );
  INV_X1 U212 ( .A(A_ns[18]), .ZN(n549) );
  OAI22_X1 U213 ( .A1(n552), .A2(n520), .B1(n553), .B2(n519), .ZN(O[1]) );
  INV_X1 U214 ( .A(A_ns[0]), .ZN(n519) );
  INV_X1 U215 ( .A(\A_s[0] ), .ZN(n520) );
  OAI221_X1 U216 ( .B1(n393), .B2(n554), .C1(n392), .C2(n555), .A(n556), .ZN(
        O[19]) );
  AOI22_X1 U217 ( .A1(A_ns[18]), .A2(n397), .B1(\A_s[18] ), .B2(n398), .ZN(
        n556) );
  INV_X1 U218 ( .A(\A_s[17] ), .ZN(n555) );
  INV_X1 U219 ( .A(A_ns[17]), .ZN(n554) );
  OAI221_X1 U220 ( .B1(n393), .B2(n557), .C1(n392), .C2(n558), .A(n559), .ZN(
        O[18]) );
  AOI22_X1 U221 ( .A1(A_ns[17]), .A2(n397), .B1(\A_s[17] ), .B2(n398), .ZN(
        n559) );
  INV_X1 U222 ( .A(\A_s[16] ), .ZN(n558) );
  INV_X1 U223 ( .A(A_ns[16]), .ZN(n557) );
  OAI221_X1 U224 ( .B1(n393), .B2(n560), .C1(n392), .C2(n561), .A(n562), .ZN(
        O[17]) );
  AOI22_X1 U225 ( .A1(A_ns[16]), .A2(n397), .B1(\A_s[16] ), .B2(n398), .ZN(
        n562) );
  INV_X1 U226 ( .A(\A_s[15] ), .ZN(n561) );
  INV_X1 U227 ( .A(A_ns[15]), .ZN(n560) );
  OAI221_X1 U228 ( .B1(n393), .B2(n563), .C1(n392), .C2(n564), .A(n565), .ZN(
        O[16]) );
  AOI22_X1 U229 ( .A1(A_ns[15]), .A2(n397), .B1(\A_s[15] ), .B2(n398), .ZN(
        n565) );
  INV_X1 U230 ( .A(\A_s[14] ), .ZN(n564) );
  INV_X1 U231 ( .A(A_ns[14]), .ZN(n563) );
  OAI221_X1 U232 ( .B1(n393), .B2(n566), .C1(n392), .C2(n567), .A(n568), .ZN(
        O[15]) );
  AOI22_X1 U233 ( .A1(A_ns[14]), .A2(n397), .B1(\A_s[14] ), .B2(n398), .ZN(
        n568) );
  INV_X1 U234 ( .A(\A_s[13] ), .ZN(n567) );
  INV_X1 U235 ( .A(A_ns[13]), .ZN(n566) );
  OAI221_X1 U236 ( .B1(n393), .B2(n569), .C1(n392), .C2(n570), .A(n571), .ZN(
        O[14]) );
  AOI22_X1 U237 ( .A1(A_ns[13]), .A2(n397), .B1(\A_s[13] ), .B2(n398), .ZN(
        n571) );
  INV_X1 U238 ( .A(\A_s[12] ), .ZN(n570) );
  INV_X1 U239 ( .A(A_ns[12]), .ZN(n569) );
  OAI221_X1 U240 ( .B1(n393), .B2(n572), .C1(n392), .C2(n573), .A(n574), .ZN(
        O[13]) );
  AOI22_X1 U241 ( .A1(A_ns[12]), .A2(n397), .B1(\A_s[12] ), .B2(n398), .ZN(
        n574) );
  INV_X1 U242 ( .A(\A_s[11] ), .ZN(n573) );
  INV_X1 U243 ( .A(A_ns[11]), .ZN(n572) );
  OAI221_X1 U244 ( .B1(n393), .B2(n575), .C1(n392), .C2(n576), .A(n577), .ZN(
        O[12]) );
  AOI22_X1 U245 ( .A1(A_ns[11]), .A2(n397), .B1(\A_s[11] ), .B2(n398), .ZN(
        n577) );
  INV_X1 U246 ( .A(\A_s[10] ), .ZN(n576) );
  INV_X1 U247 ( .A(A_ns[10]), .ZN(n575) );
  OAI221_X1 U248 ( .B1(n393), .B2(n578), .C1(n392), .C2(n579), .A(n580), .ZN(
        O[11]) );
  AOI22_X1 U249 ( .A1(A_ns[10]), .A2(n397), .B1(\A_s[10] ), .B2(n398), .ZN(
        n580) );
  INV_X1 U250 ( .A(\A_s[9] ), .ZN(n579) );
  INV_X1 U251 ( .A(A_ns[9]), .ZN(n578) );
  OAI221_X1 U252 ( .B1(n581), .B2(n393), .C1(n582), .C2(n392), .A(n583), .ZN(
        O[10]) );
  AOI22_X1 U253 ( .A1(A_ns[9]), .A2(n397), .B1(\A_s[9] ), .B2(n398), .ZN(n583)
         );
  NAND2_X1 U254 ( .A1(n584), .A2(n552), .ZN(n553) );
  NAND2_X1 U255 ( .A1(n584), .A2(n585), .ZN(n552) );
  XOR2_X1 U256 ( .A(B[17]), .B(B[18]), .Z(n584) );
  INV_X1 U257 ( .A(\A_s[8] ), .ZN(n582) );
  INV_X1 U258 ( .A(B[19]), .ZN(n585) );
  INV_X1 U259 ( .A(A_ns[8]), .ZN(n581) );
endmodule


module BOOTHENC_NBIT64_i20 ( A, A_n, A_ns, A_s, B, O, A_so, A_nso );
  input [63:0] A;
  input [63:0] A_n;
  input [63:0] A_ns;
  input [63:0] A_s;
  input [63:0] B;
  output [63:0] O;
  output [63:0] A_so;
  output [63:0] A_nso;
  wire   \A_s[61] , \A_s[60] , \A_s[59] , \A_s[58] , \A_s[57] , \A_s[56] ,
         \A_s[55] , \A_s[54] , \A_s[53] , \A_s[52] , \A_s[51] , \A_s[50] ,
         \A_s[49] , \A_s[48] , \A_s[47] , \A_s[46] , \A_s[45] , \A_s[44] ,
         \A_s[43] , \A_s[42] , \A_s[41] , \A_s[40] , \A_s[39] , \A_s[38] ,
         \A_s[37] , \A_s[36] , \A_s[35] , \A_s[34] , \A_s[33] , \A_s[32] ,
         \A_s[31] , \A_s[30] , \A_s[29] , \A_s[28] , \A_s[27] , \A_s[26] ,
         \A_s[25] , \A_s[24] , \A_s[23] , \A_s[22] , \A_s[21] , \A_s[20] ,
         \A_s[19] , \A_s[18] , \A_s[17] , \A_s[16] , \A_s[15] , \A_s[14] ,
         \A_s[13] , \A_s[12] , \A_s[11] , \A_s[10] , \A_s[9] , \A_s[8] ,
         \A_s[7] , \A_s[6] , \A_s[5] , \A_s[4] , \A_s[3] , \A_s[2] , \A_s[1] ,
         \A_s[0] , n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585;
  assign A_nso[0] = 1'b0;
  assign A_nso[1] = 1'b0;
  assign A_so[0] = 1'b0;
  assign A_so[1] = 1'b0;
  assign O[0] = 1'b0;
  assign A_nso[63] = \A_s[61] ;
  assign A_so[63] = \A_s[61] ;
  assign \A_s[61]  = A_s[61];
  assign A_nso[62] = \A_s[60] ;
  assign A_so[62] = \A_s[60] ;
  assign \A_s[60]  = A_s[60];
  assign A_nso[61] = \A_s[59] ;
  assign A_so[61] = \A_s[59] ;
  assign \A_s[59]  = A_s[59];
  assign A_nso[60] = \A_s[58] ;
  assign A_so[60] = \A_s[58] ;
  assign \A_s[58]  = A_s[58];
  assign A_nso[59] = \A_s[57] ;
  assign A_so[59] = \A_s[57] ;
  assign \A_s[57]  = A_s[57];
  assign A_nso[58] = \A_s[56] ;
  assign A_so[58] = \A_s[56] ;
  assign \A_s[56]  = A_s[56];
  assign A_nso[57] = \A_s[55] ;
  assign A_so[57] = \A_s[55] ;
  assign \A_s[55]  = A_s[55];
  assign A_nso[56] = \A_s[54] ;
  assign A_so[56] = \A_s[54] ;
  assign \A_s[54]  = A_s[54];
  assign A_nso[55] = \A_s[53] ;
  assign A_so[55] = \A_s[53] ;
  assign \A_s[53]  = A_s[53];
  assign A_nso[54] = \A_s[52] ;
  assign A_so[54] = \A_s[52] ;
  assign \A_s[52]  = A_s[52];
  assign A_nso[53] = \A_s[51] ;
  assign A_so[53] = \A_s[51] ;
  assign \A_s[51]  = A_s[51];
  assign A_nso[52] = \A_s[50] ;
  assign A_so[52] = \A_s[50] ;
  assign \A_s[50]  = A_s[50];
  assign A_nso[51] = \A_s[49] ;
  assign A_so[51] = \A_s[49] ;
  assign \A_s[49]  = A_s[49];
  assign A_nso[50] = \A_s[48] ;
  assign A_so[50] = \A_s[48] ;
  assign \A_s[48]  = A_s[48];
  assign A_nso[49] = \A_s[47] ;
  assign A_so[49] = \A_s[47] ;
  assign \A_s[47]  = A_s[47];
  assign A_nso[48] = \A_s[46] ;
  assign A_so[48] = \A_s[46] ;
  assign \A_s[46]  = A_s[46];
  assign A_nso[47] = \A_s[45] ;
  assign A_so[47] = \A_s[45] ;
  assign \A_s[45]  = A_s[45];
  assign A_nso[46] = \A_s[44] ;
  assign A_so[46] = \A_s[44] ;
  assign \A_s[44]  = A_s[44];
  assign A_nso[45] = \A_s[43] ;
  assign A_so[45] = \A_s[43] ;
  assign \A_s[43]  = A_s[43];
  assign A_nso[44] = \A_s[42] ;
  assign A_so[44] = \A_s[42] ;
  assign \A_s[42]  = A_s[42];
  assign A_nso[43] = \A_s[41] ;
  assign A_so[43] = \A_s[41] ;
  assign \A_s[41]  = A_s[41];
  assign A_nso[42] = \A_s[40] ;
  assign A_so[42] = \A_s[40] ;
  assign \A_s[40]  = A_s[40];
  assign A_nso[41] = \A_s[39] ;
  assign A_so[41] = \A_s[39] ;
  assign \A_s[39]  = A_s[39];
  assign A_nso[40] = \A_s[38] ;
  assign A_so[40] = \A_s[38] ;
  assign \A_s[38]  = A_s[38];
  assign A_nso[39] = \A_s[37] ;
  assign A_so[39] = \A_s[37] ;
  assign \A_s[37]  = A_s[37];
  assign A_nso[38] = \A_s[36] ;
  assign A_so[38] = \A_s[36] ;
  assign \A_s[36]  = A_s[36];
  assign A_nso[37] = \A_s[35] ;
  assign A_so[37] = \A_s[35] ;
  assign \A_s[35]  = A_s[35];
  assign A_nso[36] = \A_s[34] ;
  assign A_so[36] = \A_s[34] ;
  assign \A_s[34]  = A_s[34];
  assign A_nso[35] = \A_s[33] ;
  assign A_so[35] = \A_s[33] ;
  assign \A_s[33]  = A_s[33];
  assign A_nso[34] = \A_s[32] ;
  assign A_so[34] = \A_s[32] ;
  assign \A_s[32]  = A_s[32];
  assign A_nso[33] = \A_s[31] ;
  assign A_so[33] = \A_s[31] ;
  assign \A_s[31]  = A_s[31];
  assign A_nso[32] = \A_s[30] ;
  assign A_so[32] = \A_s[30] ;
  assign \A_s[30]  = A_s[30];
  assign A_nso[31] = \A_s[29] ;
  assign A_so[31] = \A_s[29] ;
  assign \A_s[29]  = A_s[29];
  assign A_nso[30] = \A_s[28] ;
  assign A_so[30] = \A_s[28] ;
  assign \A_s[28]  = A_s[28];
  assign A_nso[29] = \A_s[27] ;
  assign A_so[29] = \A_s[27] ;
  assign \A_s[27]  = A_s[27];
  assign A_nso[28] = \A_s[26] ;
  assign A_so[28] = \A_s[26] ;
  assign \A_s[26]  = A_s[26];
  assign A_nso[27] = \A_s[25] ;
  assign A_so[27] = \A_s[25] ;
  assign \A_s[25]  = A_s[25];
  assign A_nso[26] = \A_s[24] ;
  assign A_so[26] = \A_s[24] ;
  assign \A_s[24]  = A_s[24];
  assign A_nso[25] = \A_s[23] ;
  assign A_so[25] = \A_s[23] ;
  assign \A_s[23]  = A_s[23];
  assign A_nso[24] = \A_s[22] ;
  assign A_so[24] = \A_s[22] ;
  assign \A_s[22]  = A_s[22];
  assign A_nso[23] = \A_s[21] ;
  assign A_so[23] = \A_s[21] ;
  assign \A_s[21]  = A_s[21];
  assign A_nso[22] = \A_s[20] ;
  assign A_so[22] = \A_s[20] ;
  assign \A_s[20]  = A_s[20];
  assign A_nso[21] = \A_s[19] ;
  assign A_so[21] = \A_s[19] ;
  assign \A_s[19]  = A_s[19];
  assign A_nso[20] = \A_s[18] ;
  assign A_so[20] = \A_s[18] ;
  assign \A_s[18]  = A_s[18];
  assign A_nso[19] = \A_s[17] ;
  assign A_so[19] = \A_s[17] ;
  assign \A_s[17]  = A_s[17];
  assign A_nso[18] = \A_s[16] ;
  assign A_so[18] = \A_s[16] ;
  assign \A_s[16]  = A_s[16];
  assign A_nso[17] = \A_s[15] ;
  assign A_so[17] = \A_s[15] ;
  assign \A_s[15]  = A_s[15];
  assign A_nso[16] = \A_s[14] ;
  assign A_so[16] = \A_s[14] ;
  assign \A_s[14]  = A_s[14];
  assign A_nso[15] = \A_s[13] ;
  assign A_so[15] = \A_s[13] ;
  assign \A_s[13]  = A_s[13];
  assign A_nso[14] = \A_s[12] ;
  assign A_so[14] = \A_s[12] ;
  assign \A_s[12]  = A_s[12];
  assign A_nso[13] = \A_s[11] ;
  assign A_so[13] = \A_s[11] ;
  assign \A_s[11]  = A_s[11];
  assign A_nso[12] = \A_s[10] ;
  assign A_so[12] = \A_s[10] ;
  assign \A_s[10]  = A_s[10];
  assign A_nso[11] = \A_s[9] ;
  assign A_so[11] = \A_s[9] ;
  assign \A_s[9]  = A_s[9];
  assign A_nso[10] = \A_s[8] ;
  assign A_so[10] = \A_s[8] ;
  assign \A_s[8]  = A_s[8];
  assign A_nso[9] = \A_s[7] ;
  assign A_so[9] = \A_s[7] ;
  assign \A_s[7]  = A_s[7];
  assign A_nso[8] = \A_s[6] ;
  assign A_so[8] = \A_s[6] ;
  assign \A_s[6]  = A_s[6];
  assign A_nso[7] = \A_s[5] ;
  assign A_so[7] = \A_s[5] ;
  assign \A_s[5]  = A_s[5];
  assign A_nso[6] = \A_s[4] ;
  assign A_so[6] = \A_s[4] ;
  assign \A_s[4]  = A_s[4];
  assign A_nso[5] = \A_s[3] ;
  assign A_so[5] = \A_s[3] ;
  assign \A_s[3]  = A_s[3];
  assign A_nso[4] = \A_s[2] ;
  assign A_so[4] = \A_s[2] ;
  assign \A_s[2]  = A_s[2];
  assign A_nso[3] = \A_s[1] ;
  assign A_so[3] = \A_s[1] ;
  assign \A_s[1]  = A_s[1];
  assign A_nso[2] = \A_s[0] ;
  assign A_so[2] = \A_s[0] ;
  assign \A_s[0]  = A_s[0];

  AND3_X1 U2 ( .A1(B[20]), .A2(n585), .A3(B[19]), .ZN(n391) );
  INV_X4 U3 ( .A(n391), .ZN(n392) );
  INV_X4 U4 ( .A(n552), .ZN(n398) );
  OR3_X4 U5 ( .A1(B[19]), .A2(B[20]), .A3(n585), .ZN(n393) );
  INV_X4 U6 ( .A(n553), .ZN(n397) );
  OAI221_X1 U7 ( .B1(n393), .B2(n394), .C1(n392), .C2(n395), .A(n396), .ZN(
        O[9]) );
  AOI22_X1 U8 ( .A1(A_ns[8]), .A2(n397), .B1(\A_s[8] ), .B2(n398), .ZN(n396)
         );
  INV_X1 U9 ( .A(\A_s[7] ), .ZN(n395) );
  INV_X1 U10 ( .A(A_ns[7]), .ZN(n394) );
  OAI221_X1 U11 ( .B1(n393), .B2(n399), .C1(n392), .C2(n400), .A(n401), .ZN(
        O[8]) );
  AOI22_X1 U12 ( .A1(A_ns[7]), .A2(n397), .B1(\A_s[7] ), .B2(n398), .ZN(n401)
         );
  INV_X1 U13 ( .A(\A_s[6] ), .ZN(n400) );
  INV_X1 U14 ( .A(A_ns[6]), .ZN(n399) );
  OAI221_X1 U15 ( .B1(n393), .B2(n402), .C1(n392), .C2(n403), .A(n404), .ZN(
        O[7]) );
  AOI22_X1 U16 ( .A1(A_ns[6]), .A2(n397), .B1(\A_s[6] ), .B2(n398), .ZN(n404)
         );
  INV_X1 U17 ( .A(\A_s[5] ), .ZN(n403) );
  INV_X1 U18 ( .A(A_ns[5]), .ZN(n402) );
  OAI221_X1 U19 ( .B1(n393), .B2(n405), .C1(n392), .C2(n406), .A(n407), .ZN(
        O[6]) );
  AOI22_X1 U20 ( .A1(A_ns[5]), .A2(n397), .B1(\A_s[5] ), .B2(n398), .ZN(n407)
         );
  INV_X1 U21 ( .A(\A_s[4] ), .ZN(n406) );
  INV_X1 U22 ( .A(A_ns[4]), .ZN(n405) );
  OAI221_X1 U23 ( .B1(n393), .B2(n408), .C1(n392), .C2(n409), .A(n410), .ZN(
        O[63]) );
  AOI22_X1 U24 ( .A1(A_ns[62]), .A2(n397), .B1(A_s[62]), .B2(n398), .ZN(n410)
         );
  INV_X1 U25 ( .A(\A_s[61] ), .ZN(n409) );
  INV_X1 U26 ( .A(A_ns[61]), .ZN(n408) );
  OAI221_X1 U27 ( .B1(n393), .B2(n411), .C1(n392), .C2(n412), .A(n413), .ZN(
        O[62]) );
  AOI22_X1 U28 ( .A1(A_ns[61]), .A2(n397), .B1(\A_s[61] ), .B2(n398), .ZN(n413) );
  INV_X1 U29 ( .A(\A_s[60] ), .ZN(n412) );
  INV_X1 U30 ( .A(A_ns[60]), .ZN(n411) );
  OAI221_X1 U31 ( .B1(n393), .B2(n414), .C1(n392), .C2(n415), .A(n416), .ZN(
        O[61]) );
  AOI22_X1 U32 ( .A1(A_ns[60]), .A2(n397), .B1(\A_s[60] ), .B2(n398), .ZN(n416) );
  INV_X1 U33 ( .A(\A_s[59] ), .ZN(n415) );
  INV_X1 U34 ( .A(A_ns[59]), .ZN(n414) );
  OAI221_X1 U35 ( .B1(n393), .B2(n417), .C1(n392), .C2(n418), .A(n419), .ZN(
        O[60]) );
  AOI22_X1 U36 ( .A1(A_ns[59]), .A2(n397), .B1(\A_s[59] ), .B2(n398), .ZN(n419) );
  INV_X1 U37 ( .A(\A_s[58] ), .ZN(n418) );
  INV_X1 U38 ( .A(A_ns[58]), .ZN(n417) );
  OAI221_X1 U39 ( .B1(n393), .B2(n420), .C1(n392), .C2(n421), .A(n422), .ZN(
        O[5]) );
  AOI22_X1 U40 ( .A1(A_ns[4]), .A2(n397), .B1(\A_s[4] ), .B2(n398), .ZN(n422)
         );
  INV_X1 U41 ( .A(\A_s[3] ), .ZN(n421) );
  INV_X1 U42 ( .A(A_ns[3]), .ZN(n420) );
  OAI221_X1 U43 ( .B1(n393), .B2(n423), .C1(n392), .C2(n424), .A(n425), .ZN(
        O[59]) );
  AOI22_X1 U44 ( .A1(A_ns[58]), .A2(n397), .B1(\A_s[58] ), .B2(n398), .ZN(n425) );
  INV_X1 U45 ( .A(\A_s[57] ), .ZN(n424) );
  INV_X1 U46 ( .A(A_ns[57]), .ZN(n423) );
  OAI221_X1 U47 ( .B1(n393), .B2(n426), .C1(n392), .C2(n427), .A(n428), .ZN(
        O[58]) );
  AOI22_X1 U48 ( .A1(A_ns[57]), .A2(n397), .B1(\A_s[57] ), .B2(n398), .ZN(n428) );
  INV_X1 U49 ( .A(\A_s[56] ), .ZN(n427) );
  INV_X1 U50 ( .A(A_ns[56]), .ZN(n426) );
  OAI221_X1 U51 ( .B1(n393), .B2(n429), .C1(n392), .C2(n430), .A(n431), .ZN(
        O[57]) );
  AOI22_X1 U52 ( .A1(A_ns[56]), .A2(n397), .B1(\A_s[56] ), .B2(n398), .ZN(n431) );
  INV_X1 U53 ( .A(\A_s[55] ), .ZN(n430) );
  INV_X1 U54 ( .A(A_ns[55]), .ZN(n429) );
  OAI221_X1 U55 ( .B1(n393), .B2(n432), .C1(n392), .C2(n433), .A(n434), .ZN(
        O[56]) );
  AOI22_X1 U56 ( .A1(A_ns[55]), .A2(n397), .B1(\A_s[55] ), .B2(n398), .ZN(n434) );
  INV_X1 U57 ( .A(\A_s[54] ), .ZN(n433) );
  INV_X1 U58 ( .A(A_ns[54]), .ZN(n432) );
  OAI221_X1 U59 ( .B1(n393), .B2(n435), .C1(n392), .C2(n436), .A(n437), .ZN(
        O[55]) );
  AOI22_X1 U60 ( .A1(A_ns[54]), .A2(n397), .B1(\A_s[54] ), .B2(n398), .ZN(n437) );
  INV_X1 U61 ( .A(\A_s[53] ), .ZN(n436) );
  INV_X1 U62 ( .A(A_ns[53]), .ZN(n435) );
  OAI221_X1 U63 ( .B1(n393), .B2(n438), .C1(n392), .C2(n439), .A(n440), .ZN(
        O[54]) );
  AOI22_X1 U64 ( .A1(A_ns[53]), .A2(n397), .B1(\A_s[53] ), .B2(n398), .ZN(n440) );
  INV_X1 U65 ( .A(\A_s[52] ), .ZN(n439) );
  INV_X1 U66 ( .A(A_ns[52]), .ZN(n438) );
  OAI221_X1 U67 ( .B1(n393), .B2(n441), .C1(n392), .C2(n442), .A(n443), .ZN(
        O[53]) );
  AOI22_X1 U68 ( .A1(A_ns[52]), .A2(n397), .B1(\A_s[52] ), .B2(n398), .ZN(n443) );
  INV_X1 U69 ( .A(\A_s[51] ), .ZN(n442) );
  INV_X1 U70 ( .A(A_ns[51]), .ZN(n441) );
  OAI221_X1 U71 ( .B1(n393), .B2(n444), .C1(n392), .C2(n445), .A(n446), .ZN(
        O[52]) );
  AOI22_X1 U72 ( .A1(A_ns[51]), .A2(n397), .B1(\A_s[51] ), .B2(n398), .ZN(n446) );
  INV_X1 U73 ( .A(\A_s[50] ), .ZN(n445) );
  INV_X1 U74 ( .A(A_ns[50]), .ZN(n444) );
  OAI221_X1 U75 ( .B1(n393), .B2(n447), .C1(n392), .C2(n448), .A(n449), .ZN(
        O[51]) );
  AOI22_X1 U76 ( .A1(A_ns[50]), .A2(n397), .B1(\A_s[50] ), .B2(n398), .ZN(n449) );
  INV_X1 U77 ( .A(\A_s[49] ), .ZN(n448) );
  INV_X1 U78 ( .A(A_ns[49]), .ZN(n447) );
  OAI221_X1 U79 ( .B1(n393), .B2(n450), .C1(n392), .C2(n451), .A(n452), .ZN(
        O[50]) );
  AOI22_X1 U80 ( .A1(A_ns[49]), .A2(n397), .B1(\A_s[49] ), .B2(n398), .ZN(n452) );
  INV_X1 U81 ( .A(\A_s[48] ), .ZN(n451) );
  INV_X1 U82 ( .A(A_ns[48]), .ZN(n450) );
  OAI221_X1 U83 ( .B1(n393), .B2(n453), .C1(n392), .C2(n454), .A(n455), .ZN(
        O[4]) );
  AOI22_X1 U84 ( .A1(A_ns[3]), .A2(n397), .B1(\A_s[3] ), .B2(n398), .ZN(n455)
         );
  INV_X1 U85 ( .A(\A_s[2] ), .ZN(n454) );
  INV_X1 U86 ( .A(A_ns[2]), .ZN(n453) );
  OAI221_X1 U87 ( .B1(n393), .B2(n456), .C1(n392), .C2(n457), .A(n458), .ZN(
        O[49]) );
  AOI22_X1 U88 ( .A1(A_ns[48]), .A2(n397), .B1(\A_s[48] ), .B2(n398), .ZN(n458) );
  INV_X1 U89 ( .A(\A_s[47] ), .ZN(n457) );
  INV_X1 U90 ( .A(A_ns[47]), .ZN(n456) );
  OAI221_X1 U91 ( .B1(n393), .B2(n459), .C1(n392), .C2(n460), .A(n461), .ZN(
        O[48]) );
  AOI22_X1 U92 ( .A1(A_ns[47]), .A2(n397), .B1(\A_s[47] ), .B2(n398), .ZN(n461) );
  INV_X1 U93 ( .A(\A_s[46] ), .ZN(n460) );
  INV_X1 U94 ( .A(A_ns[46]), .ZN(n459) );
  OAI221_X1 U95 ( .B1(n393), .B2(n462), .C1(n392), .C2(n463), .A(n464), .ZN(
        O[47]) );
  AOI22_X1 U96 ( .A1(A_ns[46]), .A2(n397), .B1(\A_s[46] ), .B2(n398), .ZN(n464) );
  INV_X1 U97 ( .A(\A_s[45] ), .ZN(n463) );
  INV_X1 U98 ( .A(A_ns[45]), .ZN(n462) );
  OAI221_X1 U99 ( .B1(n393), .B2(n465), .C1(n392), .C2(n466), .A(n467), .ZN(
        O[46]) );
  AOI22_X1 U100 ( .A1(A_ns[45]), .A2(n397), .B1(\A_s[45] ), .B2(n398), .ZN(
        n467) );
  INV_X1 U101 ( .A(\A_s[44] ), .ZN(n466) );
  INV_X1 U102 ( .A(A_ns[44]), .ZN(n465) );
  OAI221_X1 U103 ( .B1(n393), .B2(n468), .C1(n392), .C2(n469), .A(n470), .ZN(
        O[45]) );
  AOI22_X1 U104 ( .A1(A_ns[44]), .A2(n397), .B1(\A_s[44] ), .B2(n398), .ZN(
        n470) );
  INV_X1 U105 ( .A(\A_s[43] ), .ZN(n469) );
  INV_X1 U106 ( .A(A_ns[43]), .ZN(n468) );
  OAI221_X1 U107 ( .B1(n393), .B2(n471), .C1(n392), .C2(n472), .A(n473), .ZN(
        O[44]) );
  AOI22_X1 U108 ( .A1(A_ns[43]), .A2(n397), .B1(\A_s[43] ), .B2(n398), .ZN(
        n473) );
  INV_X1 U109 ( .A(\A_s[42] ), .ZN(n472) );
  INV_X1 U110 ( .A(A_ns[42]), .ZN(n471) );
  OAI221_X1 U111 ( .B1(n393), .B2(n474), .C1(n392), .C2(n475), .A(n476), .ZN(
        O[43]) );
  AOI22_X1 U112 ( .A1(A_ns[42]), .A2(n397), .B1(\A_s[42] ), .B2(n398), .ZN(
        n476) );
  INV_X1 U113 ( .A(\A_s[41] ), .ZN(n475) );
  INV_X1 U114 ( .A(A_ns[41]), .ZN(n474) );
  OAI221_X1 U115 ( .B1(n393), .B2(n477), .C1(n392), .C2(n478), .A(n479), .ZN(
        O[42]) );
  AOI22_X1 U116 ( .A1(A_ns[41]), .A2(n397), .B1(\A_s[41] ), .B2(n398), .ZN(
        n479) );
  INV_X1 U117 ( .A(\A_s[40] ), .ZN(n478) );
  INV_X1 U118 ( .A(A_ns[40]), .ZN(n477) );
  OAI221_X1 U119 ( .B1(n393), .B2(n480), .C1(n392), .C2(n481), .A(n482), .ZN(
        O[41]) );
  AOI22_X1 U120 ( .A1(A_ns[40]), .A2(n397), .B1(\A_s[40] ), .B2(n398), .ZN(
        n482) );
  INV_X1 U121 ( .A(\A_s[39] ), .ZN(n481) );
  INV_X1 U122 ( .A(A_ns[39]), .ZN(n480) );
  OAI221_X1 U123 ( .B1(n393), .B2(n483), .C1(n392), .C2(n484), .A(n485), .ZN(
        O[40]) );
  AOI22_X1 U124 ( .A1(A_ns[39]), .A2(n397), .B1(\A_s[39] ), .B2(n398), .ZN(
        n485) );
  INV_X1 U125 ( .A(\A_s[38] ), .ZN(n484) );
  INV_X1 U126 ( .A(A_ns[38]), .ZN(n483) );
  OAI221_X1 U127 ( .B1(n393), .B2(n486), .C1(n392), .C2(n487), .A(n488), .ZN(
        O[3]) );
  AOI22_X1 U128 ( .A1(A_ns[2]), .A2(n397), .B1(\A_s[2] ), .B2(n398), .ZN(n488)
         );
  INV_X1 U129 ( .A(\A_s[1] ), .ZN(n487) );
  INV_X1 U130 ( .A(A_ns[1]), .ZN(n486) );
  OAI221_X1 U131 ( .B1(n393), .B2(n489), .C1(n392), .C2(n490), .A(n491), .ZN(
        O[39]) );
  AOI22_X1 U132 ( .A1(A_ns[38]), .A2(n397), .B1(\A_s[38] ), .B2(n398), .ZN(
        n491) );
  INV_X1 U133 ( .A(\A_s[37] ), .ZN(n490) );
  INV_X1 U134 ( .A(A_ns[37]), .ZN(n489) );
  OAI221_X1 U135 ( .B1(n393), .B2(n492), .C1(n392), .C2(n493), .A(n494), .ZN(
        O[38]) );
  AOI22_X1 U136 ( .A1(A_ns[37]), .A2(n397), .B1(\A_s[37] ), .B2(n398), .ZN(
        n494) );
  INV_X1 U137 ( .A(\A_s[36] ), .ZN(n493) );
  INV_X1 U138 ( .A(A_ns[36]), .ZN(n492) );
  OAI221_X1 U139 ( .B1(n393), .B2(n495), .C1(n392), .C2(n496), .A(n497), .ZN(
        O[37]) );
  AOI22_X1 U140 ( .A1(A_ns[36]), .A2(n397), .B1(\A_s[36] ), .B2(n398), .ZN(
        n497) );
  INV_X1 U141 ( .A(\A_s[35] ), .ZN(n496) );
  INV_X1 U142 ( .A(A_ns[35]), .ZN(n495) );
  OAI221_X1 U143 ( .B1(n393), .B2(n498), .C1(n392), .C2(n499), .A(n500), .ZN(
        O[36]) );
  AOI22_X1 U144 ( .A1(A_ns[35]), .A2(n397), .B1(\A_s[35] ), .B2(n398), .ZN(
        n500) );
  INV_X1 U145 ( .A(\A_s[34] ), .ZN(n499) );
  INV_X1 U146 ( .A(A_ns[34]), .ZN(n498) );
  OAI221_X1 U147 ( .B1(n393), .B2(n501), .C1(n392), .C2(n502), .A(n503), .ZN(
        O[35]) );
  AOI22_X1 U148 ( .A1(A_ns[34]), .A2(n397), .B1(\A_s[34] ), .B2(n398), .ZN(
        n503) );
  INV_X1 U149 ( .A(\A_s[33] ), .ZN(n502) );
  INV_X1 U150 ( .A(A_ns[33]), .ZN(n501) );
  OAI221_X1 U151 ( .B1(n393), .B2(n504), .C1(n392), .C2(n505), .A(n506), .ZN(
        O[34]) );
  AOI22_X1 U152 ( .A1(A_ns[33]), .A2(n397), .B1(\A_s[33] ), .B2(n398), .ZN(
        n506) );
  INV_X1 U153 ( .A(\A_s[32] ), .ZN(n505) );
  INV_X1 U154 ( .A(A_ns[32]), .ZN(n504) );
  OAI221_X1 U155 ( .B1(n393), .B2(n507), .C1(n392), .C2(n508), .A(n509), .ZN(
        O[33]) );
  AOI22_X1 U156 ( .A1(A_ns[32]), .A2(n397), .B1(\A_s[32] ), .B2(n398), .ZN(
        n509) );
  INV_X1 U157 ( .A(\A_s[31] ), .ZN(n508) );
  INV_X1 U158 ( .A(A_ns[31]), .ZN(n507) );
  OAI221_X1 U159 ( .B1(n393), .B2(n510), .C1(n392), .C2(n511), .A(n512), .ZN(
        O[32]) );
  AOI22_X1 U160 ( .A1(A_ns[31]), .A2(n397), .B1(\A_s[31] ), .B2(n398), .ZN(
        n512) );
  INV_X1 U161 ( .A(\A_s[30] ), .ZN(n511) );
  INV_X1 U162 ( .A(A_ns[30]), .ZN(n510) );
  OAI221_X1 U163 ( .B1(n393), .B2(n513), .C1(n392), .C2(n514), .A(n515), .ZN(
        O[31]) );
  AOI22_X1 U164 ( .A1(A_ns[30]), .A2(n397), .B1(\A_s[30] ), .B2(n398), .ZN(
        n515) );
  INV_X1 U165 ( .A(\A_s[29] ), .ZN(n514) );
  INV_X1 U166 ( .A(A_ns[29]), .ZN(n513) );
  OAI221_X1 U167 ( .B1(n393), .B2(n516), .C1(n392), .C2(n517), .A(n518), .ZN(
        O[30]) );
  AOI22_X1 U168 ( .A1(A_ns[29]), .A2(n397), .B1(\A_s[29] ), .B2(n398), .ZN(
        n518) );
  INV_X1 U169 ( .A(\A_s[28] ), .ZN(n517) );
  INV_X1 U170 ( .A(A_ns[28]), .ZN(n516) );
  OAI221_X1 U171 ( .B1(n393), .B2(n519), .C1(n392), .C2(n520), .A(n521), .ZN(
        O[2]) );
  AOI22_X1 U172 ( .A1(A_ns[1]), .A2(n397), .B1(\A_s[1] ), .B2(n398), .ZN(n521)
         );
  OAI221_X1 U173 ( .B1(n393), .B2(n522), .C1(n392), .C2(n523), .A(n524), .ZN(
        O[29]) );
  AOI22_X1 U174 ( .A1(A_ns[28]), .A2(n397), .B1(\A_s[28] ), .B2(n398), .ZN(
        n524) );
  INV_X1 U175 ( .A(\A_s[27] ), .ZN(n523) );
  INV_X1 U176 ( .A(A_ns[27]), .ZN(n522) );
  OAI221_X1 U177 ( .B1(n393), .B2(n525), .C1(n392), .C2(n526), .A(n527), .ZN(
        O[28]) );
  AOI22_X1 U178 ( .A1(A_ns[27]), .A2(n397), .B1(\A_s[27] ), .B2(n398), .ZN(
        n527) );
  INV_X1 U179 ( .A(\A_s[26] ), .ZN(n526) );
  INV_X1 U180 ( .A(A_ns[26]), .ZN(n525) );
  OAI221_X1 U181 ( .B1(n393), .B2(n528), .C1(n392), .C2(n529), .A(n530), .ZN(
        O[27]) );
  AOI22_X1 U182 ( .A1(A_ns[26]), .A2(n397), .B1(\A_s[26] ), .B2(n398), .ZN(
        n530) );
  INV_X1 U183 ( .A(\A_s[25] ), .ZN(n529) );
  INV_X1 U184 ( .A(A_ns[25]), .ZN(n528) );
  OAI221_X1 U185 ( .B1(n393), .B2(n531), .C1(n392), .C2(n532), .A(n533), .ZN(
        O[26]) );
  AOI22_X1 U186 ( .A1(A_ns[25]), .A2(n397), .B1(\A_s[25] ), .B2(n398), .ZN(
        n533) );
  INV_X1 U187 ( .A(\A_s[24] ), .ZN(n532) );
  INV_X1 U188 ( .A(A_ns[24]), .ZN(n531) );
  OAI221_X1 U189 ( .B1(n393), .B2(n534), .C1(n392), .C2(n535), .A(n536), .ZN(
        O[25]) );
  AOI22_X1 U190 ( .A1(A_ns[24]), .A2(n397), .B1(\A_s[24] ), .B2(n398), .ZN(
        n536) );
  INV_X1 U191 ( .A(\A_s[23] ), .ZN(n535) );
  INV_X1 U192 ( .A(A_ns[23]), .ZN(n534) );
  OAI221_X1 U193 ( .B1(n393), .B2(n537), .C1(n392), .C2(n538), .A(n539), .ZN(
        O[24]) );
  AOI22_X1 U194 ( .A1(A_ns[23]), .A2(n397), .B1(\A_s[23] ), .B2(n398), .ZN(
        n539) );
  INV_X1 U195 ( .A(\A_s[22] ), .ZN(n538) );
  INV_X1 U196 ( .A(A_ns[22]), .ZN(n537) );
  OAI221_X1 U197 ( .B1(n393), .B2(n540), .C1(n392), .C2(n541), .A(n542), .ZN(
        O[23]) );
  AOI22_X1 U198 ( .A1(A_ns[22]), .A2(n397), .B1(\A_s[22] ), .B2(n398), .ZN(
        n542) );
  INV_X1 U199 ( .A(\A_s[21] ), .ZN(n541) );
  INV_X1 U200 ( .A(A_ns[21]), .ZN(n540) );
  OAI221_X1 U201 ( .B1(n393), .B2(n543), .C1(n392), .C2(n544), .A(n545), .ZN(
        O[22]) );
  AOI22_X1 U202 ( .A1(A_ns[21]), .A2(n397), .B1(\A_s[21] ), .B2(n398), .ZN(
        n545) );
  INV_X1 U203 ( .A(\A_s[20] ), .ZN(n544) );
  INV_X1 U204 ( .A(A_ns[20]), .ZN(n543) );
  OAI221_X1 U205 ( .B1(n393), .B2(n546), .C1(n392), .C2(n547), .A(n548), .ZN(
        O[21]) );
  AOI22_X1 U206 ( .A1(A_ns[20]), .A2(n397), .B1(\A_s[20] ), .B2(n398), .ZN(
        n548) );
  INV_X1 U207 ( .A(\A_s[19] ), .ZN(n547) );
  INV_X1 U208 ( .A(A_ns[19]), .ZN(n546) );
  OAI221_X1 U209 ( .B1(n393), .B2(n549), .C1(n392), .C2(n550), .A(n551), .ZN(
        O[20]) );
  AOI22_X1 U210 ( .A1(A_ns[19]), .A2(n397), .B1(\A_s[19] ), .B2(n398), .ZN(
        n551) );
  INV_X1 U211 ( .A(\A_s[18] ), .ZN(n550) );
  INV_X1 U212 ( .A(A_ns[18]), .ZN(n549) );
  OAI22_X1 U213 ( .A1(n552), .A2(n520), .B1(n553), .B2(n519), .ZN(O[1]) );
  INV_X1 U214 ( .A(A_ns[0]), .ZN(n519) );
  INV_X1 U215 ( .A(\A_s[0] ), .ZN(n520) );
  OAI221_X1 U216 ( .B1(n393), .B2(n554), .C1(n392), .C2(n555), .A(n556), .ZN(
        O[19]) );
  AOI22_X1 U217 ( .A1(A_ns[18]), .A2(n397), .B1(\A_s[18] ), .B2(n398), .ZN(
        n556) );
  INV_X1 U218 ( .A(\A_s[17] ), .ZN(n555) );
  INV_X1 U219 ( .A(A_ns[17]), .ZN(n554) );
  OAI221_X1 U220 ( .B1(n393), .B2(n557), .C1(n392), .C2(n558), .A(n559), .ZN(
        O[18]) );
  AOI22_X1 U221 ( .A1(A_ns[17]), .A2(n397), .B1(\A_s[17] ), .B2(n398), .ZN(
        n559) );
  INV_X1 U222 ( .A(\A_s[16] ), .ZN(n558) );
  INV_X1 U223 ( .A(A_ns[16]), .ZN(n557) );
  OAI221_X1 U224 ( .B1(n393), .B2(n560), .C1(n392), .C2(n561), .A(n562), .ZN(
        O[17]) );
  AOI22_X1 U225 ( .A1(A_ns[16]), .A2(n397), .B1(\A_s[16] ), .B2(n398), .ZN(
        n562) );
  INV_X1 U226 ( .A(\A_s[15] ), .ZN(n561) );
  INV_X1 U227 ( .A(A_ns[15]), .ZN(n560) );
  OAI221_X1 U228 ( .B1(n393), .B2(n563), .C1(n392), .C2(n564), .A(n565), .ZN(
        O[16]) );
  AOI22_X1 U229 ( .A1(A_ns[15]), .A2(n397), .B1(\A_s[15] ), .B2(n398), .ZN(
        n565) );
  INV_X1 U230 ( .A(\A_s[14] ), .ZN(n564) );
  INV_X1 U231 ( .A(A_ns[14]), .ZN(n563) );
  OAI221_X1 U232 ( .B1(n393), .B2(n566), .C1(n392), .C2(n567), .A(n568), .ZN(
        O[15]) );
  AOI22_X1 U233 ( .A1(A_ns[14]), .A2(n397), .B1(\A_s[14] ), .B2(n398), .ZN(
        n568) );
  INV_X1 U234 ( .A(\A_s[13] ), .ZN(n567) );
  INV_X1 U235 ( .A(A_ns[13]), .ZN(n566) );
  OAI221_X1 U236 ( .B1(n393), .B2(n569), .C1(n392), .C2(n570), .A(n571), .ZN(
        O[14]) );
  AOI22_X1 U237 ( .A1(A_ns[13]), .A2(n397), .B1(\A_s[13] ), .B2(n398), .ZN(
        n571) );
  INV_X1 U238 ( .A(\A_s[12] ), .ZN(n570) );
  INV_X1 U239 ( .A(A_ns[12]), .ZN(n569) );
  OAI221_X1 U240 ( .B1(n393), .B2(n572), .C1(n392), .C2(n573), .A(n574), .ZN(
        O[13]) );
  AOI22_X1 U241 ( .A1(A_ns[12]), .A2(n397), .B1(\A_s[12] ), .B2(n398), .ZN(
        n574) );
  INV_X1 U242 ( .A(\A_s[11] ), .ZN(n573) );
  INV_X1 U243 ( .A(A_ns[11]), .ZN(n572) );
  OAI221_X1 U244 ( .B1(n393), .B2(n575), .C1(n392), .C2(n576), .A(n577), .ZN(
        O[12]) );
  AOI22_X1 U245 ( .A1(A_ns[11]), .A2(n397), .B1(\A_s[11] ), .B2(n398), .ZN(
        n577) );
  INV_X1 U246 ( .A(\A_s[10] ), .ZN(n576) );
  INV_X1 U247 ( .A(A_ns[10]), .ZN(n575) );
  OAI221_X1 U248 ( .B1(n393), .B2(n578), .C1(n392), .C2(n579), .A(n580), .ZN(
        O[11]) );
  AOI22_X1 U249 ( .A1(A_ns[10]), .A2(n397), .B1(\A_s[10] ), .B2(n398), .ZN(
        n580) );
  INV_X1 U250 ( .A(\A_s[9] ), .ZN(n579) );
  INV_X1 U251 ( .A(A_ns[9]), .ZN(n578) );
  OAI221_X1 U252 ( .B1(n581), .B2(n393), .C1(n582), .C2(n392), .A(n583), .ZN(
        O[10]) );
  AOI22_X1 U253 ( .A1(A_ns[9]), .A2(n397), .B1(\A_s[9] ), .B2(n398), .ZN(n583)
         );
  NAND2_X1 U254 ( .A1(n584), .A2(n552), .ZN(n553) );
  NAND2_X1 U255 ( .A1(n584), .A2(n585), .ZN(n552) );
  XOR2_X1 U256 ( .A(B[19]), .B(B[20]), .Z(n584) );
  INV_X1 U257 ( .A(\A_s[8] ), .ZN(n582) );
  INV_X1 U258 ( .A(B[21]), .ZN(n585) );
  INV_X1 U259 ( .A(A_ns[8]), .ZN(n581) );
endmodule


module BOOTHENC_NBIT64_i22 ( A, A_n, A_ns, A_s, B, O, A_so, A_nso );
  input [63:0] A;
  input [63:0] A_n;
  input [63:0] A_ns;
  input [63:0] A_s;
  input [63:0] B;
  output [63:0] O;
  output [63:0] A_so;
  output [63:0] A_nso;
  wire   \A_s[61] , \A_s[60] , \A_s[59] , \A_s[58] , \A_s[57] , \A_s[56] ,
         \A_s[55] , \A_s[54] , \A_s[53] , \A_s[52] , \A_s[51] , \A_s[50] ,
         \A_s[49] , \A_s[48] , \A_s[47] , \A_s[46] , \A_s[45] , \A_s[44] ,
         \A_s[43] , \A_s[42] , \A_s[41] , \A_s[40] , \A_s[39] , \A_s[38] ,
         \A_s[37] , \A_s[36] , \A_s[35] , \A_s[34] , \A_s[33] , \A_s[32] ,
         \A_s[31] , \A_s[30] , \A_s[29] , \A_s[28] , \A_s[27] , \A_s[26] ,
         \A_s[25] , \A_s[24] , \A_s[23] , \A_s[22] , \A_s[21] , \A_s[20] ,
         \A_s[19] , \A_s[18] , \A_s[17] , \A_s[16] , \A_s[15] , \A_s[14] ,
         \A_s[13] , \A_s[12] , \A_s[11] , \A_s[10] , \A_s[9] , \A_s[8] ,
         \A_s[7] , \A_s[6] , \A_s[5] , \A_s[4] , \A_s[3] , \A_s[2] , \A_s[1] ,
         \A_s[0] , n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585;
  assign A_nso[0] = 1'b0;
  assign A_nso[1] = 1'b0;
  assign A_so[0] = 1'b0;
  assign A_so[1] = 1'b0;
  assign O[0] = 1'b0;
  assign A_nso[63] = \A_s[61] ;
  assign A_so[63] = \A_s[61] ;
  assign \A_s[61]  = A_s[61];
  assign A_nso[62] = \A_s[60] ;
  assign A_so[62] = \A_s[60] ;
  assign \A_s[60]  = A_s[60];
  assign A_nso[61] = \A_s[59] ;
  assign A_so[61] = \A_s[59] ;
  assign \A_s[59]  = A_s[59];
  assign A_nso[60] = \A_s[58] ;
  assign A_so[60] = \A_s[58] ;
  assign \A_s[58]  = A_s[58];
  assign A_nso[59] = \A_s[57] ;
  assign A_so[59] = \A_s[57] ;
  assign \A_s[57]  = A_s[57];
  assign A_nso[58] = \A_s[56] ;
  assign A_so[58] = \A_s[56] ;
  assign \A_s[56]  = A_s[56];
  assign A_nso[57] = \A_s[55] ;
  assign A_so[57] = \A_s[55] ;
  assign \A_s[55]  = A_s[55];
  assign A_nso[56] = \A_s[54] ;
  assign A_so[56] = \A_s[54] ;
  assign \A_s[54]  = A_s[54];
  assign A_nso[55] = \A_s[53] ;
  assign A_so[55] = \A_s[53] ;
  assign \A_s[53]  = A_s[53];
  assign A_nso[54] = \A_s[52] ;
  assign A_so[54] = \A_s[52] ;
  assign \A_s[52]  = A_s[52];
  assign A_nso[53] = \A_s[51] ;
  assign A_so[53] = \A_s[51] ;
  assign \A_s[51]  = A_s[51];
  assign A_nso[52] = \A_s[50] ;
  assign A_so[52] = \A_s[50] ;
  assign \A_s[50]  = A_s[50];
  assign A_nso[51] = \A_s[49] ;
  assign A_so[51] = \A_s[49] ;
  assign \A_s[49]  = A_s[49];
  assign A_nso[50] = \A_s[48] ;
  assign A_so[50] = \A_s[48] ;
  assign \A_s[48]  = A_s[48];
  assign A_nso[49] = \A_s[47] ;
  assign A_so[49] = \A_s[47] ;
  assign \A_s[47]  = A_s[47];
  assign A_nso[48] = \A_s[46] ;
  assign A_so[48] = \A_s[46] ;
  assign \A_s[46]  = A_s[46];
  assign A_nso[47] = \A_s[45] ;
  assign A_so[47] = \A_s[45] ;
  assign \A_s[45]  = A_s[45];
  assign A_nso[46] = \A_s[44] ;
  assign A_so[46] = \A_s[44] ;
  assign \A_s[44]  = A_s[44];
  assign A_nso[45] = \A_s[43] ;
  assign A_so[45] = \A_s[43] ;
  assign \A_s[43]  = A_s[43];
  assign A_nso[44] = \A_s[42] ;
  assign A_so[44] = \A_s[42] ;
  assign \A_s[42]  = A_s[42];
  assign A_nso[43] = \A_s[41] ;
  assign A_so[43] = \A_s[41] ;
  assign \A_s[41]  = A_s[41];
  assign A_nso[42] = \A_s[40] ;
  assign A_so[42] = \A_s[40] ;
  assign \A_s[40]  = A_s[40];
  assign A_nso[41] = \A_s[39] ;
  assign A_so[41] = \A_s[39] ;
  assign \A_s[39]  = A_s[39];
  assign A_nso[40] = \A_s[38] ;
  assign A_so[40] = \A_s[38] ;
  assign \A_s[38]  = A_s[38];
  assign A_nso[39] = \A_s[37] ;
  assign A_so[39] = \A_s[37] ;
  assign \A_s[37]  = A_s[37];
  assign A_nso[38] = \A_s[36] ;
  assign A_so[38] = \A_s[36] ;
  assign \A_s[36]  = A_s[36];
  assign A_nso[37] = \A_s[35] ;
  assign A_so[37] = \A_s[35] ;
  assign \A_s[35]  = A_s[35];
  assign A_nso[36] = \A_s[34] ;
  assign A_so[36] = \A_s[34] ;
  assign \A_s[34]  = A_s[34];
  assign A_nso[35] = \A_s[33] ;
  assign A_so[35] = \A_s[33] ;
  assign \A_s[33]  = A_s[33];
  assign A_nso[34] = \A_s[32] ;
  assign A_so[34] = \A_s[32] ;
  assign \A_s[32]  = A_s[32];
  assign A_nso[33] = \A_s[31] ;
  assign A_so[33] = \A_s[31] ;
  assign \A_s[31]  = A_s[31];
  assign A_nso[32] = \A_s[30] ;
  assign A_so[32] = \A_s[30] ;
  assign \A_s[30]  = A_s[30];
  assign A_nso[31] = \A_s[29] ;
  assign A_so[31] = \A_s[29] ;
  assign \A_s[29]  = A_s[29];
  assign A_nso[30] = \A_s[28] ;
  assign A_so[30] = \A_s[28] ;
  assign \A_s[28]  = A_s[28];
  assign A_nso[29] = \A_s[27] ;
  assign A_so[29] = \A_s[27] ;
  assign \A_s[27]  = A_s[27];
  assign A_nso[28] = \A_s[26] ;
  assign A_so[28] = \A_s[26] ;
  assign \A_s[26]  = A_s[26];
  assign A_nso[27] = \A_s[25] ;
  assign A_so[27] = \A_s[25] ;
  assign \A_s[25]  = A_s[25];
  assign A_nso[26] = \A_s[24] ;
  assign A_so[26] = \A_s[24] ;
  assign \A_s[24]  = A_s[24];
  assign A_nso[25] = \A_s[23] ;
  assign A_so[25] = \A_s[23] ;
  assign \A_s[23]  = A_s[23];
  assign A_nso[24] = \A_s[22] ;
  assign A_so[24] = \A_s[22] ;
  assign \A_s[22]  = A_s[22];
  assign A_nso[23] = \A_s[21] ;
  assign A_so[23] = \A_s[21] ;
  assign \A_s[21]  = A_s[21];
  assign A_nso[22] = \A_s[20] ;
  assign A_so[22] = \A_s[20] ;
  assign \A_s[20]  = A_s[20];
  assign A_nso[21] = \A_s[19] ;
  assign A_so[21] = \A_s[19] ;
  assign \A_s[19]  = A_s[19];
  assign A_nso[20] = \A_s[18] ;
  assign A_so[20] = \A_s[18] ;
  assign \A_s[18]  = A_s[18];
  assign A_nso[19] = \A_s[17] ;
  assign A_so[19] = \A_s[17] ;
  assign \A_s[17]  = A_s[17];
  assign A_nso[18] = \A_s[16] ;
  assign A_so[18] = \A_s[16] ;
  assign \A_s[16]  = A_s[16];
  assign A_nso[17] = \A_s[15] ;
  assign A_so[17] = \A_s[15] ;
  assign \A_s[15]  = A_s[15];
  assign A_nso[16] = \A_s[14] ;
  assign A_so[16] = \A_s[14] ;
  assign \A_s[14]  = A_s[14];
  assign A_nso[15] = \A_s[13] ;
  assign A_so[15] = \A_s[13] ;
  assign \A_s[13]  = A_s[13];
  assign A_nso[14] = \A_s[12] ;
  assign A_so[14] = \A_s[12] ;
  assign \A_s[12]  = A_s[12];
  assign A_nso[13] = \A_s[11] ;
  assign A_so[13] = \A_s[11] ;
  assign \A_s[11]  = A_s[11];
  assign A_nso[12] = \A_s[10] ;
  assign A_so[12] = \A_s[10] ;
  assign \A_s[10]  = A_s[10];
  assign A_nso[11] = \A_s[9] ;
  assign A_so[11] = \A_s[9] ;
  assign \A_s[9]  = A_s[9];
  assign A_nso[10] = \A_s[8] ;
  assign A_so[10] = \A_s[8] ;
  assign \A_s[8]  = A_s[8];
  assign A_nso[9] = \A_s[7] ;
  assign A_so[9] = \A_s[7] ;
  assign \A_s[7]  = A_s[7];
  assign A_nso[8] = \A_s[6] ;
  assign A_so[8] = \A_s[6] ;
  assign \A_s[6]  = A_s[6];
  assign A_nso[7] = \A_s[5] ;
  assign A_so[7] = \A_s[5] ;
  assign \A_s[5]  = A_s[5];
  assign A_nso[6] = \A_s[4] ;
  assign A_so[6] = \A_s[4] ;
  assign \A_s[4]  = A_s[4];
  assign A_nso[5] = \A_s[3] ;
  assign A_so[5] = \A_s[3] ;
  assign \A_s[3]  = A_s[3];
  assign A_nso[4] = \A_s[2] ;
  assign A_so[4] = \A_s[2] ;
  assign \A_s[2]  = A_s[2];
  assign A_nso[3] = \A_s[1] ;
  assign A_so[3] = \A_s[1] ;
  assign \A_s[1]  = A_s[1];
  assign A_nso[2] = \A_s[0] ;
  assign A_so[2] = \A_s[0] ;
  assign \A_s[0]  = A_s[0];

  AND3_X1 U2 ( .A1(B[22]), .A2(n585), .A3(B[21]), .ZN(n391) );
  INV_X4 U3 ( .A(n391), .ZN(n392) );
  INV_X4 U4 ( .A(n552), .ZN(n398) );
  OR3_X4 U5 ( .A1(B[21]), .A2(B[22]), .A3(n585), .ZN(n393) );
  INV_X4 U6 ( .A(n553), .ZN(n397) );
  OAI221_X1 U7 ( .B1(n393), .B2(n394), .C1(n392), .C2(n395), .A(n396), .ZN(
        O[9]) );
  AOI22_X1 U8 ( .A1(A_ns[8]), .A2(n397), .B1(\A_s[8] ), .B2(n398), .ZN(n396)
         );
  INV_X1 U9 ( .A(\A_s[7] ), .ZN(n395) );
  INV_X1 U10 ( .A(A_ns[7]), .ZN(n394) );
  OAI221_X1 U11 ( .B1(n393), .B2(n399), .C1(n392), .C2(n400), .A(n401), .ZN(
        O[8]) );
  AOI22_X1 U12 ( .A1(A_ns[7]), .A2(n397), .B1(\A_s[7] ), .B2(n398), .ZN(n401)
         );
  INV_X1 U13 ( .A(\A_s[6] ), .ZN(n400) );
  INV_X1 U14 ( .A(A_ns[6]), .ZN(n399) );
  OAI221_X1 U15 ( .B1(n393), .B2(n402), .C1(n392), .C2(n403), .A(n404), .ZN(
        O[7]) );
  AOI22_X1 U16 ( .A1(A_ns[6]), .A2(n397), .B1(\A_s[6] ), .B2(n398), .ZN(n404)
         );
  INV_X1 U17 ( .A(\A_s[5] ), .ZN(n403) );
  INV_X1 U18 ( .A(A_ns[5]), .ZN(n402) );
  OAI221_X1 U19 ( .B1(n393), .B2(n405), .C1(n392), .C2(n406), .A(n407), .ZN(
        O[6]) );
  AOI22_X1 U20 ( .A1(A_ns[5]), .A2(n397), .B1(\A_s[5] ), .B2(n398), .ZN(n407)
         );
  INV_X1 U21 ( .A(\A_s[4] ), .ZN(n406) );
  INV_X1 U22 ( .A(A_ns[4]), .ZN(n405) );
  OAI221_X1 U23 ( .B1(n393), .B2(n408), .C1(n392), .C2(n409), .A(n410), .ZN(
        O[63]) );
  AOI22_X1 U24 ( .A1(A_ns[62]), .A2(n397), .B1(A_s[62]), .B2(n398), .ZN(n410)
         );
  INV_X1 U25 ( .A(\A_s[61] ), .ZN(n409) );
  INV_X1 U26 ( .A(A_ns[61]), .ZN(n408) );
  OAI221_X1 U27 ( .B1(n393), .B2(n411), .C1(n392), .C2(n412), .A(n413), .ZN(
        O[62]) );
  AOI22_X1 U28 ( .A1(A_ns[61]), .A2(n397), .B1(\A_s[61] ), .B2(n398), .ZN(n413) );
  INV_X1 U29 ( .A(\A_s[60] ), .ZN(n412) );
  INV_X1 U30 ( .A(A_ns[60]), .ZN(n411) );
  OAI221_X1 U31 ( .B1(n393), .B2(n414), .C1(n392), .C2(n415), .A(n416), .ZN(
        O[61]) );
  AOI22_X1 U32 ( .A1(A_ns[60]), .A2(n397), .B1(\A_s[60] ), .B2(n398), .ZN(n416) );
  INV_X1 U33 ( .A(\A_s[59] ), .ZN(n415) );
  INV_X1 U34 ( .A(A_ns[59]), .ZN(n414) );
  OAI221_X1 U35 ( .B1(n393), .B2(n417), .C1(n392), .C2(n418), .A(n419), .ZN(
        O[60]) );
  AOI22_X1 U36 ( .A1(A_ns[59]), .A2(n397), .B1(\A_s[59] ), .B2(n398), .ZN(n419) );
  INV_X1 U37 ( .A(\A_s[58] ), .ZN(n418) );
  INV_X1 U38 ( .A(A_ns[58]), .ZN(n417) );
  OAI221_X1 U39 ( .B1(n393), .B2(n420), .C1(n392), .C2(n421), .A(n422), .ZN(
        O[5]) );
  AOI22_X1 U40 ( .A1(A_ns[4]), .A2(n397), .B1(\A_s[4] ), .B2(n398), .ZN(n422)
         );
  INV_X1 U41 ( .A(\A_s[3] ), .ZN(n421) );
  INV_X1 U42 ( .A(A_ns[3]), .ZN(n420) );
  OAI221_X1 U43 ( .B1(n393), .B2(n423), .C1(n392), .C2(n424), .A(n425), .ZN(
        O[59]) );
  AOI22_X1 U44 ( .A1(A_ns[58]), .A2(n397), .B1(\A_s[58] ), .B2(n398), .ZN(n425) );
  INV_X1 U45 ( .A(\A_s[57] ), .ZN(n424) );
  INV_X1 U46 ( .A(A_ns[57]), .ZN(n423) );
  OAI221_X1 U47 ( .B1(n393), .B2(n426), .C1(n392), .C2(n427), .A(n428), .ZN(
        O[58]) );
  AOI22_X1 U48 ( .A1(A_ns[57]), .A2(n397), .B1(\A_s[57] ), .B2(n398), .ZN(n428) );
  INV_X1 U49 ( .A(\A_s[56] ), .ZN(n427) );
  INV_X1 U50 ( .A(A_ns[56]), .ZN(n426) );
  OAI221_X1 U51 ( .B1(n393), .B2(n429), .C1(n392), .C2(n430), .A(n431), .ZN(
        O[57]) );
  AOI22_X1 U52 ( .A1(A_ns[56]), .A2(n397), .B1(\A_s[56] ), .B2(n398), .ZN(n431) );
  INV_X1 U53 ( .A(\A_s[55] ), .ZN(n430) );
  INV_X1 U54 ( .A(A_ns[55]), .ZN(n429) );
  OAI221_X1 U55 ( .B1(n393), .B2(n432), .C1(n392), .C2(n433), .A(n434), .ZN(
        O[56]) );
  AOI22_X1 U56 ( .A1(A_ns[55]), .A2(n397), .B1(\A_s[55] ), .B2(n398), .ZN(n434) );
  INV_X1 U57 ( .A(\A_s[54] ), .ZN(n433) );
  INV_X1 U58 ( .A(A_ns[54]), .ZN(n432) );
  OAI221_X1 U59 ( .B1(n393), .B2(n435), .C1(n392), .C2(n436), .A(n437), .ZN(
        O[55]) );
  AOI22_X1 U60 ( .A1(A_ns[54]), .A2(n397), .B1(\A_s[54] ), .B2(n398), .ZN(n437) );
  INV_X1 U61 ( .A(\A_s[53] ), .ZN(n436) );
  INV_X1 U62 ( .A(A_ns[53]), .ZN(n435) );
  OAI221_X1 U63 ( .B1(n393), .B2(n438), .C1(n392), .C2(n439), .A(n440), .ZN(
        O[54]) );
  AOI22_X1 U64 ( .A1(A_ns[53]), .A2(n397), .B1(\A_s[53] ), .B2(n398), .ZN(n440) );
  INV_X1 U65 ( .A(\A_s[52] ), .ZN(n439) );
  INV_X1 U66 ( .A(A_ns[52]), .ZN(n438) );
  OAI221_X1 U67 ( .B1(n393), .B2(n441), .C1(n392), .C2(n442), .A(n443), .ZN(
        O[53]) );
  AOI22_X1 U68 ( .A1(A_ns[52]), .A2(n397), .B1(\A_s[52] ), .B2(n398), .ZN(n443) );
  INV_X1 U69 ( .A(\A_s[51] ), .ZN(n442) );
  INV_X1 U70 ( .A(A_ns[51]), .ZN(n441) );
  OAI221_X1 U71 ( .B1(n393), .B2(n444), .C1(n392), .C2(n445), .A(n446), .ZN(
        O[52]) );
  AOI22_X1 U72 ( .A1(A_ns[51]), .A2(n397), .B1(\A_s[51] ), .B2(n398), .ZN(n446) );
  INV_X1 U73 ( .A(\A_s[50] ), .ZN(n445) );
  INV_X1 U74 ( .A(A_ns[50]), .ZN(n444) );
  OAI221_X1 U75 ( .B1(n393), .B2(n447), .C1(n392), .C2(n448), .A(n449), .ZN(
        O[51]) );
  AOI22_X1 U76 ( .A1(A_ns[50]), .A2(n397), .B1(\A_s[50] ), .B2(n398), .ZN(n449) );
  INV_X1 U77 ( .A(\A_s[49] ), .ZN(n448) );
  INV_X1 U78 ( .A(A_ns[49]), .ZN(n447) );
  OAI221_X1 U79 ( .B1(n393), .B2(n450), .C1(n392), .C2(n451), .A(n452), .ZN(
        O[50]) );
  AOI22_X1 U80 ( .A1(A_ns[49]), .A2(n397), .B1(\A_s[49] ), .B2(n398), .ZN(n452) );
  INV_X1 U81 ( .A(\A_s[48] ), .ZN(n451) );
  INV_X1 U82 ( .A(A_ns[48]), .ZN(n450) );
  OAI221_X1 U83 ( .B1(n393), .B2(n453), .C1(n392), .C2(n454), .A(n455), .ZN(
        O[4]) );
  AOI22_X1 U84 ( .A1(A_ns[3]), .A2(n397), .B1(\A_s[3] ), .B2(n398), .ZN(n455)
         );
  INV_X1 U85 ( .A(\A_s[2] ), .ZN(n454) );
  INV_X1 U86 ( .A(A_ns[2]), .ZN(n453) );
  OAI221_X1 U87 ( .B1(n393), .B2(n456), .C1(n392), .C2(n457), .A(n458), .ZN(
        O[49]) );
  AOI22_X1 U88 ( .A1(A_ns[48]), .A2(n397), .B1(\A_s[48] ), .B2(n398), .ZN(n458) );
  INV_X1 U89 ( .A(\A_s[47] ), .ZN(n457) );
  INV_X1 U90 ( .A(A_ns[47]), .ZN(n456) );
  OAI221_X1 U91 ( .B1(n393), .B2(n459), .C1(n392), .C2(n460), .A(n461), .ZN(
        O[48]) );
  AOI22_X1 U92 ( .A1(A_ns[47]), .A2(n397), .B1(\A_s[47] ), .B2(n398), .ZN(n461) );
  INV_X1 U93 ( .A(\A_s[46] ), .ZN(n460) );
  INV_X1 U94 ( .A(A_ns[46]), .ZN(n459) );
  OAI221_X1 U95 ( .B1(n393), .B2(n462), .C1(n392), .C2(n463), .A(n464), .ZN(
        O[47]) );
  AOI22_X1 U96 ( .A1(A_ns[46]), .A2(n397), .B1(\A_s[46] ), .B2(n398), .ZN(n464) );
  INV_X1 U97 ( .A(\A_s[45] ), .ZN(n463) );
  INV_X1 U98 ( .A(A_ns[45]), .ZN(n462) );
  OAI221_X1 U99 ( .B1(n393), .B2(n465), .C1(n392), .C2(n466), .A(n467), .ZN(
        O[46]) );
  AOI22_X1 U100 ( .A1(A_ns[45]), .A2(n397), .B1(\A_s[45] ), .B2(n398), .ZN(
        n467) );
  INV_X1 U101 ( .A(\A_s[44] ), .ZN(n466) );
  INV_X1 U102 ( .A(A_ns[44]), .ZN(n465) );
  OAI221_X1 U103 ( .B1(n393), .B2(n468), .C1(n392), .C2(n469), .A(n470), .ZN(
        O[45]) );
  AOI22_X1 U104 ( .A1(A_ns[44]), .A2(n397), .B1(\A_s[44] ), .B2(n398), .ZN(
        n470) );
  INV_X1 U105 ( .A(\A_s[43] ), .ZN(n469) );
  INV_X1 U106 ( .A(A_ns[43]), .ZN(n468) );
  OAI221_X1 U107 ( .B1(n393), .B2(n471), .C1(n392), .C2(n472), .A(n473), .ZN(
        O[44]) );
  AOI22_X1 U108 ( .A1(A_ns[43]), .A2(n397), .B1(\A_s[43] ), .B2(n398), .ZN(
        n473) );
  INV_X1 U109 ( .A(\A_s[42] ), .ZN(n472) );
  INV_X1 U110 ( .A(A_ns[42]), .ZN(n471) );
  OAI221_X1 U111 ( .B1(n393), .B2(n474), .C1(n392), .C2(n475), .A(n476), .ZN(
        O[43]) );
  AOI22_X1 U112 ( .A1(A_ns[42]), .A2(n397), .B1(\A_s[42] ), .B2(n398), .ZN(
        n476) );
  INV_X1 U113 ( .A(\A_s[41] ), .ZN(n475) );
  INV_X1 U114 ( .A(A_ns[41]), .ZN(n474) );
  OAI221_X1 U115 ( .B1(n393), .B2(n477), .C1(n392), .C2(n478), .A(n479), .ZN(
        O[42]) );
  AOI22_X1 U116 ( .A1(A_ns[41]), .A2(n397), .B1(\A_s[41] ), .B2(n398), .ZN(
        n479) );
  INV_X1 U117 ( .A(\A_s[40] ), .ZN(n478) );
  INV_X1 U118 ( .A(A_ns[40]), .ZN(n477) );
  OAI221_X1 U119 ( .B1(n393), .B2(n480), .C1(n392), .C2(n481), .A(n482), .ZN(
        O[41]) );
  AOI22_X1 U120 ( .A1(A_ns[40]), .A2(n397), .B1(\A_s[40] ), .B2(n398), .ZN(
        n482) );
  INV_X1 U121 ( .A(\A_s[39] ), .ZN(n481) );
  INV_X1 U122 ( .A(A_ns[39]), .ZN(n480) );
  OAI221_X1 U123 ( .B1(n393), .B2(n483), .C1(n392), .C2(n484), .A(n485), .ZN(
        O[40]) );
  AOI22_X1 U124 ( .A1(A_ns[39]), .A2(n397), .B1(\A_s[39] ), .B2(n398), .ZN(
        n485) );
  INV_X1 U125 ( .A(\A_s[38] ), .ZN(n484) );
  INV_X1 U126 ( .A(A_ns[38]), .ZN(n483) );
  OAI221_X1 U127 ( .B1(n393), .B2(n486), .C1(n392), .C2(n487), .A(n488), .ZN(
        O[3]) );
  AOI22_X1 U128 ( .A1(A_ns[2]), .A2(n397), .B1(\A_s[2] ), .B2(n398), .ZN(n488)
         );
  INV_X1 U129 ( .A(\A_s[1] ), .ZN(n487) );
  INV_X1 U130 ( .A(A_ns[1]), .ZN(n486) );
  OAI221_X1 U131 ( .B1(n393), .B2(n489), .C1(n392), .C2(n490), .A(n491), .ZN(
        O[39]) );
  AOI22_X1 U132 ( .A1(A_ns[38]), .A2(n397), .B1(\A_s[38] ), .B2(n398), .ZN(
        n491) );
  INV_X1 U133 ( .A(\A_s[37] ), .ZN(n490) );
  INV_X1 U134 ( .A(A_ns[37]), .ZN(n489) );
  OAI221_X1 U135 ( .B1(n393), .B2(n492), .C1(n392), .C2(n493), .A(n494), .ZN(
        O[38]) );
  AOI22_X1 U136 ( .A1(A_ns[37]), .A2(n397), .B1(\A_s[37] ), .B2(n398), .ZN(
        n494) );
  INV_X1 U137 ( .A(\A_s[36] ), .ZN(n493) );
  INV_X1 U138 ( .A(A_ns[36]), .ZN(n492) );
  OAI221_X1 U139 ( .B1(n393), .B2(n495), .C1(n392), .C2(n496), .A(n497), .ZN(
        O[37]) );
  AOI22_X1 U140 ( .A1(A_ns[36]), .A2(n397), .B1(\A_s[36] ), .B2(n398), .ZN(
        n497) );
  INV_X1 U141 ( .A(\A_s[35] ), .ZN(n496) );
  INV_X1 U142 ( .A(A_ns[35]), .ZN(n495) );
  OAI221_X1 U143 ( .B1(n393), .B2(n498), .C1(n392), .C2(n499), .A(n500), .ZN(
        O[36]) );
  AOI22_X1 U144 ( .A1(A_ns[35]), .A2(n397), .B1(\A_s[35] ), .B2(n398), .ZN(
        n500) );
  INV_X1 U145 ( .A(\A_s[34] ), .ZN(n499) );
  INV_X1 U146 ( .A(A_ns[34]), .ZN(n498) );
  OAI221_X1 U147 ( .B1(n393), .B2(n501), .C1(n392), .C2(n502), .A(n503), .ZN(
        O[35]) );
  AOI22_X1 U148 ( .A1(A_ns[34]), .A2(n397), .B1(\A_s[34] ), .B2(n398), .ZN(
        n503) );
  INV_X1 U149 ( .A(\A_s[33] ), .ZN(n502) );
  INV_X1 U150 ( .A(A_ns[33]), .ZN(n501) );
  OAI221_X1 U151 ( .B1(n393), .B2(n504), .C1(n392), .C2(n505), .A(n506), .ZN(
        O[34]) );
  AOI22_X1 U152 ( .A1(A_ns[33]), .A2(n397), .B1(\A_s[33] ), .B2(n398), .ZN(
        n506) );
  INV_X1 U153 ( .A(\A_s[32] ), .ZN(n505) );
  INV_X1 U154 ( .A(A_ns[32]), .ZN(n504) );
  OAI221_X1 U155 ( .B1(n393), .B2(n507), .C1(n392), .C2(n508), .A(n509), .ZN(
        O[33]) );
  AOI22_X1 U156 ( .A1(A_ns[32]), .A2(n397), .B1(\A_s[32] ), .B2(n398), .ZN(
        n509) );
  INV_X1 U157 ( .A(\A_s[31] ), .ZN(n508) );
  INV_X1 U158 ( .A(A_ns[31]), .ZN(n507) );
  OAI221_X1 U159 ( .B1(n393), .B2(n510), .C1(n392), .C2(n511), .A(n512), .ZN(
        O[32]) );
  AOI22_X1 U160 ( .A1(A_ns[31]), .A2(n397), .B1(\A_s[31] ), .B2(n398), .ZN(
        n512) );
  INV_X1 U161 ( .A(\A_s[30] ), .ZN(n511) );
  INV_X1 U162 ( .A(A_ns[30]), .ZN(n510) );
  OAI221_X1 U163 ( .B1(n393), .B2(n513), .C1(n392), .C2(n514), .A(n515), .ZN(
        O[31]) );
  AOI22_X1 U164 ( .A1(A_ns[30]), .A2(n397), .B1(\A_s[30] ), .B2(n398), .ZN(
        n515) );
  INV_X1 U165 ( .A(\A_s[29] ), .ZN(n514) );
  INV_X1 U166 ( .A(A_ns[29]), .ZN(n513) );
  OAI221_X1 U167 ( .B1(n393), .B2(n516), .C1(n392), .C2(n517), .A(n518), .ZN(
        O[30]) );
  AOI22_X1 U168 ( .A1(A_ns[29]), .A2(n397), .B1(\A_s[29] ), .B2(n398), .ZN(
        n518) );
  INV_X1 U169 ( .A(\A_s[28] ), .ZN(n517) );
  INV_X1 U170 ( .A(A_ns[28]), .ZN(n516) );
  OAI221_X1 U171 ( .B1(n393), .B2(n519), .C1(n392), .C2(n520), .A(n521), .ZN(
        O[2]) );
  AOI22_X1 U172 ( .A1(A_ns[1]), .A2(n397), .B1(\A_s[1] ), .B2(n398), .ZN(n521)
         );
  OAI221_X1 U173 ( .B1(n393), .B2(n522), .C1(n392), .C2(n523), .A(n524), .ZN(
        O[29]) );
  AOI22_X1 U174 ( .A1(A_ns[28]), .A2(n397), .B1(\A_s[28] ), .B2(n398), .ZN(
        n524) );
  INV_X1 U175 ( .A(\A_s[27] ), .ZN(n523) );
  INV_X1 U176 ( .A(A_ns[27]), .ZN(n522) );
  OAI221_X1 U177 ( .B1(n393), .B2(n525), .C1(n392), .C2(n526), .A(n527), .ZN(
        O[28]) );
  AOI22_X1 U178 ( .A1(A_ns[27]), .A2(n397), .B1(\A_s[27] ), .B2(n398), .ZN(
        n527) );
  INV_X1 U179 ( .A(\A_s[26] ), .ZN(n526) );
  INV_X1 U180 ( .A(A_ns[26]), .ZN(n525) );
  OAI221_X1 U181 ( .B1(n393), .B2(n528), .C1(n392), .C2(n529), .A(n530), .ZN(
        O[27]) );
  AOI22_X1 U182 ( .A1(A_ns[26]), .A2(n397), .B1(\A_s[26] ), .B2(n398), .ZN(
        n530) );
  INV_X1 U183 ( .A(\A_s[25] ), .ZN(n529) );
  INV_X1 U184 ( .A(A_ns[25]), .ZN(n528) );
  OAI221_X1 U185 ( .B1(n393), .B2(n531), .C1(n392), .C2(n532), .A(n533), .ZN(
        O[26]) );
  AOI22_X1 U186 ( .A1(A_ns[25]), .A2(n397), .B1(\A_s[25] ), .B2(n398), .ZN(
        n533) );
  INV_X1 U187 ( .A(\A_s[24] ), .ZN(n532) );
  INV_X1 U188 ( .A(A_ns[24]), .ZN(n531) );
  OAI221_X1 U189 ( .B1(n393), .B2(n534), .C1(n392), .C2(n535), .A(n536), .ZN(
        O[25]) );
  AOI22_X1 U190 ( .A1(A_ns[24]), .A2(n397), .B1(\A_s[24] ), .B2(n398), .ZN(
        n536) );
  INV_X1 U191 ( .A(\A_s[23] ), .ZN(n535) );
  INV_X1 U192 ( .A(A_ns[23]), .ZN(n534) );
  OAI221_X1 U193 ( .B1(n393), .B2(n537), .C1(n392), .C2(n538), .A(n539), .ZN(
        O[24]) );
  AOI22_X1 U194 ( .A1(A_ns[23]), .A2(n397), .B1(\A_s[23] ), .B2(n398), .ZN(
        n539) );
  INV_X1 U195 ( .A(\A_s[22] ), .ZN(n538) );
  INV_X1 U196 ( .A(A_ns[22]), .ZN(n537) );
  OAI221_X1 U197 ( .B1(n393), .B2(n540), .C1(n392), .C2(n541), .A(n542), .ZN(
        O[23]) );
  AOI22_X1 U198 ( .A1(A_ns[22]), .A2(n397), .B1(\A_s[22] ), .B2(n398), .ZN(
        n542) );
  INV_X1 U199 ( .A(\A_s[21] ), .ZN(n541) );
  INV_X1 U200 ( .A(A_ns[21]), .ZN(n540) );
  OAI221_X1 U201 ( .B1(n393), .B2(n543), .C1(n392), .C2(n544), .A(n545), .ZN(
        O[22]) );
  AOI22_X1 U202 ( .A1(A_ns[21]), .A2(n397), .B1(\A_s[21] ), .B2(n398), .ZN(
        n545) );
  INV_X1 U203 ( .A(\A_s[20] ), .ZN(n544) );
  INV_X1 U204 ( .A(A_ns[20]), .ZN(n543) );
  OAI221_X1 U205 ( .B1(n393), .B2(n546), .C1(n392), .C2(n547), .A(n548), .ZN(
        O[21]) );
  AOI22_X1 U206 ( .A1(A_ns[20]), .A2(n397), .B1(\A_s[20] ), .B2(n398), .ZN(
        n548) );
  INV_X1 U207 ( .A(\A_s[19] ), .ZN(n547) );
  INV_X1 U208 ( .A(A_ns[19]), .ZN(n546) );
  OAI221_X1 U209 ( .B1(n393), .B2(n549), .C1(n392), .C2(n550), .A(n551), .ZN(
        O[20]) );
  AOI22_X1 U210 ( .A1(A_ns[19]), .A2(n397), .B1(\A_s[19] ), .B2(n398), .ZN(
        n551) );
  INV_X1 U211 ( .A(\A_s[18] ), .ZN(n550) );
  INV_X1 U212 ( .A(A_ns[18]), .ZN(n549) );
  OAI22_X1 U213 ( .A1(n552), .A2(n520), .B1(n553), .B2(n519), .ZN(O[1]) );
  INV_X1 U214 ( .A(A_ns[0]), .ZN(n519) );
  INV_X1 U215 ( .A(\A_s[0] ), .ZN(n520) );
  OAI221_X1 U216 ( .B1(n393), .B2(n554), .C1(n392), .C2(n555), .A(n556), .ZN(
        O[19]) );
  AOI22_X1 U217 ( .A1(A_ns[18]), .A2(n397), .B1(\A_s[18] ), .B2(n398), .ZN(
        n556) );
  INV_X1 U218 ( .A(\A_s[17] ), .ZN(n555) );
  INV_X1 U219 ( .A(A_ns[17]), .ZN(n554) );
  OAI221_X1 U220 ( .B1(n393), .B2(n557), .C1(n392), .C2(n558), .A(n559), .ZN(
        O[18]) );
  AOI22_X1 U221 ( .A1(A_ns[17]), .A2(n397), .B1(\A_s[17] ), .B2(n398), .ZN(
        n559) );
  INV_X1 U222 ( .A(\A_s[16] ), .ZN(n558) );
  INV_X1 U223 ( .A(A_ns[16]), .ZN(n557) );
  OAI221_X1 U224 ( .B1(n393), .B2(n560), .C1(n392), .C2(n561), .A(n562), .ZN(
        O[17]) );
  AOI22_X1 U225 ( .A1(A_ns[16]), .A2(n397), .B1(\A_s[16] ), .B2(n398), .ZN(
        n562) );
  INV_X1 U226 ( .A(\A_s[15] ), .ZN(n561) );
  INV_X1 U227 ( .A(A_ns[15]), .ZN(n560) );
  OAI221_X1 U228 ( .B1(n393), .B2(n563), .C1(n392), .C2(n564), .A(n565), .ZN(
        O[16]) );
  AOI22_X1 U229 ( .A1(A_ns[15]), .A2(n397), .B1(\A_s[15] ), .B2(n398), .ZN(
        n565) );
  INV_X1 U230 ( .A(\A_s[14] ), .ZN(n564) );
  INV_X1 U231 ( .A(A_ns[14]), .ZN(n563) );
  OAI221_X1 U232 ( .B1(n393), .B2(n566), .C1(n392), .C2(n567), .A(n568), .ZN(
        O[15]) );
  AOI22_X1 U233 ( .A1(A_ns[14]), .A2(n397), .B1(\A_s[14] ), .B2(n398), .ZN(
        n568) );
  INV_X1 U234 ( .A(\A_s[13] ), .ZN(n567) );
  INV_X1 U235 ( .A(A_ns[13]), .ZN(n566) );
  OAI221_X1 U236 ( .B1(n393), .B2(n569), .C1(n392), .C2(n570), .A(n571), .ZN(
        O[14]) );
  AOI22_X1 U237 ( .A1(A_ns[13]), .A2(n397), .B1(\A_s[13] ), .B2(n398), .ZN(
        n571) );
  INV_X1 U238 ( .A(\A_s[12] ), .ZN(n570) );
  INV_X1 U239 ( .A(A_ns[12]), .ZN(n569) );
  OAI221_X1 U240 ( .B1(n393), .B2(n572), .C1(n392), .C2(n573), .A(n574), .ZN(
        O[13]) );
  AOI22_X1 U241 ( .A1(A_ns[12]), .A2(n397), .B1(\A_s[12] ), .B2(n398), .ZN(
        n574) );
  INV_X1 U242 ( .A(\A_s[11] ), .ZN(n573) );
  INV_X1 U243 ( .A(A_ns[11]), .ZN(n572) );
  OAI221_X1 U244 ( .B1(n393), .B2(n575), .C1(n392), .C2(n576), .A(n577), .ZN(
        O[12]) );
  AOI22_X1 U245 ( .A1(A_ns[11]), .A2(n397), .B1(\A_s[11] ), .B2(n398), .ZN(
        n577) );
  INV_X1 U246 ( .A(\A_s[10] ), .ZN(n576) );
  INV_X1 U247 ( .A(A_ns[10]), .ZN(n575) );
  OAI221_X1 U248 ( .B1(n393), .B2(n578), .C1(n392), .C2(n579), .A(n580), .ZN(
        O[11]) );
  AOI22_X1 U249 ( .A1(A_ns[10]), .A2(n397), .B1(\A_s[10] ), .B2(n398), .ZN(
        n580) );
  INV_X1 U250 ( .A(\A_s[9] ), .ZN(n579) );
  INV_X1 U251 ( .A(A_ns[9]), .ZN(n578) );
  OAI221_X1 U252 ( .B1(n581), .B2(n393), .C1(n582), .C2(n392), .A(n583), .ZN(
        O[10]) );
  AOI22_X1 U253 ( .A1(A_ns[9]), .A2(n397), .B1(\A_s[9] ), .B2(n398), .ZN(n583)
         );
  NAND2_X1 U254 ( .A1(n584), .A2(n552), .ZN(n553) );
  NAND2_X1 U255 ( .A1(n584), .A2(n585), .ZN(n552) );
  XOR2_X1 U256 ( .A(B[21]), .B(B[22]), .Z(n584) );
  INV_X1 U257 ( .A(\A_s[8] ), .ZN(n582) );
  INV_X1 U258 ( .A(B[23]), .ZN(n585) );
  INV_X1 U259 ( .A(A_ns[8]), .ZN(n581) );
endmodule


module BOOTHENC_NBIT64_i24 ( A, A_n, A_ns, A_s, B, O, A_so, A_nso );
  input [63:0] A;
  input [63:0] A_n;
  input [63:0] A_ns;
  input [63:0] A_s;
  input [63:0] B;
  output [63:0] O;
  output [63:0] A_so;
  output [63:0] A_nso;
  wire   \A_s[61] , \A_s[60] , \A_s[59] , \A_s[58] , \A_s[57] , \A_s[56] ,
         \A_s[55] , \A_s[54] , \A_s[53] , \A_s[52] , \A_s[51] , \A_s[50] ,
         \A_s[49] , \A_s[48] , \A_s[47] , \A_s[46] , \A_s[45] , \A_s[44] ,
         \A_s[43] , \A_s[42] , \A_s[41] , \A_s[40] , \A_s[39] , \A_s[38] ,
         \A_s[37] , \A_s[36] , \A_s[35] , \A_s[34] , \A_s[33] , \A_s[32] ,
         \A_s[31] , \A_s[30] , \A_s[29] , \A_s[28] , \A_s[27] , \A_s[26] ,
         \A_s[25] , \A_s[24] , \A_s[23] , \A_s[22] , \A_s[21] , \A_s[20] ,
         \A_s[19] , \A_s[18] , \A_s[17] , \A_s[16] , \A_s[15] , \A_s[14] ,
         \A_s[13] , \A_s[12] , \A_s[11] , \A_s[10] , \A_s[9] , \A_s[8] ,
         \A_s[7] , \A_s[6] , \A_s[5] , \A_s[4] , \A_s[3] , \A_s[2] , \A_s[1] ,
         \A_s[0] , n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585;
  assign A_nso[0] = 1'b0;
  assign A_nso[1] = 1'b0;
  assign A_so[0] = 1'b0;
  assign A_so[1] = 1'b0;
  assign O[0] = 1'b0;
  assign A_nso[63] = \A_s[61] ;
  assign A_so[63] = \A_s[61] ;
  assign \A_s[61]  = A_s[61];
  assign A_nso[62] = \A_s[60] ;
  assign A_so[62] = \A_s[60] ;
  assign \A_s[60]  = A_s[60];
  assign A_nso[61] = \A_s[59] ;
  assign A_so[61] = \A_s[59] ;
  assign \A_s[59]  = A_s[59];
  assign A_nso[60] = \A_s[58] ;
  assign A_so[60] = \A_s[58] ;
  assign \A_s[58]  = A_s[58];
  assign A_nso[59] = \A_s[57] ;
  assign A_so[59] = \A_s[57] ;
  assign \A_s[57]  = A_s[57];
  assign A_nso[58] = \A_s[56] ;
  assign A_so[58] = \A_s[56] ;
  assign \A_s[56]  = A_s[56];
  assign A_nso[57] = \A_s[55] ;
  assign A_so[57] = \A_s[55] ;
  assign \A_s[55]  = A_s[55];
  assign A_nso[56] = \A_s[54] ;
  assign A_so[56] = \A_s[54] ;
  assign \A_s[54]  = A_s[54];
  assign A_nso[55] = \A_s[53] ;
  assign A_so[55] = \A_s[53] ;
  assign \A_s[53]  = A_s[53];
  assign A_nso[54] = \A_s[52] ;
  assign A_so[54] = \A_s[52] ;
  assign \A_s[52]  = A_s[52];
  assign A_nso[53] = \A_s[51] ;
  assign A_so[53] = \A_s[51] ;
  assign \A_s[51]  = A_s[51];
  assign A_nso[52] = \A_s[50] ;
  assign A_so[52] = \A_s[50] ;
  assign \A_s[50]  = A_s[50];
  assign A_nso[51] = \A_s[49] ;
  assign A_so[51] = \A_s[49] ;
  assign \A_s[49]  = A_s[49];
  assign A_nso[50] = \A_s[48] ;
  assign A_so[50] = \A_s[48] ;
  assign \A_s[48]  = A_s[48];
  assign A_nso[49] = \A_s[47] ;
  assign A_so[49] = \A_s[47] ;
  assign \A_s[47]  = A_s[47];
  assign A_nso[48] = \A_s[46] ;
  assign A_so[48] = \A_s[46] ;
  assign \A_s[46]  = A_s[46];
  assign A_nso[47] = \A_s[45] ;
  assign A_so[47] = \A_s[45] ;
  assign \A_s[45]  = A_s[45];
  assign A_nso[46] = \A_s[44] ;
  assign A_so[46] = \A_s[44] ;
  assign \A_s[44]  = A_s[44];
  assign A_nso[45] = \A_s[43] ;
  assign A_so[45] = \A_s[43] ;
  assign \A_s[43]  = A_s[43];
  assign A_nso[44] = \A_s[42] ;
  assign A_so[44] = \A_s[42] ;
  assign \A_s[42]  = A_s[42];
  assign A_nso[43] = \A_s[41] ;
  assign A_so[43] = \A_s[41] ;
  assign \A_s[41]  = A_s[41];
  assign A_nso[42] = \A_s[40] ;
  assign A_so[42] = \A_s[40] ;
  assign \A_s[40]  = A_s[40];
  assign A_nso[41] = \A_s[39] ;
  assign A_so[41] = \A_s[39] ;
  assign \A_s[39]  = A_s[39];
  assign A_nso[40] = \A_s[38] ;
  assign A_so[40] = \A_s[38] ;
  assign \A_s[38]  = A_s[38];
  assign A_nso[39] = \A_s[37] ;
  assign A_so[39] = \A_s[37] ;
  assign \A_s[37]  = A_s[37];
  assign A_nso[38] = \A_s[36] ;
  assign A_so[38] = \A_s[36] ;
  assign \A_s[36]  = A_s[36];
  assign A_nso[37] = \A_s[35] ;
  assign A_so[37] = \A_s[35] ;
  assign \A_s[35]  = A_s[35];
  assign A_nso[36] = \A_s[34] ;
  assign A_so[36] = \A_s[34] ;
  assign \A_s[34]  = A_s[34];
  assign A_nso[35] = \A_s[33] ;
  assign A_so[35] = \A_s[33] ;
  assign \A_s[33]  = A_s[33];
  assign A_nso[34] = \A_s[32] ;
  assign A_so[34] = \A_s[32] ;
  assign \A_s[32]  = A_s[32];
  assign A_nso[33] = \A_s[31] ;
  assign A_so[33] = \A_s[31] ;
  assign \A_s[31]  = A_s[31];
  assign A_nso[32] = \A_s[30] ;
  assign A_so[32] = \A_s[30] ;
  assign \A_s[30]  = A_s[30];
  assign A_nso[31] = \A_s[29] ;
  assign A_so[31] = \A_s[29] ;
  assign \A_s[29]  = A_s[29];
  assign A_nso[30] = \A_s[28] ;
  assign A_so[30] = \A_s[28] ;
  assign \A_s[28]  = A_s[28];
  assign A_nso[29] = \A_s[27] ;
  assign A_so[29] = \A_s[27] ;
  assign \A_s[27]  = A_s[27];
  assign A_nso[28] = \A_s[26] ;
  assign A_so[28] = \A_s[26] ;
  assign \A_s[26]  = A_s[26];
  assign A_nso[27] = \A_s[25] ;
  assign A_so[27] = \A_s[25] ;
  assign \A_s[25]  = A_s[25];
  assign A_nso[26] = \A_s[24] ;
  assign A_so[26] = \A_s[24] ;
  assign \A_s[24]  = A_s[24];
  assign A_nso[25] = \A_s[23] ;
  assign A_so[25] = \A_s[23] ;
  assign \A_s[23]  = A_s[23];
  assign A_nso[24] = \A_s[22] ;
  assign A_so[24] = \A_s[22] ;
  assign \A_s[22]  = A_s[22];
  assign A_nso[23] = \A_s[21] ;
  assign A_so[23] = \A_s[21] ;
  assign \A_s[21]  = A_s[21];
  assign A_nso[22] = \A_s[20] ;
  assign A_so[22] = \A_s[20] ;
  assign \A_s[20]  = A_s[20];
  assign A_nso[21] = \A_s[19] ;
  assign A_so[21] = \A_s[19] ;
  assign \A_s[19]  = A_s[19];
  assign A_nso[20] = \A_s[18] ;
  assign A_so[20] = \A_s[18] ;
  assign \A_s[18]  = A_s[18];
  assign A_nso[19] = \A_s[17] ;
  assign A_so[19] = \A_s[17] ;
  assign \A_s[17]  = A_s[17];
  assign A_nso[18] = \A_s[16] ;
  assign A_so[18] = \A_s[16] ;
  assign \A_s[16]  = A_s[16];
  assign A_nso[17] = \A_s[15] ;
  assign A_so[17] = \A_s[15] ;
  assign \A_s[15]  = A_s[15];
  assign A_nso[16] = \A_s[14] ;
  assign A_so[16] = \A_s[14] ;
  assign \A_s[14]  = A_s[14];
  assign A_nso[15] = \A_s[13] ;
  assign A_so[15] = \A_s[13] ;
  assign \A_s[13]  = A_s[13];
  assign A_nso[14] = \A_s[12] ;
  assign A_so[14] = \A_s[12] ;
  assign \A_s[12]  = A_s[12];
  assign A_nso[13] = \A_s[11] ;
  assign A_so[13] = \A_s[11] ;
  assign \A_s[11]  = A_s[11];
  assign A_nso[12] = \A_s[10] ;
  assign A_so[12] = \A_s[10] ;
  assign \A_s[10]  = A_s[10];
  assign A_nso[11] = \A_s[9] ;
  assign A_so[11] = \A_s[9] ;
  assign \A_s[9]  = A_s[9];
  assign A_nso[10] = \A_s[8] ;
  assign A_so[10] = \A_s[8] ;
  assign \A_s[8]  = A_s[8];
  assign A_nso[9] = \A_s[7] ;
  assign A_so[9] = \A_s[7] ;
  assign \A_s[7]  = A_s[7];
  assign A_nso[8] = \A_s[6] ;
  assign A_so[8] = \A_s[6] ;
  assign \A_s[6]  = A_s[6];
  assign A_nso[7] = \A_s[5] ;
  assign A_so[7] = \A_s[5] ;
  assign \A_s[5]  = A_s[5];
  assign A_nso[6] = \A_s[4] ;
  assign A_so[6] = \A_s[4] ;
  assign \A_s[4]  = A_s[4];
  assign A_nso[5] = \A_s[3] ;
  assign A_so[5] = \A_s[3] ;
  assign \A_s[3]  = A_s[3];
  assign A_nso[4] = \A_s[2] ;
  assign A_so[4] = \A_s[2] ;
  assign \A_s[2]  = A_s[2];
  assign A_nso[3] = \A_s[1] ;
  assign A_so[3] = \A_s[1] ;
  assign \A_s[1]  = A_s[1];
  assign A_nso[2] = \A_s[0] ;
  assign A_so[2] = \A_s[0] ;
  assign \A_s[0]  = A_s[0];

  AND3_X1 U2 ( .A1(B[24]), .A2(n585), .A3(B[23]), .ZN(n391) );
  INV_X4 U3 ( .A(n391), .ZN(n392) );
  INV_X4 U4 ( .A(n552), .ZN(n398) );
  OR3_X4 U5 ( .A1(B[23]), .A2(B[24]), .A3(n585), .ZN(n393) );
  INV_X4 U6 ( .A(n553), .ZN(n397) );
  OAI221_X1 U7 ( .B1(n393), .B2(n394), .C1(n392), .C2(n395), .A(n396), .ZN(
        O[9]) );
  AOI22_X1 U8 ( .A1(A_ns[8]), .A2(n397), .B1(\A_s[8] ), .B2(n398), .ZN(n396)
         );
  INV_X1 U9 ( .A(\A_s[7] ), .ZN(n395) );
  INV_X1 U10 ( .A(A_ns[7]), .ZN(n394) );
  OAI221_X1 U11 ( .B1(n393), .B2(n399), .C1(n392), .C2(n400), .A(n401), .ZN(
        O[8]) );
  AOI22_X1 U12 ( .A1(A_ns[7]), .A2(n397), .B1(\A_s[7] ), .B2(n398), .ZN(n401)
         );
  INV_X1 U13 ( .A(\A_s[6] ), .ZN(n400) );
  INV_X1 U14 ( .A(A_ns[6]), .ZN(n399) );
  OAI221_X1 U15 ( .B1(n393), .B2(n402), .C1(n392), .C2(n403), .A(n404), .ZN(
        O[7]) );
  AOI22_X1 U16 ( .A1(A_ns[6]), .A2(n397), .B1(\A_s[6] ), .B2(n398), .ZN(n404)
         );
  INV_X1 U17 ( .A(\A_s[5] ), .ZN(n403) );
  INV_X1 U18 ( .A(A_ns[5]), .ZN(n402) );
  OAI221_X1 U19 ( .B1(n393), .B2(n405), .C1(n392), .C2(n406), .A(n407), .ZN(
        O[6]) );
  AOI22_X1 U20 ( .A1(A_ns[5]), .A2(n397), .B1(\A_s[5] ), .B2(n398), .ZN(n407)
         );
  INV_X1 U21 ( .A(\A_s[4] ), .ZN(n406) );
  INV_X1 U22 ( .A(A_ns[4]), .ZN(n405) );
  OAI221_X1 U23 ( .B1(n393), .B2(n408), .C1(n392), .C2(n409), .A(n410), .ZN(
        O[63]) );
  AOI22_X1 U24 ( .A1(A_ns[62]), .A2(n397), .B1(A_s[62]), .B2(n398), .ZN(n410)
         );
  INV_X1 U25 ( .A(\A_s[61] ), .ZN(n409) );
  INV_X1 U26 ( .A(A_ns[61]), .ZN(n408) );
  OAI221_X1 U27 ( .B1(n393), .B2(n411), .C1(n392), .C2(n412), .A(n413), .ZN(
        O[62]) );
  AOI22_X1 U28 ( .A1(A_ns[61]), .A2(n397), .B1(\A_s[61] ), .B2(n398), .ZN(n413) );
  INV_X1 U29 ( .A(\A_s[60] ), .ZN(n412) );
  INV_X1 U30 ( .A(A_ns[60]), .ZN(n411) );
  OAI221_X1 U31 ( .B1(n393), .B2(n414), .C1(n392), .C2(n415), .A(n416), .ZN(
        O[61]) );
  AOI22_X1 U32 ( .A1(A_ns[60]), .A2(n397), .B1(\A_s[60] ), .B2(n398), .ZN(n416) );
  INV_X1 U33 ( .A(\A_s[59] ), .ZN(n415) );
  INV_X1 U34 ( .A(A_ns[59]), .ZN(n414) );
  OAI221_X1 U35 ( .B1(n393), .B2(n417), .C1(n392), .C2(n418), .A(n419), .ZN(
        O[60]) );
  AOI22_X1 U36 ( .A1(A_ns[59]), .A2(n397), .B1(\A_s[59] ), .B2(n398), .ZN(n419) );
  INV_X1 U37 ( .A(\A_s[58] ), .ZN(n418) );
  INV_X1 U38 ( .A(A_ns[58]), .ZN(n417) );
  OAI221_X1 U39 ( .B1(n393), .B2(n420), .C1(n392), .C2(n421), .A(n422), .ZN(
        O[5]) );
  AOI22_X1 U40 ( .A1(A_ns[4]), .A2(n397), .B1(\A_s[4] ), .B2(n398), .ZN(n422)
         );
  INV_X1 U41 ( .A(\A_s[3] ), .ZN(n421) );
  INV_X1 U42 ( .A(A_ns[3]), .ZN(n420) );
  OAI221_X1 U43 ( .B1(n393), .B2(n423), .C1(n392), .C2(n424), .A(n425), .ZN(
        O[59]) );
  AOI22_X1 U44 ( .A1(A_ns[58]), .A2(n397), .B1(\A_s[58] ), .B2(n398), .ZN(n425) );
  INV_X1 U45 ( .A(\A_s[57] ), .ZN(n424) );
  INV_X1 U46 ( .A(A_ns[57]), .ZN(n423) );
  OAI221_X1 U47 ( .B1(n393), .B2(n426), .C1(n392), .C2(n427), .A(n428), .ZN(
        O[58]) );
  AOI22_X1 U48 ( .A1(A_ns[57]), .A2(n397), .B1(\A_s[57] ), .B2(n398), .ZN(n428) );
  INV_X1 U49 ( .A(\A_s[56] ), .ZN(n427) );
  INV_X1 U50 ( .A(A_ns[56]), .ZN(n426) );
  OAI221_X1 U51 ( .B1(n393), .B2(n429), .C1(n392), .C2(n430), .A(n431), .ZN(
        O[57]) );
  AOI22_X1 U52 ( .A1(A_ns[56]), .A2(n397), .B1(\A_s[56] ), .B2(n398), .ZN(n431) );
  INV_X1 U53 ( .A(\A_s[55] ), .ZN(n430) );
  INV_X1 U54 ( .A(A_ns[55]), .ZN(n429) );
  OAI221_X1 U55 ( .B1(n393), .B2(n432), .C1(n392), .C2(n433), .A(n434), .ZN(
        O[56]) );
  AOI22_X1 U56 ( .A1(A_ns[55]), .A2(n397), .B1(\A_s[55] ), .B2(n398), .ZN(n434) );
  INV_X1 U57 ( .A(\A_s[54] ), .ZN(n433) );
  INV_X1 U58 ( .A(A_ns[54]), .ZN(n432) );
  OAI221_X1 U59 ( .B1(n393), .B2(n435), .C1(n392), .C2(n436), .A(n437), .ZN(
        O[55]) );
  AOI22_X1 U60 ( .A1(A_ns[54]), .A2(n397), .B1(\A_s[54] ), .B2(n398), .ZN(n437) );
  INV_X1 U61 ( .A(\A_s[53] ), .ZN(n436) );
  INV_X1 U62 ( .A(A_ns[53]), .ZN(n435) );
  OAI221_X1 U63 ( .B1(n393), .B2(n438), .C1(n392), .C2(n439), .A(n440), .ZN(
        O[54]) );
  AOI22_X1 U64 ( .A1(A_ns[53]), .A2(n397), .B1(\A_s[53] ), .B2(n398), .ZN(n440) );
  INV_X1 U65 ( .A(\A_s[52] ), .ZN(n439) );
  INV_X1 U66 ( .A(A_ns[52]), .ZN(n438) );
  OAI221_X1 U67 ( .B1(n393), .B2(n441), .C1(n392), .C2(n442), .A(n443), .ZN(
        O[53]) );
  AOI22_X1 U68 ( .A1(A_ns[52]), .A2(n397), .B1(\A_s[52] ), .B2(n398), .ZN(n443) );
  INV_X1 U69 ( .A(\A_s[51] ), .ZN(n442) );
  INV_X1 U70 ( .A(A_ns[51]), .ZN(n441) );
  OAI221_X1 U71 ( .B1(n393), .B2(n444), .C1(n392), .C2(n445), .A(n446), .ZN(
        O[52]) );
  AOI22_X1 U72 ( .A1(A_ns[51]), .A2(n397), .B1(\A_s[51] ), .B2(n398), .ZN(n446) );
  INV_X1 U73 ( .A(\A_s[50] ), .ZN(n445) );
  INV_X1 U74 ( .A(A_ns[50]), .ZN(n444) );
  OAI221_X1 U75 ( .B1(n393), .B2(n447), .C1(n392), .C2(n448), .A(n449), .ZN(
        O[51]) );
  AOI22_X1 U76 ( .A1(A_ns[50]), .A2(n397), .B1(\A_s[50] ), .B2(n398), .ZN(n449) );
  INV_X1 U77 ( .A(\A_s[49] ), .ZN(n448) );
  INV_X1 U78 ( .A(A_ns[49]), .ZN(n447) );
  OAI221_X1 U79 ( .B1(n393), .B2(n450), .C1(n392), .C2(n451), .A(n452), .ZN(
        O[50]) );
  AOI22_X1 U80 ( .A1(A_ns[49]), .A2(n397), .B1(\A_s[49] ), .B2(n398), .ZN(n452) );
  INV_X1 U81 ( .A(\A_s[48] ), .ZN(n451) );
  INV_X1 U82 ( .A(A_ns[48]), .ZN(n450) );
  OAI221_X1 U83 ( .B1(n393), .B2(n453), .C1(n392), .C2(n454), .A(n455), .ZN(
        O[4]) );
  AOI22_X1 U84 ( .A1(A_ns[3]), .A2(n397), .B1(\A_s[3] ), .B2(n398), .ZN(n455)
         );
  INV_X1 U85 ( .A(\A_s[2] ), .ZN(n454) );
  INV_X1 U86 ( .A(A_ns[2]), .ZN(n453) );
  OAI221_X1 U87 ( .B1(n393), .B2(n456), .C1(n392), .C2(n457), .A(n458), .ZN(
        O[49]) );
  AOI22_X1 U88 ( .A1(A_ns[48]), .A2(n397), .B1(\A_s[48] ), .B2(n398), .ZN(n458) );
  INV_X1 U89 ( .A(\A_s[47] ), .ZN(n457) );
  INV_X1 U90 ( .A(A_ns[47]), .ZN(n456) );
  OAI221_X1 U91 ( .B1(n393), .B2(n459), .C1(n392), .C2(n460), .A(n461), .ZN(
        O[48]) );
  AOI22_X1 U92 ( .A1(A_ns[47]), .A2(n397), .B1(\A_s[47] ), .B2(n398), .ZN(n461) );
  INV_X1 U93 ( .A(\A_s[46] ), .ZN(n460) );
  INV_X1 U94 ( .A(A_ns[46]), .ZN(n459) );
  OAI221_X1 U95 ( .B1(n393), .B2(n462), .C1(n392), .C2(n463), .A(n464), .ZN(
        O[47]) );
  AOI22_X1 U96 ( .A1(A_ns[46]), .A2(n397), .B1(\A_s[46] ), .B2(n398), .ZN(n464) );
  INV_X1 U97 ( .A(\A_s[45] ), .ZN(n463) );
  INV_X1 U98 ( .A(A_ns[45]), .ZN(n462) );
  OAI221_X1 U99 ( .B1(n393), .B2(n465), .C1(n392), .C2(n466), .A(n467), .ZN(
        O[46]) );
  AOI22_X1 U100 ( .A1(A_ns[45]), .A2(n397), .B1(\A_s[45] ), .B2(n398), .ZN(
        n467) );
  INV_X1 U101 ( .A(\A_s[44] ), .ZN(n466) );
  INV_X1 U102 ( .A(A_ns[44]), .ZN(n465) );
  OAI221_X1 U103 ( .B1(n393), .B2(n468), .C1(n392), .C2(n469), .A(n470), .ZN(
        O[45]) );
  AOI22_X1 U104 ( .A1(A_ns[44]), .A2(n397), .B1(\A_s[44] ), .B2(n398), .ZN(
        n470) );
  INV_X1 U105 ( .A(\A_s[43] ), .ZN(n469) );
  INV_X1 U106 ( .A(A_ns[43]), .ZN(n468) );
  OAI221_X1 U107 ( .B1(n393), .B2(n471), .C1(n392), .C2(n472), .A(n473), .ZN(
        O[44]) );
  AOI22_X1 U108 ( .A1(A_ns[43]), .A2(n397), .B1(\A_s[43] ), .B2(n398), .ZN(
        n473) );
  INV_X1 U109 ( .A(\A_s[42] ), .ZN(n472) );
  INV_X1 U110 ( .A(A_ns[42]), .ZN(n471) );
  OAI221_X1 U111 ( .B1(n393), .B2(n474), .C1(n392), .C2(n475), .A(n476), .ZN(
        O[43]) );
  AOI22_X1 U112 ( .A1(A_ns[42]), .A2(n397), .B1(\A_s[42] ), .B2(n398), .ZN(
        n476) );
  INV_X1 U113 ( .A(\A_s[41] ), .ZN(n475) );
  INV_X1 U114 ( .A(A_ns[41]), .ZN(n474) );
  OAI221_X1 U115 ( .B1(n393), .B2(n477), .C1(n392), .C2(n478), .A(n479), .ZN(
        O[42]) );
  AOI22_X1 U116 ( .A1(A_ns[41]), .A2(n397), .B1(\A_s[41] ), .B2(n398), .ZN(
        n479) );
  INV_X1 U117 ( .A(\A_s[40] ), .ZN(n478) );
  INV_X1 U118 ( .A(A_ns[40]), .ZN(n477) );
  OAI221_X1 U119 ( .B1(n393), .B2(n480), .C1(n392), .C2(n481), .A(n482), .ZN(
        O[41]) );
  AOI22_X1 U120 ( .A1(A_ns[40]), .A2(n397), .B1(\A_s[40] ), .B2(n398), .ZN(
        n482) );
  INV_X1 U121 ( .A(\A_s[39] ), .ZN(n481) );
  INV_X1 U122 ( .A(A_ns[39]), .ZN(n480) );
  OAI221_X1 U123 ( .B1(n393), .B2(n483), .C1(n392), .C2(n484), .A(n485), .ZN(
        O[40]) );
  AOI22_X1 U124 ( .A1(A_ns[39]), .A2(n397), .B1(\A_s[39] ), .B2(n398), .ZN(
        n485) );
  INV_X1 U125 ( .A(\A_s[38] ), .ZN(n484) );
  INV_X1 U126 ( .A(A_ns[38]), .ZN(n483) );
  OAI221_X1 U127 ( .B1(n393), .B2(n486), .C1(n392), .C2(n487), .A(n488), .ZN(
        O[3]) );
  AOI22_X1 U128 ( .A1(A_ns[2]), .A2(n397), .B1(\A_s[2] ), .B2(n398), .ZN(n488)
         );
  INV_X1 U129 ( .A(\A_s[1] ), .ZN(n487) );
  INV_X1 U130 ( .A(A_ns[1]), .ZN(n486) );
  OAI221_X1 U131 ( .B1(n393), .B2(n489), .C1(n392), .C2(n490), .A(n491), .ZN(
        O[39]) );
  AOI22_X1 U132 ( .A1(A_ns[38]), .A2(n397), .B1(\A_s[38] ), .B2(n398), .ZN(
        n491) );
  INV_X1 U133 ( .A(\A_s[37] ), .ZN(n490) );
  INV_X1 U134 ( .A(A_ns[37]), .ZN(n489) );
  OAI221_X1 U135 ( .B1(n393), .B2(n492), .C1(n392), .C2(n493), .A(n494), .ZN(
        O[38]) );
  AOI22_X1 U136 ( .A1(A_ns[37]), .A2(n397), .B1(\A_s[37] ), .B2(n398), .ZN(
        n494) );
  INV_X1 U137 ( .A(\A_s[36] ), .ZN(n493) );
  INV_X1 U138 ( .A(A_ns[36]), .ZN(n492) );
  OAI221_X1 U139 ( .B1(n393), .B2(n495), .C1(n392), .C2(n496), .A(n497), .ZN(
        O[37]) );
  AOI22_X1 U140 ( .A1(A_ns[36]), .A2(n397), .B1(\A_s[36] ), .B2(n398), .ZN(
        n497) );
  INV_X1 U141 ( .A(\A_s[35] ), .ZN(n496) );
  INV_X1 U142 ( .A(A_ns[35]), .ZN(n495) );
  OAI221_X1 U143 ( .B1(n393), .B2(n498), .C1(n392), .C2(n499), .A(n500), .ZN(
        O[36]) );
  AOI22_X1 U144 ( .A1(A_ns[35]), .A2(n397), .B1(\A_s[35] ), .B2(n398), .ZN(
        n500) );
  INV_X1 U145 ( .A(\A_s[34] ), .ZN(n499) );
  INV_X1 U146 ( .A(A_ns[34]), .ZN(n498) );
  OAI221_X1 U147 ( .B1(n393), .B2(n501), .C1(n392), .C2(n502), .A(n503), .ZN(
        O[35]) );
  AOI22_X1 U148 ( .A1(A_ns[34]), .A2(n397), .B1(\A_s[34] ), .B2(n398), .ZN(
        n503) );
  INV_X1 U149 ( .A(\A_s[33] ), .ZN(n502) );
  INV_X1 U150 ( .A(A_ns[33]), .ZN(n501) );
  OAI221_X1 U151 ( .B1(n393), .B2(n504), .C1(n392), .C2(n505), .A(n506), .ZN(
        O[34]) );
  AOI22_X1 U152 ( .A1(A_ns[33]), .A2(n397), .B1(\A_s[33] ), .B2(n398), .ZN(
        n506) );
  INV_X1 U153 ( .A(\A_s[32] ), .ZN(n505) );
  INV_X1 U154 ( .A(A_ns[32]), .ZN(n504) );
  OAI221_X1 U155 ( .B1(n393), .B2(n507), .C1(n392), .C2(n508), .A(n509), .ZN(
        O[33]) );
  AOI22_X1 U156 ( .A1(A_ns[32]), .A2(n397), .B1(\A_s[32] ), .B2(n398), .ZN(
        n509) );
  INV_X1 U157 ( .A(\A_s[31] ), .ZN(n508) );
  INV_X1 U158 ( .A(A_ns[31]), .ZN(n507) );
  OAI221_X1 U159 ( .B1(n393), .B2(n510), .C1(n392), .C2(n511), .A(n512), .ZN(
        O[32]) );
  AOI22_X1 U160 ( .A1(A_ns[31]), .A2(n397), .B1(\A_s[31] ), .B2(n398), .ZN(
        n512) );
  INV_X1 U161 ( .A(\A_s[30] ), .ZN(n511) );
  INV_X1 U162 ( .A(A_ns[30]), .ZN(n510) );
  OAI221_X1 U163 ( .B1(n393), .B2(n513), .C1(n392), .C2(n514), .A(n515), .ZN(
        O[31]) );
  AOI22_X1 U164 ( .A1(A_ns[30]), .A2(n397), .B1(\A_s[30] ), .B2(n398), .ZN(
        n515) );
  INV_X1 U165 ( .A(\A_s[29] ), .ZN(n514) );
  INV_X1 U166 ( .A(A_ns[29]), .ZN(n513) );
  OAI221_X1 U167 ( .B1(n393), .B2(n516), .C1(n392), .C2(n517), .A(n518), .ZN(
        O[30]) );
  AOI22_X1 U168 ( .A1(A_ns[29]), .A2(n397), .B1(\A_s[29] ), .B2(n398), .ZN(
        n518) );
  INV_X1 U169 ( .A(\A_s[28] ), .ZN(n517) );
  INV_X1 U170 ( .A(A_ns[28]), .ZN(n516) );
  OAI221_X1 U171 ( .B1(n393), .B2(n519), .C1(n392), .C2(n520), .A(n521), .ZN(
        O[2]) );
  AOI22_X1 U172 ( .A1(A_ns[1]), .A2(n397), .B1(\A_s[1] ), .B2(n398), .ZN(n521)
         );
  OAI221_X1 U173 ( .B1(n393), .B2(n522), .C1(n392), .C2(n523), .A(n524), .ZN(
        O[29]) );
  AOI22_X1 U174 ( .A1(A_ns[28]), .A2(n397), .B1(\A_s[28] ), .B2(n398), .ZN(
        n524) );
  INV_X1 U175 ( .A(\A_s[27] ), .ZN(n523) );
  INV_X1 U176 ( .A(A_ns[27]), .ZN(n522) );
  OAI221_X1 U177 ( .B1(n393), .B2(n525), .C1(n392), .C2(n526), .A(n527), .ZN(
        O[28]) );
  AOI22_X1 U178 ( .A1(A_ns[27]), .A2(n397), .B1(\A_s[27] ), .B2(n398), .ZN(
        n527) );
  INV_X1 U179 ( .A(\A_s[26] ), .ZN(n526) );
  INV_X1 U180 ( .A(A_ns[26]), .ZN(n525) );
  OAI221_X1 U181 ( .B1(n393), .B2(n528), .C1(n392), .C2(n529), .A(n530), .ZN(
        O[27]) );
  AOI22_X1 U182 ( .A1(A_ns[26]), .A2(n397), .B1(\A_s[26] ), .B2(n398), .ZN(
        n530) );
  INV_X1 U183 ( .A(\A_s[25] ), .ZN(n529) );
  INV_X1 U184 ( .A(A_ns[25]), .ZN(n528) );
  OAI221_X1 U185 ( .B1(n393), .B2(n531), .C1(n392), .C2(n532), .A(n533), .ZN(
        O[26]) );
  AOI22_X1 U186 ( .A1(A_ns[25]), .A2(n397), .B1(\A_s[25] ), .B2(n398), .ZN(
        n533) );
  INV_X1 U187 ( .A(\A_s[24] ), .ZN(n532) );
  INV_X1 U188 ( .A(A_ns[24]), .ZN(n531) );
  OAI221_X1 U189 ( .B1(n393), .B2(n534), .C1(n392), .C2(n535), .A(n536), .ZN(
        O[25]) );
  AOI22_X1 U190 ( .A1(A_ns[24]), .A2(n397), .B1(\A_s[24] ), .B2(n398), .ZN(
        n536) );
  INV_X1 U191 ( .A(\A_s[23] ), .ZN(n535) );
  INV_X1 U192 ( .A(A_ns[23]), .ZN(n534) );
  OAI221_X1 U193 ( .B1(n393), .B2(n537), .C1(n392), .C2(n538), .A(n539), .ZN(
        O[24]) );
  AOI22_X1 U194 ( .A1(A_ns[23]), .A2(n397), .B1(\A_s[23] ), .B2(n398), .ZN(
        n539) );
  INV_X1 U195 ( .A(\A_s[22] ), .ZN(n538) );
  INV_X1 U196 ( .A(A_ns[22]), .ZN(n537) );
  OAI221_X1 U197 ( .B1(n393), .B2(n540), .C1(n392), .C2(n541), .A(n542), .ZN(
        O[23]) );
  AOI22_X1 U198 ( .A1(A_ns[22]), .A2(n397), .B1(\A_s[22] ), .B2(n398), .ZN(
        n542) );
  INV_X1 U199 ( .A(\A_s[21] ), .ZN(n541) );
  INV_X1 U200 ( .A(A_ns[21]), .ZN(n540) );
  OAI221_X1 U201 ( .B1(n393), .B2(n543), .C1(n392), .C2(n544), .A(n545), .ZN(
        O[22]) );
  AOI22_X1 U202 ( .A1(A_ns[21]), .A2(n397), .B1(\A_s[21] ), .B2(n398), .ZN(
        n545) );
  INV_X1 U203 ( .A(\A_s[20] ), .ZN(n544) );
  INV_X1 U204 ( .A(A_ns[20]), .ZN(n543) );
  OAI221_X1 U205 ( .B1(n393), .B2(n546), .C1(n392), .C2(n547), .A(n548), .ZN(
        O[21]) );
  AOI22_X1 U206 ( .A1(A_ns[20]), .A2(n397), .B1(\A_s[20] ), .B2(n398), .ZN(
        n548) );
  INV_X1 U207 ( .A(\A_s[19] ), .ZN(n547) );
  INV_X1 U208 ( .A(A_ns[19]), .ZN(n546) );
  OAI221_X1 U209 ( .B1(n393), .B2(n549), .C1(n392), .C2(n550), .A(n551), .ZN(
        O[20]) );
  AOI22_X1 U210 ( .A1(A_ns[19]), .A2(n397), .B1(\A_s[19] ), .B2(n398), .ZN(
        n551) );
  INV_X1 U211 ( .A(\A_s[18] ), .ZN(n550) );
  INV_X1 U212 ( .A(A_ns[18]), .ZN(n549) );
  OAI22_X1 U213 ( .A1(n552), .A2(n520), .B1(n553), .B2(n519), .ZN(O[1]) );
  INV_X1 U214 ( .A(A_ns[0]), .ZN(n519) );
  INV_X1 U215 ( .A(\A_s[0] ), .ZN(n520) );
  OAI221_X1 U216 ( .B1(n393), .B2(n554), .C1(n392), .C2(n555), .A(n556), .ZN(
        O[19]) );
  AOI22_X1 U217 ( .A1(A_ns[18]), .A2(n397), .B1(\A_s[18] ), .B2(n398), .ZN(
        n556) );
  INV_X1 U218 ( .A(\A_s[17] ), .ZN(n555) );
  INV_X1 U219 ( .A(A_ns[17]), .ZN(n554) );
  OAI221_X1 U220 ( .B1(n393), .B2(n557), .C1(n392), .C2(n558), .A(n559), .ZN(
        O[18]) );
  AOI22_X1 U221 ( .A1(A_ns[17]), .A2(n397), .B1(\A_s[17] ), .B2(n398), .ZN(
        n559) );
  INV_X1 U222 ( .A(\A_s[16] ), .ZN(n558) );
  INV_X1 U223 ( .A(A_ns[16]), .ZN(n557) );
  OAI221_X1 U224 ( .B1(n393), .B2(n560), .C1(n392), .C2(n561), .A(n562), .ZN(
        O[17]) );
  AOI22_X1 U225 ( .A1(A_ns[16]), .A2(n397), .B1(\A_s[16] ), .B2(n398), .ZN(
        n562) );
  INV_X1 U226 ( .A(\A_s[15] ), .ZN(n561) );
  INV_X1 U227 ( .A(A_ns[15]), .ZN(n560) );
  OAI221_X1 U228 ( .B1(n393), .B2(n563), .C1(n392), .C2(n564), .A(n565), .ZN(
        O[16]) );
  AOI22_X1 U229 ( .A1(A_ns[15]), .A2(n397), .B1(\A_s[15] ), .B2(n398), .ZN(
        n565) );
  INV_X1 U230 ( .A(\A_s[14] ), .ZN(n564) );
  INV_X1 U231 ( .A(A_ns[14]), .ZN(n563) );
  OAI221_X1 U232 ( .B1(n393), .B2(n566), .C1(n392), .C2(n567), .A(n568), .ZN(
        O[15]) );
  AOI22_X1 U233 ( .A1(A_ns[14]), .A2(n397), .B1(\A_s[14] ), .B2(n398), .ZN(
        n568) );
  INV_X1 U234 ( .A(\A_s[13] ), .ZN(n567) );
  INV_X1 U235 ( .A(A_ns[13]), .ZN(n566) );
  OAI221_X1 U236 ( .B1(n393), .B2(n569), .C1(n392), .C2(n570), .A(n571), .ZN(
        O[14]) );
  AOI22_X1 U237 ( .A1(A_ns[13]), .A2(n397), .B1(\A_s[13] ), .B2(n398), .ZN(
        n571) );
  INV_X1 U238 ( .A(\A_s[12] ), .ZN(n570) );
  INV_X1 U239 ( .A(A_ns[12]), .ZN(n569) );
  OAI221_X1 U240 ( .B1(n393), .B2(n572), .C1(n392), .C2(n573), .A(n574), .ZN(
        O[13]) );
  AOI22_X1 U241 ( .A1(A_ns[12]), .A2(n397), .B1(\A_s[12] ), .B2(n398), .ZN(
        n574) );
  INV_X1 U242 ( .A(\A_s[11] ), .ZN(n573) );
  INV_X1 U243 ( .A(A_ns[11]), .ZN(n572) );
  OAI221_X1 U244 ( .B1(n393), .B2(n575), .C1(n392), .C2(n576), .A(n577), .ZN(
        O[12]) );
  AOI22_X1 U245 ( .A1(A_ns[11]), .A2(n397), .B1(\A_s[11] ), .B2(n398), .ZN(
        n577) );
  INV_X1 U246 ( .A(\A_s[10] ), .ZN(n576) );
  INV_X1 U247 ( .A(A_ns[10]), .ZN(n575) );
  OAI221_X1 U248 ( .B1(n393), .B2(n578), .C1(n392), .C2(n579), .A(n580), .ZN(
        O[11]) );
  AOI22_X1 U249 ( .A1(A_ns[10]), .A2(n397), .B1(\A_s[10] ), .B2(n398), .ZN(
        n580) );
  INV_X1 U250 ( .A(\A_s[9] ), .ZN(n579) );
  INV_X1 U251 ( .A(A_ns[9]), .ZN(n578) );
  OAI221_X1 U252 ( .B1(n581), .B2(n393), .C1(n582), .C2(n392), .A(n583), .ZN(
        O[10]) );
  AOI22_X1 U253 ( .A1(A_ns[9]), .A2(n397), .B1(\A_s[9] ), .B2(n398), .ZN(n583)
         );
  NAND2_X1 U254 ( .A1(n584), .A2(n552), .ZN(n553) );
  NAND2_X1 U255 ( .A1(n584), .A2(n585), .ZN(n552) );
  XOR2_X1 U256 ( .A(B[23]), .B(B[24]), .Z(n584) );
  INV_X1 U257 ( .A(\A_s[8] ), .ZN(n582) );
  INV_X1 U258 ( .A(B[25]), .ZN(n585) );
  INV_X1 U259 ( .A(A_ns[8]), .ZN(n581) );
endmodule


module BOOTHENC_NBIT64_i26 ( A, A_n, A_ns, A_s, B, O, A_so, A_nso );
  input [63:0] A;
  input [63:0] A_n;
  input [63:0] A_ns;
  input [63:0] A_s;
  input [63:0] B;
  output [63:0] O;
  output [63:0] A_so;
  output [63:0] A_nso;
  wire   \A_s[61] , \A_s[60] , \A_s[59] , \A_s[58] , \A_s[57] , \A_s[56] ,
         \A_s[55] , \A_s[54] , \A_s[53] , \A_s[52] , \A_s[51] , \A_s[50] ,
         \A_s[49] , \A_s[48] , \A_s[47] , \A_s[46] , \A_s[45] , \A_s[44] ,
         \A_s[43] , \A_s[42] , \A_s[41] , \A_s[40] , \A_s[39] , \A_s[38] ,
         \A_s[37] , \A_s[36] , \A_s[35] , \A_s[34] , \A_s[33] , \A_s[32] ,
         \A_s[31] , \A_s[30] , \A_s[29] , \A_s[28] , \A_s[27] , \A_s[26] ,
         \A_s[25] , \A_s[24] , \A_s[23] , \A_s[22] , \A_s[21] , \A_s[20] ,
         \A_s[19] , \A_s[18] , \A_s[17] , \A_s[16] , \A_s[15] , \A_s[14] ,
         \A_s[13] , \A_s[12] , \A_s[11] , \A_s[10] , \A_s[9] , \A_s[8] ,
         \A_s[7] , \A_s[6] , \A_s[5] , \A_s[4] , \A_s[3] , \A_s[2] , \A_s[1] ,
         \A_s[0] , n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585;
  assign A_nso[0] = 1'b0;
  assign A_nso[1] = 1'b0;
  assign A_so[0] = 1'b0;
  assign A_so[1] = 1'b0;
  assign O[0] = 1'b0;
  assign A_nso[63] = \A_s[61] ;
  assign A_so[63] = \A_s[61] ;
  assign \A_s[61]  = A_s[61];
  assign A_nso[62] = \A_s[60] ;
  assign A_so[62] = \A_s[60] ;
  assign \A_s[60]  = A_s[60];
  assign A_nso[61] = \A_s[59] ;
  assign A_so[61] = \A_s[59] ;
  assign \A_s[59]  = A_s[59];
  assign A_nso[60] = \A_s[58] ;
  assign A_so[60] = \A_s[58] ;
  assign \A_s[58]  = A_s[58];
  assign A_nso[59] = \A_s[57] ;
  assign A_so[59] = \A_s[57] ;
  assign \A_s[57]  = A_s[57];
  assign A_nso[58] = \A_s[56] ;
  assign A_so[58] = \A_s[56] ;
  assign \A_s[56]  = A_s[56];
  assign A_nso[57] = \A_s[55] ;
  assign A_so[57] = \A_s[55] ;
  assign \A_s[55]  = A_s[55];
  assign A_nso[56] = \A_s[54] ;
  assign A_so[56] = \A_s[54] ;
  assign \A_s[54]  = A_s[54];
  assign A_nso[55] = \A_s[53] ;
  assign A_so[55] = \A_s[53] ;
  assign \A_s[53]  = A_s[53];
  assign A_nso[54] = \A_s[52] ;
  assign A_so[54] = \A_s[52] ;
  assign \A_s[52]  = A_s[52];
  assign A_nso[53] = \A_s[51] ;
  assign A_so[53] = \A_s[51] ;
  assign \A_s[51]  = A_s[51];
  assign A_nso[52] = \A_s[50] ;
  assign A_so[52] = \A_s[50] ;
  assign \A_s[50]  = A_s[50];
  assign A_nso[51] = \A_s[49] ;
  assign A_so[51] = \A_s[49] ;
  assign \A_s[49]  = A_s[49];
  assign A_nso[50] = \A_s[48] ;
  assign A_so[50] = \A_s[48] ;
  assign \A_s[48]  = A_s[48];
  assign A_nso[49] = \A_s[47] ;
  assign A_so[49] = \A_s[47] ;
  assign \A_s[47]  = A_s[47];
  assign A_nso[48] = \A_s[46] ;
  assign A_so[48] = \A_s[46] ;
  assign \A_s[46]  = A_s[46];
  assign A_nso[47] = \A_s[45] ;
  assign A_so[47] = \A_s[45] ;
  assign \A_s[45]  = A_s[45];
  assign A_nso[46] = \A_s[44] ;
  assign A_so[46] = \A_s[44] ;
  assign \A_s[44]  = A_s[44];
  assign A_nso[45] = \A_s[43] ;
  assign A_so[45] = \A_s[43] ;
  assign \A_s[43]  = A_s[43];
  assign A_nso[44] = \A_s[42] ;
  assign A_so[44] = \A_s[42] ;
  assign \A_s[42]  = A_s[42];
  assign A_nso[43] = \A_s[41] ;
  assign A_so[43] = \A_s[41] ;
  assign \A_s[41]  = A_s[41];
  assign A_nso[42] = \A_s[40] ;
  assign A_so[42] = \A_s[40] ;
  assign \A_s[40]  = A_s[40];
  assign A_nso[41] = \A_s[39] ;
  assign A_so[41] = \A_s[39] ;
  assign \A_s[39]  = A_s[39];
  assign A_nso[40] = \A_s[38] ;
  assign A_so[40] = \A_s[38] ;
  assign \A_s[38]  = A_s[38];
  assign A_nso[39] = \A_s[37] ;
  assign A_so[39] = \A_s[37] ;
  assign \A_s[37]  = A_s[37];
  assign A_nso[38] = \A_s[36] ;
  assign A_so[38] = \A_s[36] ;
  assign \A_s[36]  = A_s[36];
  assign A_nso[37] = \A_s[35] ;
  assign A_so[37] = \A_s[35] ;
  assign \A_s[35]  = A_s[35];
  assign A_nso[36] = \A_s[34] ;
  assign A_so[36] = \A_s[34] ;
  assign \A_s[34]  = A_s[34];
  assign A_nso[35] = \A_s[33] ;
  assign A_so[35] = \A_s[33] ;
  assign \A_s[33]  = A_s[33];
  assign A_nso[34] = \A_s[32] ;
  assign A_so[34] = \A_s[32] ;
  assign \A_s[32]  = A_s[32];
  assign A_nso[33] = \A_s[31] ;
  assign A_so[33] = \A_s[31] ;
  assign \A_s[31]  = A_s[31];
  assign A_nso[32] = \A_s[30] ;
  assign A_so[32] = \A_s[30] ;
  assign \A_s[30]  = A_s[30];
  assign A_nso[31] = \A_s[29] ;
  assign A_so[31] = \A_s[29] ;
  assign \A_s[29]  = A_s[29];
  assign A_nso[30] = \A_s[28] ;
  assign A_so[30] = \A_s[28] ;
  assign \A_s[28]  = A_s[28];
  assign A_nso[29] = \A_s[27] ;
  assign A_so[29] = \A_s[27] ;
  assign \A_s[27]  = A_s[27];
  assign A_nso[28] = \A_s[26] ;
  assign A_so[28] = \A_s[26] ;
  assign \A_s[26]  = A_s[26];
  assign A_nso[27] = \A_s[25] ;
  assign A_so[27] = \A_s[25] ;
  assign \A_s[25]  = A_s[25];
  assign A_nso[26] = \A_s[24] ;
  assign A_so[26] = \A_s[24] ;
  assign \A_s[24]  = A_s[24];
  assign A_nso[25] = \A_s[23] ;
  assign A_so[25] = \A_s[23] ;
  assign \A_s[23]  = A_s[23];
  assign A_nso[24] = \A_s[22] ;
  assign A_so[24] = \A_s[22] ;
  assign \A_s[22]  = A_s[22];
  assign A_nso[23] = \A_s[21] ;
  assign A_so[23] = \A_s[21] ;
  assign \A_s[21]  = A_s[21];
  assign A_nso[22] = \A_s[20] ;
  assign A_so[22] = \A_s[20] ;
  assign \A_s[20]  = A_s[20];
  assign A_nso[21] = \A_s[19] ;
  assign A_so[21] = \A_s[19] ;
  assign \A_s[19]  = A_s[19];
  assign A_nso[20] = \A_s[18] ;
  assign A_so[20] = \A_s[18] ;
  assign \A_s[18]  = A_s[18];
  assign A_nso[19] = \A_s[17] ;
  assign A_so[19] = \A_s[17] ;
  assign \A_s[17]  = A_s[17];
  assign A_nso[18] = \A_s[16] ;
  assign A_so[18] = \A_s[16] ;
  assign \A_s[16]  = A_s[16];
  assign A_nso[17] = \A_s[15] ;
  assign A_so[17] = \A_s[15] ;
  assign \A_s[15]  = A_s[15];
  assign A_nso[16] = \A_s[14] ;
  assign A_so[16] = \A_s[14] ;
  assign \A_s[14]  = A_s[14];
  assign A_nso[15] = \A_s[13] ;
  assign A_so[15] = \A_s[13] ;
  assign \A_s[13]  = A_s[13];
  assign A_nso[14] = \A_s[12] ;
  assign A_so[14] = \A_s[12] ;
  assign \A_s[12]  = A_s[12];
  assign A_nso[13] = \A_s[11] ;
  assign A_so[13] = \A_s[11] ;
  assign \A_s[11]  = A_s[11];
  assign A_nso[12] = \A_s[10] ;
  assign A_so[12] = \A_s[10] ;
  assign \A_s[10]  = A_s[10];
  assign A_nso[11] = \A_s[9] ;
  assign A_so[11] = \A_s[9] ;
  assign \A_s[9]  = A_s[9];
  assign A_nso[10] = \A_s[8] ;
  assign A_so[10] = \A_s[8] ;
  assign \A_s[8]  = A_s[8];
  assign A_nso[9] = \A_s[7] ;
  assign A_so[9] = \A_s[7] ;
  assign \A_s[7]  = A_s[7];
  assign A_nso[8] = \A_s[6] ;
  assign A_so[8] = \A_s[6] ;
  assign \A_s[6]  = A_s[6];
  assign A_nso[7] = \A_s[5] ;
  assign A_so[7] = \A_s[5] ;
  assign \A_s[5]  = A_s[5];
  assign A_nso[6] = \A_s[4] ;
  assign A_so[6] = \A_s[4] ;
  assign \A_s[4]  = A_s[4];
  assign A_nso[5] = \A_s[3] ;
  assign A_so[5] = \A_s[3] ;
  assign \A_s[3]  = A_s[3];
  assign A_nso[4] = \A_s[2] ;
  assign A_so[4] = \A_s[2] ;
  assign \A_s[2]  = A_s[2];
  assign A_nso[3] = \A_s[1] ;
  assign A_so[3] = \A_s[1] ;
  assign \A_s[1]  = A_s[1];
  assign A_nso[2] = \A_s[0] ;
  assign A_so[2] = \A_s[0] ;
  assign \A_s[0]  = A_s[0];

  AND3_X1 U2 ( .A1(B[26]), .A2(n585), .A3(B[25]), .ZN(n391) );
  INV_X4 U3 ( .A(n391), .ZN(n392) );
  INV_X4 U4 ( .A(n552), .ZN(n398) );
  OR3_X4 U5 ( .A1(B[25]), .A2(B[26]), .A3(n585), .ZN(n393) );
  INV_X4 U6 ( .A(n553), .ZN(n397) );
  OAI221_X1 U7 ( .B1(n393), .B2(n394), .C1(n392), .C2(n395), .A(n396), .ZN(
        O[9]) );
  AOI22_X1 U8 ( .A1(A_ns[8]), .A2(n397), .B1(\A_s[8] ), .B2(n398), .ZN(n396)
         );
  INV_X1 U9 ( .A(\A_s[7] ), .ZN(n395) );
  INV_X1 U10 ( .A(A_ns[7]), .ZN(n394) );
  OAI221_X1 U11 ( .B1(n393), .B2(n399), .C1(n392), .C2(n400), .A(n401), .ZN(
        O[8]) );
  AOI22_X1 U12 ( .A1(A_ns[7]), .A2(n397), .B1(\A_s[7] ), .B2(n398), .ZN(n401)
         );
  INV_X1 U13 ( .A(\A_s[6] ), .ZN(n400) );
  INV_X1 U14 ( .A(A_ns[6]), .ZN(n399) );
  OAI221_X1 U15 ( .B1(n393), .B2(n402), .C1(n392), .C2(n403), .A(n404), .ZN(
        O[7]) );
  AOI22_X1 U16 ( .A1(A_ns[6]), .A2(n397), .B1(\A_s[6] ), .B2(n398), .ZN(n404)
         );
  INV_X1 U17 ( .A(\A_s[5] ), .ZN(n403) );
  INV_X1 U18 ( .A(A_ns[5]), .ZN(n402) );
  OAI221_X1 U19 ( .B1(n393), .B2(n405), .C1(n392), .C2(n406), .A(n407), .ZN(
        O[6]) );
  AOI22_X1 U20 ( .A1(A_ns[5]), .A2(n397), .B1(\A_s[5] ), .B2(n398), .ZN(n407)
         );
  INV_X1 U21 ( .A(\A_s[4] ), .ZN(n406) );
  INV_X1 U22 ( .A(A_ns[4]), .ZN(n405) );
  OAI221_X1 U23 ( .B1(n393), .B2(n408), .C1(n392), .C2(n409), .A(n410), .ZN(
        O[63]) );
  AOI22_X1 U24 ( .A1(A_ns[62]), .A2(n397), .B1(A_s[62]), .B2(n398), .ZN(n410)
         );
  INV_X1 U25 ( .A(\A_s[61] ), .ZN(n409) );
  INV_X1 U26 ( .A(A_ns[61]), .ZN(n408) );
  OAI221_X1 U27 ( .B1(n393), .B2(n411), .C1(n392), .C2(n412), .A(n413), .ZN(
        O[62]) );
  AOI22_X1 U28 ( .A1(A_ns[61]), .A2(n397), .B1(\A_s[61] ), .B2(n398), .ZN(n413) );
  INV_X1 U29 ( .A(\A_s[60] ), .ZN(n412) );
  INV_X1 U30 ( .A(A_ns[60]), .ZN(n411) );
  OAI221_X1 U31 ( .B1(n393), .B2(n414), .C1(n392), .C2(n415), .A(n416), .ZN(
        O[61]) );
  AOI22_X1 U32 ( .A1(A_ns[60]), .A2(n397), .B1(\A_s[60] ), .B2(n398), .ZN(n416) );
  INV_X1 U33 ( .A(\A_s[59] ), .ZN(n415) );
  INV_X1 U34 ( .A(A_ns[59]), .ZN(n414) );
  OAI221_X1 U35 ( .B1(n393), .B2(n417), .C1(n392), .C2(n418), .A(n419), .ZN(
        O[60]) );
  AOI22_X1 U36 ( .A1(A_ns[59]), .A2(n397), .B1(\A_s[59] ), .B2(n398), .ZN(n419) );
  INV_X1 U37 ( .A(\A_s[58] ), .ZN(n418) );
  INV_X1 U38 ( .A(A_ns[58]), .ZN(n417) );
  OAI221_X1 U39 ( .B1(n393), .B2(n420), .C1(n392), .C2(n421), .A(n422), .ZN(
        O[5]) );
  AOI22_X1 U40 ( .A1(A_ns[4]), .A2(n397), .B1(\A_s[4] ), .B2(n398), .ZN(n422)
         );
  INV_X1 U41 ( .A(\A_s[3] ), .ZN(n421) );
  INV_X1 U42 ( .A(A_ns[3]), .ZN(n420) );
  OAI221_X1 U43 ( .B1(n393), .B2(n423), .C1(n392), .C2(n424), .A(n425), .ZN(
        O[59]) );
  AOI22_X1 U44 ( .A1(A_ns[58]), .A2(n397), .B1(\A_s[58] ), .B2(n398), .ZN(n425) );
  INV_X1 U45 ( .A(\A_s[57] ), .ZN(n424) );
  INV_X1 U46 ( .A(A_ns[57]), .ZN(n423) );
  OAI221_X1 U47 ( .B1(n393), .B2(n426), .C1(n392), .C2(n427), .A(n428), .ZN(
        O[58]) );
  AOI22_X1 U48 ( .A1(A_ns[57]), .A2(n397), .B1(\A_s[57] ), .B2(n398), .ZN(n428) );
  INV_X1 U49 ( .A(\A_s[56] ), .ZN(n427) );
  INV_X1 U50 ( .A(A_ns[56]), .ZN(n426) );
  OAI221_X1 U51 ( .B1(n393), .B2(n429), .C1(n392), .C2(n430), .A(n431), .ZN(
        O[57]) );
  AOI22_X1 U52 ( .A1(A_ns[56]), .A2(n397), .B1(\A_s[56] ), .B2(n398), .ZN(n431) );
  INV_X1 U53 ( .A(\A_s[55] ), .ZN(n430) );
  INV_X1 U54 ( .A(A_ns[55]), .ZN(n429) );
  OAI221_X1 U55 ( .B1(n393), .B2(n432), .C1(n392), .C2(n433), .A(n434), .ZN(
        O[56]) );
  AOI22_X1 U56 ( .A1(A_ns[55]), .A2(n397), .B1(\A_s[55] ), .B2(n398), .ZN(n434) );
  INV_X1 U57 ( .A(\A_s[54] ), .ZN(n433) );
  INV_X1 U58 ( .A(A_ns[54]), .ZN(n432) );
  OAI221_X1 U59 ( .B1(n393), .B2(n435), .C1(n392), .C2(n436), .A(n437), .ZN(
        O[55]) );
  AOI22_X1 U60 ( .A1(A_ns[54]), .A2(n397), .B1(\A_s[54] ), .B2(n398), .ZN(n437) );
  INV_X1 U61 ( .A(\A_s[53] ), .ZN(n436) );
  INV_X1 U62 ( .A(A_ns[53]), .ZN(n435) );
  OAI221_X1 U63 ( .B1(n393), .B2(n438), .C1(n392), .C2(n439), .A(n440), .ZN(
        O[54]) );
  AOI22_X1 U64 ( .A1(A_ns[53]), .A2(n397), .B1(\A_s[53] ), .B2(n398), .ZN(n440) );
  INV_X1 U65 ( .A(\A_s[52] ), .ZN(n439) );
  INV_X1 U66 ( .A(A_ns[52]), .ZN(n438) );
  OAI221_X1 U67 ( .B1(n393), .B2(n441), .C1(n392), .C2(n442), .A(n443), .ZN(
        O[53]) );
  AOI22_X1 U68 ( .A1(A_ns[52]), .A2(n397), .B1(\A_s[52] ), .B2(n398), .ZN(n443) );
  INV_X1 U69 ( .A(\A_s[51] ), .ZN(n442) );
  INV_X1 U70 ( .A(A_ns[51]), .ZN(n441) );
  OAI221_X1 U71 ( .B1(n393), .B2(n444), .C1(n392), .C2(n445), .A(n446), .ZN(
        O[52]) );
  AOI22_X1 U72 ( .A1(A_ns[51]), .A2(n397), .B1(\A_s[51] ), .B2(n398), .ZN(n446) );
  INV_X1 U73 ( .A(\A_s[50] ), .ZN(n445) );
  INV_X1 U74 ( .A(A_ns[50]), .ZN(n444) );
  OAI221_X1 U75 ( .B1(n393), .B2(n447), .C1(n392), .C2(n448), .A(n449), .ZN(
        O[51]) );
  AOI22_X1 U76 ( .A1(A_ns[50]), .A2(n397), .B1(\A_s[50] ), .B2(n398), .ZN(n449) );
  INV_X1 U77 ( .A(\A_s[49] ), .ZN(n448) );
  INV_X1 U78 ( .A(A_ns[49]), .ZN(n447) );
  OAI221_X1 U79 ( .B1(n393), .B2(n450), .C1(n392), .C2(n451), .A(n452), .ZN(
        O[50]) );
  AOI22_X1 U80 ( .A1(A_ns[49]), .A2(n397), .B1(\A_s[49] ), .B2(n398), .ZN(n452) );
  INV_X1 U81 ( .A(\A_s[48] ), .ZN(n451) );
  INV_X1 U82 ( .A(A_ns[48]), .ZN(n450) );
  OAI221_X1 U83 ( .B1(n393), .B2(n453), .C1(n392), .C2(n454), .A(n455), .ZN(
        O[4]) );
  AOI22_X1 U84 ( .A1(A_ns[3]), .A2(n397), .B1(\A_s[3] ), .B2(n398), .ZN(n455)
         );
  INV_X1 U85 ( .A(\A_s[2] ), .ZN(n454) );
  INV_X1 U86 ( .A(A_ns[2]), .ZN(n453) );
  OAI221_X1 U87 ( .B1(n393), .B2(n456), .C1(n392), .C2(n457), .A(n458), .ZN(
        O[49]) );
  AOI22_X1 U88 ( .A1(A_ns[48]), .A2(n397), .B1(\A_s[48] ), .B2(n398), .ZN(n458) );
  INV_X1 U89 ( .A(\A_s[47] ), .ZN(n457) );
  INV_X1 U90 ( .A(A_ns[47]), .ZN(n456) );
  OAI221_X1 U91 ( .B1(n393), .B2(n459), .C1(n392), .C2(n460), .A(n461), .ZN(
        O[48]) );
  AOI22_X1 U92 ( .A1(A_ns[47]), .A2(n397), .B1(\A_s[47] ), .B2(n398), .ZN(n461) );
  INV_X1 U93 ( .A(\A_s[46] ), .ZN(n460) );
  INV_X1 U94 ( .A(A_ns[46]), .ZN(n459) );
  OAI221_X1 U95 ( .B1(n393), .B2(n462), .C1(n392), .C2(n463), .A(n464), .ZN(
        O[47]) );
  AOI22_X1 U96 ( .A1(A_ns[46]), .A2(n397), .B1(\A_s[46] ), .B2(n398), .ZN(n464) );
  INV_X1 U97 ( .A(\A_s[45] ), .ZN(n463) );
  INV_X1 U98 ( .A(A_ns[45]), .ZN(n462) );
  OAI221_X1 U99 ( .B1(n393), .B2(n465), .C1(n392), .C2(n466), .A(n467), .ZN(
        O[46]) );
  AOI22_X1 U100 ( .A1(A_ns[45]), .A2(n397), .B1(\A_s[45] ), .B2(n398), .ZN(
        n467) );
  INV_X1 U101 ( .A(\A_s[44] ), .ZN(n466) );
  INV_X1 U102 ( .A(A_ns[44]), .ZN(n465) );
  OAI221_X1 U103 ( .B1(n393), .B2(n468), .C1(n392), .C2(n469), .A(n470), .ZN(
        O[45]) );
  AOI22_X1 U104 ( .A1(A_ns[44]), .A2(n397), .B1(\A_s[44] ), .B2(n398), .ZN(
        n470) );
  INV_X1 U105 ( .A(\A_s[43] ), .ZN(n469) );
  INV_X1 U106 ( .A(A_ns[43]), .ZN(n468) );
  OAI221_X1 U107 ( .B1(n393), .B2(n471), .C1(n392), .C2(n472), .A(n473), .ZN(
        O[44]) );
  AOI22_X1 U108 ( .A1(A_ns[43]), .A2(n397), .B1(\A_s[43] ), .B2(n398), .ZN(
        n473) );
  INV_X1 U109 ( .A(\A_s[42] ), .ZN(n472) );
  INV_X1 U110 ( .A(A_ns[42]), .ZN(n471) );
  OAI221_X1 U111 ( .B1(n393), .B2(n474), .C1(n392), .C2(n475), .A(n476), .ZN(
        O[43]) );
  AOI22_X1 U112 ( .A1(A_ns[42]), .A2(n397), .B1(\A_s[42] ), .B2(n398), .ZN(
        n476) );
  INV_X1 U113 ( .A(\A_s[41] ), .ZN(n475) );
  INV_X1 U114 ( .A(A_ns[41]), .ZN(n474) );
  OAI221_X1 U115 ( .B1(n393), .B2(n477), .C1(n392), .C2(n478), .A(n479), .ZN(
        O[42]) );
  AOI22_X1 U116 ( .A1(A_ns[41]), .A2(n397), .B1(\A_s[41] ), .B2(n398), .ZN(
        n479) );
  INV_X1 U117 ( .A(\A_s[40] ), .ZN(n478) );
  INV_X1 U118 ( .A(A_ns[40]), .ZN(n477) );
  OAI221_X1 U119 ( .B1(n393), .B2(n480), .C1(n392), .C2(n481), .A(n482), .ZN(
        O[41]) );
  AOI22_X1 U120 ( .A1(A_ns[40]), .A2(n397), .B1(\A_s[40] ), .B2(n398), .ZN(
        n482) );
  INV_X1 U121 ( .A(\A_s[39] ), .ZN(n481) );
  INV_X1 U122 ( .A(A_ns[39]), .ZN(n480) );
  OAI221_X1 U123 ( .B1(n393), .B2(n483), .C1(n392), .C2(n484), .A(n485), .ZN(
        O[40]) );
  AOI22_X1 U124 ( .A1(A_ns[39]), .A2(n397), .B1(\A_s[39] ), .B2(n398), .ZN(
        n485) );
  INV_X1 U125 ( .A(\A_s[38] ), .ZN(n484) );
  INV_X1 U126 ( .A(A_ns[38]), .ZN(n483) );
  OAI221_X1 U127 ( .B1(n393), .B2(n486), .C1(n392), .C2(n487), .A(n488), .ZN(
        O[3]) );
  AOI22_X1 U128 ( .A1(A_ns[2]), .A2(n397), .B1(\A_s[2] ), .B2(n398), .ZN(n488)
         );
  INV_X1 U129 ( .A(\A_s[1] ), .ZN(n487) );
  INV_X1 U130 ( .A(A_ns[1]), .ZN(n486) );
  OAI221_X1 U131 ( .B1(n393), .B2(n489), .C1(n392), .C2(n490), .A(n491), .ZN(
        O[39]) );
  AOI22_X1 U132 ( .A1(A_ns[38]), .A2(n397), .B1(\A_s[38] ), .B2(n398), .ZN(
        n491) );
  INV_X1 U133 ( .A(\A_s[37] ), .ZN(n490) );
  INV_X1 U134 ( .A(A_ns[37]), .ZN(n489) );
  OAI221_X1 U135 ( .B1(n393), .B2(n492), .C1(n392), .C2(n493), .A(n494), .ZN(
        O[38]) );
  AOI22_X1 U136 ( .A1(A_ns[37]), .A2(n397), .B1(\A_s[37] ), .B2(n398), .ZN(
        n494) );
  INV_X1 U137 ( .A(\A_s[36] ), .ZN(n493) );
  INV_X1 U138 ( .A(A_ns[36]), .ZN(n492) );
  OAI221_X1 U139 ( .B1(n393), .B2(n495), .C1(n392), .C2(n496), .A(n497), .ZN(
        O[37]) );
  AOI22_X1 U140 ( .A1(A_ns[36]), .A2(n397), .B1(\A_s[36] ), .B2(n398), .ZN(
        n497) );
  INV_X1 U141 ( .A(\A_s[35] ), .ZN(n496) );
  INV_X1 U142 ( .A(A_ns[35]), .ZN(n495) );
  OAI221_X1 U143 ( .B1(n393), .B2(n498), .C1(n392), .C2(n499), .A(n500), .ZN(
        O[36]) );
  AOI22_X1 U144 ( .A1(A_ns[35]), .A2(n397), .B1(\A_s[35] ), .B2(n398), .ZN(
        n500) );
  INV_X1 U145 ( .A(\A_s[34] ), .ZN(n499) );
  INV_X1 U146 ( .A(A_ns[34]), .ZN(n498) );
  OAI221_X1 U147 ( .B1(n393), .B2(n501), .C1(n392), .C2(n502), .A(n503), .ZN(
        O[35]) );
  AOI22_X1 U148 ( .A1(A_ns[34]), .A2(n397), .B1(\A_s[34] ), .B2(n398), .ZN(
        n503) );
  INV_X1 U149 ( .A(\A_s[33] ), .ZN(n502) );
  INV_X1 U150 ( .A(A_ns[33]), .ZN(n501) );
  OAI221_X1 U151 ( .B1(n393), .B2(n504), .C1(n392), .C2(n505), .A(n506), .ZN(
        O[34]) );
  AOI22_X1 U152 ( .A1(A_ns[33]), .A2(n397), .B1(\A_s[33] ), .B2(n398), .ZN(
        n506) );
  INV_X1 U153 ( .A(\A_s[32] ), .ZN(n505) );
  INV_X1 U154 ( .A(A_ns[32]), .ZN(n504) );
  OAI221_X1 U155 ( .B1(n393), .B2(n507), .C1(n392), .C2(n508), .A(n509), .ZN(
        O[33]) );
  AOI22_X1 U156 ( .A1(A_ns[32]), .A2(n397), .B1(\A_s[32] ), .B2(n398), .ZN(
        n509) );
  INV_X1 U157 ( .A(\A_s[31] ), .ZN(n508) );
  INV_X1 U158 ( .A(A_ns[31]), .ZN(n507) );
  OAI221_X1 U159 ( .B1(n393), .B2(n510), .C1(n392), .C2(n511), .A(n512), .ZN(
        O[32]) );
  AOI22_X1 U160 ( .A1(A_ns[31]), .A2(n397), .B1(\A_s[31] ), .B2(n398), .ZN(
        n512) );
  INV_X1 U161 ( .A(\A_s[30] ), .ZN(n511) );
  INV_X1 U162 ( .A(A_ns[30]), .ZN(n510) );
  OAI221_X1 U163 ( .B1(n393), .B2(n513), .C1(n392), .C2(n514), .A(n515), .ZN(
        O[31]) );
  AOI22_X1 U164 ( .A1(A_ns[30]), .A2(n397), .B1(\A_s[30] ), .B2(n398), .ZN(
        n515) );
  INV_X1 U165 ( .A(\A_s[29] ), .ZN(n514) );
  INV_X1 U166 ( .A(A_ns[29]), .ZN(n513) );
  OAI221_X1 U167 ( .B1(n393), .B2(n516), .C1(n392), .C2(n517), .A(n518), .ZN(
        O[30]) );
  AOI22_X1 U168 ( .A1(A_ns[29]), .A2(n397), .B1(\A_s[29] ), .B2(n398), .ZN(
        n518) );
  INV_X1 U169 ( .A(\A_s[28] ), .ZN(n517) );
  INV_X1 U170 ( .A(A_ns[28]), .ZN(n516) );
  OAI221_X1 U171 ( .B1(n393), .B2(n519), .C1(n392), .C2(n520), .A(n521), .ZN(
        O[2]) );
  AOI22_X1 U172 ( .A1(A_ns[1]), .A2(n397), .B1(\A_s[1] ), .B2(n398), .ZN(n521)
         );
  OAI221_X1 U173 ( .B1(n393), .B2(n522), .C1(n392), .C2(n523), .A(n524), .ZN(
        O[29]) );
  AOI22_X1 U174 ( .A1(A_ns[28]), .A2(n397), .B1(\A_s[28] ), .B2(n398), .ZN(
        n524) );
  INV_X1 U175 ( .A(\A_s[27] ), .ZN(n523) );
  INV_X1 U176 ( .A(A_ns[27]), .ZN(n522) );
  OAI221_X1 U177 ( .B1(n393), .B2(n525), .C1(n392), .C2(n526), .A(n527), .ZN(
        O[28]) );
  AOI22_X1 U178 ( .A1(A_ns[27]), .A2(n397), .B1(\A_s[27] ), .B2(n398), .ZN(
        n527) );
  INV_X1 U179 ( .A(\A_s[26] ), .ZN(n526) );
  INV_X1 U180 ( .A(A_ns[26]), .ZN(n525) );
  OAI221_X1 U181 ( .B1(n393), .B2(n528), .C1(n392), .C2(n529), .A(n530), .ZN(
        O[27]) );
  AOI22_X1 U182 ( .A1(A_ns[26]), .A2(n397), .B1(\A_s[26] ), .B2(n398), .ZN(
        n530) );
  INV_X1 U183 ( .A(\A_s[25] ), .ZN(n529) );
  INV_X1 U184 ( .A(A_ns[25]), .ZN(n528) );
  OAI221_X1 U185 ( .B1(n393), .B2(n531), .C1(n392), .C2(n532), .A(n533), .ZN(
        O[26]) );
  AOI22_X1 U186 ( .A1(A_ns[25]), .A2(n397), .B1(\A_s[25] ), .B2(n398), .ZN(
        n533) );
  INV_X1 U187 ( .A(\A_s[24] ), .ZN(n532) );
  INV_X1 U188 ( .A(A_ns[24]), .ZN(n531) );
  OAI221_X1 U189 ( .B1(n393), .B2(n534), .C1(n392), .C2(n535), .A(n536), .ZN(
        O[25]) );
  AOI22_X1 U190 ( .A1(A_ns[24]), .A2(n397), .B1(\A_s[24] ), .B2(n398), .ZN(
        n536) );
  INV_X1 U191 ( .A(\A_s[23] ), .ZN(n535) );
  INV_X1 U192 ( .A(A_ns[23]), .ZN(n534) );
  OAI221_X1 U193 ( .B1(n393), .B2(n537), .C1(n392), .C2(n538), .A(n539), .ZN(
        O[24]) );
  AOI22_X1 U194 ( .A1(A_ns[23]), .A2(n397), .B1(\A_s[23] ), .B2(n398), .ZN(
        n539) );
  INV_X1 U195 ( .A(\A_s[22] ), .ZN(n538) );
  INV_X1 U196 ( .A(A_ns[22]), .ZN(n537) );
  OAI221_X1 U197 ( .B1(n393), .B2(n540), .C1(n392), .C2(n541), .A(n542), .ZN(
        O[23]) );
  AOI22_X1 U198 ( .A1(A_ns[22]), .A2(n397), .B1(\A_s[22] ), .B2(n398), .ZN(
        n542) );
  INV_X1 U199 ( .A(\A_s[21] ), .ZN(n541) );
  INV_X1 U200 ( .A(A_ns[21]), .ZN(n540) );
  OAI221_X1 U201 ( .B1(n393), .B2(n543), .C1(n392), .C2(n544), .A(n545), .ZN(
        O[22]) );
  AOI22_X1 U202 ( .A1(A_ns[21]), .A2(n397), .B1(\A_s[21] ), .B2(n398), .ZN(
        n545) );
  INV_X1 U203 ( .A(\A_s[20] ), .ZN(n544) );
  INV_X1 U204 ( .A(A_ns[20]), .ZN(n543) );
  OAI221_X1 U205 ( .B1(n393), .B2(n546), .C1(n392), .C2(n547), .A(n548), .ZN(
        O[21]) );
  AOI22_X1 U206 ( .A1(A_ns[20]), .A2(n397), .B1(\A_s[20] ), .B2(n398), .ZN(
        n548) );
  INV_X1 U207 ( .A(\A_s[19] ), .ZN(n547) );
  INV_X1 U208 ( .A(A_ns[19]), .ZN(n546) );
  OAI221_X1 U209 ( .B1(n393), .B2(n549), .C1(n392), .C2(n550), .A(n551), .ZN(
        O[20]) );
  AOI22_X1 U210 ( .A1(A_ns[19]), .A2(n397), .B1(\A_s[19] ), .B2(n398), .ZN(
        n551) );
  INV_X1 U211 ( .A(\A_s[18] ), .ZN(n550) );
  INV_X1 U212 ( .A(A_ns[18]), .ZN(n549) );
  OAI22_X1 U213 ( .A1(n552), .A2(n520), .B1(n553), .B2(n519), .ZN(O[1]) );
  INV_X1 U214 ( .A(A_ns[0]), .ZN(n519) );
  INV_X1 U215 ( .A(\A_s[0] ), .ZN(n520) );
  OAI221_X1 U216 ( .B1(n393), .B2(n554), .C1(n392), .C2(n555), .A(n556), .ZN(
        O[19]) );
  AOI22_X1 U217 ( .A1(A_ns[18]), .A2(n397), .B1(\A_s[18] ), .B2(n398), .ZN(
        n556) );
  INV_X1 U218 ( .A(\A_s[17] ), .ZN(n555) );
  INV_X1 U219 ( .A(A_ns[17]), .ZN(n554) );
  OAI221_X1 U220 ( .B1(n393), .B2(n557), .C1(n392), .C2(n558), .A(n559), .ZN(
        O[18]) );
  AOI22_X1 U221 ( .A1(A_ns[17]), .A2(n397), .B1(\A_s[17] ), .B2(n398), .ZN(
        n559) );
  INV_X1 U222 ( .A(\A_s[16] ), .ZN(n558) );
  INV_X1 U223 ( .A(A_ns[16]), .ZN(n557) );
  OAI221_X1 U224 ( .B1(n393), .B2(n560), .C1(n392), .C2(n561), .A(n562), .ZN(
        O[17]) );
  AOI22_X1 U225 ( .A1(A_ns[16]), .A2(n397), .B1(\A_s[16] ), .B2(n398), .ZN(
        n562) );
  INV_X1 U226 ( .A(\A_s[15] ), .ZN(n561) );
  INV_X1 U227 ( .A(A_ns[15]), .ZN(n560) );
  OAI221_X1 U228 ( .B1(n393), .B2(n563), .C1(n392), .C2(n564), .A(n565), .ZN(
        O[16]) );
  AOI22_X1 U229 ( .A1(A_ns[15]), .A2(n397), .B1(\A_s[15] ), .B2(n398), .ZN(
        n565) );
  INV_X1 U230 ( .A(\A_s[14] ), .ZN(n564) );
  INV_X1 U231 ( .A(A_ns[14]), .ZN(n563) );
  OAI221_X1 U232 ( .B1(n393), .B2(n566), .C1(n392), .C2(n567), .A(n568), .ZN(
        O[15]) );
  AOI22_X1 U233 ( .A1(A_ns[14]), .A2(n397), .B1(\A_s[14] ), .B2(n398), .ZN(
        n568) );
  INV_X1 U234 ( .A(\A_s[13] ), .ZN(n567) );
  INV_X1 U235 ( .A(A_ns[13]), .ZN(n566) );
  OAI221_X1 U236 ( .B1(n393), .B2(n569), .C1(n392), .C2(n570), .A(n571), .ZN(
        O[14]) );
  AOI22_X1 U237 ( .A1(A_ns[13]), .A2(n397), .B1(\A_s[13] ), .B2(n398), .ZN(
        n571) );
  INV_X1 U238 ( .A(\A_s[12] ), .ZN(n570) );
  INV_X1 U239 ( .A(A_ns[12]), .ZN(n569) );
  OAI221_X1 U240 ( .B1(n393), .B2(n572), .C1(n392), .C2(n573), .A(n574), .ZN(
        O[13]) );
  AOI22_X1 U241 ( .A1(A_ns[12]), .A2(n397), .B1(\A_s[12] ), .B2(n398), .ZN(
        n574) );
  INV_X1 U242 ( .A(\A_s[11] ), .ZN(n573) );
  INV_X1 U243 ( .A(A_ns[11]), .ZN(n572) );
  OAI221_X1 U244 ( .B1(n393), .B2(n575), .C1(n392), .C2(n576), .A(n577), .ZN(
        O[12]) );
  AOI22_X1 U245 ( .A1(A_ns[11]), .A2(n397), .B1(\A_s[11] ), .B2(n398), .ZN(
        n577) );
  INV_X1 U246 ( .A(\A_s[10] ), .ZN(n576) );
  INV_X1 U247 ( .A(A_ns[10]), .ZN(n575) );
  OAI221_X1 U248 ( .B1(n393), .B2(n578), .C1(n392), .C2(n579), .A(n580), .ZN(
        O[11]) );
  AOI22_X1 U249 ( .A1(A_ns[10]), .A2(n397), .B1(\A_s[10] ), .B2(n398), .ZN(
        n580) );
  INV_X1 U250 ( .A(\A_s[9] ), .ZN(n579) );
  INV_X1 U251 ( .A(A_ns[9]), .ZN(n578) );
  OAI221_X1 U252 ( .B1(n581), .B2(n393), .C1(n582), .C2(n392), .A(n583), .ZN(
        O[10]) );
  AOI22_X1 U253 ( .A1(A_ns[9]), .A2(n397), .B1(\A_s[9] ), .B2(n398), .ZN(n583)
         );
  NAND2_X1 U254 ( .A1(n584), .A2(n552), .ZN(n553) );
  NAND2_X1 U255 ( .A1(n584), .A2(n585), .ZN(n552) );
  XOR2_X1 U256 ( .A(B[25]), .B(B[26]), .Z(n584) );
  INV_X1 U257 ( .A(\A_s[8] ), .ZN(n582) );
  INV_X1 U258 ( .A(B[27]), .ZN(n585) );
  INV_X1 U259 ( .A(A_ns[8]), .ZN(n581) );
endmodule


module BOOTHENC_NBIT64_i28 ( A, A_n, A_ns, A_s, B, O, A_so, A_nso );
  input [63:0] A;
  input [63:0] A_n;
  input [63:0] A_ns;
  input [63:0] A_s;
  input [63:0] B;
  output [63:0] O;
  output [63:0] A_so;
  output [63:0] A_nso;
  wire   \A_s[61] , \A_s[60] , \A_s[59] , \A_s[58] , \A_s[57] , \A_s[56] ,
         \A_s[55] , \A_s[54] , \A_s[53] , \A_s[52] , \A_s[51] , \A_s[50] ,
         \A_s[49] , \A_s[48] , \A_s[47] , \A_s[46] , \A_s[45] , \A_s[44] ,
         \A_s[43] , \A_s[42] , \A_s[41] , \A_s[40] , \A_s[39] , \A_s[38] ,
         \A_s[37] , \A_s[36] , \A_s[35] , \A_s[34] , \A_s[33] , \A_s[32] ,
         \A_s[31] , \A_s[30] , \A_s[29] , \A_s[28] , \A_s[27] , \A_s[26] ,
         \A_s[25] , \A_s[24] , \A_s[23] , \A_s[22] , \A_s[21] , \A_s[20] ,
         \A_s[19] , \A_s[18] , \A_s[17] , \A_s[16] , \A_s[15] , \A_s[14] ,
         \A_s[13] , \A_s[12] , \A_s[11] , \A_s[10] , \A_s[9] , \A_s[8] ,
         \A_s[7] , \A_s[6] , \A_s[5] , \A_s[4] , \A_s[3] , \A_s[2] , \A_s[1] ,
         \A_s[0] , n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585;
  assign A_nso[0] = 1'b0;
  assign A_nso[1] = 1'b0;
  assign A_so[0] = 1'b0;
  assign A_so[1] = 1'b0;
  assign O[0] = 1'b0;
  assign A_nso[63] = \A_s[61] ;
  assign A_so[63] = \A_s[61] ;
  assign \A_s[61]  = A_s[61];
  assign A_nso[62] = \A_s[60] ;
  assign A_so[62] = \A_s[60] ;
  assign \A_s[60]  = A_s[60];
  assign A_nso[61] = \A_s[59] ;
  assign A_so[61] = \A_s[59] ;
  assign \A_s[59]  = A_s[59];
  assign A_nso[60] = \A_s[58] ;
  assign A_so[60] = \A_s[58] ;
  assign \A_s[58]  = A_s[58];
  assign A_nso[59] = \A_s[57] ;
  assign A_so[59] = \A_s[57] ;
  assign \A_s[57]  = A_s[57];
  assign A_nso[58] = \A_s[56] ;
  assign A_so[58] = \A_s[56] ;
  assign \A_s[56]  = A_s[56];
  assign A_nso[57] = \A_s[55] ;
  assign A_so[57] = \A_s[55] ;
  assign \A_s[55]  = A_s[55];
  assign A_nso[56] = \A_s[54] ;
  assign A_so[56] = \A_s[54] ;
  assign \A_s[54]  = A_s[54];
  assign A_nso[55] = \A_s[53] ;
  assign A_so[55] = \A_s[53] ;
  assign \A_s[53]  = A_s[53];
  assign A_nso[54] = \A_s[52] ;
  assign A_so[54] = \A_s[52] ;
  assign \A_s[52]  = A_s[52];
  assign A_nso[53] = \A_s[51] ;
  assign A_so[53] = \A_s[51] ;
  assign \A_s[51]  = A_s[51];
  assign A_nso[52] = \A_s[50] ;
  assign A_so[52] = \A_s[50] ;
  assign \A_s[50]  = A_s[50];
  assign A_nso[51] = \A_s[49] ;
  assign A_so[51] = \A_s[49] ;
  assign \A_s[49]  = A_s[49];
  assign A_nso[50] = \A_s[48] ;
  assign A_so[50] = \A_s[48] ;
  assign \A_s[48]  = A_s[48];
  assign A_nso[49] = \A_s[47] ;
  assign A_so[49] = \A_s[47] ;
  assign \A_s[47]  = A_s[47];
  assign A_nso[48] = \A_s[46] ;
  assign A_so[48] = \A_s[46] ;
  assign \A_s[46]  = A_s[46];
  assign A_nso[47] = \A_s[45] ;
  assign A_so[47] = \A_s[45] ;
  assign \A_s[45]  = A_s[45];
  assign A_nso[46] = \A_s[44] ;
  assign A_so[46] = \A_s[44] ;
  assign \A_s[44]  = A_s[44];
  assign A_nso[45] = \A_s[43] ;
  assign A_so[45] = \A_s[43] ;
  assign \A_s[43]  = A_s[43];
  assign A_nso[44] = \A_s[42] ;
  assign A_so[44] = \A_s[42] ;
  assign \A_s[42]  = A_s[42];
  assign A_nso[43] = \A_s[41] ;
  assign A_so[43] = \A_s[41] ;
  assign \A_s[41]  = A_s[41];
  assign A_nso[42] = \A_s[40] ;
  assign A_so[42] = \A_s[40] ;
  assign \A_s[40]  = A_s[40];
  assign A_nso[41] = \A_s[39] ;
  assign A_so[41] = \A_s[39] ;
  assign \A_s[39]  = A_s[39];
  assign A_nso[40] = \A_s[38] ;
  assign A_so[40] = \A_s[38] ;
  assign \A_s[38]  = A_s[38];
  assign A_nso[39] = \A_s[37] ;
  assign A_so[39] = \A_s[37] ;
  assign \A_s[37]  = A_s[37];
  assign A_nso[38] = \A_s[36] ;
  assign A_so[38] = \A_s[36] ;
  assign \A_s[36]  = A_s[36];
  assign A_nso[37] = \A_s[35] ;
  assign A_so[37] = \A_s[35] ;
  assign \A_s[35]  = A_s[35];
  assign A_nso[36] = \A_s[34] ;
  assign A_so[36] = \A_s[34] ;
  assign \A_s[34]  = A_s[34];
  assign A_nso[35] = \A_s[33] ;
  assign A_so[35] = \A_s[33] ;
  assign \A_s[33]  = A_s[33];
  assign A_nso[34] = \A_s[32] ;
  assign A_so[34] = \A_s[32] ;
  assign \A_s[32]  = A_s[32];
  assign A_nso[33] = \A_s[31] ;
  assign A_so[33] = \A_s[31] ;
  assign \A_s[31]  = A_s[31];
  assign A_nso[32] = \A_s[30] ;
  assign A_so[32] = \A_s[30] ;
  assign \A_s[30]  = A_s[30];
  assign A_nso[31] = \A_s[29] ;
  assign A_so[31] = \A_s[29] ;
  assign \A_s[29]  = A_s[29];
  assign A_nso[30] = \A_s[28] ;
  assign A_so[30] = \A_s[28] ;
  assign \A_s[28]  = A_s[28];
  assign A_nso[29] = \A_s[27] ;
  assign A_so[29] = \A_s[27] ;
  assign \A_s[27]  = A_s[27];
  assign A_nso[28] = \A_s[26] ;
  assign A_so[28] = \A_s[26] ;
  assign \A_s[26]  = A_s[26];
  assign A_nso[27] = \A_s[25] ;
  assign A_so[27] = \A_s[25] ;
  assign \A_s[25]  = A_s[25];
  assign A_nso[26] = \A_s[24] ;
  assign A_so[26] = \A_s[24] ;
  assign \A_s[24]  = A_s[24];
  assign A_nso[25] = \A_s[23] ;
  assign A_so[25] = \A_s[23] ;
  assign \A_s[23]  = A_s[23];
  assign A_nso[24] = \A_s[22] ;
  assign A_so[24] = \A_s[22] ;
  assign \A_s[22]  = A_s[22];
  assign A_nso[23] = \A_s[21] ;
  assign A_so[23] = \A_s[21] ;
  assign \A_s[21]  = A_s[21];
  assign A_nso[22] = \A_s[20] ;
  assign A_so[22] = \A_s[20] ;
  assign \A_s[20]  = A_s[20];
  assign A_nso[21] = \A_s[19] ;
  assign A_so[21] = \A_s[19] ;
  assign \A_s[19]  = A_s[19];
  assign A_nso[20] = \A_s[18] ;
  assign A_so[20] = \A_s[18] ;
  assign \A_s[18]  = A_s[18];
  assign A_nso[19] = \A_s[17] ;
  assign A_so[19] = \A_s[17] ;
  assign \A_s[17]  = A_s[17];
  assign A_nso[18] = \A_s[16] ;
  assign A_so[18] = \A_s[16] ;
  assign \A_s[16]  = A_s[16];
  assign A_nso[17] = \A_s[15] ;
  assign A_so[17] = \A_s[15] ;
  assign \A_s[15]  = A_s[15];
  assign A_nso[16] = \A_s[14] ;
  assign A_so[16] = \A_s[14] ;
  assign \A_s[14]  = A_s[14];
  assign A_nso[15] = \A_s[13] ;
  assign A_so[15] = \A_s[13] ;
  assign \A_s[13]  = A_s[13];
  assign A_nso[14] = \A_s[12] ;
  assign A_so[14] = \A_s[12] ;
  assign \A_s[12]  = A_s[12];
  assign A_nso[13] = \A_s[11] ;
  assign A_so[13] = \A_s[11] ;
  assign \A_s[11]  = A_s[11];
  assign A_nso[12] = \A_s[10] ;
  assign A_so[12] = \A_s[10] ;
  assign \A_s[10]  = A_s[10];
  assign A_nso[11] = \A_s[9] ;
  assign A_so[11] = \A_s[9] ;
  assign \A_s[9]  = A_s[9];
  assign A_nso[10] = \A_s[8] ;
  assign A_so[10] = \A_s[8] ;
  assign \A_s[8]  = A_s[8];
  assign A_nso[9] = \A_s[7] ;
  assign A_so[9] = \A_s[7] ;
  assign \A_s[7]  = A_s[7];
  assign A_nso[8] = \A_s[6] ;
  assign A_so[8] = \A_s[6] ;
  assign \A_s[6]  = A_s[6];
  assign A_nso[7] = \A_s[5] ;
  assign A_so[7] = \A_s[5] ;
  assign \A_s[5]  = A_s[5];
  assign A_nso[6] = \A_s[4] ;
  assign A_so[6] = \A_s[4] ;
  assign \A_s[4]  = A_s[4];
  assign A_nso[5] = \A_s[3] ;
  assign A_so[5] = \A_s[3] ;
  assign \A_s[3]  = A_s[3];
  assign A_nso[4] = \A_s[2] ;
  assign A_so[4] = \A_s[2] ;
  assign \A_s[2]  = A_s[2];
  assign A_nso[3] = \A_s[1] ;
  assign A_so[3] = \A_s[1] ;
  assign \A_s[1]  = A_s[1];
  assign A_nso[2] = \A_s[0] ;
  assign A_so[2] = \A_s[0] ;
  assign \A_s[0]  = A_s[0];

  AND3_X1 U2 ( .A1(B[28]), .A2(n585), .A3(B[27]), .ZN(n391) );
  INV_X4 U3 ( .A(n391), .ZN(n392) );
  INV_X4 U4 ( .A(n552), .ZN(n398) );
  OR3_X4 U5 ( .A1(B[27]), .A2(B[28]), .A3(n585), .ZN(n393) );
  INV_X4 U6 ( .A(n553), .ZN(n397) );
  OAI221_X1 U7 ( .B1(n393), .B2(n394), .C1(n392), .C2(n395), .A(n396), .ZN(
        O[9]) );
  AOI22_X1 U8 ( .A1(A_ns[8]), .A2(n397), .B1(\A_s[8] ), .B2(n398), .ZN(n396)
         );
  INV_X1 U9 ( .A(\A_s[7] ), .ZN(n395) );
  INV_X1 U10 ( .A(A_ns[7]), .ZN(n394) );
  OAI221_X1 U11 ( .B1(n393), .B2(n399), .C1(n392), .C2(n400), .A(n401), .ZN(
        O[8]) );
  AOI22_X1 U12 ( .A1(A_ns[7]), .A2(n397), .B1(\A_s[7] ), .B2(n398), .ZN(n401)
         );
  INV_X1 U13 ( .A(\A_s[6] ), .ZN(n400) );
  INV_X1 U14 ( .A(A_ns[6]), .ZN(n399) );
  OAI221_X1 U15 ( .B1(n393), .B2(n402), .C1(n392), .C2(n403), .A(n404), .ZN(
        O[7]) );
  AOI22_X1 U16 ( .A1(A_ns[6]), .A2(n397), .B1(\A_s[6] ), .B2(n398), .ZN(n404)
         );
  INV_X1 U17 ( .A(\A_s[5] ), .ZN(n403) );
  INV_X1 U18 ( .A(A_ns[5]), .ZN(n402) );
  OAI221_X1 U19 ( .B1(n393), .B2(n405), .C1(n392), .C2(n406), .A(n407), .ZN(
        O[6]) );
  AOI22_X1 U20 ( .A1(A_ns[5]), .A2(n397), .B1(\A_s[5] ), .B2(n398), .ZN(n407)
         );
  INV_X1 U21 ( .A(\A_s[4] ), .ZN(n406) );
  INV_X1 U22 ( .A(A_ns[4]), .ZN(n405) );
  OAI221_X1 U23 ( .B1(n393), .B2(n408), .C1(n392), .C2(n409), .A(n410), .ZN(
        O[63]) );
  AOI22_X1 U24 ( .A1(A_ns[62]), .A2(n397), .B1(A_s[62]), .B2(n398), .ZN(n410)
         );
  INV_X1 U25 ( .A(\A_s[61] ), .ZN(n409) );
  INV_X1 U26 ( .A(A_ns[61]), .ZN(n408) );
  OAI221_X1 U27 ( .B1(n393), .B2(n411), .C1(n392), .C2(n412), .A(n413), .ZN(
        O[62]) );
  AOI22_X1 U28 ( .A1(A_ns[61]), .A2(n397), .B1(\A_s[61] ), .B2(n398), .ZN(n413) );
  INV_X1 U29 ( .A(\A_s[60] ), .ZN(n412) );
  INV_X1 U30 ( .A(A_ns[60]), .ZN(n411) );
  OAI221_X1 U31 ( .B1(n393), .B2(n414), .C1(n392), .C2(n415), .A(n416), .ZN(
        O[61]) );
  AOI22_X1 U32 ( .A1(A_ns[60]), .A2(n397), .B1(\A_s[60] ), .B2(n398), .ZN(n416) );
  INV_X1 U33 ( .A(\A_s[59] ), .ZN(n415) );
  INV_X1 U34 ( .A(A_ns[59]), .ZN(n414) );
  OAI221_X1 U35 ( .B1(n393), .B2(n417), .C1(n392), .C2(n418), .A(n419), .ZN(
        O[60]) );
  AOI22_X1 U36 ( .A1(A_ns[59]), .A2(n397), .B1(\A_s[59] ), .B2(n398), .ZN(n419) );
  INV_X1 U37 ( .A(\A_s[58] ), .ZN(n418) );
  INV_X1 U38 ( .A(A_ns[58]), .ZN(n417) );
  OAI221_X1 U39 ( .B1(n393), .B2(n420), .C1(n392), .C2(n421), .A(n422), .ZN(
        O[5]) );
  AOI22_X1 U40 ( .A1(A_ns[4]), .A2(n397), .B1(\A_s[4] ), .B2(n398), .ZN(n422)
         );
  INV_X1 U41 ( .A(\A_s[3] ), .ZN(n421) );
  INV_X1 U42 ( .A(A_ns[3]), .ZN(n420) );
  OAI221_X1 U43 ( .B1(n393), .B2(n423), .C1(n392), .C2(n424), .A(n425), .ZN(
        O[59]) );
  AOI22_X1 U44 ( .A1(A_ns[58]), .A2(n397), .B1(\A_s[58] ), .B2(n398), .ZN(n425) );
  INV_X1 U45 ( .A(\A_s[57] ), .ZN(n424) );
  INV_X1 U46 ( .A(A_ns[57]), .ZN(n423) );
  OAI221_X1 U47 ( .B1(n393), .B2(n426), .C1(n392), .C2(n427), .A(n428), .ZN(
        O[58]) );
  AOI22_X1 U48 ( .A1(A_ns[57]), .A2(n397), .B1(\A_s[57] ), .B2(n398), .ZN(n428) );
  INV_X1 U49 ( .A(\A_s[56] ), .ZN(n427) );
  INV_X1 U50 ( .A(A_ns[56]), .ZN(n426) );
  OAI221_X1 U51 ( .B1(n393), .B2(n429), .C1(n392), .C2(n430), .A(n431), .ZN(
        O[57]) );
  AOI22_X1 U52 ( .A1(A_ns[56]), .A2(n397), .B1(\A_s[56] ), .B2(n398), .ZN(n431) );
  INV_X1 U53 ( .A(\A_s[55] ), .ZN(n430) );
  INV_X1 U54 ( .A(A_ns[55]), .ZN(n429) );
  OAI221_X1 U55 ( .B1(n393), .B2(n432), .C1(n392), .C2(n433), .A(n434), .ZN(
        O[56]) );
  AOI22_X1 U56 ( .A1(A_ns[55]), .A2(n397), .B1(\A_s[55] ), .B2(n398), .ZN(n434) );
  INV_X1 U57 ( .A(\A_s[54] ), .ZN(n433) );
  INV_X1 U58 ( .A(A_ns[54]), .ZN(n432) );
  OAI221_X1 U59 ( .B1(n393), .B2(n435), .C1(n392), .C2(n436), .A(n437), .ZN(
        O[55]) );
  AOI22_X1 U60 ( .A1(A_ns[54]), .A2(n397), .B1(\A_s[54] ), .B2(n398), .ZN(n437) );
  INV_X1 U61 ( .A(\A_s[53] ), .ZN(n436) );
  INV_X1 U62 ( .A(A_ns[53]), .ZN(n435) );
  OAI221_X1 U63 ( .B1(n393), .B2(n438), .C1(n392), .C2(n439), .A(n440), .ZN(
        O[54]) );
  AOI22_X1 U64 ( .A1(A_ns[53]), .A2(n397), .B1(\A_s[53] ), .B2(n398), .ZN(n440) );
  INV_X1 U65 ( .A(\A_s[52] ), .ZN(n439) );
  INV_X1 U66 ( .A(A_ns[52]), .ZN(n438) );
  OAI221_X1 U67 ( .B1(n393), .B2(n441), .C1(n392), .C2(n442), .A(n443), .ZN(
        O[53]) );
  AOI22_X1 U68 ( .A1(A_ns[52]), .A2(n397), .B1(\A_s[52] ), .B2(n398), .ZN(n443) );
  INV_X1 U69 ( .A(\A_s[51] ), .ZN(n442) );
  INV_X1 U70 ( .A(A_ns[51]), .ZN(n441) );
  OAI221_X1 U71 ( .B1(n393), .B2(n444), .C1(n392), .C2(n445), .A(n446), .ZN(
        O[52]) );
  AOI22_X1 U72 ( .A1(A_ns[51]), .A2(n397), .B1(\A_s[51] ), .B2(n398), .ZN(n446) );
  INV_X1 U73 ( .A(\A_s[50] ), .ZN(n445) );
  INV_X1 U74 ( .A(A_ns[50]), .ZN(n444) );
  OAI221_X1 U75 ( .B1(n393), .B2(n447), .C1(n392), .C2(n448), .A(n449), .ZN(
        O[51]) );
  AOI22_X1 U76 ( .A1(A_ns[50]), .A2(n397), .B1(\A_s[50] ), .B2(n398), .ZN(n449) );
  INV_X1 U77 ( .A(\A_s[49] ), .ZN(n448) );
  INV_X1 U78 ( .A(A_ns[49]), .ZN(n447) );
  OAI221_X1 U79 ( .B1(n393), .B2(n450), .C1(n392), .C2(n451), .A(n452), .ZN(
        O[50]) );
  AOI22_X1 U80 ( .A1(A_ns[49]), .A2(n397), .B1(\A_s[49] ), .B2(n398), .ZN(n452) );
  INV_X1 U81 ( .A(\A_s[48] ), .ZN(n451) );
  INV_X1 U82 ( .A(A_ns[48]), .ZN(n450) );
  OAI221_X1 U83 ( .B1(n393), .B2(n453), .C1(n392), .C2(n454), .A(n455), .ZN(
        O[4]) );
  AOI22_X1 U84 ( .A1(A_ns[3]), .A2(n397), .B1(\A_s[3] ), .B2(n398), .ZN(n455)
         );
  INV_X1 U85 ( .A(\A_s[2] ), .ZN(n454) );
  INV_X1 U86 ( .A(A_ns[2]), .ZN(n453) );
  OAI221_X1 U87 ( .B1(n393), .B2(n456), .C1(n392), .C2(n457), .A(n458), .ZN(
        O[49]) );
  AOI22_X1 U88 ( .A1(A_ns[48]), .A2(n397), .B1(\A_s[48] ), .B2(n398), .ZN(n458) );
  INV_X1 U89 ( .A(\A_s[47] ), .ZN(n457) );
  INV_X1 U90 ( .A(A_ns[47]), .ZN(n456) );
  OAI221_X1 U91 ( .B1(n393), .B2(n459), .C1(n392), .C2(n460), .A(n461), .ZN(
        O[48]) );
  AOI22_X1 U92 ( .A1(A_ns[47]), .A2(n397), .B1(\A_s[47] ), .B2(n398), .ZN(n461) );
  INV_X1 U93 ( .A(\A_s[46] ), .ZN(n460) );
  INV_X1 U94 ( .A(A_ns[46]), .ZN(n459) );
  OAI221_X1 U95 ( .B1(n393), .B2(n462), .C1(n392), .C2(n463), .A(n464), .ZN(
        O[47]) );
  AOI22_X1 U96 ( .A1(A_ns[46]), .A2(n397), .B1(\A_s[46] ), .B2(n398), .ZN(n464) );
  INV_X1 U97 ( .A(\A_s[45] ), .ZN(n463) );
  INV_X1 U98 ( .A(A_ns[45]), .ZN(n462) );
  OAI221_X1 U99 ( .B1(n393), .B2(n465), .C1(n392), .C2(n466), .A(n467), .ZN(
        O[46]) );
  AOI22_X1 U100 ( .A1(A_ns[45]), .A2(n397), .B1(\A_s[45] ), .B2(n398), .ZN(
        n467) );
  INV_X1 U101 ( .A(\A_s[44] ), .ZN(n466) );
  INV_X1 U102 ( .A(A_ns[44]), .ZN(n465) );
  OAI221_X1 U103 ( .B1(n393), .B2(n468), .C1(n392), .C2(n469), .A(n470), .ZN(
        O[45]) );
  AOI22_X1 U104 ( .A1(A_ns[44]), .A2(n397), .B1(\A_s[44] ), .B2(n398), .ZN(
        n470) );
  INV_X1 U105 ( .A(\A_s[43] ), .ZN(n469) );
  INV_X1 U106 ( .A(A_ns[43]), .ZN(n468) );
  OAI221_X1 U107 ( .B1(n393), .B2(n471), .C1(n392), .C2(n472), .A(n473), .ZN(
        O[44]) );
  AOI22_X1 U108 ( .A1(A_ns[43]), .A2(n397), .B1(\A_s[43] ), .B2(n398), .ZN(
        n473) );
  INV_X1 U109 ( .A(\A_s[42] ), .ZN(n472) );
  INV_X1 U110 ( .A(A_ns[42]), .ZN(n471) );
  OAI221_X1 U111 ( .B1(n393), .B2(n474), .C1(n392), .C2(n475), .A(n476), .ZN(
        O[43]) );
  AOI22_X1 U112 ( .A1(A_ns[42]), .A2(n397), .B1(\A_s[42] ), .B2(n398), .ZN(
        n476) );
  INV_X1 U113 ( .A(\A_s[41] ), .ZN(n475) );
  INV_X1 U114 ( .A(A_ns[41]), .ZN(n474) );
  OAI221_X1 U115 ( .B1(n393), .B2(n477), .C1(n392), .C2(n478), .A(n479), .ZN(
        O[42]) );
  AOI22_X1 U116 ( .A1(A_ns[41]), .A2(n397), .B1(\A_s[41] ), .B2(n398), .ZN(
        n479) );
  INV_X1 U117 ( .A(\A_s[40] ), .ZN(n478) );
  INV_X1 U118 ( .A(A_ns[40]), .ZN(n477) );
  OAI221_X1 U119 ( .B1(n393), .B2(n480), .C1(n392), .C2(n481), .A(n482), .ZN(
        O[41]) );
  AOI22_X1 U120 ( .A1(A_ns[40]), .A2(n397), .B1(\A_s[40] ), .B2(n398), .ZN(
        n482) );
  INV_X1 U121 ( .A(\A_s[39] ), .ZN(n481) );
  INV_X1 U122 ( .A(A_ns[39]), .ZN(n480) );
  OAI221_X1 U123 ( .B1(n393), .B2(n483), .C1(n392), .C2(n484), .A(n485), .ZN(
        O[40]) );
  AOI22_X1 U124 ( .A1(A_ns[39]), .A2(n397), .B1(\A_s[39] ), .B2(n398), .ZN(
        n485) );
  INV_X1 U125 ( .A(\A_s[38] ), .ZN(n484) );
  INV_X1 U126 ( .A(A_ns[38]), .ZN(n483) );
  OAI221_X1 U127 ( .B1(n393), .B2(n486), .C1(n392), .C2(n487), .A(n488), .ZN(
        O[3]) );
  AOI22_X1 U128 ( .A1(A_ns[2]), .A2(n397), .B1(\A_s[2] ), .B2(n398), .ZN(n488)
         );
  INV_X1 U129 ( .A(\A_s[1] ), .ZN(n487) );
  INV_X1 U130 ( .A(A_ns[1]), .ZN(n486) );
  OAI221_X1 U131 ( .B1(n393), .B2(n489), .C1(n392), .C2(n490), .A(n491), .ZN(
        O[39]) );
  AOI22_X1 U132 ( .A1(A_ns[38]), .A2(n397), .B1(\A_s[38] ), .B2(n398), .ZN(
        n491) );
  INV_X1 U133 ( .A(\A_s[37] ), .ZN(n490) );
  INV_X1 U134 ( .A(A_ns[37]), .ZN(n489) );
  OAI221_X1 U135 ( .B1(n393), .B2(n492), .C1(n392), .C2(n493), .A(n494), .ZN(
        O[38]) );
  AOI22_X1 U136 ( .A1(A_ns[37]), .A2(n397), .B1(\A_s[37] ), .B2(n398), .ZN(
        n494) );
  INV_X1 U137 ( .A(\A_s[36] ), .ZN(n493) );
  INV_X1 U138 ( .A(A_ns[36]), .ZN(n492) );
  OAI221_X1 U139 ( .B1(n393), .B2(n495), .C1(n392), .C2(n496), .A(n497), .ZN(
        O[37]) );
  AOI22_X1 U140 ( .A1(A_ns[36]), .A2(n397), .B1(\A_s[36] ), .B2(n398), .ZN(
        n497) );
  INV_X1 U141 ( .A(\A_s[35] ), .ZN(n496) );
  INV_X1 U142 ( .A(A_ns[35]), .ZN(n495) );
  OAI221_X1 U143 ( .B1(n393), .B2(n498), .C1(n392), .C2(n499), .A(n500), .ZN(
        O[36]) );
  AOI22_X1 U144 ( .A1(A_ns[35]), .A2(n397), .B1(\A_s[35] ), .B2(n398), .ZN(
        n500) );
  INV_X1 U145 ( .A(\A_s[34] ), .ZN(n499) );
  INV_X1 U146 ( .A(A_ns[34]), .ZN(n498) );
  OAI221_X1 U147 ( .B1(n393), .B2(n501), .C1(n392), .C2(n502), .A(n503), .ZN(
        O[35]) );
  AOI22_X1 U148 ( .A1(A_ns[34]), .A2(n397), .B1(\A_s[34] ), .B2(n398), .ZN(
        n503) );
  INV_X1 U149 ( .A(\A_s[33] ), .ZN(n502) );
  INV_X1 U150 ( .A(A_ns[33]), .ZN(n501) );
  OAI221_X1 U151 ( .B1(n393), .B2(n504), .C1(n392), .C2(n505), .A(n506), .ZN(
        O[34]) );
  AOI22_X1 U152 ( .A1(A_ns[33]), .A2(n397), .B1(\A_s[33] ), .B2(n398), .ZN(
        n506) );
  INV_X1 U153 ( .A(\A_s[32] ), .ZN(n505) );
  INV_X1 U154 ( .A(A_ns[32]), .ZN(n504) );
  OAI221_X1 U155 ( .B1(n393), .B2(n507), .C1(n392), .C2(n508), .A(n509), .ZN(
        O[33]) );
  AOI22_X1 U156 ( .A1(A_ns[32]), .A2(n397), .B1(\A_s[32] ), .B2(n398), .ZN(
        n509) );
  INV_X1 U157 ( .A(\A_s[31] ), .ZN(n508) );
  INV_X1 U158 ( .A(A_ns[31]), .ZN(n507) );
  OAI221_X1 U159 ( .B1(n393), .B2(n510), .C1(n392), .C2(n511), .A(n512), .ZN(
        O[32]) );
  AOI22_X1 U160 ( .A1(A_ns[31]), .A2(n397), .B1(\A_s[31] ), .B2(n398), .ZN(
        n512) );
  INV_X1 U161 ( .A(\A_s[30] ), .ZN(n511) );
  INV_X1 U162 ( .A(A_ns[30]), .ZN(n510) );
  OAI221_X1 U163 ( .B1(n393), .B2(n513), .C1(n392), .C2(n514), .A(n515), .ZN(
        O[31]) );
  AOI22_X1 U164 ( .A1(A_ns[30]), .A2(n397), .B1(\A_s[30] ), .B2(n398), .ZN(
        n515) );
  INV_X1 U165 ( .A(\A_s[29] ), .ZN(n514) );
  INV_X1 U166 ( .A(A_ns[29]), .ZN(n513) );
  OAI221_X1 U167 ( .B1(n393), .B2(n516), .C1(n392), .C2(n517), .A(n518), .ZN(
        O[30]) );
  AOI22_X1 U168 ( .A1(A_ns[29]), .A2(n397), .B1(\A_s[29] ), .B2(n398), .ZN(
        n518) );
  INV_X1 U169 ( .A(\A_s[28] ), .ZN(n517) );
  INV_X1 U170 ( .A(A_ns[28]), .ZN(n516) );
  OAI221_X1 U171 ( .B1(n393), .B2(n519), .C1(n392), .C2(n520), .A(n521), .ZN(
        O[2]) );
  AOI22_X1 U172 ( .A1(A_ns[1]), .A2(n397), .B1(\A_s[1] ), .B2(n398), .ZN(n521)
         );
  OAI221_X1 U173 ( .B1(n393), .B2(n522), .C1(n392), .C2(n523), .A(n524), .ZN(
        O[29]) );
  AOI22_X1 U174 ( .A1(A_ns[28]), .A2(n397), .B1(\A_s[28] ), .B2(n398), .ZN(
        n524) );
  INV_X1 U175 ( .A(\A_s[27] ), .ZN(n523) );
  INV_X1 U176 ( .A(A_ns[27]), .ZN(n522) );
  OAI221_X1 U177 ( .B1(n393), .B2(n525), .C1(n392), .C2(n526), .A(n527), .ZN(
        O[28]) );
  AOI22_X1 U178 ( .A1(A_ns[27]), .A2(n397), .B1(\A_s[27] ), .B2(n398), .ZN(
        n527) );
  INV_X1 U179 ( .A(\A_s[26] ), .ZN(n526) );
  INV_X1 U180 ( .A(A_ns[26]), .ZN(n525) );
  OAI221_X1 U181 ( .B1(n393), .B2(n528), .C1(n392), .C2(n529), .A(n530), .ZN(
        O[27]) );
  AOI22_X1 U182 ( .A1(A_ns[26]), .A2(n397), .B1(\A_s[26] ), .B2(n398), .ZN(
        n530) );
  INV_X1 U183 ( .A(\A_s[25] ), .ZN(n529) );
  INV_X1 U184 ( .A(A_ns[25]), .ZN(n528) );
  OAI221_X1 U185 ( .B1(n393), .B2(n531), .C1(n392), .C2(n532), .A(n533), .ZN(
        O[26]) );
  AOI22_X1 U186 ( .A1(A_ns[25]), .A2(n397), .B1(\A_s[25] ), .B2(n398), .ZN(
        n533) );
  INV_X1 U187 ( .A(\A_s[24] ), .ZN(n532) );
  INV_X1 U188 ( .A(A_ns[24]), .ZN(n531) );
  OAI221_X1 U189 ( .B1(n393), .B2(n534), .C1(n392), .C2(n535), .A(n536), .ZN(
        O[25]) );
  AOI22_X1 U190 ( .A1(A_ns[24]), .A2(n397), .B1(\A_s[24] ), .B2(n398), .ZN(
        n536) );
  INV_X1 U191 ( .A(\A_s[23] ), .ZN(n535) );
  INV_X1 U192 ( .A(A_ns[23]), .ZN(n534) );
  OAI221_X1 U193 ( .B1(n393), .B2(n537), .C1(n392), .C2(n538), .A(n539), .ZN(
        O[24]) );
  AOI22_X1 U194 ( .A1(A_ns[23]), .A2(n397), .B1(\A_s[23] ), .B2(n398), .ZN(
        n539) );
  INV_X1 U195 ( .A(\A_s[22] ), .ZN(n538) );
  INV_X1 U196 ( .A(A_ns[22]), .ZN(n537) );
  OAI221_X1 U197 ( .B1(n393), .B2(n540), .C1(n392), .C2(n541), .A(n542), .ZN(
        O[23]) );
  AOI22_X1 U198 ( .A1(A_ns[22]), .A2(n397), .B1(\A_s[22] ), .B2(n398), .ZN(
        n542) );
  INV_X1 U199 ( .A(\A_s[21] ), .ZN(n541) );
  INV_X1 U200 ( .A(A_ns[21]), .ZN(n540) );
  OAI221_X1 U201 ( .B1(n393), .B2(n543), .C1(n392), .C2(n544), .A(n545), .ZN(
        O[22]) );
  AOI22_X1 U202 ( .A1(A_ns[21]), .A2(n397), .B1(\A_s[21] ), .B2(n398), .ZN(
        n545) );
  INV_X1 U203 ( .A(\A_s[20] ), .ZN(n544) );
  INV_X1 U204 ( .A(A_ns[20]), .ZN(n543) );
  OAI221_X1 U205 ( .B1(n393), .B2(n546), .C1(n392), .C2(n547), .A(n548), .ZN(
        O[21]) );
  AOI22_X1 U206 ( .A1(A_ns[20]), .A2(n397), .B1(\A_s[20] ), .B2(n398), .ZN(
        n548) );
  INV_X1 U207 ( .A(\A_s[19] ), .ZN(n547) );
  INV_X1 U208 ( .A(A_ns[19]), .ZN(n546) );
  OAI221_X1 U209 ( .B1(n393), .B2(n549), .C1(n392), .C2(n550), .A(n551), .ZN(
        O[20]) );
  AOI22_X1 U210 ( .A1(A_ns[19]), .A2(n397), .B1(\A_s[19] ), .B2(n398), .ZN(
        n551) );
  INV_X1 U211 ( .A(\A_s[18] ), .ZN(n550) );
  INV_X1 U212 ( .A(A_ns[18]), .ZN(n549) );
  OAI22_X1 U213 ( .A1(n552), .A2(n520), .B1(n553), .B2(n519), .ZN(O[1]) );
  INV_X1 U214 ( .A(A_ns[0]), .ZN(n519) );
  INV_X1 U215 ( .A(\A_s[0] ), .ZN(n520) );
  OAI221_X1 U216 ( .B1(n393), .B2(n554), .C1(n392), .C2(n555), .A(n556), .ZN(
        O[19]) );
  AOI22_X1 U217 ( .A1(A_ns[18]), .A2(n397), .B1(\A_s[18] ), .B2(n398), .ZN(
        n556) );
  INV_X1 U218 ( .A(\A_s[17] ), .ZN(n555) );
  INV_X1 U219 ( .A(A_ns[17]), .ZN(n554) );
  OAI221_X1 U220 ( .B1(n393), .B2(n557), .C1(n392), .C2(n558), .A(n559), .ZN(
        O[18]) );
  AOI22_X1 U221 ( .A1(A_ns[17]), .A2(n397), .B1(\A_s[17] ), .B2(n398), .ZN(
        n559) );
  INV_X1 U222 ( .A(\A_s[16] ), .ZN(n558) );
  INV_X1 U223 ( .A(A_ns[16]), .ZN(n557) );
  OAI221_X1 U224 ( .B1(n393), .B2(n560), .C1(n392), .C2(n561), .A(n562), .ZN(
        O[17]) );
  AOI22_X1 U225 ( .A1(A_ns[16]), .A2(n397), .B1(\A_s[16] ), .B2(n398), .ZN(
        n562) );
  INV_X1 U226 ( .A(\A_s[15] ), .ZN(n561) );
  INV_X1 U227 ( .A(A_ns[15]), .ZN(n560) );
  OAI221_X1 U228 ( .B1(n393), .B2(n563), .C1(n392), .C2(n564), .A(n565), .ZN(
        O[16]) );
  AOI22_X1 U229 ( .A1(A_ns[15]), .A2(n397), .B1(\A_s[15] ), .B2(n398), .ZN(
        n565) );
  INV_X1 U230 ( .A(\A_s[14] ), .ZN(n564) );
  INV_X1 U231 ( .A(A_ns[14]), .ZN(n563) );
  OAI221_X1 U232 ( .B1(n393), .B2(n566), .C1(n392), .C2(n567), .A(n568), .ZN(
        O[15]) );
  AOI22_X1 U233 ( .A1(A_ns[14]), .A2(n397), .B1(\A_s[14] ), .B2(n398), .ZN(
        n568) );
  INV_X1 U234 ( .A(\A_s[13] ), .ZN(n567) );
  INV_X1 U235 ( .A(A_ns[13]), .ZN(n566) );
  OAI221_X1 U236 ( .B1(n393), .B2(n569), .C1(n392), .C2(n570), .A(n571), .ZN(
        O[14]) );
  AOI22_X1 U237 ( .A1(A_ns[13]), .A2(n397), .B1(\A_s[13] ), .B2(n398), .ZN(
        n571) );
  INV_X1 U238 ( .A(\A_s[12] ), .ZN(n570) );
  INV_X1 U239 ( .A(A_ns[12]), .ZN(n569) );
  OAI221_X1 U240 ( .B1(n393), .B2(n572), .C1(n392), .C2(n573), .A(n574), .ZN(
        O[13]) );
  AOI22_X1 U241 ( .A1(A_ns[12]), .A2(n397), .B1(\A_s[12] ), .B2(n398), .ZN(
        n574) );
  INV_X1 U242 ( .A(\A_s[11] ), .ZN(n573) );
  INV_X1 U243 ( .A(A_ns[11]), .ZN(n572) );
  OAI221_X1 U244 ( .B1(n393), .B2(n575), .C1(n392), .C2(n576), .A(n577), .ZN(
        O[12]) );
  AOI22_X1 U245 ( .A1(A_ns[11]), .A2(n397), .B1(\A_s[11] ), .B2(n398), .ZN(
        n577) );
  INV_X1 U246 ( .A(\A_s[10] ), .ZN(n576) );
  INV_X1 U247 ( .A(A_ns[10]), .ZN(n575) );
  OAI221_X1 U248 ( .B1(n393), .B2(n578), .C1(n392), .C2(n579), .A(n580), .ZN(
        O[11]) );
  AOI22_X1 U249 ( .A1(A_ns[10]), .A2(n397), .B1(\A_s[10] ), .B2(n398), .ZN(
        n580) );
  INV_X1 U250 ( .A(\A_s[9] ), .ZN(n579) );
  INV_X1 U251 ( .A(A_ns[9]), .ZN(n578) );
  OAI221_X1 U252 ( .B1(n581), .B2(n393), .C1(n582), .C2(n392), .A(n583), .ZN(
        O[10]) );
  AOI22_X1 U253 ( .A1(A_ns[9]), .A2(n397), .B1(\A_s[9] ), .B2(n398), .ZN(n583)
         );
  NAND2_X1 U254 ( .A1(n584), .A2(n552), .ZN(n553) );
  NAND2_X1 U255 ( .A1(n584), .A2(n585), .ZN(n552) );
  XOR2_X1 U256 ( .A(B[27]), .B(B[28]), .Z(n584) );
  INV_X1 U257 ( .A(\A_s[8] ), .ZN(n582) );
  INV_X1 U258 ( .A(B[29]), .ZN(n585) );
  INV_X1 U259 ( .A(A_ns[8]), .ZN(n581) );
endmodule


module BOOTHENC_NBIT64_i30 ( A, A_n, A_ns, A_s, B, O, A_so, A_nso );
  input [63:0] A;
  input [63:0] A_n;
  input [63:0] A_ns;
  input [63:0] A_s;
  input [63:0] B;
  output [63:0] O;
  output [63:0] A_so;
  output [63:0] A_nso;
  wire   \A_s[61] , \A_s[60] , \A_s[59] , \A_s[58] , \A_s[57] , \A_s[56] ,
         \A_s[55] , \A_s[54] , \A_s[53] , \A_s[52] , \A_s[51] , \A_s[50] ,
         \A_s[49] , \A_s[48] , \A_s[47] , \A_s[46] , \A_s[45] , \A_s[44] ,
         \A_s[43] , \A_s[42] , \A_s[41] , \A_s[40] , \A_s[39] , \A_s[38] ,
         \A_s[37] , \A_s[36] , \A_s[35] , \A_s[34] , \A_s[33] , \A_s[32] ,
         \A_s[31] , \A_s[30] , \A_s[29] , \A_s[28] , \A_s[27] , \A_s[26] ,
         \A_s[25] , \A_s[24] , \A_s[23] , \A_s[22] , \A_s[21] , \A_s[20] ,
         \A_s[19] , \A_s[18] , \A_s[17] , \A_s[16] , \A_s[15] , \A_s[14] ,
         \A_s[13] , \A_s[12] , \A_s[11] , \A_s[10] , \A_s[9] , \A_s[8] ,
         \A_s[7] , \A_s[6] , \A_s[5] , \A_s[4] , \A_s[3] , \A_s[2] , \A_s[1] ,
         \A_s[0] , n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585;
  assign A_nso[0] = 1'b0;
  assign A_nso[1] = 1'b0;
  assign A_so[0] = 1'b0;
  assign A_so[1] = 1'b0;
  assign O[0] = 1'b0;
  assign A_nso[63] = \A_s[61] ;
  assign A_so[63] = \A_s[61] ;
  assign \A_s[61]  = A_s[61];
  assign A_nso[62] = \A_s[60] ;
  assign A_so[62] = \A_s[60] ;
  assign \A_s[60]  = A_s[60];
  assign A_nso[61] = \A_s[59] ;
  assign A_so[61] = \A_s[59] ;
  assign \A_s[59]  = A_s[59];
  assign A_nso[60] = \A_s[58] ;
  assign A_so[60] = \A_s[58] ;
  assign \A_s[58]  = A_s[58];
  assign A_nso[59] = \A_s[57] ;
  assign A_so[59] = \A_s[57] ;
  assign \A_s[57]  = A_s[57];
  assign A_nso[58] = \A_s[56] ;
  assign A_so[58] = \A_s[56] ;
  assign \A_s[56]  = A_s[56];
  assign A_nso[57] = \A_s[55] ;
  assign A_so[57] = \A_s[55] ;
  assign \A_s[55]  = A_s[55];
  assign A_nso[56] = \A_s[54] ;
  assign A_so[56] = \A_s[54] ;
  assign \A_s[54]  = A_s[54];
  assign A_nso[55] = \A_s[53] ;
  assign A_so[55] = \A_s[53] ;
  assign \A_s[53]  = A_s[53];
  assign A_nso[54] = \A_s[52] ;
  assign A_so[54] = \A_s[52] ;
  assign \A_s[52]  = A_s[52];
  assign A_nso[53] = \A_s[51] ;
  assign A_so[53] = \A_s[51] ;
  assign \A_s[51]  = A_s[51];
  assign A_nso[52] = \A_s[50] ;
  assign A_so[52] = \A_s[50] ;
  assign \A_s[50]  = A_s[50];
  assign A_nso[51] = \A_s[49] ;
  assign A_so[51] = \A_s[49] ;
  assign \A_s[49]  = A_s[49];
  assign A_nso[50] = \A_s[48] ;
  assign A_so[50] = \A_s[48] ;
  assign \A_s[48]  = A_s[48];
  assign A_nso[49] = \A_s[47] ;
  assign A_so[49] = \A_s[47] ;
  assign \A_s[47]  = A_s[47];
  assign A_nso[48] = \A_s[46] ;
  assign A_so[48] = \A_s[46] ;
  assign \A_s[46]  = A_s[46];
  assign A_nso[47] = \A_s[45] ;
  assign A_so[47] = \A_s[45] ;
  assign \A_s[45]  = A_s[45];
  assign A_nso[46] = \A_s[44] ;
  assign A_so[46] = \A_s[44] ;
  assign \A_s[44]  = A_s[44];
  assign A_nso[45] = \A_s[43] ;
  assign A_so[45] = \A_s[43] ;
  assign \A_s[43]  = A_s[43];
  assign A_nso[44] = \A_s[42] ;
  assign A_so[44] = \A_s[42] ;
  assign \A_s[42]  = A_s[42];
  assign A_nso[43] = \A_s[41] ;
  assign A_so[43] = \A_s[41] ;
  assign \A_s[41]  = A_s[41];
  assign A_nso[42] = \A_s[40] ;
  assign A_so[42] = \A_s[40] ;
  assign \A_s[40]  = A_s[40];
  assign A_nso[41] = \A_s[39] ;
  assign A_so[41] = \A_s[39] ;
  assign \A_s[39]  = A_s[39];
  assign A_nso[40] = \A_s[38] ;
  assign A_so[40] = \A_s[38] ;
  assign \A_s[38]  = A_s[38];
  assign A_nso[39] = \A_s[37] ;
  assign A_so[39] = \A_s[37] ;
  assign \A_s[37]  = A_s[37];
  assign A_nso[38] = \A_s[36] ;
  assign A_so[38] = \A_s[36] ;
  assign \A_s[36]  = A_s[36];
  assign A_nso[37] = \A_s[35] ;
  assign A_so[37] = \A_s[35] ;
  assign \A_s[35]  = A_s[35];
  assign A_nso[36] = \A_s[34] ;
  assign A_so[36] = \A_s[34] ;
  assign \A_s[34]  = A_s[34];
  assign A_nso[35] = \A_s[33] ;
  assign A_so[35] = \A_s[33] ;
  assign \A_s[33]  = A_s[33];
  assign A_nso[34] = \A_s[32] ;
  assign A_so[34] = \A_s[32] ;
  assign \A_s[32]  = A_s[32];
  assign A_nso[33] = \A_s[31] ;
  assign A_so[33] = \A_s[31] ;
  assign \A_s[31]  = A_s[31];
  assign A_nso[32] = \A_s[30] ;
  assign A_so[32] = \A_s[30] ;
  assign \A_s[30]  = A_s[30];
  assign A_nso[31] = \A_s[29] ;
  assign A_so[31] = \A_s[29] ;
  assign \A_s[29]  = A_s[29];
  assign A_nso[30] = \A_s[28] ;
  assign A_so[30] = \A_s[28] ;
  assign \A_s[28]  = A_s[28];
  assign A_nso[29] = \A_s[27] ;
  assign A_so[29] = \A_s[27] ;
  assign \A_s[27]  = A_s[27];
  assign A_nso[28] = \A_s[26] ;
  assign A_so[28] = \A_s[26] ;
  assign \A_s[26]  = A_s[26];
  assign A_nso[27] = \A_s[25] ;
  assign A_so[27] = \A_s[25] ;
  assign \A_s[25]  = A_s[25];
  assign A_nso[26] = \A_s[24] ;
  assign A_so[26] = \A_s[24] ;
  assign \A_s[24]  = A_s[24];
  assign A_nso[25] = \A_s[23] ;
  assign A_so[25] = \A_s[23] ;
  assign \A_s[23]  = A_s[23];
  assign A_nso[24] = \A_s[22] ;
  assign A_so[24] = \A_s[22] ;
  assign \A_s[22]  = A_s[22];
  assign A_nso[23] = \A_s[21] ;
  assign A_so[23] = \A_s[21] ;
  assign \A_s[21]  = A_s[21];
  assign A_nso[22] = \A_s[20] ;
  assign A_so[22] = \A_s[20] ;
  assign \A_s[20]  = A_s[20];
  assign A_nso[21] = \A_s[19] ;
  assign A_so[21] = \A_s[19] ;
  assign \A_s[19]  = A_s[19];
  assign A_nso[20] = \A_s[18] ;
  assign A_so[20] = \A_s[18] ;
  assign \A_s[18]  = A_s[18];
  assign A_nso[19] = \A_s[17] ;
  assign A_so[19] = \A_s[17] ;
  assign \A_s[17]  = A_s[17];
  assign A_nso[18] = \A_s[16] ;
  assign A_so[18] = \A_s[16] ;
  assign \A_s[16]  = A_s[16];
  assign A_nso[17] = \A_s[15] ;
  assign A_so[17] = \A_s[15] ;
  assign \A_s[15]  = A_s[15];
  assign A_nso[16] = \A_s[14] ;
  assign A_so[16] = \A_s[14] ;
  assign \A_s[14]  = A_s[14];
  assign A_nso[15] = \A_s[13] ;
  assign A_so[15] = \A_s[13] ;
  assign \A_s[13]  = A_s[13];
  assign A_nso[14] = \A_s[12] ;
  assign A_so[14] = \A_s[12] ;
  assign \A_s[12]  = A_s[12];
  assign A_nso[13] = \A_s[11] ;
  assign A_so[13] = \A_s[11] ;
  assign \A_s[11]  = A_s[11];
  assign A_nso[12] = \A_s[10] ;
  assign A_so[12] = \A_s[10] ;
  assign \A_s[10]  = A_s[10];
  assign A_nso[11] = \A_s[9] ;
  assign A_so[11] = \A_s[9] ;
  assign \A_s[9]  = A_s[9];
  assign A_nso[10] = \A_s[8] ;
  assign A_so[10] = \A_s[8] ;
  assign \A_s[8]  = A_s[8];
  assign A_nso[9] = \A_s[7] ;
  assign A_so[9] = \A_s[7] ;
  assign \A_s[7]  = A_s[7];
  assign A_nso[8] = \A_s[6] ;
  assign A_so[8] = \A_s[6] ;
  assign \A_s[6]  = A_s[6];
  assign A_nso[7] = \A_s[5] ;
  assign A_so[7] = \A_s[5] ;
  assign \A_s[5]  = A_s[5];
  assign A_nso[6] = \A_s[4] ;
  assign A_so[6] = \A_s[4] ;
  assign \A_s[4]  = A_s[4];
  assign A_nso[5] = \A_s[3] ;
  assign A_so[5] = \A_s[3] ;
  assign \A_s[3]  = A_s[3];
  assign A_nso[4] = \A_s[2] ;
  assign A_so[4] = \A_s[2] ;
  assign \A_s[2]  = A_s[2];
  assign A_nso[3] = \A_s[1] ;
  assign A_so[3] = \A_s[1] ;
  assign \A_s[1]  = A_s[1];
  assign A_nso[2] = \A_s[0] ;
  assign A_so[2] = \A_s[0] ;
  assign \A_s[0]  = A_s[0];

  AND3_X1 U2 ( .A1(B[30]), .A2(n585), .A3(B[29]), .ZN(n391) );
  INV_X4 U3 ( .A(n391), .ZN(n392) );
  INV_X4 U4 ( .A(n552), .ZN(n398) );
  OR3_X4 U5 ( .A1(B[29]), .A2(B[30]), .A3(n585), .ZN(n393) );
  INV_X4 U6 ( .A(n553), .ZN(n397) );
  OAI221_X1 U7 ( .B1(n393), .B2(n394), .C1(n392), .C2(n395), .A(n396), .ZN(
        O[9]) );
  AOI22_X1 U8 ( .A1(A_ns[8]), .A2(n397), .B1(\A_s[8] ), .B2(n398), .ZN(n396)
         );
  INV_X1 U9 ( .A(\A_s[7] ), .ZN(n395) );
  INV_X1 U10 ( .A(A_ns[7]), .ZN(n394) );
  OAI221_X1 U11 ( .B1(n393), .B2(n399), .C1(n392), .C2(n400), .A(n401), .ZN(
        O[8]) );
  AOI22_X1 U12 ( .A1(A_ns[7]), .A2(n397), .B1(\A_s[7] ), .B2(n398), .ZN(n401)
         );
  INV_X1 U13 ( .A(\A_s[6] ), .ZN(n400) );
  INV_X1 U14 ( .A(A_ns[6]), .ZN(n399) );
  OAI221_X1 U15 ( .B1(n393), .B2(n402), .C1(n392), .C2(n403), .A(n404), .ZN(
        O[7]) );
  AOI22_X1 U16 ( .A1(A_ns[6]), .A2(n397), .B1(\A_s[6] ), .B2(n398), .ZN(n404)
         );
  INV_X1 U17 ( .A(\A_s[5] ), .ZN(n403) );
  INV_X1 U18 ( .A(A_ns[5]), .ZN(n402) );
  OAI221_X1 U19 ( .B1(n393), .B2(n405), .C1(n392), .C2(n406), .A(n407), .ZN(
        O[6]) );
  AOI22_X1 U20 ( .A1(A_ns[5]), .A2(n397), .B1(\A_s[5] ), .B2(n398), .ZN(n407)
         );
  INV_X1 U21 ( .A(\A_s[4] ), .ZN(n406) );
  INV_X1 U22 ( .A(A_ns[4]), .ZN(n405) );
  OAI221_X1 U23 ( .B1(n393), .B2(n408), .C1(n392), .C2(n409), .A(n410), .ZN(
        O[63]) );
  AOI22_X1 U24 ( .A1(A_ns[62]), .A2(n397), .B1(A_s[62]), .B2(n398), .ZN(n410)
         );
  INV_X1 U25 ( .A(\A_s[61] ), .ZN(n409) );
  INV_X1 U26 ( .A(A_ns[61]), .ZN(n408) );
  OAI221_X1 U27 ( .B1(n393), .B2(n411), .C1(n392), .C2(n412), .A(n413), .ZN(
        O[62]) );
  AOI22_X1 U28 ( .A1(A_ns[61]), .A2(n397), .B1(\A_s[61] ), .B2(n398), .ZN(n413) );
  INV_X1 U29 ( .A(\A_s[60] ), .ZN(n412) );
  INV_X1 U30 ( .A(A_ns[60]), .ZN(n411) );
  OAI221_X1 U31 ( .B1(n393), .B2(n414), .C1(n392), .C2(n415), .A(n416), .ZN(
        O[61]) );
  AOI22_X1 U32 ( .A1(A_ns[60]), .A2(n397), .B1(\A_s[60] ), .B2(n398), .ZN(n416) );
  INV_X1 U33 ( .A(\A_s[59] ), .ZN(n415) );
  INV_X1 U34 ( .A(A_ns[59]), .ZN(n414) );
  OAI221_X1 U35 ( .B1(n393), .B2(n417), .C1(n392), .C2(n418), .A(n419), .ZN(
        O[60]) );
  AOI22_X1 U36 ( .A1(A_ns[59]), .A2(n397), .B1(\A_s[59] ), .B2(n398), .ZN(n419) );
  INV_X1 U37 ( .A(\A_s[58] ), .ZN(n418) );
  INV_X1 U38 ( .A(A_ns[58]), .ZN(n417) );
  OAI221_X1 U39 ( .B1(n393), .B2(n420), .C1(n392), .C2(n421), .A(n422), .ZN(
        O[5]) );
  AOI22_X1 U40 ( .A1(A_ns[4]), .A2(n397), .B1(\A_s[4] ), .B2(n398), .ZN(n422)
         );
  INV_X1 U41 ( .A(\A_s[3] ), .ZN(n421) );
  INV_X1 U42 ( .A(A_ns[3]), .ZN(n420) );
  OAI221_X1 U43 ( .B1(n393), .B2(n423), .C1(n392), .C2(n424), .A(n425), .ZN(
        O[59]) );
  AOI22_X1 U44 ( .A1(A_ns[58]), .A2(n397), .B1(\A_s[58] ), .B2(n398), .ZN(n425) );
  INV_X1 U45 ( .A(\A_s[57] ), .ZN(n424) );
  INV_X1 U46 ( .A(A_ns[57]), .ZN(n423) );
  OAI221_X1 U47 ( .B1(n393), .B2(n426), .C1(n392), .C2(n427), .A(n428), .ZN(
        O[58]) );
  AOI22_X1 U48 ( .A1(A_ns[57]), .A2(n397), .B1(\A_s[57] ), .B2(n398), .ZN(n428) );
  INV_X1 U49 ( .A(\A_s[56] ), .ZN(n427) );
  INV_X1 U50 ( .A(A_ns[56]), .ZN(n426) );
  OAI221_X1 U51 ( .B1(n393), .B2(n429), .C1(n392), .C2(n430), .A(n431), .ZN(
        O[57]) );
  AOI22_X1 U52 ( .A1(A_ns[56]), .A2(n397), .B1(\A_s[56] ), .B2(n398), .ZN(n431) );
  INV_X1 U53 ( .A(\A_s[55] ), .ZN(n430) );
  INV_X1 U54 ( .A(A_ns[55]), .ZN(n429) );
  OAI221_X1 U55 ( .B1(n393), .B2(n432), .C1(n392), .C2(n433), .A(n434), .ZN(
        O[56]) );
  AOI22_X1 U56 ( .A1(A_ns[55]), .A2(n397), .B1(\A_s[55] ), .B2(n398), .ZN(n434) );
  INV_X1 U57 ( .A(\A_s[54] ), .ZN(n433) );
  INV_X1 U58 ( .A(A_ns[54]), .ZN(n432) );
  OAI221_X1 U59 ( .B1(n393), .B2(n435), .C1(n392), .C2(n436), .A(n437), .ZN(
        O[55]) );
  AOI22_X1 U60 ( .A1(A_ns[54]), .A2(n397), .B1(\A_s[54] ), .B2(n398), .ZN(n437) );
  INV_X1 U61 ( .A(\A_s[53] ), .ZN(n436) );
  INV_X1 U62 ( .A(A_ns[53]), .ZN(n435) );
  OAI221_X1 U63 ( .B1(n393), .B2(n438), .C1(n392), .C2(n439), .A(n440), .ZN(
        O[54]) );
  AOI22_X1 U64 ( .A1(A_ns[53]), .A2(n397), .B1(\A_s[53] ), .B2(n398), .ZN(n440) );
  INV_X1 U65 ( .A(\A_s[52] ), .ZN(n439) );
  INV_X1 U66 ( .A(A_ns[52]), .ZN(n438) );
  OAI221_X1 U67 ( .B1(n393), .B2(n441), .C1(n392), .C2(n442), .A(n443), .ZN(
        O[53]) );
  AOI22_X1 U68 ( .A1(A_ns[52]), .A2(n397), .B1(\A_s[52] ), .B2(n398), .ZN(n443) );
  INV_X1 U69 ( .A(\A_s[51] ), .ZN(n442) );
  INV_X1 U70 ( .A(A_ns[51]), .ZN(n441) );
  OAI221_X1 U71 ( .B1(n393), .B2(n444), .C1(n392), .C2(n445), .A(n446), .ZN(
        O[52]) );
  AOI22_X1 U72 ( .A1(A_ns[51]), .A2(n397), .B1(\A_s[51] ), .B2(n398), .ZN(n446) );
  INV_X1 U73 ( .A(\A_s[50] ), .ZN(n445) );
  INV_X1 U74 ( .A(A_ns[50]), .ZN(n444) );
  OAI221_X1 U75 ( .B1(n393), .B2(n447), .C1(n392), .C2(n448), .A(n449), .ZN(
        O[51]) );
  AOI22_X1 U76 ( .A1(A_ns[50]), .A2(n397), .B1(\A_s[50] ), .B2(n398), .ZN(n449) );
  INV_X1 U77 ( .A(\A_s[49] ), .ZN(n448) );
  INV_X1 U78 ( .A(A_ns[49]), .ZN(n447) );
  OAI221_X1 U79 ( .B1(n393), .B2(n450), .C1(n392), .C2(n451), .A(n452), .ZN(
        O[50]) );
  AOI22_X1 U80 ( .A1(A_ns[49]), .A2(n397), .B1(\A_s[49] ), .B2(n398), .ZN(n452) );
  INV_X1 U81 ( .A(\A_s[48] ), .ZN(n451) );
  INV_X1 U82 ( .A(A_ns[48]), .ZN(n450) );
  OAI221_X1 U83 ( .B1(n393), .B2(n453), .C1(n392), .C2(n454), .A(n455), .ZN(
        O[4]) );
  AOI22_X1 U84 ( .A1(A_ns[3]), .A2(n397), .B1(\A_s[3] ), .B2(n398), .ZN(n455)
         );
  INV_X1 U85 ( .A(\A_s[2] ), .ZN(n454) );
  INV_X1 U86 ( .A(A_ns[2]), .ZN(n453) );
  OAI221_X1 U87 ( .B1(n393), .B2(n456), .C1(n392), .C2(n457), .A(n458), .ZN(
        O[49]) );
  AOI22_X1 U88 ( .A1(A_ns[48]), .A2(n397), .B1(\A_s[48] ), .B2(n398), .ZN(n458) );
  INV_X1 U89 ( .A(\A_s[47] ), .ZN(n457) );
  INV_X1 U90 ( .A(A_ns[47]), .ZN(n456) );
  OAI221_X1 U91 ( .B1(n393), .B2(n459), .C1(n392), .C2(n460), .A(n461), .ZN(
        O[48]) );
  AOI22_X1 U92 ( .A1(A_ns[47]), .A2(n397), .B1(\A_s[47] ), .B2(n398), .ZN(n461) );
  INV_X1 U93 ( .A(\A_s[46] ), .ZN(n460) );
  INV_X1 U94 ( .A(A_ns[46]), .ZN(n459) );
  OAI221_X1 U95 ( .B1(n393), .B2(n462), .C1(n392), .C2(n463), .A(n464), .ZN(
        O[47]) );
  AOI22_X1 U96 ( .A1(A_ns[46]), .A2(n397), .B1(\A_s[46] ), .B2(n398), .ZN(n464) );
  INV_X1 U97 ( .A(\A_s[45] ), .ZN(n463) );
  INV_X1 U98 ( .A(A_ns[45]), .ZN(n462) );
  OAI221_X1 U99 ( .B1(n393), .B2(n465), .C1(n392), .C2(n466), .A(n467), .ZN(
        O[46]) );
  AOI22_X1 U100 ( .A1(A_ns[45]), .A2(n397), .B1(\A_s[45] ), .B2(n398), .ZN(
        n467) );
  INV_X1 U101 ( .A(\A_s[44] ), .ZN(n466) );
  INV_X1 U102 ( .A(A_ns[44]), .ZN(n465) );
  OAI221_X1 U103 ( .B1(n393), .B2(n468), .C1(n392), .C2(n469), .A(n470), .ZN(
        O[45]) );
  AOI22_X1 U104 ( .A1(A_ns[44]), .A2(n397), .B1(\A_s[44] ), .B2(n398), .ZN(
        n470) );
  INV_X1 U105 ( .A(\A_s[43] ), .ZN(n469) );
  INV_X1 U106 ( .A(A_ns[43]), .ZN(n468) );
  OAI221_X1 U107 ( .B1(n393), .B2(n471), .C1(n392), .C2(n472), .A(n473), .ZN(
        O[44]) );
  AOI22_X1 U108 ( .A1(A_ns[43]), .A2(n397), .B1(\A_s[43] ), .B2(n398), .ZN(
        n473) );
  INV_X1 U109 ( .A(\A_s[42] ), .ZN(n472) );
  INV_X1 U110 ( .A(A_ns[42]), .ZN(n471) );
  OAI221_X1 U111 ( .B1(n393), .B2(n474), .C1(n392), .C2(n475), .A(n476), .ZN(
        O[43]) );
  AOI22_X1 U112 ( .A1(A_ns[42]), .A2(n397), .B1(\A_s[42] ), .B2(n398), .ZN(
        n476) );
  INV_X1 U113 ( .A(\A_s[41] ), .ZN(n475) );
  INV_X1 U114 ( .A(A_ns[41]), .ZN(n474) );
  OAI221_X1 U115 ( .B1(n393), .B2(n477), .C1(n392), .C2(n478), .A(n479), .ZN(
        O[42]) );
  AOI22_X1 U116 ( .A1(A_ns[41]), .A2(n397), .B1(\A_s[41] ), .B2(n398), .ZN(
        n479) );
  INV_X1 U117 ( .A(\A_s[40] ), .ZN(n478) );
  INV_X1 U118 ( .A(A_ns[40]), .ZN(n477) );
  OAI221_X1 U119 ( .B1(n393), .B2(n480), .C1(n392), .C2(n481), .A(n482), .ZN(
        O[41]) );
  AOI22_X1 U120 ( .A1(A_ns[40]), .A2(n397), .B1(\A_s[40] ), .B2(n398), .ZN(
        n482) );
  INV_X1 U121 ( .A(\A_s[39] ), .ZN(n481) );
  INV_X1 U122 ( .A(A_ns[39]), .ZN(n480) );
  OAI221_X1 U123 ( .B1(n393), .B2(n483), .C1(n392), .C2(n484), .A(n485), .ZN(
        O[40]) );
  AOI22_X1 U124 ( .A1(A_ns[39]), .A2(n397), .B1(\A_s[39] ), .B2(n398), .ZN(
        n485) );
  INV_X1 U125 ( .A(\A_s[38] ), .ZN(n484) );
  INV_X1 U126 ( .A(A_ns[38]), .ZN(n483) );
  OAI221_X1 U127 ( .B1(n393), .B2(n486), .C1(n392), .C2(n487), .A(n488), .ZN(
        O[3]) );
  AOI22_X1 U128 ( .A1(A_ns[2]), .A2(n397), .B1(\A_s[2] ), .B2(n398), .ZN(n488)
         );
  INV_X1 U129 ( .A(\A_s[1] ), .ZN(n487) );
  INV_X1 U130 ( .A(A_ns[1]), .ZN(n486) );
  OAI221_X1 U131 ( .B1(n393), .B2(n489), .C1(n392), .C2(n490), .A(n491), .ZN(
        O[39]) );
  AOI22_X1 U132 ( .A1(A_ns[38]), .A2(n397), .B1(\A_s[38] ), .B2(n398), .ZN(
        n491) );
  INV_X1 U133 ( .A(\A_s[37] ), .ZN(n490) );
  INV_X1 U134 ( .A(A_ns[37]), .ZN(n489) );
  OAI221_X1 U135 ( .B1(n393), .B2(n492), .C1(n392), .C2(n493), .A(n494), .ZN(
        O[38]) );
  AOI22_X1 U136 ( .A1(A_ns[37]), .A2(n397), .B1(\A_s[37] ), .B2(n398), .ZN(
        n494) );
  INV_X1 U137 ( .A(\A_s[36] ), .ZN(n493) );
  INV_X1 U138 ( .A(A_ns[36]), .ZN(n492) );
  OAI221_X1 U139 ( .B1(n393), .B2(n495), .C1(n392), .C2(n496), .A(n497), .ZN(
        O[37]) );
  AOI22_X1 U140 ( .A1(A_ns[36]), .A2(n397), .B1(\A_s[36] ), .B2(n398), .ZN(
        n497) );
  INV_X1 U141 ( .A(\A_s[35] ), .ZN(n496) );
  INV_X1 U142 ( .A(A_ns[35]), .ZN(n495) );
  OAI221_X1 U143 ( .B1(n393), .B2(n498), .C1(n392), .C2(n499), .A(n500), .ZN(
        O[36]) );
  AOI22_X1 U144 ( .A1(A_ns[35]), .A2(n397), .B1(\A_s[35] ), .B2(n398), .ZN(
        n500) );
  INV_X1 U145 ( .A(\A_s[34] ), .ZN(n499) );
  INV_X1 U146 ( .A(A_ns[34]), .ZN(n498) );
  OAI221_X1 U147 ( .B1(n393), .B2(n501), .C1(n392), .C2(n502), .A(n503), .ZN(
        O[35]) );
  AOI22_X1 U148 ( .A1(A_ns[34]), .A2(n397), .B1(\A_s[34] ), .B2(n398), .ZN(
        n503) );
  INV_X1 U149 ( .A(\A_s[33] ), .ZN(n502) );
  INV_X1 U150 ( .A(A_ns[33]), .ZN(n501) );
  OAI221_X1 U151 ( .B1(n393), .B2(n504), .C1(n392), .C2(n505), .A(n506), .ZN(
        O[34]) );
  AOI22_X1 U152 ( .A1(A_ns[33]), .A2(n397), .B1(\A_s[33] ), .B2(n398), .ZN(
        n506) );
  INV_X1 U153 ( .A(\A_s[32] ), .ZN(n505) );
  INV_X1 U154 ( .A(A_ns[32]), .ZN(n504) );
  OAI221_X1 U155 ( .B1(n393), .B2(n507), .C1(n392), .C2(n508), .A(n509), .ZN(
        O[33]) );
  AOI22_X1 U156 ( .A1(A_ns[32]), .A2(n397), .B1(\A_s[32] ), .B2(n398), .ZN(
        n509) );
  INV_X1 U157 ( .A(\A_s[31] ), .ZN(n508) );
  INV_X1 U158 ( .A(A_ns[31]), .ZN(n507) );
  OAI221_X1 U159 ( .B1(n393), .B2(n510), .C1(n392), .C2(n511), .A(n512), .ZN(
        O[32]) );
  AOI22_X1 U160 ( .A1(A_ns[31]), .A2(n397), .B1(\A_s[31] ), .B2(n398), .ZN(
        n512) );
  INV_X1 U161 ( .A(\A_s[30] ), .ZN(n511) );
  INV_X1 U162 ( .A(A_ns[30]), .ZN(n510) );
  OAI221_X1 U163 ( .B1(n393), .B2(n513), .C1(n392), .C2(n514), .A(n515), .ZN(
        O[31]) );
  AOI22_X1 U164 ( .A1(A_ns[30]), .A2(n397), .B1(\A_s[30] ), .B2(n398), .ZN(
        n515) );
  INV_X1 U165 ( .A(\A_s[29] ), .ZN(n514) );
  INV_X1 U166 ( .A(A_ns[29]), .ZN(n513) );
  OAI221_X1 U167 ( .B1(n393), .B2(n516), .C1(n392), .C2(n517), .A(n518), .ZN(
        O[30]) );
  AOI22_X1 U168 ( .A1(A_ns[29]), .A2(n397), .B1(\A_s[29] ), .B2(n398), .ZN(
        n518) );
  INV_X1 U169 ( .A(\A_s[28] ), .ZN(n517) );
  INV_X1 U170 ( .A(A_ns[28]), .ZN(n516) );
  OAI221_X1 U171 ( .B1(n393), .B2(n519), .C1(n392), .C2(n520), .A(n521), .ZN(
        O[2]) );
  AOI22_X1 U172 ( .A1(A_ns[1]), .A2(n397), .B1(\A_s[1] ), .B2(n398), .ZN(n521)
         );
  OAI221_X1 U173 ( .B1(n393), .B2(n522), .C1(n392), .C2(n523), .A(n524), .ZN(
        O[29]) );
  AOI22_X1 U174 ( .A1(A_ns[28]), .A2(n397), .B1(\A_s[28] ), .B2(n398), .ZN(
        n524) );
  INV_X1 U175 ( .A(\A_s[27] ), .ZN(n523) );
  INV_X1 U176 ( .A(A_ns[27]), .ZN(n522) );
  OAI221_X1 U177 ( .B1(n393), .B2(n525), .C1(n392), .C2(n526), .A(n527), .ZN(
        O[28]) );
  AOI22_X1 U178 ( .A1(A_ns[27]), .A2(n397), .B1(\A_s[27] ), .B2(n398), .ZN(
        n527) );
  INV_X1 U179 ( .A(\A_s[26] ), .ZN(n526) );
  INV_X1 U180 ( .A(A_ns[26]), .ZN(n525) );
  OAI221_X1 U181 ( .B1(n393), .B2(n528), .C1(n392), .C2(n529), .A(n530), .ZN(
        O[27]) );
  AOI22_X1 U182 ( .A1(A_ns[26]), .A2(n397), .B1(\A_s[26] ), .B2(n398), .ZN(
        n530) );
  INV_X1 U183 ( .A(\A_s[25] ), .ZN(n529) );
  INV_X1 U184 ( .A(A_ns[25]), .ZN(n528) );
  OAI221_X1 U185 ( .B1(n393), .B2(n531), .C1(n392), .C2(n532), .A(n533), .ZN(
        O[26]) );
  AOI22_X1 U186 ( .A1(A_ns[25]), .A2(n397), .B1(\A_s[25] ), .B2(n398), .ZN(
        n533) );
  INV_X1 U187 ( .A(\A_s[24] ), .ZN(n532) );
  INV_X1 U188 ( .A(A_ns[24]), .ZN(n531) );
  OAI221_X1 U189 ( .B1(n393), .B2(n534), .C1(n392), .C2(n535), .A(n536), .ZN(
        O[25]) );
  AOI22_X1 U190 ( .A1(A_ns[24]), .A2(n397), .B1(\A_s[24] ), .B2(n398), .ZN(
        n536) );
  INV_X1 U191 ( .A(\A_s[23] ), .ZN(n535) );
  INV_X1 U192 ( .A(A_ns[23]), .ZN(n534) );
  OAI221_X1 U193 ( .B1(n393), .B2(n537), .C1(n392), .C2(n538), .A(n539), .ZN(
        O[24]) );
  AOI22_X1 U194 ( .A1(A_ns[23]), .A2(n397), .B1(\A_s[23] ), .B2(n398), .ZN(
        n539) );
  INV_X1 U195 ( .A(\A_s[22] ), .ZN(n538) );
  INV_X1 U196 ( .A(A_ns[22]), .ZN(n537) );
  OAI221_X1 U197 ( .B1(n393), .B2(n540), .C1(n392), .C2(n541), .A(n542), .ZN(
        O[23]) );
  AOI22_X1 U198 ( .A1(A_ns[22]), .A2(n397), .B1(\A_s[22] ), .B2(n398), .ZN(
        n542) );
  INV_X1 U199 ( .A(\A_s[21] ), .ZN(n541) );
  INV_X1 U200 ( .A(A_ns[21]), .ZN(n540) );
  OAI221_X1 U201 ( .B1(n393), .B2(n543), .C1(n392), .C2(n544), .A(n545), .ZN(
        O[22]) );
  AOI22_X1 U202 ( .A1(A_ns[21]), .A2(n397), .B1(\A_s[21] ), .B2(n398), .ZN(
        n545) );
  INV_X1 U203 ( .A(\A_s[20] ), .ZN(n544) );
  INV_X1 U204 ( .A(A_ns[20]), .ZN(n543) );
  OAI221_X1 U205 ( .B1(n393), .B2(n546), .C1(n392), .C2(n547), .A(n548), .ZN(
        O[21]) );
  AOI22_X1 U206 ( .A1(A_ns[20]), .A2(n397), .B1(\A_s[20] ), .B2(n398), .ZN(
        n548) );
  INV_X1 U207 ( .A(\A_s[19] ), .ZN(n547) );
  INV_X1 U208 ( .A(A_ns[19]), .ZN(n546) );
  OAI221_X1 U209 ( .B1(n393), .B2(n549), .C1(n392), .C2(n550), .A(n551), .ZN(
        O[20]) );
  AOI22_X1 U210 ( .A1(A_ns[19]), .A2(n397), .B1(\A_s[19] ), .B2(n398), .ZN(
        n551) );
  INV_X1 U211 ( .A(\A_s[18] ), .ZN(n550) );
  INV_X1 U212 ( .A(A_ns[18]), .ZN(n549) );
  OAI22_X1 U213 ( .A1(n552), .A2(n520), .B1(n553), .B2(n519), .ZN(O[1]) );
  INV_X1 U214 ( .A(A_ns[0]), .ZN(n519) );
  INV_X1 U215 ( .A(\A_s[0] ), .ZN(n520) );
  OAI221_X1 U216 ( .B1(n393), .B2(n554), .C1(n392), .C2(n555), .A(n556), .ZN(
        O[19]) );
  AOI22_X1 U217 ( .A1(A_ns[18]), .A2(n397), .B1(\A_s[18] ), .B2(n398), .ZN(
        n556) );
  INV_X1 U218 ( .A(\A_s[17] ), .ZN(n555) );
  INV_X1 U219 ( .A(A_ns[17]), .ZN(n554) );
  OAI221_X1 U220 ( .B1(n393), .B2(n557), .C1(n392), .C2(n558), .A(n559), .ZN(
        O[18]) );
  AOI22_X1 U221 ( .A1(A_ns[17]), .A2(n397), .B1(\A_s[17] ), .B2(n398), .ZN(
        n559) );
  INV_X1 U222 ( .A(\A_s[16] ), .ZN(n558) );
  INV_X1 U223 ( .A(A_ns[16]), .ZN(n557) );
  OAI221_X1 U224 ( .B1(n393), .B2(n560), .C1(n392), .C2(n561), .A(n562), .ZN(
        O[17]) );
  AOI22_X1 U225 ( .A1(A_ns[16]), .A2(n397), .B1(\A_s[16] ), .B2(n398), .ZN(
        n562) );
  INV_X1 U226 ( .A(\A_s[15] ), .ZN(n561) );
  INV_X1 U227 ( .A(A_ns[15]), .ZN(n560) );
  OAI221_X1 U228 ( .B1(n393), .B2(n563), .C1(n392), .C2(n564), .A(n565), .ZN(
        O[16]) );
  AOI22_X1 U229 ( .A1(A_ns[15]), .A2(n397), .B1(\A_s[15] ), .B2(n398), .ZN(
        n565) );
  INV_X1 U230 ( .A(\A_s[14] ), .ZN(n564) );
  INV_X1 U231 ( .A(A_ns[14]), .ZN(n563) );
  OAI221_X1 U232 ( .B1(n393), .B2(n566), .C1(n392), .C2(n567), .A(n568), .ZN(
        O[15]) );
  AOI22_X1 U233 ( .A1(A_ns[14]), .A2(n397), .B1(\A_s[14] ), .B2(n398), .ZN(
        n568) );
  INV_X1 U234 ( .A(\A_s[13] ), .ZN(n567) );
  INV_X1 U235 ( .A(A_ns[13]), .ZN(n566) );
  OAI221_X1 U236 ( .B1(n393), .B2(n569), .C1(n392), .C2(n570), .A(n571), .ZN(
        O[14]) );
  AOI22_X1 U237 ( .A1(A_ns[13]), .A2(n397), .B1(\A_s[13] ), .B2(n398), .ZN(
        n571) );
  INV_X1 U238 ( .A(\A_s[12] ), .ZN(n570) );
  INV_X1 U239 ( .A(A_ns[12]), .ZN(n569) );
  OAI221_X1 U240 ( .B1(n393), .B2(n572), .C1(n392), .C2(n573), .A(n574), .ZN(
        O[13]) );
  AOI22_X1 U241 ( .A1(A_ns[12]), .A2(n397), .B1(\A_s[12] ), .B2(n398), .ZN(
        n574) );
  INV_X1 U242 ( .A(\A_s[11] ), .ZN(n573) );
  INV_X1 U243 ( .A(A_ns[11]), .ZN(n572) );
  OAI221_X1 U244 ( .B1(n393), .B2(n575), .C1(n392), .C2(n576), .A(n577), .ZN(
        O[12]) );
  AOI22_X1 U245 ( .A1(A_ns[11]), .A2(n397), .B1(\A_s[11] ), .B2(n398), .ZN(
        n577) );
  INV_X1 U246 ( .A(\A_s[10] ), .ZN(n576) );
  INV_X1 U247 ( .A(A_ns[10]), .ZN(n575) );
  OAI221_X1 U248 ( .B1(n393), .B2(n578), .C1(n392), .C2(n579), .A(n580), .ZN(
        O[11]) );
  AOI22_X1 U249 ( .A1(A_ns[10]), .A2(n397), .B1(\A_s[10] ), .B2(n398), .ZN(
        n580) );
  INV_X1 U250 ( .A(\A_s[9] ), .ZN(n579) );
  INV_X1 U251 ( .A(A_ns[9]), .ZN(n578) );
  OAI221_X1 U252 ( .B1(n581), .B2(n393), .C1(n582), .C2(n392), .A(n583), .ZN(
        O[10]) );
  AOI22_X1 U253 ( .A1(A_ns[9]), .A2(n397), .B1(\A_s[9] ), .B2(n398), .ZN(n583)
         );
  NAND2_X1 U254 ( .A1(n584), .A2(n552), .ZN(n553) );
  NAND2_X1 U255 ( .A1(n584), .A2(n585), .ZN(n552) );
  XOR2_X1 U256 ( .A(B[29]), .B(B[30]), .Z(n584) );
  INV_X1 U257 ( .A(\A_s[8] ), .ZN(n582) );
  INV_X1 U258 ( .A(B[31]), .ZN(n585) );
  INV_X1 U259 ( .A(A_ns[8]), .ZN(n581) );
endmodule


module RCA_NBIT64_15_DW01_add_0 ( A, B, CI, SUM, CO );
  input [64:0] A;
  input [64:0] B;
  output [64:0] SUM;
  input CI;
  output CO;

  wire   [64:1] carry;

  FA_X1 U1_63 ( .A(A[63]), .B(B[63]), .CI(carry[63]), .CO(SUM[64]), .S(SUM[63]) );
  FA_X1 U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  FA_X1 U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  FA_X1 U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  FA_X1 U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  FA_X1 U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  FA_X1 U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  FA_X1 U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  FA_X1 U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  FA_X1 U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  FA_X1 U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  FA_X1 U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  FA_X1 U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  FA_X1 U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  FA_X1 U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  FA_X1 U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  FA_X1 U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  FA_X1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FA_X1 U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  FA_X1 U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  FA_X1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FA_X1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FA_X1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FA_X1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FA_X1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FA_X1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FA_X1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FA_X1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FA_X1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FA_X1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FA_X1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FA_X1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FA_X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(CI), .CO(carry[1]), .S(SUM[0]) );
endmodule


module RCA_NBIT64_15 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;


  RCA_NBIT64_15_DW01_add_0 add_1_root_add_81_2 ( .A({1'b0, A}), .B({1'b0, B}), 
        .CI(Ci), .SUM({Co, S}) );
endmodule


module RCA_NBIT64_29_DW01_add_0 ( A, B, CI, SUM, CO );
  input [64:0] A;
  input [64:0] B;
  output [64:0] SUM;
  input CI;
  output CO;

  wire   [64:1] carry;

  FA_X1 U1_63 ( .A(A[63]), .B(B[63]), .CI(carry[63]), .CO(SUM[64]), .S(SUM[63]) );
  FA_X1 U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  FA_X1 U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  FA_X1 U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  FA_X1 U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  FA_X1 U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  FA_X1 U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  FA_X1 U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  FA_X1 U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  FA_X1 U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  FA_X1 U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  FA_X1 U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  FA_X1 U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  FA_X1 U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  FA_X1 U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  FA_X1 U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  FA_X1 U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  FA_X1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FA_X1 U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  FA_X1 U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  FA_X1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FA_X1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FA_X1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FA_X1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FA_X1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FA_X1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FA_X1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FA_X1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FA_X1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FA_X1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FA_X1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FA_X1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FA_X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(CI), .CO(carry[1]), .S(SUM[0]) );
endmodule


module RCA_NBIT64_29 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;


  RCA_NBIT64_29_DW01_add_0 add_1_root_add_81_2 ( .A({1'b0, A}), .B({1'b0, B}), 
        .CI(Ci), .SUM({Co, S}) );
endmodule


module RCA_NBIT64_28_DW01_add_0 ( A, B, CI, SUM, CO );
  input [64:0] A;
  input [64:0] B;
  output [64:0] SUM;
  input CI;
  output CO;

  wire   [64:1] carry;

  FA_X1 U1_63 ( .A(A[63]), .B(B[63]), .CI(carry[63]), .CO(SUM[64]), .S(SUM[63]) );
  FA_X1 U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  FA_X1 U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  FA_X1 U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  FA_X1 U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  FA_X1 U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  FA_X1 U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  FA_X1 U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  FA_X1 U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  FA_X1 U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  FA_X1 U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  FA_X1 U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  FA_X1 U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  FA_X1 U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  FA_X1 U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  FA_X1 U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  FA_X1 U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  FA_X1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FA_X1 U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  FA_X1 U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  FA_X1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FA_X1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FA_X1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FA_X1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FA_X1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FA_X1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FA_X1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FA_X1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FA_X1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FA_X1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FA_X1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FA_X1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FA_X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(CI), .CO(carry[1]), .S(SUM[0]) );
endmodule


module RCA_NBIT64_28 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;


  RCA_NBIT64_28_DW01_add_0 add_1_root_add_81_2 ( .A({1'b0, A}), .B({1'b0, B}), 
        .CI(Ci), .SUM({Co, S}) );
endmodule


module RCA_NBIT64_27_DW01_add_0 ( A, B, CI, SUM, CO );
  input [64:0] A;
  input [64:0] B;
  output [64:0] SUM;
  input CI;
  output CO;

  wire   [64:1] carry;

  FA_X1 U1_63 ( .A(A[63]), .B(B[63]), .CI(carry[63]), .CO(SUM[64]), .S(SUM[63]) );
  FA_X1 U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  FA_X1 U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  FA_X1 U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  FA_X1 U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  FA_X1 U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  FA_X1 U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  FA_X1 U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  FA_X1 U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  FA_X1 U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  FA_X1 U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  FA_X1 U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  FA_X1 U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  FA_X1 U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  FA_X1 U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  FA_X1 U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  FA_X1 U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  FA_X1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FA_X1 U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  FA_X1 U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  FA_X1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FA_X1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FA_X1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FA_X1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FA_X1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FA_X1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FA_X1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FA_X1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FA_X1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FA_X1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FA_X1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FA_X1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FA_X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(CI), .CO(carry[1]), .S(SUM[0]) );
endmodule


module RCA_NBIT64_27 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;


  RCA_NBIT64_27_DW01_add_0 add_1_root_add_81_2 ( .A({1'b0, A}), .B({1'b0, B}), 
        .CI(Ci), .SUM({Co, S}) );
endmodule


module RCA_NBIT64_26_DW01_add_0 ( A, B, CI, SUM, CO );
  input [64:0] A;
  input [64:0] B;
  output [64:0] SUM;
  input CI;
  output CO;

  wire   [64:1] carry;

  FA_X1 U1_63 ( .A(A[63]), .B(B[63]), .CI(carry[63]), .CO(SUM[64]), .S(SUM[63]) );
  FA_X1 U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  FA_X1 U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  FA_X1 U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  FA_X1 U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  FA_X1 U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  FA_X1 U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  FA_X1 U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  FA_X1 U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  FA_X1 U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  FA_X1 U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  FA_X1 U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  FA_X1 U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  FA_X1 U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  FA_X1 U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  FA_X1 U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  FA_X1 U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  FA_X1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FA_X1 U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  FA_X1 U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  FA_X1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FA_X1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FA_X1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FA_X1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FA_X1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FA_X1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FA_X1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FA_X1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FA_X1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FA_X1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FA_X1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FA_X1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FA_X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(CI), .CO(carry[1]), .S(SUM[0]) );
endmodule


module RCA_NBIT64_26 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;


  RCA_NBIT64_26_DW01_add_0 add_1_root_add_81_2 ( .A({1'b0, A}), .B({1'b0, B}), 
        .CI(Ci), .SUM({Co, S}) );
endmodule


module RCA_NBIT64_25_DW01_add_0 ( A, B, CI, SUM, CO );
  input [64:0] A;
  input [64:0] B;
  output [64:0] SUM;
  input CI;
  output CO;

  wire   [64:1] carry;

  FA_X1 U1_63 ( .A(A[63]), .B(B[63]), .CI(carry[63]), .CO(SUM[64]), .S(SUM[63]) );
  FA_X1 U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  FA_X1 U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  FA_X1 U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  FA_X1 U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  FA_X1 U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  FA_X1 U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  FA_X1 U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  FA_X1 U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  FA_X1 U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  FA_X1 U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  FA_X1 U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  FA_X1 U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  FA_X1 U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  FA_X1 U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  FA_X1 U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  FA_X1 U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  FA_X1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FA_X1 U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  FA_X1 U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  FA_X1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FA_X1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FA_X1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FA_X1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FA_X1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FA_X1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FA_X1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FA_X1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FA_X1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FA_X1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FA_X1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FA_X1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FA_X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(CI), .CO(carry[1]), .S(SUM[0]) );
endmodule


module RCA_NBIT64_25 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;


  RCA_NBIT64_25_DW01_add_0 add_1_root_add_81_2 ( .A({1'b0, A}), .B({1'b0, B}), 
        .CI(Ci), .SUM({Co, S}) );
endmodule


module RCA_NBIT64_24_DW01_add_0 ( A, B, CI, SUM, CO );
  input [64:0] A;
  input [64:0] B;
  output [64:0] SUM;
  input CI;
  output CO;

  wire   [64:1] carry;

  FA_X1 U1_63 ( .A(A[63]), .B(B[63]), .CI(carry[63]), .CO(SUM[64]), .S(SUM[63]) );
  FA_X1 U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  FA_X1 U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  FA_X1 U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  FA_X1 U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  FA_X1 U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  FA_X1 U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  FA_X1 U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  FA_X1 U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  FA_X1 U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  FA_X1 U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  FA_X1 U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  FA_X1 U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  FA_X1 U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  FA_X1 U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  FA_X1 U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  FA_X1 U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  FA_X1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FA_X1 U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  FA_X1 U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  FA_X1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FA_X1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FA_X1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FA_X1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FA_X1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FA_X1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FA_X1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FA_X1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FA_X1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FA_X1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FA_X1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FA_X1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FA_X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(CI), .CO(carry[1]), .S(SUM[0]) );
endmodule


module RCA_NBIT64_24 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;


  RCA_NBIT64_24_DW01_add_0 add_1_root_add_81_2 ( .A({1'b0, A}), .B({1'b0, B}), 
        .CI(Ci), .SUM({Co, S}) );
endmodule


module RCA_NBIT64_23_DW01_add_0 ( A, B, CI, SUM, CO );
  input [64:0] A;
  input [64:0] B;
  output [64:0] SUM;
  input CI;
  output CO;

  wire   [64:1] carry;

  FA_X1 U1_63 ( .A(A[63]), .B(B[63]), .CI(carry[63]), .CO(SUM[64]), .S(SUM[63]) );
  FA_X1 U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  FA_X1 U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  FA_X1 U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  FA_X1 U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  FA_X1 U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  FA_X1 U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  FA_X1 U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  FA_X1 U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  FA_X1 U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  FA_X1 U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  FA_X1 U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  FA_X1 U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  FA_X1 U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  FA_X1 U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  FA_X1 U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  FA_X1 U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  FA_X1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FA_X1 U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  FA_X1 U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  FA_X1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FA_X1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FA_X1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FA_X1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FA_X1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FA_X1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FA_X1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FA_X1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FA_X1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FA_X1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FA_X1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FA_X1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FA_X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(CI), .CO(carry[1]), .S(SUM[0]) );
endmodule


module RCA_NBIT64_23 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;


  RCA_NBIT64_23_DW01_add_0 add_1_root_add_81_2 ( .A({1'b0, A}), .B({1'b0, B}), 
        .CI(Ci), .SUM({Co, S}) );
endmodule


module RCA_NBIT64_22_DW01_add_0 ( A, B, CI, SUM, CO );
  input [64:0] A;
  input [64:0] B;
  output [64:0] SUM;
  input CI;
  output CO;

  wire   [64:1] carry;

  FA_X1 U1_63 ( .A(A[63]), .B(B[63]), .CI(carry[63]), .CO(SUM[64]), .S(SUM[63]) );
  FA_X1 U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  FA_X1 U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  FA_X1 U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  FA_X1 U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  FA_X1 U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  FA_X1 U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  FA_X1 U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  FA_X1 U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  FA_X1 U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  FA_X1 U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  FA_X1 U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  FA_X1 U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  FA_X1 U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  FA_X1 U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  FA_X1 U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  FA_X1 U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  FA_X1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FA_X1 U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  FA_X1 U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  FA_X1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FA_X1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FA_X1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FA_X1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FA_X1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FA_X1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FA_X1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FA_X1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FA_X1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FA_X1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FA_X1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FA_X1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FA_X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(CI), .CO(carry[1]), .S(SUM[0]) );
endmodule


module RCA_NBIT64_22 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;


  RCA_NBIT64_22_DW01_add_0 add_1_root_add_81_2 ( .A({1'b0, A}), .B({1'b0, B}), 
        .CI(Ci), .SUM({Co, S}) );
endmodule


module RCA_NBIT64_21_DW01_add_0 ( A, B, CI, SUM, CO );
  input [64:0] A;
  input [64:0] B;
  output [64:0] SUM;
  input CI;
  output CO;

  wire   [64:1] carry;

  FA_X1 U1_63 ( .A(A[63]), .B(B[63]), .CI(carry[63]), .CO(SUM[64]), .S(SUM[63]) );
  FA_X1 U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  FA_X1 U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  FA_X1 U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  FA_X1 U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  FA_X1 U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  FA_X1 U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  FA_X1 U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  FA_X1 U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  FA_X1 U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  FA_X1 U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  FA_X1 U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  FA_X1 U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  FA_X1 U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  FA_X1 U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  FA_X1 U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  FA_X1 U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  FA_X1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FA_X1 U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  FA_X1 U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  FA_X1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FA_X1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FA_X1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FA_X1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FA_X1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FA_X1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FA_X1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FA_X1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FA_X1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FA_X1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FA_X1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FA_X1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FA_X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(CI), .CO(carry[1]), .S(SUM[0]) );
endmodule


module RCA_NBIT64_21 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;


  RCA_NBIT64_21_DW01_add_0 add_1_root_add_81_2 ( .A({1'b0, A}), .B({1'b0, B}), 
        .CI(Ci), .SUM({Co, S}) );
endmodule


module RCA_NBIT64_20_DW01_add_0 ( A, B, CI, SUM, CO );
  input [64:0] A;
  input [64:0] B;
  output [64:0] SUM;
  input CI;
  output CO;

  wire   [64:1] carry;

  FA_X1 U1_63 ( .A(A[63]), .B(B[63]), .CI(carry[63]), .CO(SUM[64]), .S(SUM[63]) );
  FA_X1 U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  FA_X1 U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  FA_X1 U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  FA_X1 U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  FA_X1 U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  FA_X1 U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  FA_X1 U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  FA_X1 U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  FA_X1 U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  FA_X1 U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  FA_X1 U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  FA_X1 U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  FA_X1 U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  FA_X1 U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  FA_X1 U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  FA_X1 U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  FA_X1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FA_X1 U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  FA_X1 U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  FA_X1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FA_X1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FA_X1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FA_X1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FA_X1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FA_X1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FA_X1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FA_X1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FA_X1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FA_X1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FA_X1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FA_X1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FA_X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(CI), .CO(carry[1]), .S(SUM[0]) );
endmodule


module RCA_NBIT64_20 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;


  RCA_NBIT64_20_DW01_add_0 add_1_root_add_81_2 ( .A({1'b0, A}), .B({1'b0, B}), 
        .CI(Ci), .SUM({Co, S}) );
endmodule


module RCA_NBIT64_19_DW01_add_0 ( A, B, CI, SUM, CO );
  input [64:0] A;
  input [64:0] B;
  output [64:0] SUM;
  input CI;
  output CO;

  wire   [64:1] carry;

  FA_X1 U1_63 ( .A(A[63]), .B(B[63]), .CI(carry[63]), .CO(SUM[64]), .S(SUM[63]) );
  FA_X1 U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  FA_X1 U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  FA_X1 U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  FA_X1 U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  FA_X1 U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  FA_X1 U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  FA_X1 U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  FA_X1 U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  FA_X1 U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  FA_X1 U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  FA_X1 U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  FA_X1 U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  FA_X1 U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  FA_X1 U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  FA_X1 U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  FA_X1 U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  FA_X1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FA_X1 U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  FA_X1 U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  FA_X1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FA_X1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FA_X1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FA_X1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FA_X1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FA_X1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FA_X1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FA_X1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FA_X1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FA_X1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FA_X1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FA_X1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FA_X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(CI), .CO(carry[1]), .S(SUM[0]) );
endmodule


module RCA_NBIT64_19 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;


  RCA_NBIT64_19_DW01_add_0 add_1_root_add_81_2 ( .A({1'b0, A}), .B({1'b0, B}), 
        .CI(Ci), .SUM({Co, S}) );
endmodule


module RCA_NBIT64_18_DW01_add_0 ( A, B, CI, SUM, CO );
  input [64:0] A;
  input [64:0] B;
  output [64:0] SUM;
  input CI;
  output CO;

  wire   [64:1] carry;

  FA_X1 U1_63 ( .A(A[63]), .B(B[63]), .CI(carry[63]), .CO(SUM[64]), .S(SUM[63]) );
  FA_X1 U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  FA_X1 U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  FA_X1 U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  FA_X1 U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  FA_X1 U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  FA_X1 U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  FA_X1 U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  FA_X1 U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  FA_X1 U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  FA_X1 U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  FA_X1 U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  FA_X1 U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  FA_X1 U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  FA_X1 U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  FA_X1 U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  FA_X1 U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  FA_X1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FA_X1 U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  FA_X1 U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  FA_X1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FA_X1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FA_X1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FA_X1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FA_X1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FA_X1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FA_X1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FA_X1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FA_X1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FA_X1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FA_X1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FA_X1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FA_X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(CI), .CO(carry[1]), .S(SUM[0]) );
endmodule


module RCA_NBIT64_18 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;


  RCA_NBIT64_18_DW01_add_0 add_1_root_add_81_2 ( .A({1'b0, A}), .B({1'b0, B}), 
        .CI(Ci), .SUM({Co, S}) );
endmodule


module RCA_NBIT64_17_DW01_add_0 ( A, B, CI, SUM, CO );
  input [64:0] A;
  input [64:0] B;
  output [64:0] SUM;
  input CI;
  output CO;

  wire   [64:1] carry;

  FA_X1 U1_63 ( .A(A[63]), .B(B[63]), .CI(carry[63]), .CO(SUM[64]), .S(SUM[63]) );
  FA_X1 U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  FA_X1 U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  FA_X1 U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  FA_X1 U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  FA_X1 U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  FA_X1 U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  FA_X1 U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  FA_X1 U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  FA_X1 U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  FA_X1 U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  FA_X1 U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  FA_X1 U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  FA_X1 U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  FA_X1 U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  FA_X1 U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  FA_X1 U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  FA_X1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FA_X1 U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  FA_X1 U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  FA_X1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FA_X1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FA_X1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FA_X1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FA_X1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FA_X1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FA_X1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FA_X1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FA_X1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FA_X1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FA_X1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FA_X1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FA_X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(CI), .CO(carry[1]), .S(SUM[0]) );
endmodule


module RCA_NBIT64_17 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;


  RCA_NBIT64_17_DW01_add_0 add_1_root_add_81_2 ( .A({1'b0, A}), .B({1'b0, B}), 
        .CI(Ci), .SUM({Co, S}) );
endmodule


module RCA_NBIT64_16_DW01_add_0 ( A, B, CI, SUM, CO );
  input [64:0] A;
  input [64:0] B;
  output [64:0] SUM;
  input CI;
  output CO;

  wire   [64:1] carry;

  FA_X1 U1_63 ( .A(A[63]), .B(B[63]), .CI(carry[63]), .CO(SUM[64]), .S(SUM[63]) );
  FA_X1 U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  FA_X1 U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  FA_X1 U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  FA_X1 U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  FA_X1 U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  FA_X1 U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  FA_X1 U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  FA_X1 U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  FA_X1 U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  FA_X1 U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  FA_X1 U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  FA_X1 U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  FA_X1 U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  FA_X1 U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  FA_X1 U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  FA_X1 U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  FA_X1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FA_X1 U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  FA_X1 U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  FA_X1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FA_X1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  FA_X1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FA_X1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  FA_X1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  FA_X1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FA_X1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  FA_X1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  FA_X1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  FA_X1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FA_X1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FA_X1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  FA_X1 U1_0 ( .A(A[0]), .B(B[0]), .CI(CI), .CO(carry[1]), .S(SUM[0]) );
endmodule


module RCA_NBIT64_16 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;


  RCA_NBIT64_16_DW01_add_0 add_1_root_add_81_2 ( .A({1'b0, A}), .B({1'b0, B}), 
        .CI(Ci), .SUM({Co, S}) );
endmodule


module BOOTHMUL_NBIT32_1_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n96, n97, n98, n99, n101, n102, n103, n104, n105, n106, n107,
         n108, n110, n111, n112, n114, n115, n116, n118, n119, n120, n122,
         n123, n94, n100, n109, n113, n117, n121, n124, n125, n126;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U42 ( .A(n97), .B(B[9]), .Z(DIFF[9]) );
  XOR2_X1 U43 ( .A(n99), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U45 ( .A(n101), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U46 ( .A(n103), .B(B[3]), .Z(DIFF[3]) );
  XOR2_X1 U47 ( .A(n96), .B(B[30]), .Z(DIFF[30]) );
  XOR2_X1 U48 ( .A(n106), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U50 ( .A(n108), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U51 ( .A(n110), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U53 ( .A(n112), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U54 ( .A(B[1]), .B(\B[0] ), .Z(DIFF[1]) );
  XOR2_X1 U55 ( .A(n114), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U57 ( .A(n116), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U58 ( .A(n118), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U60 ( .A(n120), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U61 ( .A(n122), .B(B[11]), .Z(DIFF[11]) );
  XOR2_X1 U1 ( .A(n100), .B(B[31]), .Z(n94) );
  INV_X2 U2 ( .A(n94), .ZN(DIFF[31]) );
  NOR2_X1 U3 ( .A1(n96), .A2(B[30]), .ZN(n100) );
  NOR3_X1 U4 ( .A1(B[27]), .A2(B[28]), .A3(n106), .ZN(n104) );
  NAND2_X1 U5 ( .A1(n104), .A2(n126), .ZN(n96) );
  INV_X1 U6 ( .A(B[29]), .ZN(n126) );
  OR3_X1 U7 ( .A1(B[25]), .A2(B[26]), .A3(n108), .ZN(n106) );
  OR3_X1 U8 ( .A1(B[1]), .A2(B[2]), .A3(\B[0] ), .ZN(n103) );
  OR3_X1 U9 ( .A1(B[5]), .A2(B[6]), .A3(n101), .ZN(n99) );
  OR3_X1 U10 ( .A1(B[10]), .A2(B[9]), .A3(n97), .ZN(n122) );
  OR3_X1 U11 ( .A1(B[13]), .A2(B[14]), .A3(n120), .ZN(n118) );
  OR3_X1 U12 ( .A1(B[17]), .A2(B[18]), .A3(n116), .ZN(n114) );
  OR3_X1 U13 ( .A1(B[21]), .A2(B[22]), .A3(n112), .ZN(n110) );
  OR3_X1 U14 ( .A1(B[3]), .A2(B[4]), .A3(n103), .ZN(n101) );
  OR3_X1 U15 ( .A1(B[7]), .A2(B[8]), .A3(n99), .ZN(n97) );
  OR3_X1 U16 ( .A1(B[11]), .A2(B[12]), .A3(n122), .ZN(n120) );
  OR3_X1 U17 ( .A1(B[15]), .A2(B[16]), .A3(n118), .ZN(n116) );
  OR3_X1 U18 ( .A1(B[19]), .A2(B[20]), .A3(n114), .ZN(n112) );
  OR3_X1 U19 ( .A1(B[23]), .A2(B[24]), .A3(n110), .ZN(n108) );
  XNOR2_X1 U20 ( .A(n104), .B(B[29]), .ZN(DIFF[29]) );
  XNOR2_X1 U21 ( .A(n109), .B(B[6]), .ZN(DIFF[6]) );
  NOR2_X1 U22 ( .A1(n101), .A2(B[5]), .ZN(n109) );
  XNOR2_X1 U23 ( .A(n113), .B(B[10]), .ZN(DIFF[10]) );
  NOR2_X1 U24 ( .A1(n97), .A2(B[9]), .ZN(n113) );
  XNOR2_X1 U25 ( .A(n117), .B(B[14]), .ZN(DIFF[14]) );
  NOR2_X1 U26 ( .A1(n120), .A2(B[13]), .ZN(n117) );
  XNOR2_X1 U27 ( .A(n121), .B(B[18]), .ZN(DIFF[18]) );
  NOR2_X1 U28 ( .A1(n116), .A2(B[17]), .ZN(n121) );
  XNOR2_X1 U29 ( .A(n124), .B(B[22]), .ZN(DIFF[22]) );
  NOR2_X1 U30 ( .A1(n112), .A2(B[21]), .ZN(n124) );
  XNOR2_X1 U31 ( .A(n125), .B(B[26]), .ZN(DIFF[26]) );
  NOR2_X1 U32 ( .A1(n108), .A2(B[25]), .ZN(n125) );
  XNOR2_X1 U33 ( .A(B[2]), .B(n105), .ZN(DIFF[2]) );
  NOR2_X1 U34 ( .A1(\B[0] ), .A2(B[1]), .ZN(n105) );
  XNOR2_X1 U35 ( .A(B[4]), .B(n102), .ZN(DIFF[4]) );
  NOR2_X1 U36 ( .A1(B[3]), .A2(n103), .ZN(n102) );
  XNOR2_X1 U37 ( .A(B[12]), .B(n123), .ZN(DIFF[12]) );
  NOR2_X1 U38 ( .A1(B[11]), .A2(n122), .ZN(n123) );
  XNOR2_X1 U39 ( .A(B[16]), .B(n119), .ZN(DIFF[16]) );
  NOR2_X1 U40 ( .A1(B[15]), .A2(n118), .ZN(n119) );
  XNOR2_X1 U41 ( .A(B[20]), .B(n115), .ZN(DIFF[20]) );
  NOR2_X1 U44 ( .A1(B[19]), .A2(n114), .ZN(n115) );
  XNOR2_X1 U49 ( .A(B[24]), .B(n111), .ZN(DIFF[24]) );
  NOR2_X1 U52 ( .A1(B[23]), .A2(n110), .ZN(n111) );
  XNOR2_X1 U56 ( .A(B[28]), .B(n107), .ZN(DIFF[28]) );
  NOR2_X1 U59 ( .A1(B[27]), .A2(n106), .ZN(n107) );
  XNOR2_X1 U62 ( .A(B[8]), .B(n98), .ZN(DIFF[8]) );
  NOR2_X1 U63 ( .A1(B[7]), .A2(n99), .ZN(n98) );
endmodule


module BOOTHMUL_NBIT32_1 ( A, B, S );
  input [31:0] A;
  input [31:0] B;
  output [63:0] S;
  wire   A_n_63;
  wire   [30:0] A_n;
  wire   [1023:64] SHIFT;
  wire   [1023:64] SHIFT_n;
  wire   [1023:0] OTMP;
  wire   [895:0] PTMP;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72;

  BOOTHENC_NBIT64_i0 BOOTHENC_I_1 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .A_n({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .A_ns({A_n_63, A_n_63, A_n_63, A_n_63, 
        A_n_63, A_n_63, A_n_63, A_n_63, A_n_63, A_n_63, A_n_63, A_n_63, A_n_63, 
        A_n_63, A_n_63, A_n_63, A_n_63, A_n_63, A_n_63, A_n_63, A_n_63, A_n_63, 
        A_n_63, A_n_63, A_n_63, A_n_63, A_n_63, A_n_63, A_n_63, A_n_63, A_n_63, 
        A_n_63, A_n_63, A_n}), .A_s({A[31], A[31], A[31], A[31], A[31], A[31], 
        A[31], A[31], A[31], A[31], A[31], A[31], A[31], A[31], A[31], A[31], 
        A[31], A[31], A[31], A[31], A[31], A[31], A[31], A[31], A[31], A[31], 
        A[31], A[31], A[31], A[31], A[31], A[31], A}), .B({B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B}), 
        .O(OTMP[63:0]), .A_so({SHIFT[127:65], SYNOPSYS_UNCONNECTED__0}), 
        .A_nso({SHIFT_n[127:65], SYNOPSYS_UNCONNECTED__1}) );
  BOOTHENC_NBIT64_i2 BOOTHENC_I_2 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .A_n({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .A_ns({SHIFT_n[127:65], 1'b0}), .A_s({
        SHIFT[127:65], 1'b0}), .B({B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B}), .O({OTMP[127:65], 
        SYNOPSYS_UNCONNECTED__2}), .A_so({SHIFT[191:130], 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4}), .A_nso({
        SHIFT_n[191:130], SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6})
         );
  BOOTHENC_NBIT64_i4 BOOTHENC_I_3 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .A_n({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .A_ns({SHIFT_n[191:130], 1'b0, 1'b0}), .A_s(
        {SHIFT[191:130], 1'b0, 1'b0}), .B({B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B}), .O({
        OTMP[191:129], SYNOPSYS_UNCONNECTED__7}), .A_so({SHIFT[255:194], 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9}), .A_nso({
        SHIFT_n[255:194], SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11})
         );
  BOOTHENC_NBIT64_i6 BOOTHENC_I_4 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .A_n({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .A_ns({SHIFT_n[255:194], 1'b0, 1'b0}), .A_s(
        {SHIFT[255:194], 1'b0, 1'b0}), .B({B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B}), .O({
        OTMP[255:193], SYNOPSYS_UNCONNECTED__12}), .A_so({SHIFT[319:258], 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14}), .A_nso({
        SHIFT_n[319:258], SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16})
         );
  BOOTHENC_NBIT64_i8 BOOTHENC_I_5 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .A_n({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .A_ns({SHIFT_n[319:258], 1'b0, 1'b0}), .A_s(
        {SHIFT[319:258], 1'b0, 1'b0}), .B({B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B}), .O({
        OTMP[319:257], SYNOPSYS_UNCONNECTED__17}), .A_so({SHIFT[383:322], 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19}), .A_nso({
        SHIFT_n[383:322], SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21})
         );
  BOOTHENC_NBIT64_i10 BOOTHENC_I_6 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .A_n({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .A_ns({SHIFT_n[383:322], 1'b0, 1'b0}), .A_s(
        {SHIFT[383:322], 1'b0, 1'b0}), .B({B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B}), .O({
        OTMP[383:321], SYNOPSYS_UNCONNECTED__22}), .A_so({SHIFT[447:386], 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24}), .A_nso({
        SHIFT_n[447:386], SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26})
         );
  BOOTHENC_NBIT64_i12 BOOTHENC_I_7 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .A_n({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .A_ns({SHIFT_n[447:386], 1'b0, 1'b0}), .A_s(
        {SHIFT[447:386], 1'b0, 1'b0}), .B({B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B}), .O({
        OTMP[447:385], SYNOPSYS_UNCONNECTED__27}), .A_so({SHIFT[511:450], 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29}), .A_nso({
        SHIFT_n[511:450], SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31})
         );
  BOOTHENC_NBIT64_i14 BOOTHENC_I_8 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .A_n({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .A_ns({SHIFT_n[511:450], 1'b0, 1'b0}), .A_s(
        {SHIFT[511:450], 1'b0, 1'b0}), .B({B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B}), .O({
        OTMP[511:449], SYNOPSYS_UNCONNECTED__32}), .A_so({SHIFT[575:514], 
        SYNOPSYS_UNCONNECTED__33, SYNOPSYS_UNCONNECTED__34}), .A_nso({
        SHIFT_n[575:514], SYNOPSYS_UNCONNECTED__35, SYNOPSYS_UNCONNECTED__36})
         );
  BOOTHENC_NBIT64_i16 BOOTHENC_I_9 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .A_n({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .A_ns({SHIFT_n[575:514], 1'b0, 1'b0}), .A_s(
        {SHIFT[575:514], 1'b0, 1'b0}), .B({B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B}), .O({
        OTMP[575:513], SYNOPSYS_UNCONNECTED__37}), .A_so({SHIFT[639:578], 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39}), .A_nso({
        SHIFT_n[639:578], SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41})
         );
  BOOTHENC_NBIT64_i18 BOOTHENC_I_10 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .A_n({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .A_ns({SHIFT_n[639:578], 1'b0, 1'b0}), .A_s(
        {SHIFT[639:578], 1'b0, 1'b0}), .B({B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B}), .O({
        OTMP[639:577], SYNOPSYS_UNCONNECTED__42}), .A_so({SHIFT[703:642], 
        SYNOPSYS_UNCONNECTED__43, SYNOPSYS_UNCONNECTED__44}), .A_nso({
        SHIFT_n[703:642], SYNOPSYS_UNCONNECTED__45, SYNOPSYS_UNCONNECTED__46})
         );
  BOOTHENC_NBIT64_i20 BOOTHENC_I_11 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .A_n({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .A_ns({SHIFT_n[703:642], 1'b0, 1'b0}), .A_s(
        {SHIFT[703:642], 1'b0, 1'b0}), .B({B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B}), .O({
        OTMP[703:641], SYNOPSYS_UNCONNECTED__47}), .A_so({SHIFT[767:706], 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49}), .A_nso({
        SHIFT_n[767:706], SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51})
         );
  BOOTHENC_NBIT64_i22 BOOTHENC_I_12 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .A_n({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .A_ns({SHIFT_n[767:706], 1'b0, 1'b0}), .A_s(
        {SHIFT[767:706], 1'b0, 1'b0}), .B({B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B}), .O({
        OTMP[767:705], SYNOPSYS_UNCONNECTED__52}), .A_so({SHIFT[831:770], 
        SYNOPSYS_UNCONNECTED__53, SYNOPSYS_UNCONNECTED__54}), .A_nso({
        SHIFT_n[831:770], SYNOPSYS_UNCONNECTED__55, SYNOPSYS_UNCONNECTED__56})
         );
  BOOTHENC_NBIT64_i24 BOOTHENC_I_13 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .A_n({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .A_ns({SHIFT_n[831:770], 1'b0, 1'b0}), .A_s(
        {SHIFT[831:770], 1'b0, 1'b0}), .B({B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B}), .O({
        OTMP[831:769], SYNOPSYS_UNCONNECTED__57}), .A_so({SHIFT[895:834], 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59}), .A_nso({
        SHIFT_n[895:834], SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61})
         );
  BOOTHENC_NBIT64_i26 BOOTHENC_I_14 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .A_n({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .A_ns({SHIFT_n[895:834], 1'b0, 1'b0}), .A_s(
        {SHIFT[895:834], 1'b0, 1'b0}), .B({B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B}), .O({
        OTMP[895:833], SYNOPSYS_UNCONNECTED__62}), .A_so({SHIFT[959:898], 
        SYNOPSYS_UNCONNECTED__63, SYNOPSYS_UNCONNECTED__64}), .A_nso({
        SHIFT_n[959:898], SYNOPSYS_UNCONNECTED__65, SYNOPSYS_UNCONNECTED__66})
         );
  BOOTHENC_NBIT64_i28 BOOTHENC_I_15 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .A_n({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .A_ns({SHIFT_n[959:898], 1'b0, 1'b0}), .A_s(
        {SHIFT[959:898], 1'b0, 1'b0}), .B({B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B}), .O({
        OTMP[959:897], SYNOPSYS_UNCONNECTED__67}), .A_so({SHIFT[1023:962], 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69}), .A_nso({
        SHIFT_n[1023:962], SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71}) );
  BOOTHENC_NBIT64_i30 BOOTHENC_I_16 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .A_n({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .A_ns({SHIFT_n[1023:962], 1'b0, 1'b0}), 
        .A_s({SHIFT[1023:962], 1'b0, 1'b0}), .B({B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], 
        B[31], B[31], B[31], B[31], B[31], B[31], B[31], B[31], B}), .O({
        OTMP[1023:961], SYNOPSYS_UNCONNECTED__72}) );
  RCA_NBIT64_15 ADDER2_2 ( .A(OTMP[63:0]), .B({OTMP[127:65], 1'b0}), .Ci(1'b0), 
        .S(PTMP[63:0]) );
  RCA_NBIT64_29 ADDERI_3 ( .A(PTMP[63:0]), .B({OTMP[191:129], 1'b0}), .Ci(1'b0), .S(PTMP[127:64]) );
  RCA_NBIT64_28 ADDERI_4 ( .A(PTMP[127:64]), .B({OTMP[255:193], 1'b0}), .Ci(
        1'b0), .S(PTMP[191:128]) );
  RCA_NBIT64_27 ADDERI_5 ( .A(PTMP[191:128]), .B({OTMP[319:257], 1'b0}), .Ci(
        1'b0), .S(PTMP[255:192]) );
  RCA_NBIT64_26 ADDERI_6 ( .A(PTMP[255:192]), .B({OTMP[383:321], 1'b0}), .Ci(
        1'b0), .S(PTMP[319:256]) );
  RCA_NBIT64_25 ADDERI_7 ( .A(PTMP[319:256]), .B({OTMP[447:385], 1'b0}), .Ci(
        1'b0), .S(PTMP[383:320]) );
  RCA_NBIT64_24 ADDERI_8 ( .A(PTMP[383:320]), .B({OTMP[511:449], 1'b0}), .Ci(
        1'b0), .S(PTMP[447:384]) );
  RCA_NBIT64_23 ADDERI_9 ( .A(PTMP[447:384]), .B({OTMP[575:513], 1'b0}), .Ci(
        1'b0), .S(PTMP[511:448]) );
  RCA_NBIT64_22 ADDERI_10 ( .A(PTMP[511:448]), .B({OTMP[639:577], 1'b0}), .Ci(
        1'b0), .S(PTMP[575:512]) );
  RCA_NBIT64_21 ADDERI_11 ( .A(PTMP[575:512]), .B({OTMP[703:641], 1'b0}), .Ci(
        1'b0), .S(PTMP[639:576]) );
  RCA_NBIT64_20 ADDERI_12 ( .A(PTMP[639:576]), .B({OTMP[767:705], 1'b0}), .Ci(
        1'b0), .S(PTMP[703:640]) );
  RCA_NBIT64_19 ADDERI_13 ( .A(PTMP[703:640]), .B({OTMP[831:769], 1'b0}), .Ci(
        1'b0), .S(PTMP[767:704]) );
  RCA_NBIT64_18 ADDERI_14 ( .A(PTMP[767:704]), .B({OTMP[895:833], 1'b0}), .Ci(
        1'b0), .S(PTMP[831:768]) );
  RCA_NBIT64_17 ADDERI_15 ( .A(PTMP[831:768]), .B({OTMP[959:897], 1'b0}), .Ci(
        1'b0), .S(PTMP[895:832]) );
  RCA_NBIT64_16 ADDERI_16 ( .A(PTMP[895:832]), .B({OTMP[1023:961], 1'b0}), 
        .Ci(1'b0), .S(S) );
  BOOTHMUL_NBIT32_1_DW01_sub_0 sub_82 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF({A_n_63, A_n}) );
endmodule

