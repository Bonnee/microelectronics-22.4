
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_BOOTHMUL_NBIT32 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_BOOTHMUL_NBIT32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHMUL_NBIT32_DW01_sub_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end BOOTHMUL_NBIT32_DW01_sub_0;

architecture SYN_rpl of BOOTHMUL_NBIT32_DW01_sub_0 is

   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, DIFF_27_port,
      DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, DIFF_22_port, 
      DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, DIFF_17_port, 
      DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, DIFF_12_port, 
      DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, DIFF_7_port, 
      DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, DIFF_2_port, 
      DIFF_1_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
      n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29
      , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
      n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58
      , n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, 
      n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93 : std_logic;

begin
   DIFF <= ( DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, 
      DIFF_2_port, DIFF_1_port, B(0) );
   
   U1 : AND2_X1 port map( A1 => n63, A2 => n30, ZN => n1);
   U2 : INV_X4 port map( A => n31, ZN => DIFF_31_port);
   U3 : XNOR2_X1 port map( A => n92, B => n93, ZN => n61);
   U4 : XNOR2_X1 port map( A => n91, B => n2, ZN => n60);
   U5 : XNOR2_X1 port map( A => n90, B => n3, ZN => n59);
   U6 : XNOR2_X1 port map( A => n89, B => n4, ZN => n58);
   U7 : XNOR2_X1 port map( A => n88, B => n5, ZN => n57);
   U8 : XNOR2_X1 port map( A => n87, B => n6, ZN => n56);
   U9 : XNOR2_X1 port map( A => n86, B => n7, ZN => n55);
   U10 : XNOR2_X1 port map( A => n85, B => n8, ZN => n54);
   U11 : XNOR2_X1 port map( A => n84, B => n9, ZN => n53);
   U12 : XNOR2_X1 port map( A => n83, B => n10, ZN => n52);
   U13 : XNOR2_X1 port map( A => n82, B => n11, ZN => n51);
   U14 : XNOR2_X1 port map( A => n81, B => n12, ZN => n50);
   U15 : XNOR2_X1 port map( A => n80, B => n13, ZN => n49);
   U16 : XNOR2_X1 port map( A => n79, B => n14, ZN => n48);
   U17 : XNOR2_X1 port map( A => n78, B => n15, ZN => n47);
   U18 : XNOR2_X1 port map( A => n77, B => n16, ZN => n46);
   U19 : XNOR2_X1 port map( A => n76, B => n17, ZN => n45);
   U20 : XNOR2_X1 port map( A => n75, B => n18, ZN => n44);
   U21 : XNOR2_X1 port map( A => n74, B => n19, ZN => n43);
   U22 : XNOR2_X1 port map( A => n73, B => n20, ZN => n42);
   U23 : XNOR2_X1 port map( A => n72, B => n21, ZN => n41);
   U24 : XNOR2_X1 port map( A => n71, B => n22, ZN => n40);
   U25 : XNOR2_X1 port map( A => n70, B => n23, ZN => n39);
   U26 : XNOR2_X1 port map( A => n69, B => n24, ZN => n38);
   U27 : XNOR2_X1 port map( A => n68, B => n25, ZN => n37);
   U28 : XNOR2_X1 port map( A => n67, B => n26, ZN => n36);
   U29 : XNOR2_X1 port map( A => n66, B => n27, ZN => n35);
   U30 : XNOR2_X1 port map( A => n65, B => n28, ZN => n34);
   U31 : XNOR2_X1 port map( A => n63, B => n30, ZN => n32);
   U32 : XNOR2_X1 port map( A => n64, B => n29, ZN => n33);
   U33 : AND2_X1 port map( A1 => n92, A2 => n93, ZN => n2);
   U34 : AND2_X1 port map( A1 => n91, A2 => n2, ZN => n3);
   U35 : AND2_X1 port map( A1 => n90, A2 => n3, ZN => n4);
   U36 : AND2_X1 port map( A1 => n89, A2 => n4, ZN => n5);
   U37 : AND2_X1 port map( A1 => n88, A2 => n5, ZN => n6);
   U38 : AND2_X1 port map( A1 => n87, A2 => n6, ZN => n7);
   U39 : AND2_X1 port map( A1 => n86, A2 => n7, ZN => n8);
   U40 : AND2_X1 port map( A1 => n85, A2 => n8, ZN => n9);
   U41 : AND2_X1 port map( A1 => n84, A2 => n9, ZN => n10);
   U42 : AND2_X1 port map( A1 => n83, A2 => n10, ZN => n11);
   U43 : AND2_X1 port map( A1 => n82, A2 => n11, ZN => n12);
   U44 : AND2_X1 port map( A1 => n81, A2 => n12, ZN => n13);
   U45 : AND2_X1 port map( A1 => n80, A2 => n13, ZN => n14);
   U46 : AND2_X1 port map( A1 => n79, A2 => n14, ZN => n15);
   U47 : AND2_X1 port map( A1 => n78, A2 => n15, ZN => n16);
   U48 : AND2_X1 port map( A1 => n77, A2 => n16, ZN => n17);
   U49 : AND2_X1 port map( A1 => n76, A2 => n17, ZN => n18);
   U50 : AND2_X1 port map( A1 => n75, A2 => n18, ZN => n19);
   U51 : AND2_X1 port map( A1 => n74, A2 => n19, ZN => n20);
   U52 : AND2_X1 port map( A1 => n73, A2 => n20, ZN => n21);
   U53 : AND2_X1 port map( A1 => n72, A2 => n21, ZN => n22);
   U54 : AND2_X1 port map( A1 => n71, A2 => n22, ZN => n23);
   U55 : AND2_X1 port map( A1 => n70, A2 => n23, ZN => n24);
   U56 : AND2_X1 port map( A1 => n69, A2 => n24, ZN => n25);
   U57 : AND2_X1 port map( A1 => n68, A2 => n25, ZN => n26);
   U58 : AND2_X1 port map( A1 => n67, A2 => n26, ZN => n27);
   U59 : AND2_X1 port map( A1 => n66, A2 => n27, ZN => n28);
   U60 : AND2_X1 port map( A1 => n65, A2 => n28, ZN => n29);
   U61 : AND2_X1 port map( A1 => n64, A2 => n29, ZN => n30);
   U62 : XNOR2_X1 port map( A => n62, B => n1, ZN => n31);
   U63 : INV_X1 port map( A => B(31), ZN => n62);
   U64 : INV_X1 port map( A => B(0), ZN => n93);
   U65 : INV_X1 port map( A => B(1), ZN => n92);
   U66 : INV_X1 port map( A => B(2), ZN => n91);
   U67 : INV_X1 port map( A => B(3), ZN => n90);
   U68 : INV_X1 port map( A => B(4), ZN => n89);
   U69 : INV_X1 port map( A => B(5), ZN => n88);
   U70 : INV_X1 port map( A => B(6), ZN => n87);
   U71 : INV_X1 port map( A => B(7), ZN => n86);
   U72 : INV_X1 port map( A => B(8), ZN => n85);
   U73 : INV_X1 port map( A => B(9), ZN => n84);
   U74 : INV_X1 port map( A => B(10), ZN => n83);
   U75 : INV_X1 port map( A => B(11), ZN => n82);
   U76 : INV_X1 port map( A => B(12), ZN => n81);
   U77 : INV_X1 port map( A => B(13), ZN => n80);
   U78 : INV_X1 port map( A => B(14), ZN => n79);
   U79 : INV_X1 port map( A => B(15), ZN => n78);
   U80 : INV_X1 port map( A => B(16), ZN => n77);
   U81 : INV_X1 port map( A => B(17), ZN => n76);
   U82 : INV_X1 port map( A => B(18), ZN => n75);
   U83 : INV_X1 port map( A => B(19), ZN => n74);
   U84 : INV_X1 port map( A => B(20), ZN => n73);
   U85 : INV_X1 port map( A => B(21), ZN => n72);
   U86 : INV_X1 port map( A => B(22), ZN => n71);
   U87 : INV_X1 port map( A => B(23), ZN => n70);
   U88 : INV_X1 port map( A => B(24), ZN => n69);
   U89 : INV_X1 port map( A => B(25), ZN => n68);
   U90 : INV_X1 port map( A => B(26), ZN => n67);
   U91 : INV_X1 port map( A => B(27), ZN => n66);
   U92 : INV_X1 port map( A => B(28), ZN => n65);
   U93 : INV_X1 port map( A => B(29), ZN => n64);
   U94 : INV_X1 port map( A => B(30), ZN => n63);
   U95 : INV_X2 port map( A => n32, ZN => DIFF_30_port);
   U96 : INV_X2 port map( A => n33, ZN => DIFF_29_port);
   U97 : INV_X2 port map( A => n34, ZN => DIFF_28_port);
   U98 : INV_X2 port map( A => n35, ZN => DIFF_27_port);
   U99 : INV_X2 port map( A => n36, ZN => DIFF_26_port);
   U100 : INV_X2 port map( A => n37, ZN => DIFF_25_port);
   U101 : INV_X2 port map( A => n38, ZN => DIFF_24_port);
   U102 : INV_X2 port map( A => n39, ZN => DIFF_23_port);
   U103 : INV_X2 port map( A => n40, ZN => DIFF_22_port);
   U104 : INV_X2 port map( A => n41, ZN => DIFF_21_port);
   U105 : INV_X2 port map( A => n42, ZN => DIFF_20_port);
   U106 : INV_X2 port map( A => n43, ZN => DIFF_19_port);
   U107 : INV_X2 port map( A => n44, ZN => DIFF_18_port);
   U108 : INV_X2 port map( A => n45, ZN => DIFF_17_port);
   U109 : INV_X2 port map( A => n46, ZN => DIFF_16_port);
   U110 : INV_X2 port map( A => n47, ZN => DIFF_15_port);
   U111 : INV_X2 port map( A => n48, ZN => DIFF_14_port);
   U112 : INV_X2 port map( A => n49, ZN => DIFF_13_port);
   U113 : INV_X2 port map( A => n50, ZN => DIFF_12_port);
   U114 : INV_X2 port map( A => n51, ZN => DIFF_11_port);
   U115 : INV_X2 port map( A => n52, ZN => DIFF_10_port);
   U116 : INV_X2 port map( A => n53, ZN => DIFF_9_port);
   U117 : INV_X2 port map( A => n54, ZN => DIFF_8_port);
   U118 : INV_X2 port map( A => n55, ZN => DIFF_7_port);
   U119 : INV_X2 port map( A => n56, ZN => DIFF_6_port);
   U120 : INV_X2 port map( A => n57, ZN => DIFF_5_port);
   U121 : INV_X2 port map( A => n58, ZN => DIFF_4_port);
   U122 : INV_X2 port map( A => n59, ZN => DIFF_3_port);
   U123 : INV_X2 port map( A => n60, ZN => DIFF_2_port);
   U124 : INV_X2 port map( A => n61, ZN => DIFF_1_port);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT64_DW01_add_0 is

   port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (63 downto 0);  CO : out std_logic);

end RCA_NBIT64_DW01_add_0;

architecture SYN_rpl of RCA_NBIT64_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_29_port, carry_28_port, carry_27_port, carry_26_port, 
      carry_25_port, carry_24_port, carry_23_port, carry_22_port, carry_21_port
      , carry_20_port, carry_19_port, carry_18_port, carry_17_port, 
      carry_16_port, carry_15_port, carry_14_port, carry_13_port, carry_12_port
      , carry_11_port, carry_10_port, carry_9_port, carry_8_port, carry_7_port,
      carry_6_port, carry_5_port, carry_4_port, carry_3_port, carry_2_port, n1,
      n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, 
      n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, 
      n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, 
      n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, 
      n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, 
      n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, 
      n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, 
      n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, 
      n753, n754, n755, n756, n757, n758, n759, n760, n761, n614, n615, n616, 
      n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, 
      n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, 
      n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, 
      n653, n654, n655, n656 : std_logic;

begin
   
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U140 : XOR2_X1 port map( A => n657, B => n658, Z => SUM(63));
   U141 : XOR2_X1 port map( A => n666, B => n667, Z => SUM(61));
   U142 : XOR2_X1 port map( A => n617, B => n672, Z => SUM(59));
   U143 : XOR2_X1 port map( A => n675, B => n673, Z => SUM(58));
   U144 : XOR2_X1 port map( A => n618, B => B(58), Z => n675);
   U145 : XOR2_X1 port map( A => n677, B => n678, Z => SUM(57));
   U146 : XOR2_X1 port map( A => B(57), B => A(57), Z => n678);
   U147 : XOR2_X1 port map( A => n681, B => n621, Z => SUM(56));
   U148 : XOR2_X1 port map( A => n620, B => B(56), Z => n681);
   U149 : XOR2_X1 port map( A => n682, B => n684, Z => SUM(55));
   U150 : XOR2_X1 port map( A => n690, B => n624, Z => SUM(53));
   U151 : XOR2_X1 port map( A => n691, B => n693, Z => SUM(52));
   U152 : XOR2_X1 port map( A => n625, B => B(52), Z => n693);
   U153 : XOR2_X1 port map( A => n697, B => n699, Z => SUM(50));
   U154 : XOR2_X1 port map( A => n703, B => n705, Z => SUM(48));
   U155 : XOR2_X1 port map( A => n712, B => n714, Z => SUM(45));
   U156 : XOR2_X1 port map( A => B(45), B => A(45), Z => n714);
   U157 : XOR2_X1 port map( A => n718, B => n720, Z => SUM(43));
   U158 : XOR2_X1 port map( A => B(43), B => A(43), Z => n720);
   U159 : XOR2_X1 port map( A => n638, B => n723, Z => SUM(42));
   U160 : XOR2_X1 port map( A => n724, B => n726, Z => SUM(41));
   U161 : XOR2_X1 port map( A => B(41), B => A(41), Z => n726);
   U162 : XOR2_X1 port map( A => n641, B => n729, Z => SUM(40));
   U163 : XOR2_X1 port map( A => B(40), B => A(40), Z => n729);
   U164 : XOR2_X1 port map( A => n730, B => n732, Z => SUM(39));
   U165 : XOR2_X1 port map( A => B(39), B => A(39), Z => n732);
   U166 : XOR2_X1 port map( A => n643, B => n735, Z => SUM(38));
   U167 : XOR2_X1 port map( A => B(38), B => A(38), Z => n735);
   U168 : XOR2_X1 port map( A => n736, B => n738, Z => SUM(37));
   U169 : XOR2_X1 port map( A => B(37), B => A(37), Z => n738);
   U170 : XOR2_X1 port map( A => n646, B => n741, Z => SUM(36));
   U171 : XOR2_X1 port map( A => B(36), B => A(36), Z => n741);
   U172 : XOR2_X1 port map( A => n742, B => n744, Z => SUM(35));
   U173 : XOR2_X1 port map( A => B(35), B => A(35), Z => n744);
   U174 : XOR2_X1 port map( A => n649, B => n747, Z => SUM(34));
   U175 : XOR2_X1 port map( A => B(34), B => A(34), Z => n747);
   U176 : XOR2_X1 port map( A => n748, B => n750, Z => SUM(33));
   U177 : XOR2_X1 port map( A => B(33), B => A(33), Z => n750);
   U178 : XOR2_X1 port map( A => n652, B => n753, Z => SUM(32));
   U179 : XOR2_X1 port map( A => n653, B => n755, Z => SUM(31));
   U180 : XOR2_X1 port map( A => B(31), B => A(31), Z => n755);
   U181 : XOR2_X1 port map( A => n654, B => n758, Z => SUM(30));
   U182 : XOR2_X1 port map( A => B(30), B => A(30), Z => n758);
   U183 : XOR2_X1 port map( A => A(29), B => n761, Z => SUM(29));
   U184 : XOR2_X1 port map( A => carry_29_port, B => B(29), Z => n761);
   U185 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : INV_X1 port map( A => A(32), ZN => n651);
   U2 : INV_X1 port map( A => n727, ZN => n641);
   U3 : INV_X1 port map( A => A(42), ZN => n637);
   U4 : INV_X1 port map( A => A(46), ZN => n631);
   U5 : INV_X1 port map( A => n751, ZN => n652);
   U6 : INV_X1 port map( A => A(52), ZN => n625);
   U7 : INV_X1 port map( A => A(56), ZN => n620);
   U8 : INV_X1 port map( A => n715, ZN => n635);
   U9 : INV_X1 port map( A => A(58), ZN => n618);
   U10 : INV_X1 port map( A => n745, ZN => n649);
   U11 : INV_X1 port map( A => n739, ZN => n646);
   U12 : INV_X1 port map( A => n680, ZN => n621);
   U13 : INV_X1 port map( A => n689, ZN => n624);
   U14 : INV_X1 port map( A => n721, ZN => n638);
   U15 : INV_X1 port map( A => n733, ZN => n643);
   U16 : INV_X1 port map( A => n671, ZN => n617);
   U17 : OAI22_X1 port map( A1 => A(54), A2 => n685, B1 => B(54), B2 => n686, 
                           ZN => n682);
   U18 : AND2_X1 port map( A1 => n685, A2 => A(54), ZN => n686);
   U19 : OAI22_X1 port map( A1 => A(60), A2 => n665, B1 => B(60), B2 => n668, 
                           ZN => n666);
   U20 : AND2_X1 port map( A1 => A(60), A2 => n665, ZN => n668);
   U21 : AOI22_X1 port map( A1 => A(57), A2 => B(57), B1 => n676, B2 => n677, 
                           ZN => n673);
   U22 : OR2_X1 port map( A1 => B(57), A2 => A(57), ZN => n676);
   U23 : OAI22_X1 port map( A1 => A(31), A2 => n653, B1 => B(31), B2 => n754, 
                           ZN => n751);
   U24 : AND2_X1 port map( A1 => n653, A2 => A(31), ZN => n754);
   U25 : OAI22_X1 port map( A1 => n706, A2 => B(47), B1 => A(47), B2 => n707, 
                           ZN => n703);
   U26 : AND2_X1 port map( A1 => n707, A2 => A(47), ZN => n706);
   U27 : OAI22_X1 port map( A1 => n700, A2 => B(49), B1 => A(49), B2 => n701, 
                           ZN => n697);
   U28 : AND2_X1 port map( A1 => n701, A2 => A(49), ZN => n700);
   U29 : OAI22_X1 port map( A1 => n694, A2 => B(51), B1 => A(51), B2 => n695, 
                           ZN => n691);
   U30 : AND2_X1 port map( A1 => n695, A2 => A(51), ZN => n694);
   U31 : AOI21_X1 port map( B1 => n617, B2 => n616, A => n670, ZN => n665);
   U32 : INV_X1 port map( A => A(59), ZN => n616);
   U33 : AOI21_X1 port map( B1 => n671, B2 => A(59), A => B(59), ZN => n670);
   U34 : AOI22_X1 port map( A1 => n730, A2 => A(39), B1 => n731, B2 => B(39), 
                           ZN => n727);
   U35 : OR2_X1 port map( A1 => A(39), A2 => n730, ZN => n731);
   U36 : OAI21_X1 port map( B1 => A(45), B2 => n712, A => n633, ZN => n709);
   U37 : INV_X1 port map( A => n713, ZN => n633);
   U38 : AOI21_X1 port map( B1 => n712, B2 => A(45), A => B(45), ZN => n713);
   U39 : AOI21_X1 port map( B1 => n623, B2 => n624, A => n688, ZN => n685);
   U40 : INV_X1 port map( A => A(53), ZN => n623);
   U41 : AOI21_X1 port map( B1 => n689, B2 => A(53), A => B(53), ZN => n688);
   U42 : AOI21_X1 port map( B1 => n631, B2 => n709, A => n710, ZN => n707);
   U43 : AOI21_X1 port map( B1 => n632, B2 => A(46), A => B(46), ZN => n710);
   U44 : INV_X1 port map( A => n709, ZN => n632);
   U45 : OAI21_X1 port map( B1 => n703, B2 => n629, A => n704, ZN => n701);
   U46 : INV_X1 port map( A => A(48), ZN => n629);
   U47 : OAI21_X1 port map( B1 => n630, B2 => A(48), A => B(48), ZN => n704);
   U48 : INV_X1 port map( A => n703, ZN => n630);
   U49 : OAI21_X1 port map( B1 => n697, B2 => n627, A => n698, ZN => n695);
   U50 : INV_X1 port map( A => A(50), ZN => n627);
   U51 : OAI21_X1 port map( B1 => n628, B2 => A(50), A => B(50), ZN => n698);
   U52 : INV_X1 port map( A => n697, ZN => n628);
   U53 : AOI21_X1 port map( B1 => n640, B2 => n727, A => n728, ZN => n724);
   U54 : INV_X1 port map( A => A(40), ZN => n640);
   U55 : AOI21_X1 port map( B1 => n641, B2 => A(40), A => B(40), ZN => n728);
   U56 : OAI21_X1 port map( B1 => n751, B2 => n651, A => n752, ZN => n748);
   U57 : OAI21_X1 port map( B1 => n652, B2 => A(32), A => B(32), ZN => n752);
   U58 : OAI21_X1 port map( B1 => n745, B2 => n648, A => n746, ZN => n742);
   U59 : INV_X1 port map( A => A(34), ZN => n648);
   U60 : OAI21_X1 port map( B1 => n649, B2 => A(34), A => B(34), ZN => n746);
   U61 : OAI21_X1 port map( B1 => n739, B2 => n645, A => n740, ZN => n736);
   U62 : INV_X1 port map( A => A(36), ZN => n645);
   U63 : OAI21_X1 port map( B1 => n646, B2 => A(36), A => B(36), ZN => n740);
   U64 : OAI21_X1 port map( B1 => n721, B2 => n637, A => n722, ZN => n718);
   U65 : OAI21_X1 port map( B1 => n638, B2 => A(42), A => B(42), ZN => n722);
   U66 : OAI21_X1 port map( B1 => n715, B2 => n634, A => n716, ZN => n712);
   U67 : INV_X1 port map( A => A(44), ZN => n634);
   U68 : OAI21_X1 port map( B1 => n635, B2 => A(44), A => B(44), ZN => n716);
   U69 : AOI21_X1 port map( B1 => n618, B2 => n673, A => n674, ZN => n671);
   U70 : AOI21_X1 port map( B1 => n619, B2 => A(58), A => B(58), ZN => n674);
   U71 : INV_X1 port map( A => n673, ZN => n619);
   U72 : OAI21_X1 port map( B1 => n733, B2 => n642, A => n734, ZN => n730);
   U73 : INV_X1 port map( A => A(38), ZN => n642);
   U74 : OAI21_X1 port map( B1 => n643, B2 => A(38), A => B(38), ZN => n734);
   U75 : OAI21_X1 port map( B1 => n691, B2 => n625, A => n692, ZN => n689);
   U76 : OAI21_X1 port map( B1 => n626, B2 => A(52), A => B(52), ZN => n692);
   U77 : INV_X1 port map( A => n691, ZN => n626);
   U78 : OAI21_X1 port map( B1 => n682, B2 => n656, A => n683, ZN => n680);
   U79 : INV_X1 port map( A => B(55), ZN => n656);
   U80 : OAI21_X1 port map( B1 => n622, B2 => B(55), A => A(55), ZN => n683);
   U81 : INV_X1 port map( A => n682, ZN => n622);
   U82 : OAI21_X1 port map( B1 => A(33), B2 => n748, A => n650, ZN => n745);
   U83 : INV_X1 port map( A => n749, ZN => n650);
   U84 : AOI21_X1 port map( B1 => n748, B2 => A(33), A => B(33), ZN => n749);
   U85 : OAI21_X1 port map( B1 => A(35), B2 => n742, A => n647, ZN => n739);
   U86 : INV_X1 port map( A => n743, ZN => n647);
   U87 : AOI21_X1 port map( B1 => n742, B2 => A(35), A => B(35), ZN => n743);
   U88 : OAI21_X1 port map( B1 => A(43), B2 => n718, A => n636, ZN => n715);
   U89 : INV_X1 port map( A => n719, ZN => n636);
   U90 : AOI21_X1 port map( B1 => n718, B2 => A(43), A => B(43), ZN => n719);
   U91 : OAI21_X1 port map( B1 => n724, B2 => A(41), A => n639, ZN => n721);
   U92 : INV_X1 port map( A => n725, ZN => n639);
   U93 : AOI21_X1 port map( B1 => n724, B2 => A(41), A => B(41), ZN => n725);
   U94 : OAI21_X1 port map( B1 => A(37), B2 => n736, A => n644, ZN => n733);
   U95 : INV_X1 port map( A => n737, ZN => n644);
   U96 : AOI21_X1 port map( B1 => n736, B2 => A(37), A => B(37), ZN => n737);
   U97 : OAI21_X1 port map( B1 => n621, B2 => n620, A => n679, ZN => n677);
   U98 : OAI21_X1 port map( B1 => A(56), B2 => n680, A => B(56), ZN => n679);
   U99 : NAND2_X1 port map( A1 => n662, A2 => n663, ZN => n660);
   U100 : OAI21_X1 port map( B1 => B(61), B2 => n614, A => A(61), ZN => n662);
   U101 : OAI211_X1 port map( C1 => A(60), C2 => B(60), A => n615, B => B(61), 
                           ZN => n663);
   U102 : INV_X1 port map( A => n666, ZN => n614);
   U103 : XNOR2_X1 port map( A => A(61), B => B(61), ZN => n667);
   U104 : XNOR2_X1 port map( A => B(55), B => A(55), ZN => n684);
   U105 : XNOR2_X1 port map( A => A(48), B => B(48), ZN => n705);
   U106 : XNOR2_X1 port map( A => A(50), B => B(50), ZN => n699);
   U107 : XNOR2_X1 port map( A => A(59), B => B(59), ZN => n672);
   U108 : XNOR2_X1 port map( A => B(32), B => n651, ZN => n753);
   U109 : XNOR2_X1 port map( A => B(42), B => n637, ZN => n723);
   U110 : XNOR2_X1 port map( A => B(63), B => A(63), ZN => n658);
   U111 : OAI22_X1 port map( A1 => n659, A2 => n660, B1 => B(62), B2 => A(62), 
                           ZN => n657);
   U112 : XNOR2_X1 port map( A => n661, B => n660, ZN => SUM(62));
   U113 : XNOR2_X1 port map( A => A(62), B => B(62), ZN => n661);
   U114 : XNOR2_X1 port map( A => n702, B => n701, ZN => SUM(49));
   U115 : XNOR2_X1 port map( A => A(49), B => B(49), ZN => n702);
   U116 : XNOR2_X1 port map( A => n696, B => n695, ZN => SUM(51));
   U117 : XNOR2_X1 port map( A => A(51), B => B(51), ZN => n696);
   U118 : XNOR2_X1 port map( A => A(53), B => B(53), ZN => n690);
   U119 : XNOR2_X1 port map( A => n665, B => n669, ZN => SUM(60));
   U120 : XNOR2_X1 port map( A => A(60), B => B(60), ZN => n669);
   U121 : XNOR2_X1 port map( A => n707, B => n708, ZN => SUM(47));
   U122 : XNOR2_X1 port map( A => A(47), B => B(47), ZN => n708);
   U123 : XNOR2_X1 port map( A => n635, B => n717, ZN => SUM(44));
   U124 : XNOR2_X1 port map( A => A(44), B => B(44), ZN => n717);
   U125 : XNOR2_X1 port map( A => n685, B => n687, ZN => SUM(54));
   U126 : XNOR2_X1 port map( A => A(54), B => B(54), ZN => n687);
   U127 : XNOR2_X1 port map( A => n709, B => n711, ZN => SUM(46));
   U128 : XNOR2_X1 port map( A => B(46), B => n631, ZN => n711);
   U129 : INV_X1 port map( A => n759, ZN => n654);
   U130 : OAI21_X1 port map( B1 => B(29), B2 => A(29), A => n655, ZN => n759);
   U131 : INV_X1 port map( A => n760, ZN => n655);
   U132 : AOI21_X1 port map( B1 => A(29), B2 => B(29), A => carry_29_port, ZN 
                           => n760);
   U133 : INV_X1 port map( A => n756, ZN => n653);
   U134 : OAI22_X1 port map( A1 => A(30), A2 => n654, B1 => B(30), B2 => n757, 
                           ZN => n756);
   U135 : AND2_X1 port map( A1 => n654, A2 => A(30), ZN => n757);
   U136 : AND2_X1 port map( A1 => A(62), A2 => B(62), ZN => n659);
   U137 : INV_X1 port map( A => n664, ZN => n615);
   U138 : AOI21_X1 port map( B1 => A(60), B2 => B(60), A => n665, ZN => n664);
   U139 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT62_DW01_add_0 is

   port( A, B : in std_logic_vector (61 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (61 downto 0);  CO : out std_logic);

end RCA_NBIT62_DW01_add_0;

architecture SYN_rpl of RCA_NBIT62_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_28_port, carry_27_port, carry_26_port, carry_25_port, 
      carry_24_port, carry_23_port, carry_22_port, carry_21_port, carry_20_port
      , carry_19_port, carry_18_port, carry_17_port, carry_16_port, 
      carry_15_port, carry_14_port, carry_13_port, carry_12_port, carry_11_port
      , carry_10_port, carry_9_port, carry_8_port, carry_7_port, carry_6_port, 
      carry_5_port, carry_4_port, carry_3_port, carry_2_port, n1, carry_59_port
      , carry_58_port, n556, n557, n558, n559, n560, n561, n562, n563, n564, 
      n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, 
      n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, 
      n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, 
      n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, 
      n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, 
      n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, 
      n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, 
      n649, n650, n651, n652, n653, n654, n509, n510, n511, n512, n513, n514, 
      n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, 
      n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, 
      n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, 
      n551, n552, n553, n554, n555 : std_logic;

begin
   
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U1_57 : FA_X1 port map( A => A(57), B => B(57), CI => n654, CO => 
                           carry_58_port, S => SUM(57));
   U1_58 : FA_X1 port map( A => A(58), B => B(58), CI => carry_58_port, CO => 
                           carry_59_port, S => SUM(58));
   U142 : XOR2_X1 port map( A => B(61), B => A(61), Z => n559);
   U143 : XOR2_X1 port map( A => n509, B => n561, Z => SUM(60));
   U144 : XOR2_X1 port map( A => B(60), B => A(60), Z => n561);
   U145 : XOR2_X1 port map( A => A(59), B => n564, Z => SUM(59));
   U146 : XOR2_X1 port map( A => carry_59_port, B => B(59), Z => n564);
   U147 : XOR2_X1 port map( A => n556, B => n565, Z => SUM(56));
   U148 : XOR2_X1 port map( A => n511, B => B(56), Z => n565);
   U149 : XOR2_X1 port map( A => n569, B => n571, Z => SUM(54));
   U150 : XOR2_X1 port map( A => n514, B => B(54), Z => n571);
   U151 : XOR2_X1 port map( A => n572, B => n576, Z => SUM(53));
   U152 : XOR2_X1 port map( A => B(53), B => A(53), Z => n576);
   U153 : XOR2_X1 port map( A => n578, B => n581, Z => SUM(52));
   U154 : XOR2_X1 port map( A => B(52), B => A(52), Z => n581);
   U155 : XOR2_X1 port map( A => n579, B => n583, Z => SUM(51));
   U156 : XOR2_X1 port map( A => B(51), B => A(51), Z => n583);
   U157 : XOR2_X1 port map( A => n519, B => n586, Z => SUM(50));
   U158 : XOR2_X1 port map( A => B(50), B => A(50), Z => n586);
   U159 : XOR2_X1 port map( A => n590, B => n592, Z => SUM(48));
   U160 : XOR2_X1 port map( A => n614, B => n616, Z => SUM(40));
   U161 : XOR2_X1 port map( A => n618, B => n619, Z => SUM(39));
   U162 : XOR2_X1 port map( A => n621, B => n622, Z => SUM(38));
   U163 : XOR2_X1 port map( A => n626, B => n628, Z => SUM(36));
   U164 : XOR2_X1 port map( A => n629, B => n631, Z => SUM(35));
   U165 : XOR2_X1 port map( A => B(35), B => A(35), Z => n631);
   U166 : XOR2_X1 port map( A => n632, B => n634, Z => SUM(34));
   U167 : XOR2_X1 port map( A => n540, B => B(34), Z => n634);
   U168 : XOR2_X1 port map( A => n635, B => n637, Z => SUM(33));
   U169 : XOR2_X1 port map( A => B(33), B => A(33), Z => n637);
   U170 : XOR2_X1 port map( A => n639, B => n644, Z => SUM(32));
   U171 : XOR2_X1 port map( A => n543, B => B(32), Z => n644);
   U172 : XOR2_X1 port map( A => n645, B => n646, Z => SUM(31));
   U173 : XOR2_X1 port map( A => n554, B => A(31), Z => n646);
   U174 : XOR2_X1 port map( A => n547, B => n648, Z => SUM(30));
   U175 : XOR2_X1 port map( A => B(30), B => A(30), Z => n648);
   U176 : XOR2_X1 port map( A => n549, B => n650, Z => SUM(29));
   U177 : XOR2_X1 port map( A => B(29), B => A(29), Z => n650);
   U178 : XOR2_X1 port map( A => A(28), B => n653, Z => SUM(28));
   U179 : XOR2_X1 port map( A => carry_28_port, B => B(28), Z => n653);
   U180 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : OAI21_X1 port map( B1 => A(30), B2 => n547, A => n647, ZN => n645);
   U2 : OAI21_X1 port map( B1 => n643, B2 => n546, A => n555, ZN => n647);
   U3 : OAI21_X1 port map( B1 => n577, B2 => n552, A => n574, ZN => n572);
   U4 : AND2_X1 port map( A1 => n516, A2 => n575, ZN => n577);
   U5 : NOR2_X1 port map( A1 => n579, A2 => A(51), ZN => n580);
   U6 : OAI21_X1 port map( B1 => A(31), B2 => n545, A => n641, ZN => n639);
   U7 : INV_X1 port map( A => n645, ZN => n545);
   U8 : INV_X1 port map( A => A(30), ZN => n546);
   U9 : NOR2_X1 port map( A1 => n547, A2 => A(30), ZN => n642);
   U10 : NAND2_X1 port map( A1 => A(52), A2 => n578, ZN => n574);
   U11 : INV_X1 port map( A => A(44), ZN => n527);
   U12 : INV_X1 port map( A => n643, ZN => n547);
   U13 : INV_X1 port map( A => A(42), ZN => n530);
   U14 : INV_X1 port map( A => A(46), ZN => n524);
   U15 : INV_X1 port map( A => A(56), ZN => n511);
   U16 : INV_X1 port map( A => A(31), ZN => n544);
   U17 : INV_X1 port map( A => A(52), ZN => n516);
   U18 : INV_X1 port map( A => A(34), ZN => n540);
   U19 : INV_X1 port map( A => A(32), ZN => n543);
   U20 : INV_X1 port map( A => n584, ZN => n519);
   U21 : XNOR2_X1 port map( A => A(48), B => B(48), ZN => n592);
   U22 : XNOR2_X1 port map( A => n558, B => n559, ZN => SUM(61));
   U23 : OAI22_X1 port map( A1 => n560, A2 => B(60), B1 => n509, B2 => A(60), 
                           ZN => n558);
   U24 : AND2_X1 port map( A1 => A(60), A2 => n509, ZN => n560);
   U25 : XNOR2_X1 port map( A => A(40), B => B(40), ZN => n616);
   U26 : XNOR2_X1 port map( A => A(38), B => B(38), ZN => n622);
   U27 : XNOR2_X1 port map( A => A(36), B => B(36), ZN => n628);
   U28 : OAI22_X1 port map( A1 => n535, A2 => A(39), B1 => B(39), B2 => n617, 
                           ZN => n614);
   U29 : AND2_X1 port map( A1 => n535, A2 => A(39), ZN => n617);
   U30 : INV_X1 port map( A => n618, ZN => n535);
   U31 : XNOR2_X1 port map( A => A(39), B => B(39), ZN => n619);
   U32 : OAI22_X1 port map( A1 => n569, A2 => n514, B1 => n570, B2 => n551, ZN 
                           => n566);
   U33 : AND2_X1 port map( A1 => n569, A2 => n514, ZN => n570);
   U34 : INV_X1 port map( A => B(54), ZN => n551);
   U35 : OAI22_X1 port map( A1 => A(53), A2 => n572, B1 => B(53), B2 => n573, 
                           ZN => n569);
   U36 : AOI221_X1 port map( B1 => n574, B2 => n552, C1 => n575, C2 => n516, A 
                           => n515, ZN => n573);
   U37 : INV_X1 port map( A => A(53), ZN => n515);
   U38 : OAI22_X1 port map( A1 => A(37), A2 => n623, B1 => B(37), B2 => n624, 
                           ZN => n621);
   U39 : AND2_X1 port map( A1 => n623, A2 => A(37), ZN => n624);
   U40 : OAI22_X1 port map( A1 => n638, A2 => n553, B1 => n639, B2 => n543, ZN 
                           => n635);
   U41 : AOI21_X1 port map( B1 => n640, B2 => n641, A => A(32), ZN => n638);
   U42 : INV_X1 port map( A => B(32), ZN => n553);
   U43 : OAI221_X1 port map( B1 => n642, B2 => n555, C1 => n643, C2 => n546, A 
                           => n544, ZN => n640);
   U44 : OAI22_X1 port map( A1 => n536, A2 => B(38), B1 => n620, B2 => A(38), 
                           ZN => n618);
   U45 : AND2_X1 port map( A1 => n536, A2 => B(38), ZN => n620);
   U46 : INV_X1 port map( A => n621, ZN => n536);
   U47 : OAI21_X1 port map( B1 => n584, B2 => n518, A => n585, ZN => n579);
   U48 : INV_X1 port map( A => A(50), ZN => n518);
   U49 : OAI21_X1 port map( B1 => A(50), B2 => n519, A => B(50), ZN => n585);
   U50 : AOI21_X1 port map( B1 => n605, B2 => A(43), A => n529, ZN => n602);
   U51 : INV_X1 port map( A => n606, ZN => n529);
   U52 : OAI21_X1 port map( B1 => n605, B2 => A(43), A => B(43), ZN => n606);
   U53 : AOI21_X1 port map( B1 => n599, B2 => A(45), A => n526, ZN => n596);
   U54 : INV_X1 port map( A => n600, ZN => n526);
   U55 : OAI21_X1 port map( B1 => n599, B2 => A(45), A => B(45), ZN => n600);
   U56 : AOI21_X1 port map( B1 => n611, B2 => A(41), A => n532, ZN => n608);
   U57 : INV_X1 port map( A => n612, ZN => n532);
   U58 : OAI21_X1 port map( B1 => A(41), B2 => n611, A => B(41), ZN => n612);
   U59 : AOI21_X1 port map( B1 => n530, B2 => n608, A => n609, ZN => n605);
   U60 : AOI21_X1 port map( B1 => n531, B2 => A(42), A => B(42), ZN => n609);
   U61 : INV_X1 port map( A => n608, ZN => n531);
   U62 : AOI21_X1 port map( B1 => n527, B2 => n602, A => n603, ZN => n599);
   U63 : AOI21_X1 port map( B1 => n528, B2 => A(44), A => B(44), ZN => n603);
   U64 : INV_X1 port map( A => n602, ZN => n528);
   U65 : AOI21_X1 port map( B1 => n524, B2 => n596, A => n597, ZN => n593);
   U66 : AOI21_X1 port map( B1 => n525, B2 => A(46), A => B(46), ZN => n597);
   U67 : INV_X1 port map( A => n596, ZN => n525);
   U68 : OAI21_X1 port map( B1 => n614, B2 => n533, A => n615, ZN => n611);
   U69 : INV_X1 port map( A => A(40), ZN => n533);
   U70 : OAI21_X1 port map( B1 => n534, B2 => A(40), A => B(40), ZN => n615);
   U71 : INV_X1 port map( A => n614, ZN => n534);
   U72 : OAI21_X1 port map( B1 => n590, B2 => n521, A => n591, ZN => n587);
   U73 : INV_X1 port map( A => A(48), ZN => n521);
   U74 : OAI21_X1 port map( B1 => A(48), B2 => n522, A => B(48), ZN => n591);
   U75 : INV_X1 port map( A => n590, ZN => n522);
   U76 : XNOR2_X1 port map( A => n602, B => n604, ZN => SUM(44));
   U77 : XNOR2_X1 port map( A => B(44), B => n527, ZN => n604);
   U78 : AOI21_X1 port map( B1 => n537, B2 => n626, A => n627, ZN => n623);
   U79 : INV_X1 port map( A => A(36), ZN => n537);
   U80 : AOI21_X1 port map( B1 => n538, B2 => A(36), A => B(36), ZN => n627);
   U81 : INV_X1 port map( A => n626, ZN => n538);
   U82 : AOI22_X1 port map( A1 => n579, A2 => A(51), B1 => n517, B2 => B(51), 
                           ZN => n575);
   U83 : INV_X1 port map( A => n580, ZN => n517);
   U84 : XNOR2_X1 port map( A => n613, B => n611, ZN => SUM(41));
   U85 : XNOR2_X1 port map( A => A(41), B => B(41), ZN => n613);
   U86 : OAI21_X1 port map( B1 => A(29), B2 => n549, A => n548, ZN => n643);
   U87 : INV_X1 port map( A => n649, ZN => n548);
   U88 : AOI21_X1 port map( B1 => n549, B2 => A(29), A => B(29), ZN => n649);
   U89 : XNOR2_X1 port map( A => n589, B => n587, ZN => SUM(49));
   U90 : XNOR2_X1 port map( A => A(49), B => B(49), ZN => n589);
   U91 : XNOR2_X1 port map( A => n623, B => n625, ZN => SUM(37));
   U92 : XNOR2_X1 port map( A => A(37), B => B(37), ZN => n625);
   U93 : XNOR2_X1 port map( A => n605, B => n607, ZN => SUM(43));
   U94 : XNOR2_X1 port map( A => A(43), B => B(43), ZN => n607);
   U95 : XNOR2_X1 port map( A => n599, B => n601, ZN => SUM(45));
   U96 : XNOR2_X1 port map( A => A(45), B => B(45), ZN => n601);
   U97 : XNOR2_X1 port map( A => n593, B => n595, ZN => SUM(47));
   U98 : XNOR2_X1 port map( A => A(47), B => B(47), ZN => n595);
   U99 : OAI21_X1 port map( B1 => A(35), B2 => n629, A => n539, ZN => n626);
   U100 : INV_X1 port map( A => n630, ZN => n539);
   U101 : AOI21_X1 port map( B1 => n629, B2 => A(35), A => B(35), ZN => n630);
   U102 : OAI21_X1 port map( B1 => n632, B2 => n540, A => n633, ZN => n629);
   U103 : OAI21_X1 port map( B1 => n541, B2 => A(34), A => B(34), ZN => n633);
   U104 : INV_X1 port map( A => n632, ZN => n541);
   U105 : OAI21_X1 port map( B1 => A(33), B2 => n635, A => n542, ZN => n632);
   U106 : INV_X1 port map( A => n636, ZN => n542);
   U107 : AOI21_X1 port map( B1 => n635, B2 => A(33), A => B(33), ZN => n636);
   U108 : OAI21_X1 port map( B1 => A(55), B2 => n566, A => n513, ZN => n556);
   U109 : INV_X1 port map( A => n567, ZN => n513);
   U110 : AOI21_X1 port map( B1 => n566, B2 => A(55), A => B(55), ZN => n567);
   U111 : OAI21_X1 port map( B1 => n593, B2 => A(47), A => n523, ZN => n590);
   U112 : INV_X1 port map( A => n594, ZN => n523);
   U113 : AOI21_X1 port map( B1 => n593, B2 => A(47), A => B(47), ZN => n594);
   U114 : XNOR2_X1 port map( A => n568, B => n566, ZN => SUM(55));
   U115 : XNOR2_X1 port map( A => A(55), B => B(55), ZN => n568);
   U116 : AOI21_X1 port map( B1 => n587, B2 => A(49), A => n520, ZN => n584);
   U117 : INV_X1 port map( A => n588, ZN => n520);
   U118 : OAI21_X1 port map( B1 => A(49), B2 => n587, A => B(49), ZN => n588);
   U119 : OAI21_X1 port map( B1 => n512, B2 => A(56), A => B(56), ZN => n557);
   U120 : INV_X1 port map( A => n556, ZN => n512);
   U121 : XNOR2_X1 port map( A => n596, B => n598, ZN => SUM(46));
   U122 : XNOR2_X1 port map( A => B(46), B => n524, ZN => n598);
   U123 : OAI21_X1 port map( B1 => n645, B2 => n544, A => n554, ZN => n641);
   U124 : XNOR2_X1 port map( A => n608, B => n610, ZN => SUM(42));
   U125 : XNOR2_X1 port map( A => B(42), B => n530, ZN => n610);
   U126 : INV_X1 port map( A => B(52), ZN => n552);
   U127 : INV_X1 port map( A => B(30), ZN => n555);
   U128 : NOR2_X1 port map( A1 => n580, A2 => n582, ZN => n578);
   U129 : AOI21_X1 port map( B1 => n579, B2 => A(51), A => B(51), ZN => n582);
   U130 : INV_X1 port map( A => n562, ZN => n509);
   U131 : OAI21_X1 port map( B1 => B(59), B2 => A(59), A => n510, ZN => n562);
   U132 : INV_X1 port map( A => n563, ZN => n510);
   U133 : AOI21_X1 port map( B1 => A(59), B2 => B(59), A => carry_59_port, ZN 
                           => n563);
   U134 : OAI21_X1 port map( B1 => n556, B2 => n511, A => n557, ZN => n654);
   U135 : INV_X1 port map( A => n651, ZN => n549);
   U136 : AOI21_X1 port map( B1 => A(28), B2 => B(28), A => n550, ZN => n651);
   U137 : INV_X1 port map( A => n652, ZN => n550);
   U138 : OAI21_X1 port map( B1 => A(28), B2 => B(28), A => carry_28_port, ZN 
                           => n652);
   U139 : INV_X1 port map( A => A(54), ZN => n514);
   U140 : INV_X1 port map( A => B(31), ZN => n554);
   U141 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT60_DW01_add_0 is

   port( A, B : in std_logic_vector (59 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (59 downto 0);  CO : out std_logic);

end RCA_NBIT60_DW01_add_0;

architecture SYN_rpl of RCA_NBIT60_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_30_port, carry_26_port, carry_25_port, carry_24_port, 
      carry_23_port, carry_22_port, carry_21_port, carry_20_port, carry_19_port
      , carry_18_port, carry_17_port, carry_16_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_10_port
      , carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, n1, n477, n478, n479, n480, 
      n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, 
      n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, 
      n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, 
      n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, 
      n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, 
      n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, 
      n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, 
      n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476 : std_logic;

begin
   
   U1_29 : FA_X1 port map( A => B(29), B => n472, CI => A(29), CO => 
                           carry_30_port, S => SUM(29));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U144 : XOR2_X1 port map( A => B(59), B => A(59), Z => n481);
   U145 : XOR2_X1 port map( A => n483, B => n484, Z => SUM(58));
   U146 : XOR2_X1 port map( A => B(58), B => A(58), Z => n484);
   U147 : XOR2_X1 port map( A => n488, B => n490, Z => SUM(56));
   U148 : XOR2_X1 port map( A => B(56), B => A(56), Z => n490);
   U149 : XOR2_X1 port map( A => n494, B => n496, Z => SUM(54));
   U150 : XOR2_X1 port map( A => B(54), B => A(54), Z => n496);
   U151 : XOR2_X1 port map( A => B(53), B => A(53), Z => n499);
   U152 : XOR2_X1 port map( A => B(52), B => A(52), Z => n502);
   U153 : XOR2_X1 port map( A => n506, B => n507, Z => SUM(51));
   U154 : XOR2_X1 port map( A => n509, B => n508, Z => SUM(50));
   U155 : XOR2_X1 port map( A => n451, B => B(46), Z => n521);
   U156 : XOR2_X1 port map( A => n455, B => n527, Z => SUM(44));
   U157 : XOR2_X1 port map( A => B(44), B => A(44), Z => n527);
   U158 : XOR2_X1 port map( A => n457, B => B(42), Z => n533);
   U159 : XOR2_X1 port map( A => n546, B => n548, Z => SUM(37));
   U160 : XOR2_X1 port map( A => B(37), B => A(37), Z => n548);
   U161 : XOR2_X1 port map( A => n555, B => n556, Z => SUM(35));
   U162 : XOR2_X1 port map( A => B(34), B => A(34), Z => n558);
   U163 : XOR2_X1 port map( A => B(33), B => A(33), Z => n561);
   U164 : XOR2_X1 port map( A => B(32), B => A(32), Z => n564);
   U165 : XOR2_X1 port map( A => B(31), B => A(31), Z => n567);
   U166 : XOR2_X1 port map( A => A(30), B => n569, Z => SUM(30));
   U167 : XOR2_X1 port map( A => carry_30_port, B => B(30), Z => n569);
   U168 : XOR2_X1 port map( A => n478, B => n570, Z => SUM(28));
   U169 : XOR2_X1 port map( A => B(28), B => A(28), Z => n570);
   U170 : XOR2_X1 port map( A => B(27), B => A(27), Z => n573);
   U171 : XOR2_X1 port map( A => carry_26_port, B => n574, Z => SUM(26));
   U172 : XOR2_X1 port map( A => A(26), B => B(26), Z => n574);
   U173 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : NOR2_X1 port map( A1 => n554, A2 => n553, ZN => n555);
   U2 : XNOR2_X1 port map( A => n476, B => A(35), ZN => n556);
   U3 : NOR2_X1 port map( A1 => n467, A2 => A(34), ZN => n553);
   U4 : NAND2_X1 port map( A1 => n508, A2 => n446, ZN => n504);
   U5 : INV_X1 port map( A => n531, ZN => n458);
   U6 : INV_X1 port map( A => A(38), ZN => n461);
   U7 : INV_X1 port map( A => A(36), ZN => n464);
   U8 : INV_X1 port map( A => n557, ZN => n467);
   U9 : INV_X1 port map( A => n491, ZN => n441);
   U10 : INV_X1 port map( A => n513, ZN => n449);
   U11 : INV_X1 port map( A => A(42), ZN => n457);
   U12 : INV_X1 port map( A => A(50), ZN => n446);
   U13 : INV_X1 port map( A => n519, ZN => n452);
   U14 : INV_X1 port map( A => n485, ZN => n437);
   U15 : INV_X1 port map( A => A(46), ZN => n451);
   U16 : INV_X1 port map( A => n525, ZN => n455);
   U17 : NAND2_X1 port map( A1 => n505, A2 => n504, ZN => n506);
   U18 : XNOR2_X1 port map( A => A(51), B => B(51), ZN => n507);
   U19 : XNOR2_X1 port map( A => n480, B => n481, ZN => SUM(59));
   U20 : OAI22_X1 port map( A1 => n482, A2 => B(58), B1 => n483, B2 => A(58), 
                           ZN => n480);
   U21 : AND2_X1 port map( A1 => A(58), A2 => n483, ZN => n482);
   U22 : XNOR2_X1 port map( A => A(50), B => B(50), ZN => n509);
   U23 : OAI22_X1 port map( A1 => A(52), A2 => n444, B1 => B(52), B2 => n500, 
                           ZN => n497);
   U24 : AND2_X1 port map( A1 => n444, A2 => A(52), ZN => n500);
   U25 : INV_X1 port map( A => n501, ZN => n444);
   U26 : AOI21_X1 port map( B1 => A(35), B2 => B(35), A => n552, ZN => n549);
   U27 : AOI211_X1 port map( C1 => n466, C2 => n476, A => n553, B => n554, ZN 
                           => n552);
   U28 : INV_X1 port map( A => A(35), ZN => n466);
   U29 : OAI22_X1 port map( A1 => A(54), A2 => n494, B1 => B(54), B2 => n495, 
                           ZN => n491);
   U30 : AND2_X1 port map( A1 => n494, A2 => A(54), ZN => n495);
   U31 : OAI22_X1 port map( A1 => n534, A2 => A(41), B1 => n459, B2 => B(41), 
                           ZN => n531);
   U32 : AND2_X1 port map( A1 => n459, A2 => B(41), ZN => n534);
   U33 : AOI21_X1 port map( B1 => A(51), B2 => B(51), A => n445, ZN => n501);
   U34 : INV_X1 port map( A => n503, ZN => n445);
   U35 : OAI211_X1 port map( C1 => A(51), C2 => B(51), A => n504, B => n505, ZN
                           => n503);
   U36 : AOI22_X1 port map( A1 => n574, A2 => carry_26_port, B1 => A(26), B2 =>
                           B(26), ZN => n571);
   U37 : AOI21_X1 port map( B1 => A(30), B2 => B(30), A => n471, ZN => n566);
   U38 : INV_X1 port map( A => n568, ZN => n471);
   U39 : OAI21_X1 port map( B1 => A(30), B2 => B(30), A => carry_30_port, ZN =>
                           n568);
   U40 : AOI21_X1 port map( B1 => n546, B2 => A(37), A => n463, ZN => n543);
   U41 : INV_X1 port map( A => n547, ZN => n463);
   U42 : OAI21_X1 port map( B1 => n546, B2 => A(37), A => B(37), ZN => n547);
   U43 : AOI21_X1 port map( B1 => n454, B2 => n525, A => n526, ZN => n522);
   U44 : INV_X1 port map( A => A(44), ZN => n454);
   U45 : AOI21_X1 port map( B1 => n455, B2 => A(44), A => B(44), ZN => n526);
   U46 : AOI21_X1 port map( B1 => n448, B2 => n513, A => n514, ZN => n510);
   U47 : INV_X1 port map( A => A(48), ZN => n448);
   U48 : AOI21_X1 port map( B1 => n449, B2 => A(48), A => B(48), ZN => n514);
   U49 : AOI22_X1 port map( A1 => n470, A2 => A(31), B1 => n565, B2 => B(31), 
                           ZN => n563);
   U50 : OR2_X1 port map( A1 => A(31), A2 => n470, ZN => n565);
   U51 : INV_X1 port map( A => n566, ZN => n470);
   U52 : AOI22_X1 port map( A1 => n469, A2 => A(32), B1 => n562, B2 => B(32), 
                           ZN => n560);
   U53 : OR2_X1 port map( A1 => A(32), A2 => n469, ZN => n562);
   U54 : INV_X1 port map( A => n563, ZN => n469);
   U55 : AOI22_X1 port map( A1 => n468, A2 => A(33), B1 => n559, B2 => B(33), 
                           ZN => n557);
   U56 : OR2_X1 port map( A1 => A(33), A2 => n468, ZN => n559);
   U57 : INV_X1 port map( A => n560, ZN => n468);
   U58 : OAI21_X1 port map( B1 => n531, B2 => n457, A => n532, ZN => n528);
   U59 : OAI21_X1 port map( B1 => A(42), B2 => n458, A => B(42), ZN => n532);
   U60 : OAI21_X1 port map( B1 => n519, B2 => n451, A => n520, ZN => n516);
   U61 : OAI21_X1 port map( B1 => n452, B2 => A(46), A => B(46), ZN => n520);
   U62 : XNOR2_X1 port map( A => n530, B => n528, ZN => SUM(43));
   U63 : XNOR2_X1 port map( A => A(43), B => B(43), ZN => n530);
   U64 : XNOR2_X1 port map( A => n518, B => n516, ZN => SUM(47));
   U65 : XNOR2_X1 port map( A => A(47), B => B(47), ZN => n518);
   U66 : XNOR2_X1 port map( A => n522, B => n524, ZN => SUM(45));
   U67 : XNOR2_X1 port map( A => A(45), B => B(45), ZN => n524);
   U68 : XNOR2_X1 port map( A => n549, B => n551, ZN => SUM(36));
   U69 : XNOR2_X1 port map( A => B(36), B => n464, ZN => n551);
   U70 : XNOR2_X1 port map( A => n459, B => n535, ZN => SUM(41));
   U71 : XNOR2_X1 port map( A => A(41), B => B(41), ZN => n535);
   U72 : XNOR2_X1 port map( A => n510, B => n512, ZN => SUM(49));
   U73 : XNOR2_X1 port map( A => A(49), B => B(49), ZN => n512);
   U74 : XNOR2_X1 port map( A => n441, B => n493, ZN => SUM(55));
   U75 : XNOR2_X1 port map( A => A(55), B => B(55), ZN => n493);
   U76 : XNOR2_X1 port map( A => n460, B => n538, ZN => SUM(40));
   U77 : XNOR2_X1 port map( A => A(40), B => B(40), ZN => n538);
   U78 : XNOR2_X1 port map( A => n449, B => n515, ZN => SUM(48));
   U79 : XNOR2_X1 port map( A => A(48), B => B(48), ZN => n515);
   U80 : AOI21_X1 port map( B1 => n461, B2 => n543, A => n544, ZN => n540);
   U81 : AOI21_X1 port map( B1 => n462, B2 => A(38), A => B(38), ZN => n544);
   U82 : INV_X1 port map( A => n543, ZN => n462);
   U83 : AOI21_X1 port map( B1 => n467, B2 => A(34), A => B(34), ZN => n554);
   U84 : AOI21_X1 port map( B1 => n510, B2 => A(49), A => n447, ZN => n508);
   U85 : INV_X1 port map( A => n511, ZN => n447);
   U86 : OAI21_X1 port map( B1 => n510, B2 => A(49), A => B(49), ZN => n511);
   U87 : AOI21_X1 port map( B1 => n464, B2 => n549, A => n550, ZN => n546);
   U88 : AOI21_X1 port map( B1 => n465, B2 => A(36), A => B(36), ZN => n550);
   U89 : INV_X1 port map( A => n549, ZN => n465);
   U90 : XNOR2_X1 port map( A => n540, B => n542, ZN => SUM(39));
   U91 : XNOR2_X1 port map( A => A(39), B => B(39), ZN => n542);
   U92 : XNOR2_X1 port map( A => n560, B => n561, ZN => SUM(33));
   U93 : XNOR2_X1 port map( A => n497, B => n499, ZN => SUM(53));
   U94 : XNOR2_X1 port map( A => n566, B => n567, ZN => SUM(31));
   U95 : XNOR2_X1 port map( A => n501, B => n502, ZN => SUM(52));
   U96 : OAI21_X1 port map( B1 => n491, B2 => n440, A => n492, ZN => n488);
   U97 : INV_X1 port map( A => A(55), ZN => n440);
   U98 : OAI21_X1 port map( B1 => n441, B2 => A(55), A => B(55), ZN => n492);
   U99 : XNOR2_X1 port map( A => A(57), B => B(57), ZN => n487);
   U100 : AOI21_X1 port map( B1 => n528, B2 => A(43), A => n456, ZN => n525);
   U101 : INV_X1 port map( A => n529, ZN => n456);
   U102 : OAI21_X1 port map( B1 => A(43), B2 => n528, A => B(43), ZN => n529);
   U103 : OAI21_X1 port map( B1 => n497, B2 => n442, A => n498, ZN => n494);
   U104 : INV_X1 port map( A => A(53), ZN => n442);
   U105 : OAI21_X1 port map( B1 => n443, B2 => A(53), A => B(53), ZN => n498);
   U106 : INV_X1 port map( A => n497, ZN => n443);
   U107 : AOI22_X1 port map( A1 => n478, A2 => A(28), B1 => n479, B2 => B(28), 
                           ZN => n477);
   U108 : OR2_X1 port map( A1 => A(28), A2 => n478, ZN => n479);
   U109 : XNOR2_X1 port map( A => n543, B => n545, ZN => SUM(38));
   U110 : XNOR2_X1 port map( A => B(38), B => n461, ZN => n545);
   U111 : OAI21_X1 port map( B1 => n571, B2 => n473, A => n572, ZN => n478);
   U112 : INV_X1 port map( A => A(27), ZN => n473);
   U113 : OAI21_X1 port map( B1 => A(27), B2 => n474, A => B(27), ZN => n572);
   U114 : INV_X1 port map( A => n571, ZN => n474);
   U115 : OAI21_X1 port map( B1 => n485, B2 => n439, A => n486, ZN => n483);
   U116 : INV_X1 port map( A => A(57), ZN => n439);
   U117 : OAI21_X1 port map( B1 => n437, B2 => A(57), A => B(57), ZN => n486);
   U118 : XNOR2_X1 port map( A => n557, B => n558, ZN => SUM(34));
   U119 : OAI21_X1 port map( B1 => A(47), B2 => n516, A => n450, ZN => n513);
   U120 : INV_X1 port map( A => n517, ZN => n450);
   U121 : AOI21_X1 port map( B1 => n516, B2 => A(47), A => B(47), ZN => n517);
   U122 : XNOR2_X1 port map( A => n458, B => n533, ZN => SUM(42));
   U123 : XNOR2_X1 port map( A => n452, B => n521, ZN => SUM(46));
   U124 : XNOR2_X1 port map( A => n563, B => n564, ZN => SUM(32));
   U125 : OAI21_X1 port map( B1 => A(45), B2 => n522, A => n453, ZN => n519);
   U126 : INV_X1 port map( A => n523, ZN => n453);
   U127 : AOI21_X1 port map( B1 => n522, B2 => A(45), A => B(45), ZN => n523);
   U128 : OAI21_X1 port map( B1 => A(56), B2 => n488, A => n438, ZN => n485);
   U129 : INV_X1 port map( A => n489, ZN => n438);
   U130 : AOI21_X1 port map( B1 => n488, B2 => A(56), A => B(56), ZN => n489);
   U131 : OAI21_X1 port map( B1 => n508, B2 => n446, A => n475, ZN => n505);
   U132 : INV_X1 port map( A => B(50), ZN => n475);
   U133 : INV_X1 port map( A => B(35), ZN => n476);
   U134 : INV_X1 port map( A => n477, ZN => n472);
   U135 : XNOR2_X1 port map( A => n571, B => n573, ZN => SUM(27));
   U136 : INV_X1 port map( A => n539, ZN => n460);
   U137 : OAI22_X1 port map( A1 => A(39), A2 => n540, B1 => B(39), B2 => n541, 
                           ZN => n539);
   U138 : AND2_X1 port map( A1 => n540, A2 => A(39), ZN => n541);
   U139 : INV_X1 port map( A => n536, ZN => n459);
   U140 : OAI22_X1 port map( A1 => A(40), A2 => n460, B1 => B(40), B2 => n537, 
                           ZN => n536);
   U141 : AND2_X1 port map( A1 => n460, A2 => A(40), ZN => n537);
   U142 : XNOR2_X1 port map( A => n437, B => n487, ZN => SUM(57));
   U143 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT58_DW01_add_0 is

   port( A, B : in std_logic_vector (57 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (57 downto 0);  CO : out std_logic);

end RCA_NBIT58_DW01_add_0;

architecture SYN_rpl of RCA_NBIT58_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_24_port, carry_23_port, carry_22_port, carry_21_port, 
      carry_20_port, carry_19_port, carry_18_port, carry_17_port, carry_16_port
      , carry_15_port, carry_14_port, carry_13_port, carry_12_port, 
      carry_11_port, carry_10_port, carry_9_port, carry_8_port, carry_7_port, 
      carry_6_port, carry_5_port, carry_4_port, carry_3_port, carry_2_port, n1,
      n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, 
      n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, 
      n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, 
      n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, 
      n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, 
      n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, 
      n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, 
      n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, 
      n686, n687, n688, n689, n690, n546, n547, n548, n549, n550, n551, n552, 
      n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, 
      n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, 
      n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, 
      n589 : std_logic;

begin
   
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U141 : XOR2_X1 port map( A => n603, B => n604, Z => SUM(53));
   U142 : XOR2_X1 port map( A => B(53), B => A(53), Z => n604);
   U143 : XOR2_X1 port map( A => n608, B => n610, Z => SUM(51));
   U144 : XOR2_X1 port map( A => B(51), B => A(51), Z => n610);
   U145 : XOR2_X1 port map( A => B(50), B => A(50), Z => n613);
   U146 : XOR2_X1 port map( A => n614, B => n616, Z => SUM(49));
   U147 : XOR2_X1 port map( A => B(49), B => A(49), Z => n616);
   U148 : XOR2_X1 port map( A => B(48), B => A(48), Z => n619);
   U149 : XOR2_X1 port map( A => n620, B => n622, Z => SUM(47));
   U150 : XOR2_X1 port map( A => B(47), B => A(47), Z => n622);
   U151 : XOR2_X1 port map( A => B(46), B => A(46), Z => n625);
   U152 : XOR2_X1 port map( A => B(45), B => A(45), Z => n628);
   U153 : XOR2_X1 port map( A => n629, B => n631, Z => SUM(44));
   U154 : XOR2_X1 port map( A => B(44), B => A(44), Z => n631);
   U155 : XOR2_X1 port map( A => n635, B => n637, Z => SUM(42));
   U156 : XOR2_X1 port map( A => B(42), B => A(42), Z => n637);
   U157 : XOR2_X1 port map( A => n641, B => n643, Z => SUM(40));
   U158 : XOR2_X1 port map( A => B(40), B => A(40), Z => n643);
   U159 : XOR2_X1 port map( A => n647, B => n649, Z => SUM(38));
   U160 : XOR2_X1 port map( A => B(38), B => A(38), Z => n649);
   U161 : XOR2_X1 port map( A => A(37), B => B(37), Z => n652);
   U162 : XOR2_X1 port map( A => n653, B => n655, Z => SUM(36));
   U163 : XOR2_X1 port map( A => B(36), B => A(36), Z => n655);
   U164 : XOR2_X1 port map( A => B(35), B => A(35), Z => n658);
   U165 : XOR2_X1 port map( A => n659, B => n661, Z => SUM(34));
   U166 : XOR2_X1 port map( A => B(34), B => A(34), Z => n661);
   U167 : XOR2_X1 port map( A => B(33), B => A(33), Z => n664);
   U168 : XOR2_X1 port map( A => n665, B => n667, Z => SUM(32));
   U169 : XOR2_X1 port map( A => B(32), B => A(32), Z => n667);
   U170 : XOR2_X1 port map( A => B(31), B => A(31), Z => n670);
   U171 : XOR2_X1 port map( A => n671, B => n673, Z => SUM(30));
   U172 : XOR2_X1 port map( A => B(30), B => A(30), Z => n673);
   U173 : XOR2_X1 port map( A => B(29), B => A(29), Z => n676);
   U174 : XOR2_X1 port map( A => n677, B => n679, Z => SUM(28));
   U175 : XOR2_X1 port map( A => B(28), B => A(28), Z => n679);
   U176 : XOR2_X1 port map( A => B(27), B => A(27), Z => n682);
   U177 : XOR2_X1 port map( A => B(26), B => A(26), Z => n685);
   U178 : XOR2_X1 port map( A => B(25), B => A(25), Z => n688);
   U179 : XOR2_X1 port map( A => A(24), B => n690, Z => SUM(24));
   U180 : XOR2_X1 port map( A => carry_24_port, B => B(24), Z => n690);
   U181 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : NOR3_X1 port map( A1 => n601, A2 => A(54), A3 => n549, ZN => n598);
   U2 : OAI21_X1 port map( B1 => n601, B2 => n549, A => A(54), ZN => n599);
   U3 : INV_X1 port map( A => A(41), ZN => n564);
   U4 : INV_X1 port map( A => n592, ZN => n546);
   U5 : INV_X1 port map( A => A(39), ZN => n566);
   U6 : INV_X1 port map( A => A(52), ZN => n550);
   U7 : INV_X1 port map( A => A(43), ZN => n562);
   U8 : AND2_X1 port map( A1 => A(53), A2 => n603, ZN => n601);
   U9 : XNOR2_X1 port map( A => n590, B => n591, ZN => SUM(57));
   U10 : OAI21_X1 port map( B1 => n548, B2 => n592, A => n593, ZN => n591);
   U11 : XNOR2_X1 port map( A => B(57), B => A(57), ZN => n590);
   U12 : INV_X1 port map( A => A(56), ZN => n548);
   U13 : OAI22_X1 port map( A1 => A(26), A2 => n586, B1 => B(26), B2 => n683, 
                           ZN => n680);
   U14 : AND2_X1 port map( A1 => n586, A2 => A(26), ZN => n683);
   U15 : INV_X1 port map( A => n684, ZN => n586);
   U16 : OAI22_X1 port map( A1 => A(25), A2 => n587, B1 => B(25), B2 => n686, 
                           ZN => n684);
   U17 : AND2_X1 port map( A1 => n587, A2 => A(25), ZN => n686);
   U18 : INV_X1 port map( A => n687, ZN => n587);
   U19 : AOI22_X1 port map( A1 => n641, A2 => A(40), B1 => n642, B2 => B(40), 
                           ZN => n638);
   U20 : OR2_X1 port map( A1 => n641, A2 => A(40), ZN => n642);
   U21 : AOI22_X1 port map( A1 => n635, A2 => A(42), B1 => n636, B2 => B(42), 
                           ZN => n632);
   U22 : OR2_X1 port map( A1 => n635, A2 => A(42), ZN => n636);
   U23 : AOI22_X1 port map( A1 => n561, A2 => A(45), B1 => n626, B2 => B(45), 
                           ZN => n623);
   U24 : OR2_X1 port map( A1 => A(45), A2 => n561, ZN => n626);
   U25 : INV_X1 port map( A => n627, ZN => n561);
   U26 : AOI21_X1 port map( B1 => n647, B2 => A(38), A => n568, ZN => n644);
   U27 : INV_X1 port map( A => n648, ZN => n568);
   U28 : OAI21_X1 port map( B1 => A(38), B2 => n647, A => B(38), ZN => n648);
   U29 : XNOR2_X1 port map( A => B(54), B => n600, ZN => SUM(54));
   U30 : NAND2_X1 port map( A1 => n599, A2 => n547, ZN => n600);
   U31 : INV_X1 port map( A => n598, ZN => n547);
   U32 : AOI21_X1 port map( B1 => n653, B2 => A(36), A => n570, ZN => n650);
   U33 : INV_X1 port map( A => n654, ZN => n570);
   U34 : OAI21_X1 port map( B1 => A(36), B2 => n653, A => B(36), ZN => n654);
   U35 : AOI21_X1 port map( B1 => n665, B2 => A(32), A => n576, ZN => n662);
   U36 : INV_X1 port map( A => n666, ZN => n576);
   U37 : OAI21_X1 port map( B1 => A(32), B2 => n665, A => B(32), ZN => n666);
   U38 : AOI21_X1 port map( B1 => n677, B2 => A(28), A => n583, ZN => n674);
   U39 : INV_X1 port map( A => n678, ZN => n583);
   U40 : OAI21_X1 port map( B1 => A(28), B2 => n677, A => B(28), ZN => n678);
   U41 : AOI21_X1 port map( B1 => n671, B2 => A(30), A => n580, ZN => n668);
   U42 : INV_X1 port map( A => n672, ZN => n580);
   U43 : OAI21_X1 port map( B1 => A(30), B2 => n671, A => B(30), ZN => n672);
   U44 : AOI21_X1 port map( B1 => n659, B2 => A(34), A => n573, ZN => n656);
   U45 : INV_X1 port map( A => n660, ZN => n573);
   U46 : OAI21_X1 port map( B1 => A(34), B2 => n659, A => B(34), ZN => n660);
   U47 : AOI21_X1 port map( B1 => n620, B2 => A(47), A => n558, ZN => n617);
   U48 : INV_X1 port map( A => n621, ZN => n558);
   U49 : OAI21_X1 port map( B1 => A(47), B2 => n620, A => B(47), ZN => n621);
   U50 : AOI21_X1 port map( B1 => n608, B2 => A(51), A => n552, ZN => n605);
   U51 : INV_X1 port map( A => n609, ZN => n552);
   U52 : OAI21_X1 port map( B1 => A(51), B2 => n608, A => B(51), ZN => n609);
   U53 : AOI21_X1 port map( B1 => n614, B2 => A(49), A => n555, ZN => n611);
   U54 : INV_X1 port map( A => n615, ZN => n555);
   U55 : OAI21_X1 port map( B1 => A(49), B2 => n614, A => B(49), ZN => n615);
   U56 : AOI22_X1 port map( A1 => n629, A2 => A(44), B1 => n630, B2 => B(44), 
                           ZN => n627);
   U57 : OR2_X1 port map( A1 => n629, A2 => A(44), ZN => n630);
   U58 : XNOR2_X1 port map( A => n656, B => n658, ZN => SUM(35));
   U59 : AOI22_X1 port map( A1 => n595, A2 => A(55), B1 => n596, B2 => B(55), 
                           ZN => n592);
   U60 : OR2_X1 port map( A1 => A(55), A2 => n595, ZN => n596);
   U61 : XNOR2_X1 port map( A => n617, B => n619, ZN => SUM(48));
   U62 : XNOR2_X1 port map( A => n632, B => n634, ZN => SUM(43));
   U63 : XNOR2_X1 port map( A => B(43), B => n562, ZN => n634);
   U64 : XNOR2_X1 port map( A => n597, B => n595, ZN => SUM(55));
   U65 : XNOR2_X1 port map( A => A(55), B => B(55), ZN => n597);
   U66 : XNOR2_X1 port map( A => n627, B => n628, ZN => SUM(45));
   U67 : OAI21_X1 port map( B1 => n598, B2 => n578, A => n599, ZN => n595);
   U68 : INV_X1 port map( A => B(54), ZN => n578);
   U69 : XNOR2_X1 port map( A => n650, B => n652, ZN => SUM(37));
   U70 : XNOR2_X1 port map( A => n594, B => n546, ZN => SUM(56));
   U71 : XNOR2_X1 port map( A => A(56), B => B(56), ZN => n594);
   U72 : XNOR2_X1 port map( A => n644, B => n646, ZN => SUM(39));
   U73 : XNOR2_X1 port map( A => B(39), B => n566, ZN => n646);
   U74 : XNOR2_X1 port map( A => n680, B => n682, ZN => SUM(27));
   U75 : OAI21_X1 port map( B1 => n623, B2 => n559, A => n624, ZN => n620);
   U76 : INV_X1 port map( A => A(46), ZN => n559);
   U77 : OAI21_X1 port map( B1 => A(46), B2 => n560, A => B(46), ZN => n624);
   U78 : INV_X1 port map( A => n623, ZN => n560);
   U79 : OAI21_X1 port map( B1 => n680, B2 => n584, A => n681, ZN => n677);
   U80 : INV_X1 port map( A => A(27), ZN => n584);
   U81 : OAI21_X1 port map( B1 => A(27), B2 => n585, A => B(27), ZN => n681);
   U82 : INV_X1 port map( A => n680, ZN => n585);
   U83 : OAI21_X1 port map( B1 => n650, B2 => n589, A => n651, ZN => n647);
   U84 : INV_X1 port map( A => B(37), ZN => n589);
   U85 : OAI21_X1 port map( B1 => B(37), B2 => n569, A => A(37), ZN => n651);
   U86 : INV_X1 port map( A => n650, ZN => n569);
   U87 : OAI21_X1 port map( B1 => n674, B2 => n581, A => n675, ZN => n671);
   U88 : INV_X1 port map( A => A(29), ZN => n581);
   U89 : OAI21_X1 port map( B1 => A(29), B2 => n582, A => B(29), ZN => n675);
   U90 : INV_X1 port map( A => n674, ZN => n582);
   U91 : OAI21_X1 port map( B1 => n668, B2 => n577, A => n669, ZN => n665);
   U92 : INV_X1 port map( A => A(31), ZN => n577);
   U93 : OAI21_X1 port map( B1 => A(31), B2 => n579, A => B(31), ZN => n669);
   U94 : INV_X1 port map( A => n668, ZN => n579);
   U95 : OAI21_X1 port map( B1 => n662, B2 => n574, A => n663, ZN => n659);
   U96 : INV_X1 port map( A => A(33), ZN => n574);
   U97 : OAI21_X1 port map( B1 => A(33), B2 => n575, A => B(33), ZN => n663);
   U98 : INV_X1 port map( A => n662, ZN => n575);
   U99 : OAI21_X1 port map( B1 => n656, B2 => n571, A => n657, ZN => n653);
   U100 : INV_X1 port map( A => A(35), ZN => n571);
   U101 : OAI21_X1 port map( B1 => A(35), B2 => n572, A => B(35), ZN => n657);
   U102 : INV_X1 port map( A => n656, ZN => n572);
   U103 : OAI21_X1 port map( B1 => n617, B2 => n556, A => n618, ZN => n614);
   U104 : INV_X1 port map( A => A(48), ZN => n556);
   U105 : OAI21_X1 port map( B1 => A(48), B2 => n557, A => B(48), ZN => n618);
   U106 : INV_X1 port map( A => n617, ZN => n557);
   U107 : AOI21_X1 port map( B1 => n564, B2 => n638, A => n639, ZN => n635);
   U108 : AOI21_X1 port map( B1 => n565, B2 => A(41), A => B(41), ZN => n639);
   U109 : INV_X1 port map( A => n638, ZN => n565);
   U110 : AOI21_X1 port map( B1 => n562, B2 => n632, A => n633, ZN => n629);
   U111 : AOI21_X1 port map( B1 => n563, B2 => A(43), A => B(43), ZN => n633);
   U112 : INV_X1 port map( A => n632, ZN => n563);
   U113 : OAI21_X1 port map( B1 => n611, B2 => n553, A => n612, ZN => n608);
   U114 : INV_X1 port map( A => A(50), ZN => n553);
   U115 : OAI21_X1 port map( B1 => A(50), B2 => n554, A => B(50), ZN => n612);
   U116 : INV_X1 port map( A => n611, ZN => n554);
   U117 : AOI21_X1 port map( B1 => n566, B2 => n644, A => n645, ZN => n641);
   U118 : AOI21_X1 port map( B1 => n567, B2 => A(39), A => B(39), ZN => n645);
   U119 : INV_X1 port map( A => n644, ZN => n567);
   U120 : XNOR2_X1 port map( A => n668, B => n670, ZN => SUM(31));
   U121 : XNOR2_X1 port map( A => n662, B => n664, ZN => SUM(33));
   U122 : XNOR2_X1 port map( A => n605, B => n607, ZN => SUM(52));
   U123 : XNOR2_X1 port map( A => B(52), B => n550, ZN => n607);
   U124 : OAI21_X1 port map( B1 => B(24), B2 => A(24), A => n588, ZN => n687);
   U125 : INV_X1 port map( A => n689, ZN => n588);
   U126 : AOI21_X1 port map( B1 => A(24), B2 => B(24), A => carry_24_port, ZN 
                           => n689);
   U127 : XNOR2_X1 port map( A => n638, B => n640, ZN => SUM(41));
   U128 : XNOR2_X1 port map( A => B(41), B => n564, ZN => n640);
   U129 : OAI21_X1 port map( B1 => n605, B2 => n550, A => n606, ZN => n603);
   U130 : OAI21_X1 port map( B1 => A(52), B2 => n551, A => B(52), ZN => n606);
   U131 : INV_X1 port map( A => n605, ZN => n551);
   U132 : XNOR2_X1 port map( A => n611, B => n613, ZN => SUM(50));
   U133 : OAI21_X1 port map( B1 => n546, B2 => A(56), A => B(56), ZN => n593);
   U134 : XNOR2_X1 port map( A => n623, B => n625, ZN => SUM(46));
   U135 : XNOR2_X1 port map( A => n684, B => n685, ZN => SUM(26));
   U136 : XNOR2_X1 port map( A => n674, B => n676, ZN => SUM(29));
   U137 : XNOR2_X1 port map( A => n687, B => n688, ZN => SUM(25));
   U138 : INV_X1 port map( A => n602, ZN => n549);
   U139 : OAI21_X1 port map( B1 => A(53), B2 => n603, A => B(53), ZN => n602);
   U140 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT56_DW01_add_0 is

   port( A, B : in std_logic_vector (55 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (55 downto 0);  CO : out std_logic);

end RCA_NBIT56_DW01_add_0;

architecture SYN_rpl of RCA_NBIT56_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_25_port, carry_22_port, carry_21_port, carry_20_port, 
      carry_19_port, carry_18_port, carry_17_port, carry_16_port, carry_15_port
      , carry_14_port, carry_13_port, carry_12_port, carry_11_port, 
      carry_10_port, carry_9_port, carry_8_port, carry_7_port, carry_6_port, 
      carry_5_port, carry_4_port, carry_3_port, carry_2_port, n1, n523, n524, 
      n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, 
      n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, 
      n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, 
      n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, 
      n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, 
      n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, 
      n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, 
      n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, 
      n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, 
      n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, 
      n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, 
      n519, n520, n521, n522 : std_logic;

begin
   
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => n521, CO => 
                           carry_25_port, S => SUM(24));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U125 : XOR2_X1 port map( A => B(55), B => A(55), Z => n526);
   U126 : XOR2_X1 port map( A => n483, B => n528, Z => SUM(54));
   U127 : XOR2_X1 port map( A => B(54), B => A(54), Z => n528);
   U128 : XOR2_X1 port map( A => n530, B => n532, Z => SUM(53));
   U129 : XOR2_X1 port map( A => B(53), B => A(53), Z => n532);
   U130 : XOR2_X1 port map( A => n485, B => n535, Z => SUM(52));
   U131 : XOR2_X1 port map( A => B(52), B => A(52), Z => n535);
   U132 : XOR2_X1 port map( A => n486, B => n537, Z => SUM(51));
   U133 : XOR2_X1 port map( A => B(51), B => A(51), Z => n537);
   U134 : XOR2_X1 port map( A => n487, B => n540, Z => SUM(50));
   U135 : XOR2_X1 port map( A => B(50), B => A(50), Z => n540);
   U136 : XOR2_X1 port map( A => n517, B => n547, Z => SUM(48));
   U137 : NAND3_X1 port map( A1 => n548, A2 => n489, A3 => A(48), ZN => n546);
   U138 : XOR2_X1 port map( A => n550, B => n551, Z => SUM(47));
   U139 : XOR2_X1 port map( A => B(47), B => A(47), Z => n551);
   U140 : XOR2_X1 port map( A => B(46), B => n555, Z => SUM(46));
   U141 : XOR2_X1 port map( A => n491, B => n558, Z => SUM(45));
   U142 : XOR2_X1 port map( A => B(44), B => A(44), Z => n561);
   U143 : XOR2_X1 port map( A => n565, B => n567, Z => SUM(42));
   U144 : XOR2_X1 port map( A => n575, B => n577, Z => SUM(39));
   U145 : XOR2_X1 port map( A => n581, B => n583, Z => SUM(37));
   U146 : XOR2_X1 port map( A => n584, B => n586, Z => SUM(36));
   U147 : XOR2_X1 port map( A => B(36), B => A(36), Z => n586);
   U148 : XOR2_X1 port map( A => n507, B => n589, Z => SUM(35));
   U149 : XOR2_X1 port map( A => B(35), B => A(35), Z => n589);
   U150 : XOR2_X1 port map( A => n590, B => n592, Z => SUM(34));
   U151 : XOR2_X1 port map( A => B(34), B => A(34), Z => n592);
   U152 : XOR2_X1 port map( A => n509, B => n595, Z => SUM(33));
   U153 : XOR2_X1 port map( A => B(33), B => A(33), Z => n595);
   U154 : XOR2_X1 port map( A => n596, B => n598, Z => SUM(32));
   U155 : XOR2_X1 port map( A => B(32), B => A(32), Z => n598);
   U156 : XOR2_X1 port map( A => n512, B => n601, Z => SUM(31));
   U157 : XOR2_X1 port map( A => B(31), B => A(31), Z => n601);
   U158 : XOR2_X1 port map( A => n602, B => n604, Z => SUM(30));
   U159 : XOR2_X1 port map( A => B(30), B => A(30), Z => n604);
   U160 : XOR2_X1 port map( A => n514, B => n607, Z => SUM(29));
   U161 : XOR2_X1 port map( A => B(29), B => A(29), Z => n607);
   U162 : XOR2_X1 port map( A => n608, B => n610, Z => SUM(28));
   U163 : XOR2_X1 port map( A => B(28), B => A(28), Z => n610);
   U164 : XOR2_X1 port map( A => n518, B => n613, Z => SUM(27));
   U165 : XOR2_X1 port map( A => n519, B => n615, Z => SUM(26));
   U166 : XOR2_X1 port map( A => B(26), B => A(26), Z => n615);
   U167 : XOR2_X1 port map( A => A(25), B => n618, Z => SUM(25));
   U168 : XOR2_X1 port map( A => carry_25_port, B => B(25), Z => n618);
   U169 : XOR2_X1 port map( A => n522, B => n524, Z => SUM(23));
   U170 : XOR2_X1 port map( A => A(23), B => B(23), Z => n524);
   U171 : XOR2_X1 port map( A => carry_22_port, B => n620, Z => SUM(22));
   U172 : XOR2_X1 port map( A => A(22), B => B(22), Z => n620);
   U173 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : AOI21_X1 port map( B1 => n548, B2 => n489, A => A(48), ZN => n545);
   U2 : NOR2_X1 port map( A1 => n554, A2 => A(46), ZN => n553);
   U3 : NOR2_X1 port map( A1 => n498, A2 => n571, ZN => n568);
   U4 : INV_X1 port map( A => A(45), ZN => n490);
   U5 : NAND2_X1 port map( A1 => n571, A2 => n498, ZN => n569);
   U6 : INV_X1 port map( A => A(27), ZN => n516);
   U7 : INV_X1 port map( A => n599, ZN => n512);
   U8 : INV_X1 port map( A => n587, ZN => n507);
   U9 : INV_X1 port map( A => n533, ZN => n485);
   U10 : INV_X1 port map( A => n611, ZN => n518);
   U11 : INV_X1 port map( A => n593, ZN => n509);
   U12 : INV_X1 port map( A => n605, ZN => n514);
   U13 : INV_X1 port map( A => n556, ZN => n491);
   U14 : OR2_X1 port map( A1 => A(47), A2 => n550, ZN => n548);
   U15 : XNOR2_X1 port map( A => n525, B => n526, ZN => SUM(55));
   U16 : OAI22_X1 port map( A1 => n527, A2 => B(54), B1 => n483, B2 => A(54), 
                           ZN => n525);
   U17 : AND2_X1 port map( A1 => A(54), A2 => n483, ZN => n527);
   U18 : AOI21_X1 port map( B1 => A(46), B2 => n554, A => n553, ZN => n555);
   U19 : XNOR2_X1 port map( A => B(27), B => n516, ZN => n613);
   U20 : NAND2_X1 port map( A1 => n546, A2 => n488, ZN => n547);
   U21 : INV_X1 port map( A => n545, ZN => n488);
   U22 : XNOR2_X1 port map( A => B(45), B => n490, ZN => n558);
   U23 : XNOR2_X1 port map( A => A(42), B => B(42), ZN => n567);
   U24 : XNOR2_X1 port map( A => A(39), B => B(39), ZN => n577);
   U25 : OAI22_X1 port map( A1 => A(26), A2 => n519, B1 => B(26), B2 => n614, 
                           ZN => n611);
   U26 : AND2_X1 port map( A1 => n519, A2 => A(26), ZN => n614);
   U27 : OAI21_X1 port map( B1 => B(38), B2 => n578, A => n502, ZN => n575);
   U28 : INV_X1 port map( A => n579, ZN => n502);
   U29 : AOI21_X1 port map( B1 => n578, B2 => B(38), A => A(38), ZN => n579);
   U30 : XNOR2_X1 port map( A => A(37), B => B(37), ZN => n583);
   U31 : AOI21_X1 port map( B1 => n503, B2 => n581, A => n582, ZN => n578);
   U32 : INV_X1 port map( A => A(37), ZN => n503);
   U33 : AOI21_X1 port map( B1 => n504, B2 => A(37), A => B(37), ZN => n582);
   U34 : INV_X1 port map( A => n581, ZN => n504);
   U35 : OAI21_X1 port map( B1 => n575, B2 => n500, A => n576, ZN => n572);
   U36 : INV_X1 port map( A => A(39), ZN => n500);
   U37 : OAI21_X1 port map( B1 => n501, B2 => A(39), A => B(39), ZN => n576);
   U38 : INV_X1 port map( A => n575, ZN => n501);
   U39 : OAI21_X1 port map( B1 => n565, B2 => n495, A => n566, ZN => n562);
   U40 : INV_X1 port map( A => A(42), ZN => n495);
   U41 : OAI21_X1 port map( B1 => A(42), B2 => n496, A => B(42), ZN => n566);
   U42 : INV_X1 port map( A => n565, ZN => n496);
   U43 : OAI21_X1 port map( B1 => n568, B2 => B(41), A => n569, ZN => n565);
   U44 : XNOR2_X1 port map( A => B(41), B => n570, ZN => SUM(41));
   U45 : NAND2_X1 port map( A1 => n497, A2 => n569, ZN => n570);
   U46 : INV_X1 port map( A => n568, ZN => n497);
   U47 : AOI22_X1 port map( A1 => n602, A2 => A(30), B1 => n603, B2 => B(30), 
                           ZN => n599);
   U48 : OR2_X1 port map( A1 => n602, A2 => A(30), ZN => n603);
   U49 : AOI22_X1 port map( A1 => n590, A2 => A(34), B1 => n591, B2 => B(34), 
                           ZN => n587);
   U50 : OR2_X1 port map( A1 => n590, A2 => A(34), ZN => n591);
   U51 : AOI22_X1 port map( A1 => n486, A2 => A(51), B1 => n536, B2 => B(51), 
                           ZN => n533);
   U52 : OR2_X1 port map( A1 => A(51), A2 => n486, ZN => n536);
   U53 : AOI21_X1 port map( B1 => n506, B2 => n587, A => n588, ZN => n584);
   U54 : INV_X1 port map( A => A(35), ZN => n506);
   U55 : AOI21_X1 port map( B1 => n507, B2 => A(35), A => B(35), ZN => n588);
   U56 : AOI21_X1 port map( B1 => n511, B2 => n599, A => n600, ZN => n596);
   U57 : INV_X1 port map( A => A(31), ZN => n511);
   U58 : AOI21_X1 port map( B1 => n512, B2 => A(31), A => B(31), ZN => n600);
   U59 : OAI21_X1 port map( B1 => n556, B2 => n490, A => n557, ZN => n554);
   U60 : OAI21_X1 port map( B1 => A(45), B2 => n491, A => B(45), ZN => n557);
   U61 : OAI21_X1 port map( B1 => n545, B2 => n517, A => n546, ZN => n542);
   U62 : XNOR2_X1 port map( A => n544, B => n542, ZN => SUM(49));
   U63 : XNOR2_X1 port map( A => A(49), B => B(49), ZN => n544);
   U64 : XNOR2_X1 port map( A => n578, B => n580, ZN => SUM(38));
   U65 : XNOR2_X1 port map( A => B(38), B => A(38), ZN => n580);
   U66 : OAI21_X1 port map( B1 => A(36), B2 => n584, A => n505, ZN => n581);
   U67 : INV_X1 port map( A => n585, ZN => n505);
   U68 : AOI21_X1 port map( B1 => n584, B2 => A(36), A => B(36), ZN => n585);
   U69 : OAI21_X1 port map( B1 => n611, B2 => n516, A => n612, ZN => n608);
   U70 : OAI21_X1 port map( B1 => A(27), B2 => n518, A => B(27), ZN => n612);
   U71 : AOI21_X1 port map( B1 => n484, B2 => n533, A => n534, ZN => n530);
   U72 : INV_X1 port map( A => A(52), ZN => n484);
   U73 : AOI21_X1 port map( B1 => n485, B2 => A(52), A => B(52), ZN => n534);
   U74 : AOI21_X1 port map( B1 => n513, B2 => n605, A => n606, ZN => n602);
   U75 : INV_X1 port map( A => A(29), ZN => n513);
   U76 : AOI21_X1 port map( B1 => n514, B2 => A(29), A => B(29), ZN => n606);
   U77 : AOI21_X1 port map( B1 => n508, B2 => n593, A => n594, ZN => n590);
   U78 : INV_X1 port map( A => A(33), ZN => n508);
   U79 : AOI21_X1 port map( B1 => n509, B2 => A(33), A => B(33), ZN => n594);
   U80 : AOI21_X1 port map( B1 => n562, B2 => A(43), A => n494, ZN => n560);
   U81 : INV_X1 port map( A => n563, ZN => n494);
   U82 : OAI21_X1 port map( B1 => A(43), B2 => n562, A => B(43), ZN => n563);
   U83 : XNOR2_X1 port map( A => n574, B => n572, ZN => SUM(40));
   U84 : XNOR2_X1 port map( A => A(40), B => B(40), ZN => n574);
   U85 : AOI22_X1 port map( A1 => B(23), A2 => A(23), B1 => n522, B2 => n524, 
                           ZN => n523);
   U86 : XNOR2_X1 port map( A => n560, B => n561, ZN => SUM(44));
   U87 : AOI21_X1 port map( B1 => n596, B2 => A(32), A => n510, ZN => n593);
   U88 : INV_X1 port map( A => n597, ZN => n510);
   U89 : OAI21_X1 port map( B1 => n596, B2 => A(32), A => B(32), ZN => n597);
   U90 : AOI21_X1 port map( B1 => n608, B2 => A(28), A => n515, ZN => n605);
   U91 : INV_X1 port map( A => n609, ZN => n515);
   U92 : OAI21_X1 port map( B1 => A(28), B2 => n608, A => B(28), ZN => n609);
   U93 : AOI21_X1 port map( B1 => n572, B2 => A(40), A => n499, ZN => n571);
   U94 : INV_X1 port map( A => n573, ZN => n499);
   U95 : OAI21_X1 port map( B1 => A(40), B2 => n572, A => B(40), ZN => n573);
   U96 : AOI21_X1 port map( B1 => n493, B2 => A(44), A => n492, ZN => n556);
   U97 : INV_X1 port map( A => n559, ZN => n492);
   U98 : OAI21_X1 port map( B1 => A(44), B2 => n493, A => B(44), ZN => n559);
   U99 : INV_X1 port map( A => n560, ZN => n493);
   U100 : XNOR2_X1 port map( A => n564, B => n562, ZN => SUM(43));
   U101 : XNOR2_X1 port map( A => A(43), B => B(43), ZN => n564);
   U102 : NOR2_X1 port map( A1 => n552, A2 => n553, ZN => n550);
   U103 : AOI21_X1 port map( B1 => n554, B2 => A(46), A => B(46), ZN => n552);
   U104 : INV_X1 port map( A => n523, ZN => n521);
   U105 : INV_X1 port map( A => n616, ZN => n519);
   U106 : OAI21_X1 port map( B1 => B(25), B2 => A(25), A => n520, ZN => n616);
   U107 : INV_X1 port map( A => n617, ZN => n520);
   U108 : AOI21_X1 port map( B1 => A(25), B2 => B(25), A => carry_25_port, ZN 
                           => n617);
   U109 : INV_X1 port map( A => n541, ZN => n487);
   U110 : AOI22_X1 port map( A1 => n542, A2 => A(49), B1 => n543, B2 => B(49), 
                           ZN => n541);
   U111 : OR2_X1 port map( A1 => A(49), A2 => n542, ZN => n543);
   U112 : INV_X1 port map( A => n529, ZN => n483);
   U113 : AOI22_X1 port map( A1 => n530, A2 => A(53), B1 => n531, B2 => B(53), 
                           ZN => n529);
   U114 : OR2_X1 port map( A1 => n530, A2 => A(53), ZN => n531);
   U115 : INV_X1 port map( A => n538, ZN => n486);
   U116 : AOI22_X1 port map( A1 => n487, A2 => A(50), B1 => n539, B2 => B(50), 
                           ZN => n538);
   U117 : OR2_X1 port map( A1 => A(50), A2 => n487, ZN => n539);
   U118 : INV_X1 port map( A => n549, ZN => n489);
   U119 : AOI21_X1 port map( B1 => n550, B2 => A(47), A => B(47), ZN => n549);
   U120 : INV_X1 port map( A => A(41), ZN => n498);
   U121 : INV_X1 port map( A => n619, ZN => n522);
   U122 : AOI22_X1 port map( A1 => n620, A2 => carry_22_port, B1 => A(22), B2 
                           => B(22), ZN => n619);
   U123 : INV_X1 port map( A => B(48), ZN => n517);
   U124 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT54_DW01_add_0 is

   port( A, B : in std_logic_vector (53 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (53 downto 0);  CO : out std_logic);

end RCA_NBIT54_DW01_add_0;

architecture SYN_rpl of RCA_NBIT54_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_51_port, carry_16_port, carry_15_port, carry_14_port, 
      carry_13_port, carry_12_port, carry_11_port, carry_10_port, carry_9_port,
      carry_8_port, carry_7_port, carry_6_port, carry_5_port, carry_4_port, 
      carry_3_port, carry_2_port, n1, carry_49_port, carry_48_port, 
      carry_47_port, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561
      , n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
      n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, 
      n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, 
      n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, 
      n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, 
      n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, 
      n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, 
      n646, n647, n648, n649, n650, n651, n652, n507, n508, n509, n510, n511, 
      n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, 
      n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, 
      n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, 
      n548, n549, n550, n551 : std_logic;

begin
   
   U1_50 : FA_X1 port map( A => A(50), B => B(50), CI => n509, CO => 
                           carry_51_port, S => SUM(50));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U1_48 : FA_X1 port map( A => B(48), B => carry_48_port, CI => A(48), CO => 
                           carry_49_port, S => SUM(48));
   U1_47 : FA_X1 port map( A => A(47), B => B(47), CI => carry_47_port, CO => 
                           carry_48_port, S => SUM(47));
   U141 : XOR2_X1 port map( A => n556, B => n557, Z => SUM(53));
   U142 : XOR2_X1 port map( A => B(53), B => A(53), Z => n557);
   U143 : XOR2_X1 port map( A => carry_51_port, B => n561, Z => SUM(51));
   U144 : XOR2_X1 port map( A => A(51), B => B(51), Z => n561);
   U145 : XOR2_X1 port map( A => carry_49_port, B => n553, Z => SUM(49));
   U146 : XOR2_X1 port map( A => A(49), B => B(49), Z => n553);
   U147 : XOR2_X1 port map( A => n563, B => n565, Z => SUM(45));
   U148 : XOR2_X1 port map( A => B(45), B => A(45), Z => n565);
   U149 : XOR2_X1 port map( A => B(44), B => A(44), Z => n568);
   U150 : XOR2_X1 port map( A => n569, B => n571, Z => SUM(43));
   U151 : XOR2_X1 port map( A => B(43), B => A(43), Z => n571);
   U152 : XOR2_X1 port map( A => B(42), B => A(42), Z => n574);
   U153 : XOR2_X1 port map( A => n575, B => n577, Z => SUM(41));
   U154 : XOR2_X1 port map( A => B(41), B => A(41), Z => n577);
   U155 : XOR2_X1 port map( A => n585, B => n587, Z => SUM(38));
   U156 : XOR2_X1 port map( A => B(38), B => A(38), Z => n587);
   U157 : XOR2_X1 port map( A => B(37), B => A(37), Z => n590);
   U158 : XOR2_X1 port map( A => n591, B => n593, Z => SUM(36));
   U159 : XOR2_X1 port map( A => B(36), B => A(36), Z => n593);
   U160 : XOR2_X1 port map( A => B(35), B => A(35), Z => n596);
   U161 : XOR2_X1 port map( A => n597, B => n599, Z => SUM(34));
   U162 : XOR2_X1 port map( A => B(34), B => A(34), Z => n599);
   U163 : XOR2_X1 port map( A => B(33), B => A(33), Z => n602);
   U164 : XOR2_X1 port map( A => n603, B => n605, Z => SUM(32));
   U165 : XOR2_X1 port map( A => B(32), B => A(32), Z => n605);
   U166 : XOR2_X1 port map( A => B(31), B => A(31), Z => n608);
   U167 : XOR2_X1 port map( A => n609, B => n611, Z => SUM(30));
   U168 : XOR2_X1 port map( A => B(30), B => A(30), Z => n611);
   U169 : XOR2_X1 port map( A => B(29), B => A(29), Z => n614);
   U170 : XOR2_X1 port map( A => n615, B => n617, Z => SUM(28));
   U171 : XOR2_X1 port map( A => B(28), B => A(28), Z => n617);
   U172 : XOR2_X1 port map( A => B(27), B => A(27), Z => n620);
   U173 : XOR2_X1 port map( A => n621, B => n623, Z => SUM(26));
   U174 : XOR2_X1 port map( A => B(26), B => A(26), Z => n623);
   U175 : XOR2_X1 port map( A => B(24), B => A(24), Z => n629);
   U176 : XOR2_X1 port map( A => n630, B => n632, Z => SUM(23));
   U177 : XOR2_X1 port map( A => B(23), B => A(23), Z => n632);
   U178 : XOR2_X1 port map( A => B(22), B => A(22), Z => n635);
   U179 : XOR2_X1 port map( A => n545, B => n638, Z => SUM(21));
   U180 : XOR2_X1 port map( A => B(18), B => A(18), Z => n647);
   U181 : XOR2_X1 port map( A => B(17), B => A(17), Z => n650);
   U182 : XOR2_X1 port map( A => A(16), B => n652, Z => SUM(16));
   U183 : XOR2_X1 port map( A => carry_16_port, B => B(16), Z => n652);
   U184 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : INV_X1 port map( A => A(52), ZN => n508);
   U2 : NAND2_X1 port map( A1 => A(40), A2 => n580, ZN => n579);
   U3 : INV_X1 port map( A => A(25), ZN => n538);
   U4 : INV_X1 port map( A => A(19), ZN => n547);
   U5 : INV_X1 port map( A => A(39), ZN => n519);
   U6 : INV_X1 port map( A => A(21), ZN => n543);
   U7 : INV_X1 port map( A => A(46), ZN => n510);
   U8 : INV_X1 port map( A => n558, ZN => n507);
   U9 : INV_X1 port map( A => n634, ZN => n542);
   U10 : INV_X1 port map( A => n636, ZN => n545);
   U11 : OAI21_X1 port map( B1 => n558, B2 => n508, A => n559, ZN => n556);
   U12 : OAI21_X1 port map( B1 => A(52), B2 => n507, A => B(52), ZN => n559);
   U13 : AOI22_X1 port map( A1 => n540, A2 => A(24), B1 => n627, B2 => B(24), 
                           ZN => n624);
   U14 : OR2_X1 port map( A1 => A(24), A2 => n540, ZN => n627);
   U15 : INV_X1 port map( A => n628, ZN => n540);
   U16 : AOI22_X1 port map( A1 => n561, A2 => carry_51_port, B1 => A(51), B2 =>
                           B(51), ZN => n558);
   U17 : AOI22_X1 port map( A1 => n621, A2 => A(26), B1 => n622, B2 => B(26), 
                           ZN => n618);
   U18 : OR2_X1 port map( A1 => n621, A2 => A(26), ZN => n622);
   U19 : AOI22_X1 port map( A1 => n615, A2 => A(28), B1 => n616, B2 => B(28), 
                           ZN => n612);
   U20 : OR2_X1 port map( A1 => A(28), A2 => n615, ZN => n616);
   U21 : XNOR2_X1 port map( A => B(40), B => n581, ZN => SUM(40));
   U22 : OAI21_X1 port map( B1 => A(40), B2 => n580, A => n579, ZN => n581);
   U23 : OAI22_X1 port map( A1 => A(18), A2 => n549, B1 => B(18), B2 => n645, 
                           ZN => n642);
   U24 : AND2_X1 port map( A1 => n549, A2 => A(18), ZN => n645);
   U25 : INV_X1 port map( A => n646, ZN => n549);
   U26 : AOI21_X1 port map( B1 => n569, B2 => A(43), A => n515, ZN => n566);
   U27 : INV_X1 port map( A => n570, ZN => n515);
   U28 : OAI21_X1 port map( B1 => A(43), B2 => n569, A => B(43), ZN => n570);
   U29 : AOI21_X1 port map( B1 => n575, B2 => A(41), A => n518, ZN => n572);
   U30 : INV_X1 port map( A => n576, ZN => n518);
   U31 : OAI21_X1 port map( B1 => A(41), B2 => n575, A => B(41), ZN => n576);
   U32 : AOI21_X1 port map( B1 => n609, B2 => A(30), A => n533, ZN => n606);
   U33 : INV_X1 port map( A => n610, ZN => n533);
   U34 : OAI21_X1 port map( B1 => A(30), B2 => n609, A => B(30), ZN => n610);
   U35 : AOI21_X1 port map( B1 => n603, B2 => A(32), A => n530, ZN => n600);
   U36 : INV_X1 port map( A => n604, ZN => n530);
   U37 : OAI21_X1 port map( B1 => A(32), B2 => n603, A => B(32), ZN => n604);
   U38 : AOI21_X1 port map( B1 => n597, B2 => A(34), A => n527, ZN => n594);
   U39 : INV_X1 port map( A => n598, ZN => n527);
   U40 : OAI21_X1 port map( B1 => A(34), B2 => n597, A => B(34), ZN => n598);
   U41 : AOI21_X1 port map( B1 => n563, B2 => A(45), A => n512, ZN => n554);
   U42 : INV_X1 port map( A => n564, ZN => n512);
   U43 : OAI21_X1 port map( B1 => A(45), B2 => n563, A => B(45), ZN => n564);
   U44 : AOI21_X1 port map( B1 => n591, B2 => A(36), A => n524, ZN => n588);
   U45 : INV_X1 port map( A => n592, ZN => n524);
   U46 : OAI21_X1 port map( B1 => A(36), B2 => n591, A => B(36), ZN => n592);
   U47 : AOI21_X1 port map( B1 => n585, B2 => A(38), A => n521, ZN => n582);
   U48 : INV_X1 port map( A => n586, ZN => n521);
   U49 : OAI21_X1 port map( B1 => A(38), B2 => n585, A => B(38), ZN => n586);
   U50 : AOI21_X1 port map( B1 => n547, B2 => n642, A => n643, ZN => n639);
   U51 : AOI21_X1 port map( B1 => n548, B2 => A(19), A => B(19), ZN => n643);
   U52 : INV_X1 port map( A => n642, ZN => n548);
   U53 : AOI22_X1 port map( A1 => n630, A2 => A(23), B1 => n631, B2 => B(23), 
                           ZN => n628);
   U54 : OR2_X1 port map( A1 => A(23), A2 => n630, ZN => n631);
   U55 : XNOR2_X1 port map( A => n588, B => n590, ZN => SUM(37));
   U56 : XNOR2_X1 port map( A => n582, B => n584, ZN => SUM(39));
   U57 : XNOR2_X1 port map( A => B(39), B => n519, ZN => n584);
   U58 : XNOR2_X1 port map( A => n572, B => n574, ZN => SUM(42));
   U59 : XNOR2_X1 port map( A => n554, B => n562, ZN => SUM(46));
   U60 : XNOR2_X1 port map( A => B(46), B => n510, ZN => n562);
   U61 : OAI21_X1 port map( B1 => n582, B2 => n519, A => n583, ZN => n580);
   U62 : OAI21_X1 port map( B1 => A(39), B2 => n520, A => B(39), ZN => n583);
   U63 : INV_X1 port map( A => n582, ZN => n520);
   U64 : XNOR2_X1 port map( A => n558, B => n560, ZN => SUM(52));
   U65 : XNOR2_X1 port map( A => B(52), B => n508, ZN => n560);
   U66 : XNOR2_X1 port map( A => n612, B => n614, ZN => SUM(29));
   U67 : XNOR2_X1 port map( A => n606, B => n608, ZN => SUM(31));
   U68 : XNOR2_X1 port map( A => n600, B => n602, ZN => SUM(33));
   U69 : XNOR2_X1 port map( A => n594, B => n596, ZN => SUM(35));
   U70 : XNOR2_X1 port map( A => n566, B => n568, ZN => SUM(44));
   U71 : OAI22_X1 port map( A1 => A(17), A2 => n550, B1 => B(17), B2 => n648, 
                           ZN => n646);
   U72 : AND2_X1 port map( A1 => n550, A2 => A(17), ZN => n648);
   U73 : INV_X1 port map( A => n649, ZN => n550);
   U74 : XNOR2_X1 port map( A => n624, B => n626, ZN => SUM(25));
   U75 : XNOR2_X1 port map( A => B(25), B => n538, ZN => n626);
   U76 : OAI21_X1 port map( B1 => n612, B2 => n534, A => n613, ZN => n609);
   U77 : INV_X1 port map( A => A(29), ZN => n534);
   U78 : OAI21_X1 port map( B1 => A(29), B2 => n535, A => B(29), ZN => n613);
   U79 : INV_X1 port map( A => n612, ZN => n535);
   U80 : OAI21_X1 port map( B1 => n606, B2 => n531, A => n607, ZN => n603);
   U81 : INV_X1 port map( A => A(31), ZN => n531);
   U82 : OAI21_X1 port map( B1 => A(31), B2 => n532, A => B(31), ZN => n607);
   U83 : INV_X1 port map( A => n606, ZN => n532);
   U84 : OAI21_X1 port map( B1 => n600, B2 => n528, A => n601, ZN => n597);
   U85 : INV_X1 port map( A => A(33), ZN => n528);
   U86 : OAI21_X1 port map( B1 => A(33), B2 => n529, A => B(33), ZN => n601);
   U87 : INV_X1 port map( A => n600, ZN => n529);
   U88 : OAI21_X1 port map( B1 => n594, B2 => n525, A => n595, ZN => n591);
   U89 : INV_X1 port map( A => A(35), ZN => n525);
   U90 : OAI21_X1 port map( B1 => A(35), B2 => n526, A => B(35), ZN => n595);
   U91 : INV_X1 port map( A => n594, ZN => n526);
   U92 : OAI21_X1 port map( B1 => n588, B2 => n522, A => n589, ZN => n585);
   U93 : INV_X1 port map( A => A(37), ZN => n522);
   U94 : OAI21_X1 port map( B1 => A(37), B2 => n523, A => B(37), ZN => n589);
   U95 : INV_X1 port map( A => n588, ZN => n523);
   U96 : OAI21_X1 port map( B1 => n572, B2 => n516, A => n573, ZN => n569);
   U97 : INV_X1 port map( A => A(42), ZN => n516);
   U98 : OAI21_X1 port map( B1 => A(42), B2 => n517, A => B(42), ZN => n573);
   U99 : INV_X1 port map( A => n572, ZN => n517);
   U100 : OAI21_X1 port map( B1 => n566, B2 => n513, A => n567, ZN => n563);
   U101 : INV_X1 port map( A => A(44), ZN => n513);
   U102 : OAI21_X1 port map( B1 => A(44), B2 => n514, A => B(44), ZN => n567);
   U103 : INV_X1 port map( A => n566, ZN => n514);
   U104 : OAI21_X1 port map( B1 => n578, B2 => n544, A => n579, ZN => n575);
   U105 : NOR2_X1 port map( A1 => A(40), A2 => n580, ZN => n578);
   U106 : INV_X1 port map( A => B(40), ZN => n544);
   U107 : AOI21_X1 port map( B1 => n538, B2 => n624, A => n625, ZN => n621);
   U108 : AOI21_X1 port map( B1 => n539, B2 => A(25), A => B(25), ZN => n625);
   U109 : INV_X1 port map( A => n624, ZN => n539);
   U110 : AOI22_X1 port map( A1 => B(49), A2 => A(49), B1 => n553, B2 => 
                           carry_49_port, ZN => n552);
   U111 : OAI21_X1 port map( B1 => B(16), B2 => A(16), A => n551, ZN => n649);
   U112 : INV_X1 port map( A => n651, ZN => n551);
   U113 : AOI21_X1 port map( B1 => A(16), B2 => B(16), A => carry_16_port, ZN 
                           => n651);
   U114 : OAI21_X1 port map( B1 => n618, B2 => n536, A => n619, ZN => n615);
   U115 : INV_X1 port map( A => A(27), ZN => n536);
   U116 : OAI21_X1 port map( B1 => A(27), B2 => n537, A => B(27), ZN => n619);
   U117 : INV_X1 port map( A => n618, ZN => n537);
   U118 : OAI21_X1 port map( B1 => n542, B2 => n541, A => n633, ZN => n630);
   U119 : INV_X1 port map( A => A(22), ZN => n541);
   U120 : OAI21_X1 port map( B1 => A(22), B2 => n634, A => B(22), ZN => n633);
   U121 : XNOR2_X1 port map( A => B(21), B => n543, ZN => n638);
   U122 : XNOR2_X1 port map( A => n618, B => n620, ZN => SUM(27));
   U123 : OAI21_X1 port map( B1 => A(46), B2 => n511, A => B(46), ZN => n555);
   U124 : INV_X1 port map( A => n554, ZN => n511);
   U125 : OAI21_X1 port map( B1 => n636, B2 => n543, A => n637, ZN => n634);
   U126 : OAI21_X1 port map( B1 => A(21), B2 => n545, A => B(21), ZN => n637);
   U127 : AOI21_X1 port map( B1 => n639, B2 => A(20), A => n546, ZN => n636);
   U128 : INV_X1 port map( A => n640, ZN => n546);
   U129 : OAI21_X1 port map( B1 => n639, B2 => A(20), A => B(20), ZN => n640);
   U130 : XNOR2_X1 port map( A => n542, B => n635, ZN => SUM(22));
   U131 : INV_X1 port map( A => n552, ZN => n509);
   U132 : XNOR2_X1 port map( A => n628, B => n629, ZN => SUM(24));
   U133 : OAI21_X1 port map( B1 => n554, B2 => n510, A => n555, ZN => 
                           carry_47_port);
   U134 : XNOR2_X1 port map( A => n649, B => n650, ZN => SUM(17));
   U135 : XNOR2_X1 port map( A => n646, B => n647, ZN => SUM(18));
   U136 : XNOR2_X1 port map( A => n642, B => n644, ZN => SUM(19));
   U137 : XNOR2_X1 port map( A => B(19), B => n547, ZN => n644);
   U138 : XNOR2_X1 port map( A => n639, B => n641, ZN => SUM(20));
   U139 : XNOR2_X1 port map( A => A(20), B => B(20), ZN => n641);
   U140 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT52_DW01_add_0 is

   port( A, B : in std_logic_vector (51 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (51 downto 0);  CO : out std_logic);

end RCA_NBIT52_DW01_add_0;

architecture SYN_rpl of RCA_NBIT52_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_18_port, carry_17_port, carry_16_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_10_port
      , carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, n1, n542, n543, n544, n545, 
      n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, 
      n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, 
      n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, 
      n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, 
      n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, 
      n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, 
      n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, 
      n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, 
      n642, n643, n644, n497, n498, n499, n500, n501, n502, n503, n504, n505, 
      n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, 
      n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, 
      n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541 : 
      std_logic;

begin
   
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U134 : XOR2_X1 port map( A => n542, B => n543, Z => SUM(51));
   U135 : XOR2_X1 port map( A => n546, B => n545, Z => SUM(50));
   U136 : XOR2_X1 port map( A => n547, B => n498, Z => SUM(49));
   U137 : XOR2_X1 port map( A => A(49), B => B(49), Z => n547);
   U138 : XOR2_X1 port map( A => n552, B => n554, Z => SUM(47));
   U139 : XOR2_X1 port map( A => n558, B => n560, Z => SUM(45));
   U140 : XOR2_X1 port map( A => n564, B => n566, Z => SUM(43));
   U141 : XOR2_X1 port map( A => n570, B => n571, Z => SUM(42));
   U142 : XOR2_X1 port map( A => B(42), B => A(42), Z => n571);
   U143 : XOR2_X1 port map( A => n572, B => n573, Z => SUM(41));
   U144 : XOR2_X1 port map( A => B(41), B => A(41), Z => n573);
   U145 : XOR2_X1 port map( A => n579, B => n580, Z => SUM(40));
   U146 : XOR2_X1 port map( A => B(40), B => A(40), Z => n580);
   U147 : XOR2_X1 port map( A => n577, B => n581, Z => SUM(39));
   U148 : XOR2_X1 port map( A => B(39), B => A(39), Z => n581);
   U149 : XOR2_X1 port map( A => n512, B => n584, Z => SUM(38));
   U150 : XOR2_X1 port map( A => B(38), B => A(38), Z => n584);
   U151 : XOR2_X1 port map( A => n513, B => n586, Z => SUM(37));
   U152 : XOR2_X1 port map( A => B(37), B => A(37), Z => n586);
   U153 : XOR2_X1 port map( A => n588, B => n590, Z => SUM(36));
   U154 : XOR2_X1 port map( A => B(36), B => A(36), Z => n590);
   U155 : XOR2_X1 port map( A => n515, B => n593, Z => SUM(35));
   U156 : XOR2_X1 port map( A => B(35), B => A(35), Z => n593);
   U157 : XOR2_X1 port map( A => n594, B => n596, Z => SUM(34));
   U158 : XOR2_X1 port map( A => B(34), B => A(34), Z => n596);
   U159 : XOR2_X1 port map( A => n518, B => n599, Z => SUM(33));
   U160 : XOR2_X1 port map( A => B(33), B => A(33), Z => n599);
   U161 : XOR2_X1 port map( A => n600, B => n602, Z => SUM(32));
   U162 : XOR2_X1 port map( A => B(32), B => A(32), Z => n602);
   U163 : XOR2_X1 port map( A => n521, B => n605, Z => SUM(31));
   U164 : XOR2_X1 port map( A => n606, B => n608, Z => SUM(30));
   U165 : XOR2_X1 port map( A => B(30), B => A(30), Z => n608);
   U166 : XOR2_X1 port map( A => n541, B => n611, Z => SUM(29));
   U167 : XOR2_X1 port map( A => n526, B => n615, Z => SUM(28));
   U168 : XOR2_X1 port map( A => B(28), B => A(28), Z => n615);
   U169 : XOR2_X1 port map( A => n616, B => n618, Z => SUM(27));
   U170 : XOR2_X1 port map( A => B(27), B => A(27), Z => n618);
   U171 : XOR2_X1 port map( A => n528, B => n621, Z => SUM(26));
   U172 : XOR2_X1 port map( A => B(26), B => A(26), Z => n621);
   U173 : XOR2_X1 port map( A => n622, B => n624, Z => SUM(25));
   U174 : XOR2_X1 port map( A => B(25), B => A(25), Z => n624);
   U175 : XOR2_X1 port map( A => n626, B => n627, Z => SUM(24));
   U176 : XOR2_X1 port map( A => n533, B => n630, Z => SUM(23));
   U177 : XOR2_X1 port map( A => n631, B => n633, Z => SUM(22));
   U178 : XOR2_X1 port map( A => B(22), B => A(22), Z => n633);
   U179 : XOR2_X1 port map( A => n536, B => n636, Z => SUM(21));
   U180 : XOR2_X1 port map( A => n539, B => n642, Z => SUM(19));
   U181 : XOR2_X1 port map( A => B(19), B => A(19), Z => n642);
   U182 : XOR2_X1 port map( A => A(18), B => n644, Z => SUM(18));
   U183 : XOR2_X1 port map( A => carry_18_port, B => B(18), Z => n644);
   U184 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : INV_X1 port map( A => n578, ZN => n510);
   U2 : NOR2_X1 port map( A1 => A(29), A2 => n612, ZN => n609);
   U3 : NAND2_X1 port map( A1 => A(39), A2 => n577, ZN => n578);
   U4 : NAND2_X1 port map( A1 => A(20), A2 => n637, ZN => n638);
   U5 : NAND2_X1 port map( A1 => A(41), A2 => n572, ZN => n568);
   U6 : INV_X1 port map( A => A(31), ZN => n520);
   U7 : INV_X1 port map( A => A(24), ZN => n530);
   U8 : INV_X1 port map( A => n545, ZN => n497);
   U9 : NAND2_X1 port map( A1 => A(29), A2 => n612, ZN => n610);
   U10 : INV_X1 port map( A => A(23), ZN => n532);
   U11 : INV_X1 port map( A => A(21), ZN => n535);
   U12 : INV_X1 port map( A => n619, ZN => n528);
   U13 : INV_X1 port map( A => n613, ZN => n526);
   U14 : INV_X1 port map( A => n582, ZN => n512);
   U15 : INV_X1 port map( A => n634, ZN => n536);
   U16 : INV_X1 port map( A => n628, ZN => n533);
   U17 : INV_X1 port map( A => n591, ZN => n515);
   U18 : INV_X1 port map( A => n640, ZN => n539);
   U19 : OR2_X1 port map( A1 => n497, A2 => A(50), ZN => n544);
   U20 : INV_X1 port map( A => n576, ZN => n509);
   U21 : INV_X1 port map( A => n603, ZN => n521);
   U22 : INV_X1 port map( A => n597, ZN => n518);
   U23 : XNOR2_X1 port map( A => B(51), B => A(51), ZN => n542);
   U24 : AOI22_X1 port map( A1 => B(50), A2 => n544, B1 => A(50), B2 => n497, 
                           ZN => n543);
   U25 : NAND2_X1 port map( A1 => n576, A2 => n578, ZN => n579);
   U26 : XNOR2_X1 port map( A => A(43), B => B(43), ZN => n566);
   U27 : XNOR2_X1 port map( A => B(45), B => A(45), ZN => n560);
   U28 : XNOR2_X1 port map( A => B(31), B => n520, ZN => n605);
   U29 : NAND2_X1 port map( A1 => n569, A2 => n568, ZN => n570);
   U30 : NAND2_X1 port map( A1 => n523, A2 => n610, ZN => n611);
   U31 : INV_X1 port map( A => n609, ZN => n523);
   U32 : XNOR2_X1 port map( A => B(24), B => n530, ZN => n627);
   U33 : XNOR2_X1 port map( A => B(23), B => n532, ZN => n630);
   U34 : OAI22_X1 port map( A1 => A(20), A2 => n637, B1 => B(20), B2 => n537, 
                           ZN => n634);
   U35 : INV_X1 port map( A => n638, ZN => n537);
   U36 : XNOR2_X1 port map( A => B(21), B => n535, ZN => n636);
   U37 : XNOR2_X1 port map( A => B(20), B => n639, ZN => SUM(20));
   U38 : OAI21_X1 port map( B1 => A(20), B2 => n637, A => n638, ZN => n639);
   U39 : AOI21_X1 port map( B1 => n511, B2 => n582, A => n583, ZN => n577);
   U40 : INV_X1 port map( A => A(38), ZN => n511);
   U41 : AOI21_X1 port map( B1 => n512, B2 => A(38), A => B(38), ZN => n583);
   U42 : OAI21_X1 port map( B1 => B(42), B2 => A(42), A => n567, ZN => n564);
   U43 : OAI211_X1 port map( C1 => n507, C2 => n529, A => n568, B => n569, ZN 
                           => n567);
   U44 : INV_X1 port map( A => A(42), ZN => n507);
   U45 : INV_X1 port map( A => B(42), ZN => n529);
   U46 : AOI21_X1 port map( B1 => n500, B2 => n552, A => n553, ZN => n549);
   U47 : INV_X1 port map( A => A(47), ZN => n500);
   U48 : AOI21_X1 port map( B1 => n501, B2 => A(47), A => B(47), ZN => n553);
   U49 : INV_X1 port map( A => n552, ZN => n501);
   U50 : AOI21_X1 port map( B1 => n538, B2 => n640, A => n641, ZN => n637);
   U51 : INV_X1 port map( A => A(19), ZN => n538);
   U52 : AOI21_X1 port map( B1 => n539, B2 => A(19), A => B(19), ZN => n641);
   U53 : OAI21_X1 port map( B1 => n564, B2 => n505, A => n565, ZN => n561);
   U54 : INV_X1 port map( A => A(43), ZN => n505);
   U55 : OAI21_X1 port map( B1 => n506, B2 => A(43), A => B(43), ZN => n565);
   U56 : INV_X1 port map( A => n564, ZN => n506);
   U57 : OAI21_X1 port map( B1 => n558, B2 => n525, A => n559, ZN => n555);
   U58 : INV_X1 port map( A => B(45), ZN => n525);
   U59 : OAI21_X1 port map( B1 => n503, B2 => B(45), A => A(45), ZN => n559);
   U60 : INV_X1 port map( A => n558, ZN => n503);
   U61 : AOI22_X1 port map( A1 => n622, A2 => A(25), B1 => n623, B2 => B(25), 
                           ZN => n619);
   U62 : OR2_X1 port map( A1 => A(25), A2 => n622, ZN => n623);
   U63 : AOI22_X1 port map( A1 => n616, A2 => A(27), B1 => n617, B2 => B(27), 
                           ZN => n613);
   U64 : OR2_X1 port map( A1 => n616, A2 => A(27), ZN => n617);
   U65 : AOI22_X1 port map( A1 => n513, A2 => A(37), B1 => n585, B2 => B(37), 
                           ZN => n582);
   U66 : OR2_X1 port map( A1 => A(37), A2 => n513, ZN => n585);
   U67 : AOI21_X1 port map( B1 => n508, B2 => n574, A => n575, ZN => n572);
   U68 : INV_X1 port map( A => A(40), ZN => n508);
   U69 : NOR3_X1 port map( A1 => n509, A2 => B(40), A3 => n510, ZN => n575);
   U70 : OAI221_X1 port map( B1 => n510, B2 => B(39), C1 => n577, C2 => A(39), 
                           A => B(40), ZN => n574);
   U71 : AOI22_X1 port map( A1 => B(49), A2 => A(49), B1 => n498, B2 => n547, 
                           ZN => n545);
   U72 : XNOR2_X1 port map( A => n563, B => n561, ZN => SUM(44));
   U73 : XNOR2_X1 port map( A => A(44), B => B(44), ZN => n563);
   U74 : OAI21_X1 port map( B1 => A(46), B2 => n555, A => n502, ZN => n552);
   U75 : INV_X1 port map( A => n556, ZN => n502);
   U76 : AOI21_X1 port map( B1 => n555, B2 => A(46), A => B(46), ZN => n556);
   U77 : OAI21_X1 port map( B1 => n628, B2 => n532, A => n629, ZN => n626);
   U78 : OAI21_X1 port map( B1 => n533, B2 => A(23), A => B(23), ZN => n629);
   U79 : OAI21_X1 port map( B1 => n634, B2 => n535, A => n635, ZN => n631);
   U80 : OAI21_X1 port map( B1 => n536, B2 => A(21), A => B(21), ZN => n635);
   U81 : OAI21_X1 port map( B1 => A(44), B2 => n561, A => n504, ZN => n558);
   U82 : INV_X1 port map( A => n562, ZN => n504);
   U83 : AOI21_X1 port map( B1 => n561, B2 => A(44), A => B(44), ZN => n562);
   U84 : OAI21_X1 port map( B1 => n609, B2 => n541, A => n610, ZN => n606);
   U85 : OAI21_X1 port map( B1 => n597, B2 => n517, A => n598, ZN => n594);
   U86 : INV_X1 port map( A => A(33), ZN => n517);
   U87 : OAI21_X1 port map( B1 => n518, B2 => A(33), A => B(33), ZN => n598);
   U88 : OAI21_X1 port map( B1 => n603, B2 => n520, A => n604, ZN => n600);
   U89 : OAI21_X1 port map( B1 => n521, B2 => A(31), A => B(31), ZN => n604);
   U90 : AOI21_X1 port map( B1 => n527, B2 => n619, A => n620, ZN => n616);
   U91 : INV_X1 port map( A => A(26), ZN => n527);
   U92 : AOI21_X1 port map( B1 => n528, B2 => A(26), A => B(26), ZN => n620);
   U93 : OAI21_X1 port map( B1 => n577, B2 => A(39), A => B(39), ZN => n576);
   U94 : AOI21_X1 port map( B1 => A(18), B2 => B(18), A => n540, ZN => n640);
   U95 : INV_X1 port map( A => n643, ZN => n540);
   U96 : OAI21_X1 port map( B1 => A(18), B2 => B(18), A => carry_18_port, ZN =>
                           n643);
   U97 : AOI21_X1 port map( B1 => n524, B2 => n613, A => n614, ZN => n612);
   U98 : INV_X1 port map( A => A(28), ZN => n524);
   U99 : AOI21_X1 port map( B1 => n526, B2 => A(28), A => B(28), ZN => n614);
   U100 : OAI21_X1 port map( B1 => A(41), B2 => n572, A => B(41), ZN => n569);
   U101 : OAI21_X1 port map( B1 => n591, B2 => n514, A => n592, ZN => n588);
   U102 : INV_X1 port map( A => A(35), ZN => n514);
   U103 : OAI21_X1 port map( B1 => n515, B2 => A(35), A => B(35), ZN => n592);
   U104 : OAI21_X1 port map( B1 => n531, B2 => n530, A => n625, ZN => n622);
   U105 : INV_X1 port map( A => n626, ZN => n531);
   U106 : OAI21_X1 port map( B1 => A(24), B2 => n626, A => B(24), ZN => n625);
   U107 : OAI21_X1 port map( B1 => A(34), B2 => n594, A => n516, ZN => n591);
   U108 : INV_X1 port map( A => n595, ZN => n516);
   U109 : AOI21_X1 port map( B1 => n594, B2 => A(34), A => B(34), ZN => n595);
   U110 : XNOR2_X1 port map( A => n557, B => n555, ZN => SUM(46));
   U111 : XNOR2_X1 port map( A => A(46), B => B(46), ZN => n557);
   U112 : OAI21_X1 port map( B1 => A(22), B2 => n631, A => n534, ZN => n628);
   U113 : INV_X1 port map( A => n632, ZN => n534);
   U114 : AOI21_X1 port map( B1 => n631, B2 => A(22), A => B(22), ZN => n632);
   U115 : OAI21_X1 port map( B1 => A(32), B2 => n600, A => n519, ZN => n597);
   U116 : INV_X1 port map( A => n601, ZN => n519);
   U117 : AOI21_X1 port map( B1 => n600, B2 => A(32), A => B(32), ZN => n601);
   U118 : XNOR2_X1 port map( A => A(47), B => B(47), ZN => n554);
   U119 : OAI21_X1 port map( B1 => A(30), B2 => n606, A => n522, ZN => n603);
   U120 : INV_X1 port map( A => n607, ZN => n522);
   U121 : AOI21_X1 port map( B1 => n606, B2 => A(30), A => B(30), ZN => n607);
   U122 : XNOR2_X1 port map( A => A(50), B => B(50), ZN => n546);
   U123 : XNOR2_X1 port map( A => n549, B => n551, ZN => SUM(48));
   U124 : XNOR2_X1 port map( A => A(48), B => B(48), ZN => n551);
   U125 : INV_X1 port map( A => n587, ZN => n513);
   U126 : AOI22_X1 port map( A1 => n588, A2 => A(36), B1 => n589, B2 => B(36), 
                           ZN => n587);
   U127 : OR2_X1 port map( A1 => A(36), A2 => n588, ZN => n589);
   U128 : INV_X1 port map( A => n548, ZN => n498);
   U129 : AOI21_X1 port map( B1 => n549, B2 => A(48), A => n499, ZN => n548);
   U130 : INV_X1 port map( A => n550, ZN => n499);
   U131 : OAI21_X1 port map( B1 => n549, B2 => A(48), A => B(48), ZN => n550);
   U132 : INV_X1 port map( A => B(29), ZN => n541);
   U133 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT50_DW01_add_0 is

   port( A, B : in std_logic_vector (49 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (49 downto 0);  CO : out std_logic);

end RCA_NBIT50_DW01_add_0;

architecture SYN_rpl of RCA_NBIT50_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_15_port, carry_14_port, carry_13_port, carry_12_port, 
      carry_11_port, carry_10_port, carry_9_port, carry_8_port, carry_7_port, 
      carry_6_port, carry_5_port, carry_4_port, carry_3_port, carry_2_port, n1,
      carry_44_port, carry_16_port, carry_43_port, carry_42_port, net76696, 
      n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, 
      n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, 
      n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, 
      n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, 
      n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, 
      n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, 
      n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, 
      n550, n551, n552, n553, n554, n555, n426, n427, n428, n429, n430, n431, 
      n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, 
      n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, 
      n456, n457, n458, n459, n460, n461, n462, n463, n464, n465 : std_logic;

begin
   
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_44 : FA_X1 port map( A => A(44), B => B(44), CI => carry_44_port, CO => 
                           net76696, S => SUM(44));
   U1_41 : FA_X1 port map( A => B(41), B => A(41), CI => n430, CO => 
                           carry_42_port, S => SUM(41));
   U1_43 : FA_X1 port map( A => A(43), B => B(43), CI => carry_43_port, CO => 
                           carry_44_port, S => SUM(43));
   U1_42 : FA_X1 port map( A => A(42), B => B(42), CI => carry_42_port, CO => 
                           carry_43_port, S => SUM(42));
   U129 : XOR2_X1 port map( A => n469, B => n470, Z => SUM(49));
   U130 : XOR2_X1 port map( A => B(46), B => A(46), Z => n479);
   U131 : XOR2_X1 port map( A => A(45), B => n481, Z => SUM(45));
   U132 : XOR2_X1 port map( A => net76696, B => B(45), Z => n481);
   U133 : XOR2_X1 port map( A => n467, B => n482, Z => SUM(40));
   U134 : XOR2_X1 port map( A => B(40), B => A(40), Z => n482);
   U135 : XOR2_X1 port map( A => n433, B => n485, Z => SUM(39));
   U136 : XOR2_X1 port map( A => B(39), B => A(39), Z => n485);
   U137 : XOR2_X1 port map( A => n435, B => B(37), Z => n491);
   U138 : XOR2_X1 port map( A => n493, B => n494, Z => SUM(36));
   U139 : XOR2_X1 port map( A => B(36), B => A(36), Z => n494);
   U140 : XOR2_X1 port map( A => B(35), B => A(35), Z => n497);
   U141 : XOR2_X1 port map( A => B(34), B => n500, Z => SUM(34));
   U142 : XOR2_X1 port map( A => B(33), B => A(33), Z => n504);
   U143 : XOR2_X1 port map( A => B(32), B => A(32), Z => n507);
   U144 : XOR2_X1 port map( A => n510, B => n511, Z => SUM(31));
   U145 : XOR2_X1 port map( A => n518, B => n520, Z => SUM(28));
   U146 : XOR2_X1 port map( A => B(28), B => A(28), Z => n520);
   U147 : XOR2_X1 port map( A => n524, B => n526, Z => SUM(26));
   U148 : XOR2_X1 port map( A => B(26), B => A(26), Z => n526);
   U149 : XOR2_X1 port map( A => n527, B => n529, Z => SUM(25));
   U150 : XOR2_X1 port map( A => n451, B => B(25), Z => n529);
   U151 : XOR2_X1 port map( A => n530, B => n532, Z => SUM(24));
   U152 : XOR2_X1 port map( A => B(24), B => A(24), Z => n532);
   U153 : XOR2_X1 port map( A => B(23), B => A(23), Z => n535);
   U154 : XOR2_X1 port map( A => n536, B => n538, Z => SUM(22));
   U155 : XOR2_X1 port map( A => B(22), B => A(22), Z => n538);
   U156 : XOR2_X1 port map( A => n542, B => n544, Z => SUM(20));
   U157 : XOR2_X1 port map( A => B(20), B => A(20), Z => n544);
   U158 : XOR2_X1 port map( A => n548, B => n550, Z => SUM(18));
   U159 : XOR2_X1 port map( A => B(18), B => A(18), Z => n550);
   U160 : XOR2_X1 port map( A => A(16), B => n555, Z => SUM(16));
   U161 : XOR2_X1 port map( A => carry_16_port, B => B(16), Z => n555);
   U162 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : NOR2_X1 port map( A1 => A(34), A2 => n440, ZN => n499);
   U2 : INV_X1 port map( A => n489, ZN => n436);
   U3 : INV_X1 port map( A => A(17), ZN => n463);
   U4 : INV_X1 port map( A => n545, ZN => n461);
   U5 : INV_X1 port map( A => n539, ZN => n458);
   U6 : INV_X1 port map( A => n521, ZN => n449);
   U7 : INV_X1 port map( A => A(25), ZN => n451);
   U8 : INV_X1 port map( A => A(37), ZN => n435);
   U9 : INV_X1 port map( A => n515, ZN => n446);
   U10 : OR2_X1 port map( A1 => A(30), A2 => n512, ZN => n509);
   U11 : INV_X1 port map( A => n483, ZN => n433);
   U12 : AND2_X1 port map( A1 => n426, A2 => A(48), ZN => n471);
   U13 : XNOR2_X1 port map( A => B(49), B => A(49), ZN => n470);
   U14 : OAI22_X1 port map( A1 => A(48), A2 => n426, B1 => B(48), B2 => n471, 
                           ZN => n469);
   U15 : AOI21_X1 port map( B1 => A(34), B2 => n440, A => n499, ZN => n500);
   U16 : NAND2_X1 port map( A1 => n444, A2 => n509, ZN => n510);
   U17 : XNOR2_X1 port map( A => A(31), B => B(31), ZN => n511);
   U18 : OAI22_X1 port map( A1 => A(32), A2 => n442, B1 => B(32), B2 => n505, 
                           ZN => n503);
   U19 : AND2_X1 port map( A1 => n442, A2 => A(32), ZN => n505);
   U20 : INV_X1 port map( A => n506, ZN => n442);
   U21 : AOI21_X1 port map( B1 => A(31), B2 => B(31), A => n443, ZN => n506);
   U22 : INV_X1 port map( A => n508, ZN => n443);
   U23 : OAI211_X1 port map( C1 => A(31), C2 => B(31), A => n509, B => n444, ZN
                           => n508);
   U24 : AOI21_X1 port map( B1 => A(16), B2 => B(16), A => n465, ZN => n551);
   U25 : INV_X1 port map( A => n554, ZN => n465);
   U26 : OAI21_X1 port map( B1 => A(16), B2 => B(16), A => carry_16_port, ZN =>
                           n554);
   U27 : OAI21_X1 port map( B1 => n498, B2 => B(34), A => n439, ZN => n495);
   U28 : INV_X1 port map( A => n499, ZN => n439);
   U29 : AND2_X1 port map( A1 => n440, A2 => A(34), ZN => n498);
   U30 : OAI22_X1 port map( A1 => n492, A2 => B(36), B1 => A(36), B2 => n493, 
                           ZN => n489);
   U31 : AND2_X1 port map( A1 => n493, A2 => A(36), ZN => n492);
   U32 : OAI21_X1 port map( B1 => n489, B2 => n435, A => n490, ZN => n486);
   U33 : OAI21_X1 port map( B1 => n436, B2 => A(37), A => B(37), ZN => n490);
   U34 : XNOR2_X1 port map( A => n426, B => n472, ZN => SUM(48));
   U35 : XNOR2_X1 port map( A => A(48), B => B(48), ZN => n472);
   U36 : XNOR2_X1 port map( A => n427, B => n475, ZN => SUM(47));
   U37 : XNOR2_X1 port map( A => A(47), B => B(47), ZN => n475);
   U38 : XNOR2_X1 port map( A => n478, B => n479, ZN => SUM(46));
   U39 : OAI21_X1 port map( B1 => A(22), B2 => n536, A => n456, ZN => n533);
   U40 : INV_X1 port map( A => n537, ZN => n456);
   U41 : AOI21_X1 port map( B1 => n536, B2 => A(22), A => B(22), ZN => n537);
   U42 : AOI21_X1 port map( B1 => n445, B2 => n515, A => n516, ZN => n512);
   U43 : INV_X1 port map( A => A(29), ZN => n445);
   U44 : AOI21_X1 port map( B1 => n446, B2 => A(29), A => B(29), ZN => n516);
   U45 : AOI21_X1 port map( B1 => n463, B2 => n551, A => n552, ZN => n548);
   U46 : AOI21_X1 port map( B1 => n464, B2 => A(17), A => B(17), ZN => n552);
   U47 : INV_X1 port map( A => n551, ZN => n464);
   U48 : OAI21_X1 port map( B1 => A(45), B2 => B(45), A => n429, ZN => n478);
   U49 : INV_X1 port map( A => n480, ZN => n429);
   U50 : AOI21_X1 port map( B1 => A(45), B2 => B(45), A => net76696, ZN => n480
                           );
   U51 : XNOR2_X1 port map( A => n488, B => n486, ZN => SUM(38));
   U52 : XNOR2_X1 port map( A => A(38), B => B(38), ZN => n488);
   U53 : XNOR2_X1 port map( A => n495, B => n497, ZN => SUM(35));
   U54 : XNOR2_X1 port map( A => n461, B => n547, ZN => SUM(19));
   U55 : XNOR2_X1 port map( A => A(19), B => B(19), ZN => n547);
   U56 : XNOR2_X1 port map( A => n506, B => n507, ZN => SUM(32));
   U57 : XNOR2_X1 port map( A => n503, B => n504, ZN => SUM(33));
   U58 : XNOR2_X1 port map( A => n512, B => n514, ZN => SUM(30));
   U59 : XNOR2_X1 port map( A => A(30), B => B(30), ZN => n514);
   U60 : OAI21_X1 port map( B1 => n533, B2 => n454, A => n534, ZN => n530);
   U61 : INV_X1 port map( A => A(23), ZN => n454);
   U62 : OAI21_X1 port map( B1 => n455, B2 => A(23), A => B(23), ZN => n534);
   U63 : INV_X1 port map( A => n533, ZN => n455);
   U64 : OAI21_X1 port map( B1 => n545, B2 => n460, A => n546, ZN => n542);
   U65 : INV_X1 port map( A => A(19), ZN => n460);
   U66 : OAI21_X1 port map( B1 => n461, B2 => A(19), A => B(19), ZN => n546);
   U67 : OAI21_X1 port map( B1 => n539, B2 => n457, A => n540, ZN => n536);
   U68 : INV_X1 port map( A => A(21), ZN => n457);
   U69 : OAI21_X1 port map( B1 => n458, B2 => A(21), A => B(21), ZN => n540);
   U70 : OAI21_X1 port map( B1 => n521, B2 => n448, A => n522, ZN => n518);
   U71 : INV_X1 port map( A => A(27), ZN => n448);
   U72 : OAI21_X1 port map( B1 => n449, B2 => A(27), A => B(27), ZN => n522);
   U73 : OAI21_X1 port map( B1 => n527, B2 => n451, A => n528, ZN => n524);
   U74 : OAI21_X1 port map( B1 => n452, B2 => A(25), A => B(25), ZN => n528);
   U75 : INV_X1 port map( A => n527, ZN => n452);
   U76 : OAI21_X1 port map( B1 => A(24), B2 => n530, A => n453, ZN => n527);
   U77 : INV_X1 port map( A => n531, ZN => n453);
   U78 : AOI21_X1 port map( B1 => n530, B2 => A(24), A => B(24), ZN => n531);
   U79 : OAI21_X1 port map( B1 => n483, B2 => n432, A => n484, ZN => n467);
   U80 : INV_X1 port map( A => A(39), ZN => n432);
   U81 : OAI21_X1 port map( B1 => A(39), B2 => n433, A => B(39), ZN => n484);
   U82 : XNOR2_X1 port map( A => n449, B => n523, ZN => SUM(27));
   U83 : XNOR2_X1 port map( A => A(27), B => B(27), ZN => n523);
   U84 : XNOR2_X1 port map( A => n436, B => n491, ZN => SUM(37));
   U85 : OAI21_X1 port map( B1 => n495, B2 => n437, A => n496, ZN => n493);
   U86 : INV_X1 port map( A => A(35), ZN => n437);
   U87 : OAI21_X1 port map( B1 => n438, B2 => A(35), A => B(35), ZN => n496);
   U88 : INV_X1 port map( A => n495, ZN => n438);
   U89 : AOI21_X1 port map( B1 => n486, B2 => A(38), A => n434, ZN => n483);
   U90 : INV_X1 port map( A => n487, ZN => n434);
   U91 : OAI21_X1 port map( B1 => A(38), B2 => n486, A => B(38), ZN => n487);
   U92 : XNOR2_X1 port map( A => n533, B => n535, ZN => SUM(23));
   U93 : XNOR2_X1 port map( A => n458, B => n541, ZN => SUM(21));
   U94 : XNOR2_X1 port map( A => A(21), B => B(21), ZN => n541);
   U95 : OAI21_X1 port map( B1 => A(28), B2 => n518, A => n447, ZN => n515);
   U96 : INV_X1 port map( A => n519, ZN => n447);
   U97 : AOI21_X1 port map( B1 => n518, B2 => A(28), A => B(28), ZN => n519);
   U98 : XNOR2_X1 port map( A => n446, B => n517, ZN => SUM(29));
   U99 : XNOR2_X1 port map( A => A(29), B => B(29), ZN => n517);
   U100 : OAI21_X1 port map( B1 => A(26), B2 => n524, A => n450, ZN => n521);
   U101 : INV_X1 port map( A => n525, ZN => n450);
   U102 : AOI21_X1 port map( B1 => n524, B2 => A(26), A => B(26), ZN => n525);
   U103 : OAI21_X1 port map( B1 => A(20), B2 => n542, A => n459, ZN => n539);
   U104 : INV_X1 port map( A => n543, ZN => n459);
   U105 : AOI21_X1 port map( B1 => n542, B2 => A(20), A => B(20), ZN => n543);
   U106 : OAI21_X1 port map( B1 => A(18), B2 => n548, A => n462, ZN => n545);
   U107 : INV_X1 port map( A => n549, ZN => n462);
   U108 : AOI21_X1 port map( B1 => n548, B2 => A(18), A => B(18), ZN => n549);
   U109 : AOI21_X1 port map( B1 => n467, B2 => A(40), A => n431, ZN => n466);
   U110 : INV_X1 port map( A => n468, ZN => n431);
   U111 : OAI21_X1 port map( B1 => A(40), B2 => n467, A => B(40), ZN => n468);
   U112 : XNOR2_X1 port map( A => n551, B => n553, ZN => SUM(17));
   U113 : XNOR2_X1 port map( A => B(17), B => n463, ZN => n553);
   U114 : INV_X1 port map( A => n476, ZN => n427);
   U115 : OAI22_X1 port map( A1 => n477, A2 => B(46), B1 => n428, B2 => A(46), 
                           ZN => n476);
   U116 : AND2_X1 port map( A1 => n428, A2 => A(46), ZN => n477);
   U117 : INV_X1 port map( A => n478, ZN => n428);
   U118 : INV_X1 port map( A => n473, ZN => n426);
   U119 : OAI22_X1 port map( A1 => A(47), A2 => n427, B1 => B(47), B2 => n474, 
                           ZN => n473);
   U120 : AND2_X1 port map( A1 => n427, A2 => A(47), ZN => n474);
   U121 : INV_X1 port map( A => n466, ZN => n430);
   U122 : INV_X1 port map( A => n501, ZN => n440);
   U123 : OAI22_X1 port map( A1 => A(33), A2 => n441, B1 => B(33), B2 => n502, 
                           ZN => n501);
   U124 : AND2_X1 port map( A1 => n441, A2 => A(33), ZN => n502);
   U125 : INV_X1 port map( A => n503, ZN => n441);
   U126 : INV_X1 port map( A => n513, ZN => n444);
   U127 : AOI21_X1 port map( B1 => n512, B2 => A(30), A => B(30), ZN => n513);
   U128 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT48_DW01_add_0 is

   port( A, B : in std_logic_vector (47 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (47 downto 0);  CO : out std_logic);

end RCA_NBIT48_DW01_add_0;

architecture SYN_rpl of RCA_NBIT48_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_14_port, carry_13_port, carry_12_port, carry_11_port, 
      carry_10_port, carry_9_port, carry_8_port, carry_7_port, carry_6_port, 
      carry_5_port, carry_4_port, carry_3_port, carry_2_port, n1, n510, n511, 
      n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, 
      n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, 
      n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, 
      n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, 
      n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, 
      n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, 
      n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, 
      n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, 
      n608, n609, n610, n611, n612, n613, n463, n464, n465, n466, n467, n468, 
      n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, 
      n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, 
      n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, 
      n505, n506, n507, n508, n509 : std_logic;

begin
   
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U139 : XOR2_X1 port map( A => B(47), B => A(47), Z => n511);
   U140 : XOR2_X1 port map( A => n512, B => n514, Z => SUM(46));
   U141 : XOR2_X1 port map( A => B(46), B => A(46), Z => n514);
   U142 : XOR2_X1 port map( A => n516, B => n517, Z => SUM(45));
   U143 : XOR2_X1 port map( A => B(45), B => A(45), Z => n517);
   U144 : XOR2_X1 port map( A => n467, B => n520, Z => SUM(44));
   U145 : XOR2_X1 port map( A => B(44), B => A(44), Z => n520);
   U146 : XOR2_X1 port map( A => n521, B => n523, Z => SUM(43));
   U147 : XOR2_X1 port map( A => B(43), B => A(43), Z => n523);
   U148 : XOR2_X1 port map( A => n470, B => n526, Z => SUM(42));
   U149 : XOR2_X1 port map( A => B(42), B => A(42), Z => n526);
   U150 : XOR2_X1 port map( A => n527, B => n529, Z => SUM(41));
   U151 : XOR2_X1 port map( A => B(41), B => A(41), Z => n529);
   U152 : XOR2_X1 port map( A => n476, B => n538, Z => SUM(38));
   U153 : XOR2_X1 port map( A => B(38), B => A(38), Z => n538);
   U154 : XOR2_X1 port map( A => n494, B => n542, Z => SUM(37));
   U155 : XOR2_X1 port map( A => B(36), B => A(36), Z => n545);
   U156 : NAND3_X1 port map( A1 => n551, A2 => n480, A3 => A(34), ZN => n550);
   U157 : XOR2_X1 port map( A => n552, B => n553, Z => SUM(34));
   U158 : XOR2_X1 port map( A => A(34), B => n497, Z => n553);
   U159 : XOR2_X1 port map( A => n481, B => n555, Z => SUM(33));
   U160 : XOR2_X1 port map( A => B(33), B => A(33), Z => n555);
   U161 : XOR2_X1 port map( A => n560, B => n562, Z => SUM(31));
   U162 : XOR2_X1 port map( A => n490, B => n574, Z => SUM(27));
   U163 : XOR2_X1 port map( A => B(27), B => A(27), Z => n574);
   U164 : XOR2_X1 port map( A => n575, B => n577, Z => SUM(26));
   U165 : XOR2_X1 port map( A => B(26), B => A(26), Z => n577);
   U166 : XOR2_X1 port map( A => n580, B => n578, Z => SUM(25));
   U167 : XOR2_X1 port map( A => n492, B => B(25), Z => n580);
   U168 : XOR2_X1 port map( A => n584, B => n586, Z => SUM(23));
   U169 : XOR2_X1 port map( A => n495, B => B(23), Z => n586);
   U170 : XOR2_X1 port map( A => n590, B => n591, Z => SUM(22));
   U171 : XOR2_X1 port map( A => B(22), B => A(22), Z => n591);
   U172 : XOR2_X1 port map( A => n498, B => n592, Z => SUM(21));
   U173 : XOR2_X1 port map( A => B(21), B => A(21), Z => n592);
   U174 : XOR2_X1 port map( A => n595, B => n596, Z => SUM(20));
   U175 : XOR2_X1 port map( A => B(20), B => A(20), Z => n596);
   U176 : XOR2_X1 port map( A => n598, B => n599, Z => SUM(19));
   U177 : XOR2_X1 port map( A => B(19), B => A(19), Z => n599);
   U178 : XOR2_X1 port map( A => n502, B => n602, Z => SUM(18));
   U179 : XOR2_X1 port map( A => n603, B => n605, Z => SUM(17));
   U180 : XOR2_X1 port map( A => B(17), B => A(17), Z => n605);
   U181 : XOR2_X1 port map( A => n505, B => n608, Z => SUM(16));
   U182 : XOR2_X1 port map( A => B(16), B => A(16), Z => n608);
   U183 : XOR2_X1 port map( A => n506, B => n610, Z => SUM(15));
   U184 : XOR2_X1 port map( A => B(15), B => A(15), Z => n610);
   U185 : XOR2_X1 port map( A => A(14), B => n613, Z => SUM(14));
   U186 : XOR2_X1 port map( A => carry_14_port, B => B(14), Z => n613);
   U187 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : NAND2_X1 port map( A1 => n541, A2 => n477, ZN => n540);
   U2 : INV_X1 port map( A => A(18), ZN => n501);
   U3 : OR2_X1 port map( A1 => n481, A2 => A(33), ZN => n551);
   U4 : INV_X1 port map( A => A(40), ZN => n472);
   U5 : INV_X1 port map( A => A(29), ZN => n486);
   U6 : INV_X1 port map( A => n606, ZN => n505);
   U7 : INV_X1 port map( A => A(25), ZN => n492);
   U8 : INV_X1 port map( A => n572, ZN => n490);
   U9 : INV_X1 port map( A => n600, ZN => n502);
   U10 : INV_X1 port map( A => n524, ZN => n470);
   U11 : INV_X1 port map( A => n518, ZN => n467);
   U12 : INV_X1 port map( A => n536, ZN => n476);
   U13 : XNOR2_X1 port map( A => n510, B => n511, ZN => SUM(47));
   U14 : AOI21_X1 port map( B1 => n512, B2 => A(46), A => n463, ZN => n510);
   U15 : INV_X1 port map( A => n513, ZN => n463);
   U16 : XNOR2_X1 port map( A => A(31), B => B(31), ZN => n562);
   U17 : XNOR2_X1 port map( A => B(18), B => n501, ZN => n602);
   U18 : NAND2_X1 port map( A1 => n589, A2 => n588, ZN => n590);
   U19 : NAND2_X1 port map( A1 => n480, A2 => n551, ZN => n552);
   U20 : OAI22_X1 port map( A1 => n584, A2 => n495, B1 => n585, B2 => n508, ZN 
                           => n581);
   U21 : AND2_X1 port map( A1 => n584, A2 => n495, ZN => n585);
   U22 : INV_X1 port map( A => B(23), ZN => n508);
   U23 : OAI21_X1 port map( B1 => n541, B2 => n477, A => n540, ZN => n542);
   U24 : AOI22_X1 port map( A1 => n581, A2 => A(24), B1 => n582, B2 => B(24), 
                           ZN => n578);
   U25 : OR2_X1 port map( A1 => A(24), A2 => n581, ZN => n582);
   U26 : AOI22_X1 port map( A1 => n478, A2 => A(36), B1 => n543, B2 => B(36), 
                           ZN => n541);
   U27 : OR2_X1 port map( A1 => A(36), A2 => n478, ZN => n543);
   U28 : INV_X1 port map( A => n544, ZN => n478);
   U29 : AOI21_X1 port map( B1 => n569, B2 => A(28), A => n488, ZN => n566);
   U30 : INV_X1 port map( A => n570, ZN => n488);
   U31 : OAI21_X1 port map( B1 => n569, B2 => A(28), A => B(28), ZN => n570);
   U32 : AOI21_X1 port map( B1 => n533, B2 => A(39), A => n474, ZN => n530);
   U33 : INV_X1 port map( A => n534, ZN => n474);
   U34 : OAI21_X1 port map( B1 => n533, B2 => A(39), A => B(39), ZN => n534);
   U35 : AOI21_X1 port map( B1 => n486, B2 => n566, A => n567, ZN => n563);
   U36 : AOI21_X1 port map( B1 => n487, B2 => A(29), A => B(29), ZN => n567);
   U37 : INV_X1 port map( A => n566, ZN => n487);
   U38 : AOI21_X1 port map( B1 => n572, B2 => n489, A => n573, ZN => n569);
   U39 : INV_X1 port map( A => A(27), ZN => n489);
   U40 : AOI21_X1 port map( B1 => n490, B2 => A(27), A => B(27), ZN => n573);
   U41 : AOI21_X1 port map( B1 => n475, B2 => n536, A => n537, ZN => n533);
   U42 : INV_X1 port map( A => A(38), ZN => n475);
   U43 : AOI21_X1 port map( B1 => n476, B2 => A(38), A => B(38), ZN => n537);
   U44 : OAI21_X1 port map( B1 => n560, B2 => n483, A => n561, ZN => n557);
   U45 : INV_X1 port map( A => A(31), ZN => n483);
   U46 : OAI21_X1 port map( B1 => n484, B2 => A(31), A => B(31), ZN => n561);
   U47 : INV_X1 port map( A => n560, ZN => n484);
   U48 : OAI21_X1 port map( B1 => n549, B2 => n497, A => n550, ZN => n546);
   U49 : AOI221_X1 port map( B1 => A(33), B2 => n481, C1 => B(33), C2 => n551, 
                           A => A(34), ZN => n549);
   U50 : OAI21_X1 port map( B1 => n563, B2 => B(30), A => n485, ZN => n560);
   U51 : INV_X1 port map( A => n564, ZN => n485);
   U52 : AOI21_X1 port map( B1 => n563, B2 => B(30), A => A(30), ZN => n564);
   U53 : XNOR2_X1 port map( A => n566, B => n568, ZN => SUM(29));
   U54 : XNOR2_X1 port map( A => B(29), B => n486, ZN => n568);
   U55 : OAI21_X1 port map( B1 => B(22), B2 => A(22), A => n587, ZN => n584);
   U56 : OAI211_X1 port map( C1 => n496, C2 => n509, A => n588, B => n589, ZN 
                           => n587);
   U57 : INV_X1 port map( A => A(22), ZN => n496);
   U58 : INV_X1 port map( A => B(22), ZN => n509);
   U59 : AOI21_X1 port map( B1 => n492, B2 => n578, A => n579, ZN => n575);
   U60 : AOI21_X1 port map( B1 => n493, B2 => A(25), A => B(25), ZN => n579);
   U61 : INV_X1 port map( A => n578, ZN => n493);
   U62 : AOI22_X1 port map( A1 => n506, A2 => A(15), B1 => n609, B2 => B(15), 
                           ZN => n606);
   U63 : OR2_X1 port map( A1 => A(15), A2 => n506, ZN => n609);
   U64 : AOI21_X1 port map( B1 => n501, B2 => n600, A => n601, ZN => n598);
   U65 : AOI21_X1 port map( B1 => n502, B2 => A(18), A => B(18), ZN => n601);
   U66 : AOI21_X1 port map( B1 => n504, B2 => n606, A => n607, ZN => n603);
   U67 : INV_X1 port map( A => A(16), ZN => n504);
   U68 : AOI21_X1 port map( B1 => n505, B2 => A(16), A => B(16), ZN => n607);
   U69 : AOI21_X1 port map( B1 => n464, B2 => n465, A => n515, ZN => n512);
   U70 : INV_X1 port map( A => n516, ZN => n465);
   U71 : INV_X1 port map( A => A(45), ZN => n464);
   U72 : AOI21_X1 port map( B1 => n516, B2 => A(45), A => B(45), ZN => n515);
   U73 : OAI21_X1 port map( B1 => B(21), B2 => n498, A => A(21), ZN => n589);
   U74 : XNOR2_X1 port map( A => n563, B => n565, ZN => SUM(30));
   U75 : XNOR2_X1 port map( A => A(30), B => B(30), ZN => n565);
   U76 : XNOR2_X1 port map( A => n583, B => n581, ZN => SUM(24));
   U77 : XNOR2_X1 port map( A => A(24), B => B(24), ZN => n583);
   U78 : XNOR2_X1 port map( A => n548, B => n546, ZN => SUM(35));
   U79 : XNOR2_X1 port map( A => A(35), B => B(35), ZN => n548);
   U80 : XNOR2_X1 port map( A => n569, B => n571, ZN => SUM(28));
   U81 : XNOR2_X1 port map( A => A(28), B => B(28), ZN => n571);
   U82 : XNOR2_X1 port map( A => n530, B => n532, ZN => SUM(40));
   U83 : XNOR2_X1 port map( A => B(40), B => n472, ZN => n532);
   U84 : XNOR2_X1 port map( A => n533, B => n535, ZN => SUM(39));
   U85 : XNOR2_X1 port map( A => A(39), B => B(39), ZN => n535);
   U86 : OAI21_X1 port map( B1 => n530, B2 => n472, A => n531, ZN => n527);
   U87 : OAI21_X1 port map( B1 => A(40), B2 => n473, A => B(40), ZN => n531);
   U88 : INV_X1 port map( A => n530, ZN => n473);
   U89 : OAI21_X1 port map( B1 => n524, B2 => n469, A => n525, ZN => n521);
   U90 : INV_X1 port map( A => A(42), ZN => n469);
   U91 : OAI21_X1 port map( B1 => n470, B2 => A(42), A => B(42), ZN => n525);
   U92 : OAI21_X1 port map( B1 => n518, B2 => n466, A => n519, ZN => n516);
   U93 : INV_X1 port map( A => A(44), ZN => n466);
   U94 : OAI21_X1 port map( B1 => n467, B2 => A(44), A => B(44), ZN => n519);
   U95 : AOI21_X1 port map( B1 => n603, B2 => A(17), A => n503, ZN => n600);
   U96 : INV_X1 port map( A => n604, ZN => n503);
   U97 : OAI21_X1 port map( B1 => n603, B2 => A(17), A => B(17), ZN => n604);
   U98 : XNOR2_X1 port map( A => n559, B => n557, ZN => SUM(32));
   U99 : XNOR2_X1 port map( A => A(32), B => B(32), ZN => n559);
   U100 : XNOR2_X1 port map( A => n544, B => n545, ZN => SUM(36));
   U101 : OAI21_X1 port map( B1 => A(35), B2 => n546, A => n479, ZN => n544);
   U102 : INV_X1 port map( A => n547, ZN => n479);
   U103 : AOI21_X1 port map( B1 => n546, B2 => A(35), A => B(35), ZN => n547);
   U104 : OAI21_X1 port map( B1 => A(26), B2 => n575, A => n491, ZN => n572);
   U105 : INV_X1 port map( A => n576, ZN => n491);
   U106 : AOI21_X1 port map( B1 => n575, B2 => A(26), A => B(26), ZN => n576);
   U107 : OAI21_X1 port map( B1 => A(41), B2 => n527, A => n471, ZN => n524);
   U108 : INV_X1 port map( A => n528, ZN => n471);
   U109 : AOI21_X1 port map( B1 => n527, B2 => A(41), A => B(41), ZN => n528);
   U110 : OAI21_X1 port map( B1 => A(43), B2 => n521, A => n468, ZN => n518);
   U111 : INV_X1 port map( A => n522, ZN => n468);
   U112 : AOI21_X1 port map( B1 => n521, B2 => A(43), A => B(43), ZN => n522);
   U113 : NAND2_X1 port map( A1 => B(21), A2 => n498, ZN => n588);
   U114 : OAI21_X1 port map( B1 => n500, B2 => n499, A => n597, ZN => n595);
   U115 : INV_X1 port map( A => n598, ZN => n500);
   U116 : INV_X1 port map( A => A(19), ZN => n499);
   U117 : OAI21_X1 port map( B1 => n598, B2 => A(19), A => B(19), ZN => n597);
   U118 : OAI21_X1 port map( B1 => n512, B2 => A(46), A => B(46), ZN => n513);
   U119 : INV_X1 port map( A => n556, ZN => n481);
   U120 : AOI21_X1 port map( B1 => n557, B2 => A(32), A => n482, ZN => n556);
   U121 : INV_X1 port map( A => n558, ZN => n482);
   U122 : OAI21_X1 port map( B1 => A(32), B2 => n557, A => B(32), ZN => n558);
   U123 : INV_X1 port map( A => n593, ZN => n498);
   U124 : OAI22_X1 port map( A1 => A(20), A2 => B(20), B1 => n594, B2 => n595, 
                           ZN => n593);
   U125 : AND2_X1 port map( A1 => A(20), A2 => B(20), ZN => n594);
   U126 : INV_X1 port map( A => A(37), ZN => n477);
   U127 : NAND2_X1 port map( A1 => n539, A2 => n540, ZN => n536);
   U128 : OAI21_X1 port map( B1 => n541, B2 => n477, A => n494, ZN => n539);
   U129 : INV_X1 port map( A => n611, ZN => n506);
   U130 : AOI21_X1 port map( B1 => A(14), B2 => B(14), A => n507, ZN => n611);
   U131 : INV_X1 port map( A => n612, ZN => n507);
   U132 : OAI21_X1 port map( B1 => A(14), B2 => B(14), A => carry_14_port, ZN 
                           => n612);
   U133 : INV_X1 port map( A => A(23), ZN => n495);
   U134 : INV_X1 port map( A => n554, ZN => n480);
   U135 : AOI21_X1 port map( B1 => n481, B2 => A(33), A => B(33), ZN => n554);
   U136 : INV_X1 port map( A => B(34), ZN => n497);
   U137 : INV_X1 port map( A => B(37), ZN => n494);
   U138 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT46_DW01_add_0 is

   port( A, B : in std_logic_vector (45 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (45 downto 0);  CO : out std_logic);

end RCA_NBIT46_DW01_add_0;

architecture SYN_rpl of RCA_NBIT46_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_12_port, carry_11_port, carry_10_port, carry_9_port, 
      carry_8_port, carry_7_port, carry_6_port, carry_5_port, carry_4_port, 
      carry_3_port, carry_2_port, n1, n525, n526, n527, n528, n529, n530, n531,
      n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, 
      n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, 
      n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, 
      n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, 
      n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, 
      n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, 
      n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, 
      n616, n617, n618, n619, n620, n621, n622, n623, n624, n482, n483, n484, 
      n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, 
      n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, 
      n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, 
      n521, n522, n523, n524 : std_logic;

begin
   
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U136 : XOR2_X1 port map( A => B(45), B => A(45), Z => n526);
   U137 : XOR2_X1 port map( A => n527, B => n529, Z => SUM(44));
   U138 : XOR2_X1 port map( A => B(44), B => A(44), Z => n529);
   U139 : XOR2_X1 port map( A => B(43), B => A(43), Z => n532);
   U140 : XOR2_X1 port map( A => n533, B => n535, Z => SUM(42));
   U141 : XOR2_X1 port map( A => B(42), B => A(42), Z => n535);
   U142 : XOR2_X1 port map( A => B(41), B => A(41), Z => n538);
   U143 : XOR2_X1 port map( A => n539, B => n541, Z => SUM(40));
   U144 : XOR2_X1 port map( A => B(40), B => A(40), Z => n541);
   U145 : XOR2_X1 port map( A => B(39), B => A(39), Z => n544);
   U146 : XOR2_X1 port map( A => n545, B => n547, Z => SUM(38));
   U147 : XOR2_X1 port map( A => B(38), B => A(38), Z => n547);
   U148 : XOR2_X1 port map( A => B(37), B => A(37), Z => n550);
   U149 : XOR2_X1 port map( A => n551, B => n553, Z => SUM(36));
   U150 : XOR2_X1 port map( A => B(36), B => A(36), Z => n553);
   U151 : XOR2_X1 port map( A => B(35), B => A(35), Z => n556);
   U152 : XOR2_X1 port map( A => n557, B => n559, Z => SUM(34));
   U153 : XOR2_X1 port map( A => B(34), B => A(34), Z => n559);
   U154 : XOR2_X1 port map( A => B(33), B => A(33), Z => n562);
   U155 : XOR2_X1 port map( A => n563, B => n565, Z => SUM(32));
   U156 : XOR2_X1 port map( A => B(32), B => A(32), Z => n565);
   U157 : XOR2_X1 port map( A => B(31), B => A(31), Z => n568);
   U158 : XOR2_X1 port map( A => n569, B => n571, Z => SUM(30));
   U159 : XOR2_X1 port map( A => B(30), B => A(30), Z => n571);
   U160 : XOR2_X1 port map( A => B(29), B => A(29), Z => n574);
   U161 : XOR2_X1 port map( A => n575, B => n577, Z => SUM(28));
   U162 : XOR2_X1 port map( A => B(28), B => A(28), Z => n577);
   U163 : XOR2_X1 port map( A => B(26), B => A(26), Z => n583);
   U164 : XOR2_X1 port map( A => B(25), B => A(25), Z => n586);
   U165 : XOR2_X1 port map( A => n587, B => n589, Z => SUM(24));
   U166 : XOR2_X1 port map( A => B(24), B => A(24), Z => n589);
   U167 : XOR2_X1 port map( A => B(22), B => A(22), Z => n595);
   U168 : XOR2_X1 port map( A => B(21), B => A(21), Z => n598);
   U169 : XOR2_X1 port map( A => n599, B => n601, Z => SUM(20));
   U170 : XOR2_X1 port map( A => B(20), B => A(20), Z => n601);
   U171 : XOR2_X1 port map( A => n605, B => n607, Z => SUM(18));
   U172 : XOR2_X1 port map( A => B(18), B => A(18), Z => n607);
   U173 : XOR2_X1 port map( A => n518, B => n610, Z => SUM(17));
   U174 : XOR2_X1 port map( A => B(17), B => A(17), Z => n610);
   U175 : XOR2_X1 port map( A => B(14), B => A(14), Z => n619);
   U176 : XOR2_X1 port map( A => B(13), B => A(13), Z => n622);
   U177 : XOR2_X1 port map( A => A(12), B => n624, Z => SUM(12));
   U178 : XOR2_X1 port map( A => carry_12_port, B => B(12), Z => n624);
   U179 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : INV_X1 port map( A => A(15), ZN => n520);
   U2 : INV_X1 port map( A => A(19), ZN => n514);
   U3 : INV_X1 port map( A => A(23), ZN => n510);
   U4 : INV_X1 port map( A => A(27), ZN => n505);
   U5 : INV_X1 port map( A => n579, ZN => n506);
   U6 : INV_X1 port map( A => n608, ZN => n518);
   U7 : XNOR2_X1 port map( A => n525, B => n526, ZN => SUM(45));
   U8 : AOI21_X1 port map( B1 => n527, B2 => A(44), A => n482, ZN => n525);
   U9 : INV_X1 port map( A => n528, ZN => n482);
   U10 : OAI22_X1 port map( A1 => A(14), A2 => n522, B1 => B(14), B2 => n617, 
                           ZN => n614);
   U11 : AND2_X1 port map( A1 => n522, A2 => A(14), ZN => n617);
   U12 : INV_X1 port map( A => n618, ZN => n522);
   U13 : AOI22_X1 port map( A1 => n512, A2 => A(22), B1 => n593, B2 => B(22), 
                           ZN => n590);
   U14 : OR2_X1 port map( A1 => A(22), A2 => n512, ZN => n593);
   U15 : INV_X1 port map( A => n594, ZN => n512);
   U16 : OAI22_X1 port map( A1 => A(13), A2 => n523, B1 => B(13), B2 => n620, 
                           ZN => n618);
   U17 : AND2_X1 port map( A1 => n523, A2 => A(13), ZN => n620);
   U18 : INV_X1 port map( A => n621, ZN => n523);
   U19 : AOI22_X1 port map( A1 => n509, A2 => A(25), B1 => n584, B2 => B(25), 
                           ZN => n581);
   U20 : OR2_X1 port map( A1 => A(25), A2 => n509, ZN => n584);
   U21 : INV_X1 port map( A => n585, ZN => n509);
   U22 : AOI22_X1 port map( A1 => n575, A2 => A(28), B1 => n576, B2 => B(28), 
                           ZN => n572);
   U23 : OR2_X1 port map( A1 => n575, A2 => A(28), ZN => n576);
   U24 : AOI22_X1 port map( A1 => n569, A2 => A(30), B1 => n570, B2 => B(30), 
                           ZN => n566);
   U25 : OR2_X1 port map( A1 => A(30), A2 => n569, ZN => n570);
   U26 : AOI21_X1 port map( B1 => n605, B2 => A(18), A => n516, ZN => n602);
   U27 : INV_X1 port map( A => n606, ZN => n516);
   U28 : OAI21_X1 port map( B1 => A(18), B2 => n605, A => B(18), ZN => n606);
   U29 : AOI21_X1 port map( B1 => n551, B2 => A(36), A => n494, ZN => n548);
   U30 : INV_X1 port map( A => n552, ZN => n494);
   U31 : OAI21_X1 port map( B1 => A(36), B2 => n551, A => B(36), ZN => n552);
   U32 : AOI21_X1 port map( B1 => n563, B2 => A(32), A => n500, ZN => n560);
   U33 : INV_X1 port map( A => n564, ZN => n500);
   U34 : OAI21_X1 port map( B1 => A(32), B2 => n563, A => B(32), ZN => n564);
   U35 : AOI21_X1 port map( B1 => n545, B2 => A(38), A => n491, ZN => n542);
   U36 : INV_X1 port map( A => n546, ZN => n491);
   U37 : OAI21_X1 port map( B1 => A(38), B2 => n545, A => B(38), ZN => n546);
   U38 : AOI21_X1 port map( B1 => n539, B2 => A(40), A => n488, ZN => n536);
   U39 : INV_X1 port map( A => n540, ZN => n488);
   U40 : OAI21_X1 port map( B1 => A(40), B2 => n539, A => B(40), ZN => n540);
   U41 : AOI21_X1 port map( B1 => n533, B2 => A(42), A => n484, ZN => n530);
   U42 : INV_X1 port map( A => n534, ZN => n484);
   U43 : OAI21_X1 port map( B1 => A(42), B2 => n533, A => B(42), ZN => n534);
   U44 : AOI21_X1 port map( B1 => n557, B2 => A(34), A => n497, ZN => n554);
   U45 : INV_X1 port map( A => n558, ZN => n497);
   U46 : OAI21_X1 port map( B1 => A(34), B2 => n557, A => B(34), ZN => n558);
   U47 : AOI21_X1 port map( B1 => n520, B2 => n614, A => n615, ZN => n611);
   U48 : AOI21_X1 port map( B1 => n521, B2 => A(15), A => B(15), ZN => n615);
   U49 : INV_X1 port map( A => n614, ZN => n521);
   U50 : XNOR2_X1 port map( A => n560, B => n562, ZN => SUM(33));
   U51 : XNOR2_X1 port map( A => n542, B => n544, ZN => SUM(39));
   U52 : XNOR2_X1 port map( A => n566, B => n568, ZN => SUM(31));
   U53 : XNOR2_X1 port map( A => n554, B => n556, ZN => SUM(35));
   U54 : AOI22_X1 port map( A1 => n599, A2 => A(20), B1 => n600, B2 => B(20), 
                           ZN => n597);
   U55 : OR2_X1 port map( A1 => n599, A2 => A(20), ZN => n600);
   U56 : AOI22_X1 port map( A1 => n513, A2 => A(21), B1 => n596, B2 => B(21), 
                           ZN => n594);
   U57 : OR2_X1 port map( A1 => A(21), A2 => n513, ZN => n596);
   U58 : INV_X1 port map( A => n597, ZN => n513);
   U59 : AOI22_X1 port map( A1 => n587, A2 => A(24), B1 => n588, B2 => B(24), 
                           ZN => n585);
   U60 : OR2_X1 port map( A1 => n587, A2 => A(24), ZN => n588);
   U61 : OAI21_X1 port map( B1 => B(12), B2 => A(12), A => n524, ZN => n621);
   U62 : INV_X1 port map( A => n623, ZN => n524);
   U63 : AOI21_X1 port map( B1 => A(12), B2 => B(12), A => carry_12_port, ZN =>
                           n623);
   U64 : XNOR2_X1 port map( A => n611, B => n613, ZN => SUM(16));
   U65 : XNOR2_X1 port map( A => A(16), B => B(16), ZN => n613);
   U66 : XNOR2_X1 port map( A => n506, B => n580, ZN => SUM(27));
   U67 : XNOR2_X1 port map( A => B(27), B => n505, ZN => n580);
   U68 : XNOR2_X1 port map( A => n581, B => n583, ZN => SUM(26));
   U69 : XNOR2_X1 port map( A => n594, B => n595, ZN => SUM(22));
   U70 : XNOR2_X1 port map( A => n536, B => n538, ZN => SUM(41));
   U71 : XNOR2_X1 port map( A => n530, B => n532, ZN => SUM(43));
   U72 : XNOR2_X1 port map( A => n602, B => n604, ZN => SUM(19));
   U73 : XNOR2_X1 port map( A => B(19), B => n514, ZN => n604);
   U74 : OAI21_X1 port map( B1 => n566, B2 => n501, A => n567, ZN => n563);
   U75 : INV_X1 port map( A => A(31), ZN => n501);
   U76 : OAI21_X1 port map( B1 => A(31), B2 => n502, A => B(31), ZN => n567);
   U77 : INV_X1 port map( A => n566, ZN => n502);
   U78 : OAI21_X1 port map( B1 => n560, B2 => n498, A => n561, ZN => n557);
   U79 : INV_X1 port map( A => A(33), ZN => n498);
   U80 : OAI21_X1 port map( B1 => A(33), B2 => n499, A => B(33), ZN => n561);
   U81 : INV_X1 port map( A => n560, ZN => n499);
   U82 : XNOR2_X1 port map( A => n618, B => n619, ZN => SUM(14));
   U83 : OAI21_X1 port map( B1 => n554, B2 => n495, A => n555, ZN => n551);
   U84 : INV_X1 port map( A => A(35), ZN => n495);
   U85 : OAI21_X1 port map( B1 => A(35), B2 => n496, A => B(35), ZN => n555);
   U86 : INV_X1 port map( A => n554, ZN => n496);
   U87 : OAI21_X1 port map( B1 => n548, B2 => n492, A => n549, ZN => n545);
   U88 : INV_X1 port map( A => A(37), ZN => n492);
   U89 : OAI21_X1 port map( B1 => A(37), B2 => n493, A => B(37), ZN => n549);
   U90 : INV_X1 port map( A => n548, ZN => n493);
   U91 : OAI21_X1 port map( B1 => n542, B2 => n489, A => n543, ZN => n539);
   U92 : INV_X1 port map( A => A(39), ZN => n489);
   U93 : OAI21_X1 port map( B1 => A(39), B2 => n490, A => B(39), ZN => n543);
   U94 : INV_X1 port map( A => n542, ZN => n490);
   U95 : OAI21_X1 port map( B1 => n536, B2 => n486, A => n537, ZN => n533);
   U96 : INV_X1 port map( A => A(41), ZN => n486);
   U97 : OAI21_X1 port map( B1 => A(41), B2 => n487, A => B(41), ZN => n537);
   U98 : INV_X1 port map( A => n536, ZN => n487);
   U99 : OAI21_X1 port map( B1 => n530, B2 => n485, A => n531, ZN => n527);
   U100 : INV_X1 port map( A => A(43), ZN => n485);
   U101 : OAI21_X1 port map( B1 => A(43), B2 => n483, A => B(43), ZN => n531);
   U102 : INV_X1 port map( A => n530, ZN => n483);
   U103 : OAI21_X1 port map( B1 => n608, B2 => n517, A => n609, ZN => n605);
   U104 : INV_X1 port map( A => A(17), ZN => n517);
   U105 : OAI21_X1 port map( B1 => A(17), B2 => n518, A => B(17), ZN => n609);
   U106 : AOI21_X1 port map( B1 => n510, B2 => n590, A => n591, ZN => n587);
   U107 : AOI21_X1 port map( B1 => n511, B2 => A(23), A => B(23), ZN => n591);
   U108 : INV_X1 port map( A => n590, ZN => n511);
   U109 : AOI21_X1 port map( B1 => n514, B2 => n602, A => n603, ZN => n599);
   U110 : AOI21_X1 port map( B1 => n515, B2 => A(19), A => B(19), ZN => n603);
   U111 : INV_X1 port map( A => n602, ZN => n515);
   U112 : AOI21_X1 port map( B1 => n505, B2 => n506, A => n578, ZN => n575);
   U113 : AOI21_X1 port map( B1 => n579, B2 => A(27), A => B(27), ZN => n578);
   U114 : XNOR2_X1 port map( A => n614, B => n616, ZN => SUM(15));
   U115 : XNOR2_X1 port map( A => B(15), B => n520, ZN => n616);
   U116 : AOI21_X1 port map( B1 => n611, B2 => A(16), A => n519, ZN => n608);
   U117 : INV_X1 port map( A => n612, ZN => n519);
   U118 : OAI21_X1 port map( B1 => n611, B2 => A(16), A => B(16), ZN => n612);
   U119 : OAI21_X1 port map( B1 => n572, B2 => n503, A => n573, ZN => n569);
   U120 : INV_X1 port map( A => A(29), ZN => n503);
   U121 : OAI21_X1 port map( B1 => A(29), B2 => n504, A => B(29), ZN => n573);
   U122 : INV_X1 port map( A => n572, ZN => n504);
   U123 : XNOR2_X1 port map( A => n572, B => n574, ZN => SUM(29));
   U124 : XNOR2_X1 port map( A => n585, B => n586, ZN => SUM(25));
   U125 : OAI21_X1 port map( B1 => n581, B2 => n507, A => n582, ZN => n579);
   U126 : INV_X1 port map( A => A(26), ZN => n507);
   U127 : OAI21_X1 port map( B1 => A(26), B2 => n508, A => B(26), ZN => n582);
   U128 : INV_X1 port map( A => n581, ZN => n508);
   U129 : XNOR2_X1 port map( A => n597, B => n598, ZN => SUM(21));
   U130 : OAI21_X1 port map( B1 => A(44), B2 => n527, A => B(44), ZN => n528);
   U131 : XNOR2_X1 port map( A => n548, B => n550, ZN => SUM(37));
   U132 : XNOR2_X1 port map( A => n590, B => n592, ZN => SUM(23));
   U133 : XNOR2_X1 port map( A => B(23), B => n510, ZN => n592);
   U134 : XNOR2_X1 port map( A => n621, B => n622, ZN => SUM(13));
   U135 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT44_DW01_add_0 is

   port( A, B : in std_logic_vector (43 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (43 downto 0);  CO : out std_logic);

end RCA_NBIT44_DW01_add_0;

architecture SYN_rpl of RCA_NBIT44_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal n1, carry_9_port, carry_8_port, carry_7_port, carry_6_port, 
      carry_5_port, carry_4_port, carry_3_port, carry_2_port, carry_10_port, 
      carry_14_port, carry_13_port, n523, n524, n525, n526, n527, n528, n529, 
      n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, 
      n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, 
      n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, 
      n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, 
      n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, 
      n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, 
      n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, 
      n614, n615, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, 
      n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, 
      n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, 
      n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522 : 
      std_logic;

begin
   
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => n521, CO => 
                           carry_13_port, S => SUM(12));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U134 : XOR2_X1 port map( A => B(43), B => A(43), Z => n526);
   U135 : XOR2_X1 port map( A => n530, B => n532, Z => SUM(41));
   U136 : XOR2_X1 port map( A => n536, B => n538, Z => SUM(39));
   U137 : XOR2_X1 port map( A => n542, B => n544, Z => SUM(37));
   U138 : XOR2_X1 port map( A => n550, B => n551, Z => SUM(35));
   U139 : XOR2_X1 port map( A => n491, B => n557, Z => SUM(33));
   U140 : XOR2_X1 port map( A => n493, B => n560, Z => SUM(32));
   U141 : XOR2_X1 port map( A => n561, B => n563, Z => SUM(31));
   U142 : XOR2_X1 port map( A => B(31), B => A(31), Z => n563);
   U143 : XOR2_X1 port map( A => n496, B => n566, Z => SUM(30));
   U144 : XOR2_X1 port map( A => B(29), B => A(29), Z => n569);
   U145 : XOR2_X1 port map( A => n504, B => n581, Z => SUM(25));
   U146 : XOR2_X1 port map( A => B(25), B => A(25), Z => n581);
   U147 : XOR2_X1 port map( A => n582, B => n584, Z => SUM(24));
   U148 : XOR2_X1 port map( A => B(24), B => A(24), Z => n584);
   U149 : XOR2_X1 port map( A => n507, B => n587, Z => SUM(23));
   U150 : XOR2_X1 port map( A => B(23), B => A(23), Z => n587);
   U151 : XOR2_X1 port map( A => n588, B => n590, Z => SUM(22));
   U152 : XOR2_X1 port map( A => B(22), B => A(22), Z => n590);
   U153 : XOR2_X1 port map( A => n510, B => n593, Z => SUM(21));
   U154 : XOR2_X1 port map( A => n594, B => n596, Z => SUM(20));
   U155 : XOR2_X1 port map( A => B(20), B => A(20), Z => n596);
   U156 : XOR2_X1 port map( A => n597, B => n599, Z => SUM(19));
   U157 : XOR2_X1 port map( A => n512, B => B(19), Z => n599);
   U158 : XOR2_X1 port map( A => n600, B => n602, Z => SUM(18));
   U159 : XOR2_X1 port map( A => B(18), B => A(18), Z => n602);
   U160 : XOR2_X1 port map( A => n603, B => n605, Z => SUM(17));
   U161 : XOR2_X1 port map( A => n515, B => B(17), Z => n605);
   U162 : XOR2_X1 port map( A => n606, B => n608, Z => SUM(16));
   U163 : XOR2_X1 port map( A => B(16), B => A(16), Z => n608);
   U164 : XOR2_X1 port map( A => n519, B => n611, Z => SUM(15));
   U165 : XOR2_X1 port map( A => B(15), B => A(15), Z => n611);
   U166 : XOR2_X1 port map( A => A(14), B => n613, Z => SUM(14));
   U167 : XOR2_X1 port map( A => carry_14_port, B => B(14), Z => n613);
   U168 : XOR2_X1 port map( A => n522, B => n524, Z => SUM(11));
   U169 : XOR2_X1 port map( A => A(11), B => B(11), Z => n524);
   U170 : XOR2_X1 port map( A => carry_10_port, B => n615, Z => SUM(10));
   U171 : XOR2_X1 port map( A => A(10), B => B(10), Z => n615);
   U172 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : NAND2_X1 port map( A1 => n547, A2 => n487, ZN => n546);
   U2 : INV_X1 port map( A => A(32), ZN => n492);
   U3 : INV_X1 port map( A => A(21), ZN => n509);
   U4 : INV_X1 port map( A => A(27), ZN => n500);
   U5 : INV_X1 port map( A => A(17), ZN => n515);
   U6 : INV_X1 port map( A => A(19), ZN => n512);
   U7 : INV_X1 port map( A => n609, ZN => n519);
   U8 : INV_X1 port map( A => n579, ZN => n504);
   U9 : INV_X1 port map( A => n558, ZN => n493);
   U10 : INV_X1 port map( A => n556, ZN => n491);
   U11 : INV_X1 port map( A => n591, ZN => n510);
   U12 : INV_X1 port map( A => n585, ZN => n507);
   U13 : INV_X1 port map( A => n564, ZN => n496);
   U14 : XNOR2_X1 port map( A => n525, B => n526, ZN => SUM(43));
   U15 : AOI21_X1 port map( B1 => n527, B2 => A(42), A => n478, ZN => n525);
   U16 : INV_X1 port map( A => n528, ZN => n478);
   U17 : XNOR2_X1 port map( A => B(32), B => n492, ZN => n560);
   U18 : XNOR2_X1 port map( A => A(33), B => B(33), ZN => n557);
   U19 : XNOR2_X1 port map( A => A(35), B => B(35), ZN => n551);
   U20 : XNOR2_X1 port map( A => A(37), B => B(37), ZN => n544);
   U21 : XNOR2_X1 port map( A => A(39), B => B(39), ZN => n538);
   U22 : XNOR2_X1 port map( A => A(41), B => B(41), ZN => n532);
   U23 : XNOR2_X1 port map( A => B(21), B => n509, ZN => n593);
   U24 : XNOR2_X1 port map( A => B(30), B => n495, ZN => n566);
   U25 : AOI21_X1 port map( B1 => n576, B2 => A(26), A => n502, ZN => n573);
   U26 : INV_X1 port map( A => n577, ZN => n502);
   U27 : OAI21_X1 port map( B1 => n576, B2 => A(26), A => B(26), ZN => n577);
   U28 : OAI22_X1 port map( A1 => n552, A2 => A(34), B1 => n553, B2 => B(34), 
                           ZN => n550);
   U29 : AND2_X1 port map( A1 => n552, A2 => A(34), ZN => n553);
   U30 : XNOR2_X1 port map( A => B(36), B => n548, ZN => SUM(36));
   U31 : OAI21_X1 port map( B1 => n547, B2 => n487, A => n546, ZN => n548);
   U32 : AOI21_X1 port map( B1 => n500, B2 => n573, A => n574, ZN => n570);
   U33 : AOI21_X1 port map( B1 => n501, B2 => A(27), A => B(27), ZN => n574);
   U34 : INV_X1 port map( A => n573, ZN => n501);
   U35 : AOI21_X1 port map( B1 => n579, B2 => n503, A => n580, ZN => n576);
   U36 : INV_X1 port map( A => A(25), ZN => n503);
   U37 : AOI21_X1 port map( B1 => n504, B2 => A(25), A => B(25), ZN => n580);
   U38 : OAI21_X1 port map( B1 => n542, B2 => n485, A => n543, ZN => n539);
   U39 : INV_X1 port map( A => A(37), ZN => n485);
   U40 : OAI21_X1 port map( B1 => A(37), B2 => n486, A => B(37), ZN => n543);
   U41 : INV_X1 port map( A => n542, ZN => n486);
   U42 : OAI21_X1 port map( B1 => n530, B2 => n479, A => n531, ZN => n527);
   U43 : INV_X1 port map( A => A(41), ZN => n479);
   U44 : OAI21_X1 port map( B1 => n480, B2 => A(41), A => B(41), ZN => n531);
   U45 : INV_X1 port map( A => n530, ZN => n480);
   U46 : OAI21_X1 port map( B1 => n536, B2 => n482, A => n537, ZN => n533);
   U47 : INV_X1 port map( A => A(39), ZN => n482);
   U48 : OAI21_X1 port map( B1 => n483, B2 => A(39), A => B(39), ZN => n537);
   U49 : INV_X1 port map( A => n536, ZN => n483);
   U50 : AOI21_X1 port map( B1 => n489, B2 => A(35), A => n488, ZN => n547);
   U51 : INV_X1 port map( A => n549, ZN => n488);
   U52 : OAI21_X1 port map( B1 => n489, B2 => A(35), A => B(35), ZN => n549);
   U53 : INV_X1 port map( A => n550, ZN => n489);
   U54 : AOI21_X1 port map( B1 => A(14), B2 => B(14), A => n520, ZN => n609);
   U55 : INV_X1 port map( A => n612, ZN => n520);
   U56 : OAI21_X1 port map( B1 => A(14), B2 => B(14), A => carry_14_port, ZN =>
                           n612);
   U57 : OAI21_X1 port map( B1 => n545, B2 => B(36), A => n546, ZN => n542);
   U58 : NOR2_X1 port map( A1 => n547, A2 => n487, ZN => n545);
   U59 : AOI21_X1 port map( B1 => n490, B2 => n491, A => n555, ZN => n552);
   U60 : INV_X1 port map( A => A(33), ZN => n490);
   U61 : AOI21_X1 port map( B1 => n556, B2 => A(33), A => B(33), ZN => n555);
   U62 : AOI21_X1 port map( B1 => n518, B2 => n609, A => n610, ZN => n606);
   U63 : INV_X1 port map( A => A(15), ZN => n518);
   U64 : AOI21_X1 port map( B1 => n519, B2 => A(15), A => B(15), ZN => n610);
   U65 : XNOR2_X1 port map( A => n529, B => n527, ZN => SUM(42));
   U66 : XNOR2_X1 port map( A => A(42), B => B(42), ZN => n529);
   U67 : XNOR2_X1 port map( A => n541, B => n539, ZN => SUM(38));
   U68 : XNOR2_X1 port map( A => A(38), B => B(38), ZN => n541);
   U69 : XNOR2_X1 port map( A => n535, B => n533, ZN => SUM(40));
   U70 : XNOR2_X1 port map( A => A(40), B => B(40), ZN => n535);
   U71 : XNOR2_X1 port map( A => n552, B => n554, ZN => SUM(34));
   U72 : XNOR2_X1 port map( A => A(34), B => B(34), ZN => n554);
   U73 : XNOR2_X1 port map( A => n568, B => n569, ZN => SUM(29));
   U74 : XNOR2_X1 port map( A => n576, B => n578, ZN => SUM(26));
   U75 : XNOR2_X1 port map( A => A(26), B => B(26), ZN => n578);
   U76 : OAI21_X1 port map( B1 => n603, B2 => n515, A => n604, ZN => n600);
   U77 : OAI21_X1 port map( B1 => n516, B2 => A(17), A => B(17), ZN => n604);
   U78 : INV_X1 port map( A => n603, ZN => n516);
   U79 : OAI21_X1 port map( B1 => n597, B2 => n512, A => n598, ZN => n594);
   U80 : OAI21_X1 port map( B1 => n513, B2 => A(19), A => B(19), ZN => n598);
   U81 : INV_X1 port map( A => n597, ZN => n513);
   U82 : OAI21_X1 port map( B1 => A(40), B2 => n533, A => n481, ZN => n530);
   U83 : INV_X1 port map( A => n534, ZN => n481);
   U84 : AOI21_X1 port map( B1 => n533, B2 => A(40), A => B(40), ZN => n534);
   U85 : OAI21_X1 port map( B1 => A(38), B2 => n539, A => n484, ZN => n536);
   U86 : INV_X1 port map( A => n540, ZN => n484);
   U87 : AOI21_X1 port map( B1 => n539, B2 => A(38), A => B(38), ZN => n540);
   U88 : OAI21_X1 port map( B1 => A(18), B2 => n600, A => n514, ZN => n597);
   U89 : INV_X1 port map( A => n601, ZN => n514);
   U90 : AOI21_X1 port map( B1 => n600, B2 => A(18), A => B(18), ZN => n601);
   U91 : OAI21_X1 port map( B1 => A(16), B2 => n606, A => n517, ZN => n603);
   U92 : INV_X1 port map( A => n607, ZN => n517);
   U93 : AOI21_X1 port map( B1 => n606, B2 => A(16), A => B(16), ZN => n607);
   U94 : OAI21_X1 port map( B1 => n591, B2 => n509, A => n592, ZN => n588);
   U95 : OAI21_X1 port map( B1 => n510, B2 => A(21), A => B(21), ZN => n592);
   U96 : OAI21_X1 port map( B1 => n564, B2 => n495, A => n565, ZN => n561);
   U97 : OAI21_X1 port map( B1 => n496, B2 => A(30), A => B(30), ZN => n565);
   U98 : OAI21_X1 port map( B1 => n585, B2 => n506, A => n586, ZN => n582);
   U99 : INV_X1 port map( A => A(23), ZN => n506);
   U100 : OAI21_X1 port map( B1 => n507, B2 => A(23), A => B(23), ZN => n586);
   U101 : AOI21_X1 port map( B1 => n570, B2 => A(28), A => n499, ZN => n568);
   U102 : INV_X1 port map( A => n571, ZN => n499);
   U103 : OAI21_X1 port map( B1 => n570, B2 => A(28), A => B(28), ZN => n571);
   U104 : XNOR2_X1 port map( A => n570, B => n572, ZN => SUM(28));
   U105 : XNOR2_X1 port map( A => A(28), B => B(28), ZN => n572);
   U106 : AOI21_X1 port map( B1 => n558, B2 => n492, A => n559, ZN => n556);
   U107 : AOI21_X1 port map( B1 => n493, B2 => A(32), A => B(32), ZN => n559);
   U108 : AOI22_X1 port map( A1 => B(11), A2 => A(11), B1 => n522, B2 => n524, 
                           ZN => n523);
   U109 : XNOR2_X1 port map( A => n573, B => n575, ZN => SUM(27));
   U110 : XNOR2_X1 port map( A => B(27), B => n500, ZN => n575);
   U111 : OAI21_X1 port map( B1 => A(24), B2 => n582, A => n505, ZN => n579);
   U112 : INV_X1 port map( A => n583, ZN => n505);
   U113 : AOI21_X1 port map( B1 => n582, B2 => A(24), A => B(24), ZN => n583);
   U114 : OAI21_X1 port map( B1 => A(31), B2 => n561, A => n494, ZN => n558);
   U115 : INV_X1 port map( A => n562, ZN => n494);
   U116 : AOI21_X1 port map( B1 => n561, B2 => A(31), A => B(31), ZN => n562);
   U117 : OAI21_X1 port map( B1 => A(29), B2 => n498, A => n497, ZN => n564);
   U118 : INV_X1 port map( A => n567, ZN => n497);
   U119 : AOI21_X1 port map( B1 => n498, B2 => A(29), A => B(29), ZN => n567);
   U120 : INV_X1 port map( A => n568, ZN => n498);
   U121 : OAI21_X1 port map( B1 => A(22), B2 => n588, A => n508, ZN => n585);
   U122 : INV_X1 port map( A => n589, ZN => n508);
   U123 : AOI21_X1 port map( B1 => n588, B2 => A(22), A => B(22), ZN => n589);
   U124 : OAI21_X1 port map( B1 => A(20), B2 => n594, A => n511, ZN => n591);
   U125 : INV_X1 port map( A => n595, ZN => n511);
   U126 : AOI21_X1 port map( B1 => n594, B2 => A(20), A => B(20), ZN => n595);
   U127 : OAI21_X1 port map( B1 => A(42), B2 => n527, A => B(42), ZN => n528);
   U128 : INV_X1 port map( A => A(36), ZN => n487);
   U129 : INV_X1 port map( A => n523, ZN => n521);
   U130 : INV_X1 port map( A => A(30), ZN => n495);
   U131 : INV_X1 port map( A => n614, ZN => n522);
   U132 : AOI22_X1 port map( A1 => n615, A2 => carry_10_port, B1 => A(10), B2 
                           => B(10), ZN => n614);
   U133 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT42_DW01_add_0 is

   port( A, B : in std_logic_vector (41 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (41 downto 0);  CO : out std_logic);

end RCA_NBIT42_DW01_add_0;

architecture SYN_rpl of RCA_NBIT42_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_39_port, carry_38_port, carry_37_port, carry_36_port, 
      carry_35_port, carry_32_port, carry_31_port, carry_30_port, carry_29_port
      , carry_28_port, carry_26_port, carry_23_port, carry_22_port, n389, n390,
      n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n351, n352, n353, n354, 
      n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, 
      n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, 
      n379, n380, n381, n382, n383, n384, n385, n386, n387, n388 : std_logic;

begin
   
   U1_38 : FA_X1 port map( A => A(38), B => B(38), CI => carry_38_port, CO => 
                           carry_39_port, S => SUM(38));
   U1_37 : FA_X1 port map( A => A(37), B => B(37), CI => carry_37_port, CO => 
                           carry_38_port, S => SUM(37));
   U1_36 : FA_X1 port map( A => A(36), B => B(36), CI => carry_36_port, CO => 
                           carry_37_port, S => SUM(36));
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => carry_35_port, CO => 
                           carry_36_port, S => SUM(35));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => n360, CO => 
                           carry_22_port, S => SUM(21));
   U1_22 : FA_X1 port map( A => B(22), B => A(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => n470, CO => 
                           carry_26_port, S => SUM(25));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => n358, CO => 
                           carry_28_port, S => SUM(27));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U100 : XOR2_X1 port map( A => n378, B => n398, Z => SUM(9));
   U101 : XOR2_X1 port map( A => B(9), B => A(9), Z => n398);
   U102 : XOR2_X1 port map( A => n399, B => n400, Z => SUM(8));
   U103 : XOR2_X1 port map( A => B(8), B => A(8), Z => n400);
   U104 : XOR2_X1 port map( A => n380, B => n401, Z => SUM(7));
   U105 : XOR2_X1 port map( A => B(7), B => A(7), Z => n401);
   U106 : XOR2_X1 port map( A => n402, B => n403, Z => SUM(6));
   U107 : XOR2_X1 port map( A => B(6), B => A(6), Z => n403);
   U108 : XOR2_X1 port map( A => n383, B => n404, Z => SUM(5));
   U109 : XOR2_X1 port map( A => B(5), B => A(5), Z => n404);
   U110 : XOR2_X1 port map( A => n405, B => n406, Z => SUM(4));
   U111 : XOR2_X1 port map( A => B(4), B => A(4), Z => n406);
   U112 : XOR2_X1 port map( A => B(41), B => A(41), Z => n408);
   U113 : XOR2_X1 port map( A => n410, B => n411, Z => SUM(40));
   U114 : XOR2_X1 port map( A => B(40), B => A(40), Z => n411);
   U115 : XOR2_X1 port map( A => n386, B => n413, Z => SUM(3));
   U116 : XOR2_X1 port map( A => B(3), B => A(3), Z => n413);
   U117 : XOR2_X1 port map( A => A(39), B => n414, Z => SUM(39));
   U118 : XOR2_X1 port map( A => carry_39_port, B => B(39), Z => n414);
   U119 : XOR2_X1 port map( A => n356, B => n418, Z => SUM(33));
   U120 : XOR2_X1 port map( A => A(32), B => n420, Z => SUM(32));
   U121 : XOR2_X1 port map( A => carry_32_port, B => B(32), Z => n420);
   U122 : XOR2_X1 port map( A => n421, B => n422, Z => SUM(2));
   U123 : XOR2_X1 port map( A => B(2), B => A(2), Z => n422);
   U124 : XOR2_X1 port map( A => carry_26_port, B => n390, Z => SUM(26));
   U125 : XOR2_X1 port map( A => A(26), B => B(26), Z => n390);
   U126 : XOR2_X1 port map( A => n392, B => n391, Z => SUM(24));
   U127 : XOR2_X1 port map( A => n359, B => B(24), Z => n392);
   U128 : XOR2_X1 port map( A => carry_23_port, B => n423, Z => SUM(23));
   U129 : XOR2_X1 port map( A => A(23), B => B(23), Z => n423);
   U130 : XOR2_X1 port map( A => n427, B => n428, Z => SUM(1));
   U131 : XOR2_X1 port map( A => B(1), B => A(1), Z => n428);
   U132 : XOR2_X1 port map( A => n425, B => n429, Z => SUM(19));
   U133 : XOR2_X1 port map( A => n430, B => n432, Z => SUM(18));
   U134 : XOR2_X1 port map( A => B(18), B => A(18), Z => n432);
   U135 : XOR2_X1 port map( A => n367, B => n435, Z => SUM(17));
   U136 : XOR2_X1 port map( A => B(17), B => A(17), Z => n435);
   U137 : XOR2_X1 port map( A => n436, B => n438, Z => SUM(16));
   U138 : XOR2_X1 port map( A => B(16), B => A(16), Z => n438);
   U139 : XOR2_X1 port map( A => n370, B => n441, Z => SUM(15));
   U140 : XOR2_X1 port map( A => B(15), B => A(15), Z => n441);
   U141 : XOR2_X1 port map( A => n442, B => n444, Z => SUM(14));
   U142 : XOR2_X1 port map( A => B(14), B => A(14), Z => n444);
   U143 : XOR2_X1 port map( A => n372, B => n447, Z => SUM(13));
   U144 : XOR2_X1 port map( A => B(13), B => A(13), Z => n447);
   U145 : XOR2_X1 port map( A => n448, B => n450, Z => SUM(12));
   U146 : XOR2_X1 port map( A => B(12), B => A(12), Z => n450);
   U147 : XOR2_X1 port map( A => n375, B => n453, Z => SUM(11));
   U148 : XOR2_X1 port map( A => B(11), B => A(11), Z => n453);
   U149 : XOR2_X1 port map( A => n454, B => n456, Z => SUM(10));
   U150 : XOR2_X1 port map( A => B(10), B => A(10), Z => n456);
   U151 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : INV_X1 port map( A => A(34), ZN => n353);
   U2 : INV_X1 port map( A => n416, ZN => n356);
   U3 : INV_X1 port map( A => n439, ZN => n370);
   U4 : INV_X1 port map( A => n397, ZN => n354);
   U5 : INV_X1 port map( A => n457, ZN => n378);
   U6 : INV_X1 port map( A => n445, ZN => n372);
   U7 : INV_X1 port map( A => n433, ZN => n367);
   U8 : INV_X1 port map( A => n460, ZN => n380);
   U9 : INV_X1 port map( A => n451, ZN => n375);
   U10 : INV_X1 port map( A => n466, ZN => n386);
   U11 : INV_X1 port map( A => n463, ZN => n383);
   U12 : XNOR2_X1 port map( A => n407, B => n408, ZN => SUM(41));
   U13 : OAI22_X1 port map( A1 => n409, A2 => B(40), B1 => n410, B2 => A(40), 
                           ZN => n407);
   U14 : AND2_X1 port map( A1 => A(40), A2 => n410, ZN => n409);
   U15 : XNOR2_X1 port map( A => B(33), B => n355, ZN => n418);
   U16 : XNOR2_X1 port map( A => A(19), B => B(19), ZN => n429);
   U17 : AOI21_X1 port map( B1 => n425, B2 => n362, A => n426, ZN => n394);
   U18 : INV_X1 port map( A => A(19), ZN => n362);
   U19 : AOI21_X1 port map( B1 => n363, B2 => A(19), A => B(19), ZN => n426);
   U20 : INV_X1 port map( A => n425, ZN => n363);
   U21 : AOI22_X1 port map( A1 => n442, A2 => A(14), B1 => n443, B2 => B(14), 
                           ZN => n439);
   U22 : OR2_X1 port map( A1 => n442, A2 => A(14), ZN => n443);
   U23 : AOI21_X1 port map( B1 => n365, B2 => n433, A => n434, ZN => n430);
   U24 : INV_X1 port map( A => A(17), ZN => n365);
   U25 : AOI21_X1 port map( B1 => n367, B2 => A(17), A => B(17), ZN => n434);
   U26 : AOI21_X1 port map( B1 => n369, B2 => n439, A => n440, ZN => n436);
   U27 : INV_X1 port map( A => A(15), ZN => n369);
   U28 : AOI21_X1 port map( B1 => n370, B2 => A(15), A => B(15), ZN => n440);
   U29 : AOI21_X1 port map( B1 => n377, B2 => n457, A => n458, ZN => n454);
   U30 : INV_X1 port map( A => A(9), ZN => n377);
   U31 : AOI21_X1 port map( B1 => n378, B2 => A(9), A => B(9), ZN => n458);
   U32 : AOI21_X1 port map( B1 => n374, B2 => n451, A => n452, ZN => n448);
   U33 : INV_X1 port map( A => A(11), ZN => n374);
   U34 : AOI21_X1 port map( B1 => n375, B2 => A(11), A => B(11), ZN => n452);
   U35 : AOI21_X1 port map( B1 => n385, B2 => n466, A => n467, ZN => n405);
   U36 : INV_X1 port map( A => A(3), ZN => n385);
   U37 : AOI21_X1 port map( B1 => n386, B2 => A(3), A => B(3), ZN => n467);
   U38 : AOI21_X1 port map( B1 => n382, B2 => n463, A => n464, ZN => n402);
   U39 : INV_X1 port map( A => A(5), ZN => n382);
   U40 : AOI21_X1 port map( B1 => n383, B2 => A(5), A => B(5), ZN => n464);
   U41 : OAI21_X1 port map( B1 => B(32), B2 => A(32), A => n357, ZN => n416);
   U42 : INV_X1 port map( A => n419, ZN => n357);
   U43 : AOI21_X1 port map( B1 => A(32), B2 => B(32), A => carry_32_port, ZN =>
                           n419);
   U44 : XNOR2_X1 port map( A => n354, B => n415, ZN => SUM(34));
   U45 : XNOR2_X1 port map( A => B(34), B => n353, ZN => n415);
   U46 : XNOR2_X1 port map( A => n394, B => n424, ZN => SUM(20));
   U47 : XNOR2_X1 port map( A => A(20), B => B(20), ZN => n424);
   U48 : AOI22_X1 port map( A1 => n399, A2 => A(8), B1 => n459, B2 => B(8), ZN 
                           => n457);
   U49 : OR2_X1 port map( A1 => n399, A2 => A(8), ZN => n459);
   U50 : AOI22_X1 port map( A1 => B(23), A2 => A(23), B1 => n423, B2 => 
                           carry_23_port, ZN => n391);
   U51 : OAI21_X1 port map( B1 => A(18), B2 => n430, A => n364, ZN => n425);
   U52 : INV_X1 port map( A => n431, ZN => n364);
   U53 : AOI21_X1 port map( B1 => n430, B2 => A(18), A => B(18), ZN => n431);
   U54 : AOI21_X1 port map( B1 => n371, B2 => n445, A => n446, ZN => n442);
   U55 : INV_X1 port map( A => A(13), ZN => n371);
   U56 : AOI21_X1 port map( B1 => n372, B2 => A(13), A => B(13), ZN => n446);
   U57 : AOI21_X1 port map( B1 => n379, B2 => n460, A => n461, ZN => n399);
   U58 : INV_X1 port map( A => A(7), ZN => n379);
   U59 : AOI21_X1 port map( B1 => n380, B2 => A(7), A => B(7), ZN => n461);
   U60 : AOI22_X1 port map( A1 => n421, A2 => A(2), B1 => n468, B2 => B(2), ZN 
                           => n466);
   U61 : OR2_X1 port map( A1 => A(2), A2 => n421, ZN => n468);
   U62 : AOI21_X1 port map( B1 => n402, B2 => A(6), A => n381, ZN => n460);
   U63 : INV_X1 port map( A => n462, ZN => n381);
   U64 : OAI21_X1 port map( B1 => n402, B2 => A(6), A => B(6), ZN => n462);
   U65 : AOI21_X1 port map( B1 => n448, B2 => A(12), A => n373, ZN => n445);
   U66 : INV_X1 port map( A => n449, ZN => n373);
   U67 : OAI21_X1 port map( B1 => n448, B2 => A(12), A => B(12), ZN => n449);
   U68 : AOI21_X1 port map( B1 => n454, B2 => A(10), A => n376, ZN => n451);
   U69 : INV_X1 port map( A => n455, ZN => n376);
   U70 : OAI21_X1 port map( B1 => n454, B2 => A(10), A => B(10), ZN => n455);
   U71 : AOI21_X1 port map( B1 => n405, B2 => A(4), A => n384, ZN => n463);
   U72 : INV_X1 port map( A => n465, ZN => n384);
   U73 : OAI21_X1 port map( B1 => n405, B2 => A(4), A => B(4), ZN => n465);
   U74 : AOI21_X1 port map( B1 => n436, B2 => A(16), A => n368, ZN => n433);
   U75 : INV_X1 port map( A => n437, ZN => n368);
   U76 : OAI21_X1 port map( B1 => n436, B2 => A(16), A => B(16), ZN => n437);
   U77 : OAI21_X1 port map( B1 => n352, B2 => n351, A => n412, ZN => n410);
   U78 : INV_X1 port map( A => B(39), ZN => n351);
   U79 : INV_X1 port map( A => A(39), ZN => n352);
   U80 : OAI21_X1 port map( B1 => A(39), B2 => B(39), A => carry_39_port, ZN =>
                           n412);
   U81 : OAI21_X1 port map( B1 => n416, B2 => n355, A => n417, ZN => n397);
   U82 : OAI21_X1 port map( B1 => n356, B2 => A(33), A => B(33), ZN => n417);
   U83 : AOI21_X1 port map( B1 => n394, B2 => A(20), A => n361, ZN => n393);
   U84 : INV_X1 port map( A => n395, ZN => n361);
   U85 : OAI21_X1 port map( B1 => n394, B2 => A(20), A => B(20), ZN => n395);
   U86 : OAI22_X1 port map( A1 => n366, A2 => n359, B1 => n391, B2 => n392, ZN 
                           => n470);
   U87 : INV_X1 port map( A => B(24), ZN => n366);
   U88 : INV_X1 port map( A => n393, ZN => n360);
   U89 : INV_X1 port map( A => n389, ZN => n358);
   U90 : AOI22_X1 port map( A1 => B(26), A2 => A(26), B1 => n390, B2 => 
                           carry_26_port, ZN => n389);
   U91 : OAI21_X1 port map( B1 => n354, B2 => n353, A => n396, ZN => 
                           carry_35_port);
   U92 : OAI21_X1 port map( B1 => A(34), B2 => n397, A => B(34), ZN => n396);
   U93 : INV_X1 port map( A => A(33), ZN => n355);
   U94 : INV_X1 port map( A => A(24), ZN => n359);
   U95 : OAI21_X1 port map( B1 => n387, B2 => n388, A => n469, ZN => n421);
   U96 : INV_X1 port map( A => B(1), ZN => n388);
   U97 : INV_X1 port map( A => A(1), ZN => n387);
   U98 : OAI211_X1 port map( C1 => A(1), C2 => B(1), A => A(0), B => B(0), ZN 
                           => n469);
   U99 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n427);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT40_DW01_add_0 is

   port( A, B : in std_logic_vector (39 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (39 downto 0);  CO : out std_logic);

end RCA_NBIT40_DW01_add_0;

architecture SYN_rpl of RCA_NBIT40_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_39_port, carry_38_port, carry_37_port, carry_36_port, 
      carry_34_port, carry_33_port, carry_30_port, carry_29_port, carry_28_port
      , carry_6_port, carry_5_port, carry_4_port, carry_3_port, carry_2_port, 
      n1, n268, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, 
      n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, 
      n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, 
      n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, 
      n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, 
      n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, 
      n428, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, 
      n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, 
      n349, n350, n351, n352, n353, n354, n355, n356, n357 : std_logic;

begin
   
   U1_38 : FA_X1 port map( A => A(38), B => B(38), CI => carry_38_port, CO => 
                           carry_39_port, S => SUM(38));
   U1_37 : FA_X1 port map( A => A(37), B => B(37), CI => carry_37_port, CO => 
                           carry_38_port, S => SUM(37));
   U1_36 : FA_X1 port map( A => A(36), B => B(36), CI => carry_36_port, CO => 
                           carry_37_port, S => SUM(36));
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => n326, CO => 
                           carry_36_port, S => SUM(35));
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1_32 : FA_X1 port map( A => B(32), B => n268, CI => A(32), CO => 
                           carry_33_port, S => SUM(32));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => n328, CO => 
                           carry_28_port, S => SUM(27));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U86 : XOR2_X1 port map( A => n353, B => n365, Z => SUM(9));
   U87 : XOR2_X1 port map( A => B(9), B => A(9), Z => n365);
   U88 : XOR2_X1 port map( A => n366, B => n367, Z => SUM(8));
   U89 : XOR2_X1 port map( A => B(8), B => A(8), Z => n367);
   U90 : XOR2_X1 port map( A => n356, B => n368, Z => SUM(7));
   U91 : XOR2_X1 port map( A => A(6), B => n369, Z => SUM(6));
   U92 : XOR2_X1 port map( A => carry_6_port, B => B(6), Z => n369);
   U93 : XOR2_X1 port map( A => A(39), B => n370, Z => SUM(39));
   U94 : XOR2_X1 port map( A => carry_39_port, B => B(39), Z => n370);
   U95 : XOR2_X1 port map( A => carry_34_port, B => n361, Z => SUM(34));
   U96 : XOR2_X1 port map( A => A(34), B => B(34), Z => n361);
   U97 : XOR2_X1 port map( A => n359, B => n358, Z => SUM(31));
   U98 : XOR2_X1 port map( A => n327, B => B(31), Z => n359);
   U99 : XOR2_X1 port map( A => carry_30_port, B => n371, Z => SUM(30));
   U100 : XOR2_X1 port map( A => A(30), B => B(30), Z => n371);
   U101 : XOR2_X1 port map( A => B(26), B => A(26), Z => n372);
   U102 : XOR2_X1 port map( A => n376, B => n377, Z => SUM(25));
   U103 : XOR2_X1 port map( A => B(25), B => A(25), Z => n377);
   U104 : XOR2_X1 port map( A => n381, B => n382, Z => SUM(24));
   U105 : XOR2_X1 port map( A => B(24), B => A(24), Z => n382);
   U106 : XOR2_X1 port map( A => n385, B => n387, Z => SUM(22));
   U107 : XOR2_X1 port map( A => B(22), B => A(22), Z => n387);
   U108 : XOR2_X1 port map( A => n390, B => n388, Z => SUM(21));
   U109 : XOR2_X1 port map( A => n333, B => B(21), Z => n390);
   U110 : XOR2_X1 port map( A => n391, B => n392, Z => SUM(20));
   U111 : XOR2_X1 port map( A => A(20), B => B(20), Z => n392);
   U112 : XOR2_X1 port map( A => n336, B => n395, Z => SUM(19));
   U113 : XOR2_X1 port map( A => B(19), B => A(19), Z => n395);
   U114 : XOR2_X1 port map( A => n397, B => n398, Z => SUM(18));
   U115 : XOR2_X1 port map( A => n399, B => n401, Z => SUM(17));
   U116 : XOR2_X1 port map( A => B(17), B => A(17), Z => n401);
   U117 : XOR2_X1 port map( A => n343, B => n404, Z => SUM(16));
   U118 : XOR2_X1 port map( A => B(16), B => A(16), Z => n404);
   U119 : XOR2_X1 port map( A => n344, B => n406, Z => SUM(15));
   U120 : XOR2_X1 port map( A => B(15), B => A(15), Z => n406);
   U121 : XOR2_X1 port map( A => n408, B => n410, Z => SUM(14));
   U122 : XOR2_X1 port map( A => B(14), B => A(14), Z => n410);
   U123 : XOR2_X1 port map( A => n347, B => n413, Z => SUM(13));
   U124 : XOR2_X1 port map( A => B(13), B => A(13), Z => n413);
   U125 : XOR2_X1 port map( A => n414, B => n416, Z => SUM(12));
   U126 : XOR2_X1 port map( A => B(12), B => A(12), Z => n416);
   U127 : XOR2_X1 port map( A => n350, B => n419, Z => SUM(11));
   U128 : XOR2_X1 port map( A => B(11), B => A(11), Z => n419);
   U129 : XOR2_X1 port map( A => n420, B => n422, Z => SUM(10));
   U130 : XOR2_X1 port map( A => A(10), B => B(10), Z => n422);
   U131 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : XNOR2_X1 port map( A => n380, B => n384, ZN => SUM(23));
   U2 : XNOR2_X1 port map( A => n338, B => A(23), ZN => n384);
   U3 : NOR2_X1 port map( A1 => n381, A2 => A(24), ZN => n374);
   U4 : NOR2_X1 port map( A1 => n374, A2 => n375, ZN => n376);
   U5 : INV_X1 port map( A => A(7), ZN => n355);
   U6 : INV_X1 port map( A => n426, ZN => n356);
   U7 : INV_X1 port map( A => n417, ZN => n350);
   U8 : INV_X1 port map( A => n402, ZN => n343);
   U9 : INV_X1 port map( A => n423, ZN => n353);
   U10 : INV_X1 port map( A => n411, ZN => n347);
   U11 : INV_X1 port map( A => n393, ZN => n336);
   U12 : XNOR2_X1 port map( A => B(7), B => n355, ZN => n368);
   U13 : XNOR2_X1 port map( A => A(18), B => B(18), ZN => n398);
   U14 : AOI22_X1 port map( A1 => n385, A2 => A(22), B1 => n386, B2 => B(22), 
                           ZN => n380);
   U15 : OR2_X1 port map( A1 => A(22), A2 => n385, ZN => n386);
   U16 : OAI22_X1 port map( A1 => n388, A2 => n333, B1 => n389, B2 => n342, ZN 
                           => n385);
   U17 : AND2_X1 port map( A1 => n333, A2 => n388, ZN => n389);
   U18 : INV_X1 port map( A => B(21), ZN => n342);
   U19 : AOI21_X1 port map( B1 => A(25), B2 => B(25), A => n373, ZN => n364);
   U20 : AOI211_X1 port map( C1 => n331, C2 => n334, A => n374, B => n375, ZN 
                           => n373);
   U21 : INV_X1 port map( A => A(25), ZN => n331);
   U22 : INV_X1 port map( A => B(25), ZN => n334);
   U23 : AOI22_X1 port map( A1 => B(20), A2 => A(20), B1 => n391, B2 => n392, 
                           ZN => n388);
   U24 : AOI22_X1 port map( A1 => n344, A2 => A(15), B1 => n405, B2 => B(15), 
                           ZN => n402);
   U25 : OR2_X1 port map( A1 => n344, A2 => A(15), ZN => n405);
   U26 : AOI21_X1 port map( B1 => n341, B2 => n402, A => n403, ZN => n399);
   U27 : INV_X1 port map( A => A(16), ZN => n341);
   U28 : AOI21_X1 port map( B1 => n343, B2 => A(16), A => B(16), ZN => n403);
   U29 : OAI21_X1 port map( B1 => B(6), B2 => A(6), A => n357, ZN => n426);
   U30 : INV_X1 port map( A => n428, ZN => n357);
   U31 : AOI21_X1 port map( B1 => A(6), B2 => B(6), A => carry_6_port, ZN => 
                           n428);
   U32 : OAI21_X1 port map( B1 => B(10), B2 => n420, A => n351, ZN => n417);
   U33 : INV_X1 port map( A => n421, ZN => n351);
   U34 : AOI21_X1 port map( B1 => n420, B2 => B(10), A => A(10), ZN => n421);
   U35 : OAI21_X1 port map( B1 => n426, B2 => n355, A => n427, ZN => n366);
   U36 : OAI21_X1 port map( B1 => n356, B2 => A(7), A => B(7), ZN => n427);
   U37 : OAI21_X1 port map( B1 => n417, B2 => n349, A => n418, ZN => n414);
   U38 : INV_X1 port map( A => A(11), ZN => n349);
   U39 : OAI21_X1 port map( B1 => n350, B2 => A(11), A => B(11), ZN => n418);
   U40 : AOI21_X1 port map( B1 => A(24), B2 => n378, A => B(24), ZN => n375);
   U41 : AOI22_X1 port map( A1 => n338, A2 => n332, B1 => n379, B2 => n380, ZN 
                           => n378);
   U42 : INV_X1 port map( A => A(23), ZN => n332);
   U43 : AOI22_X1 port map( A1 => B(30), A2 => A(30), B1 => n371, B2 => 
                           carry_30_port, ZN => n358);
   U44 : OAI21_X1 port map( B1 => n423, B2 => n352, A => n424, ZN => n420);
   U45 : INV_X1 port map( A => A(9), ZN => n352);
   U46 : OAI21_X1 port map( B1 => n353, B2 => A(9), A => B(9), ZN => n424);
   U47 : OAI21_X1 port map( B1 => n411, B2 => n346, A => n412, ZN => n408);
   U48 : INV_X1 port map( A => A(13), ZN => n346);
   U49 : OAI21_X1 port map( B1 => n347, B2 => A(13), A => B(13), ZN => n412);
   U50 : AOI21_X1 port map( B1 => n339, B2 => A(18), A => n337, ZN => n393);
   U51 : INV_X1 port map( A => n396, ZN => n337);
   U52 : OAI21_X1 port map( B1 => n339, B2 => A(18), A => B(18), ZN => n396);
   U53 : INV_X1 port map( A => n397, ZN => n339);
   U54 : AOI22_X1 port map( A1 => n330, A2 => A(26), B1 => n363, B2 => B(26), 
                           ZN => n362);
   U55 : OR2_X1 port map( A1 => A(26), A2 => n330, ZN => n363);
   U56 : INV_X1 port map( A => n364, ZN => n330);
   U57 : OAI21_X1 port map( B1 => A(12), B2 => n414, A => n348, ZN => n411);
   U58 : INV_X1 port map( A => n415, ZN => n348);
   U59 : AOI21_X1 port map( B1 => n414, B2 => A(12), A => B(12), ZN => n415);
   U60 : OAI21_X1 port map( B1 => A(8), B2 => n366, A => n354, ZN => n423);
   U61 : INV_X1 port map( A => n425, ZN => n354);
   U62 : AOI21_X1 port map( B1 => n366, B2 => A(8), A => B(8), ZN => n425);
   U63 : XNOR2_X1 port map( A => n364, B => n372, ZN => SUM(26));
   U64 : OAI21_X1 port map( B1 => n380, B2 => n383, A => n379, ZN => n381);
   U65 : NOR2_X1 port map( A1 => A(23), A2 => B(23), ZN => n383);
   U66 : NAND2_X1 port map( A1 => B(23), A2 => A(23), ZN => n379);
   U67 : OAI21_X1 port map( B1 => n399, B2 => A(17), A => n340, ZN => n397);
   U68 : INV_X1 port map( A => n400, ZN => n340);
   U69 : AOI21_X1 port map( B1 => n399, B2 => A(17), A => B(17), ZN => n400);
   U70 : OAI21_X1 port map( B1 => n393, B2 => n335, A => n394, ZN => n391);
   U71 : INV_X1 port map( A => A(19), ZN => n335);
   U72 : OAI21_X1 port map( B1 => A(19), B2 => n336, A => B(19), ZN => n394);
   U73 : INV_X1 port map( A => B(23), ZN => n338);
   U74 : INV_X1 port map( A => n362, ZN => n328);
   U75 : OAI22_X1 port map( A1 => n329, A2 => n327, B1 => n358, B2 => n359, ZN 
                           => n268);
   U76 : INV_X1 port map( A => B(31), ZN => n329);
   U77 : INV_X1 port map( A => n360, ZN => n326);
   U78 : AOI22_X1 port map( A1 => B(34), A2 => A(34), B1 => n361, B2 => 
                           carry_34_port, ZN => n360);
   U79 : INV_X1 port map( A => n407, ZN => n344);
   U80 : OAI21_X1 port map( B1 => A(14), B2 => n408, A => n345, ZN => n407);
   U81 : INV_X1 port map( A => n409, ZN => n345);
   U82 : AOI21_X1 port map( B1 => n408, B2 => A(14), A => B(14), ZN => n409);
   U83 : INV_X1 port map( A => A(21), ZN => n333);
   U84 : INV_X1 port map( A => A(31), ZN => n327);
   U85 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT38_DW01_add_0 is

   port( A, B : in std_logic_vector (37 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (37 downto 0);  CO : out std_logic);

end RCA_NBIT38_DW01_add_0;

architecture SYN_rpl of RCA_NBIT38_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_36_port, carry_34_port, carry_33_port, carry_4_port, 
      carry_3_port, carry_2_port, n1, n435, n436, n437, n438, n439, n440, n441,
      n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, 
      n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, 
      n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, 
      n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, 
      n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, 
      n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, 
      n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, 
      n526, n527, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434 : std_logic;

begin
   
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => n393, CO => 
                           carry_36_port, S => SUM(35));
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => n394, CO => 
                           carry_33_port, S => SUM(32));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U131 : XOR2_X1 port map( A => B(9), B => A(9), Z => n441);
   U132 : XOR2_X1 port map( A => n442, B => n443, Z => SUM(8));
   U133 : XOR2_X1 port map( A => B(8), B => A(8), Z => n443);
   U134 : XOR2_X1 port map( A => n446, B => n447, Z => SUM(6));
   U135 : XOR2_X1 port map( A => B(6), B => A(6), Z => n447);
   U136 : XOR2_X1 port map( A => B(5), B => A(5), Z => n449);
   U137 : XOR2_X1 port map( A => A(4), B => n450, Z => SUM(4));
   U138 : XOR2_X1 port map( A => carry_4_port, B => B(4), Z => n450);
   U139 : XOR2_X1 port map( A => n451, B => n452, Z => SUM(37));
   U140 : XOR2_X1 port map( A => carry_36_port, B => n453, Z => SUM(36));
   U141 : XOR2_X1 port map( A => A(36), B => B(36), Z => n453);
   U142 : XOR2_X1 port map( A => carry_34_port, B => n436, Z => SUM(34));
   U143 : XOR2_X1 port map( A => A(34), B => B(34), Z => n436);
   U144 : XOR2_X1 port map( A => B(31), B => A(31), Z => n454);
   U145 : XOR2_X1 port map( A => B(30), B => A(30), Z => n457);
   U146 : XOR2_X1 port map( A => n458, B => n460, Z => SUM(29));
   U147 : XOR2_X1 port map( A => B(29), B => A(29), Z => n460);
   U148 : XOR2_X1 port map( A => B(27), B => A(27), Z => n466);
   U149 : XOR2_X1 port map( A => n467, B => n469, Z => SUM(26));
   U150 : XOR2_X1 port map( A => B(26), B => A(26), Z => n469);
   U151 : XOR2_X1 port map( A => n403, B => n472, Z => SUM(25));
   U152 : XOR2_X1 port map( A => B(25), B => A(25), Z => n472);
   U153 : XOR2_X1 port map( A => n479, B => n481, Z => SUM(22));
   U154 : XOR2_X1 port map( A => B(22), B => A(22), Z => n481);
   U155 : XOR2_X1 port map( A => n489, B => n491, Z => SUM(19));
   U156 : XOR2_X1 port map( A => B(19), B => A(19), Z => n491);
   U157 : XOR2_X1 port map( A => n492, B => n494, Z => SUM(18));
   U158 : NAND3_X1 port map( A1 => n499, A2 => n413, A3 => n498, ZN => n496);
   U159 : XOR2_X1 port map( A => n500, B => n501, Z => SUM(16));
   U160 : XOR2_X1 port map( A => B(16), B => A(16), Z => n501);
   U161 : XOR2_X1 port map( A => n502, B => n504, Z => SUM(15));
   U162 : NAND3_X1 port map( A1 => A(14), A2 => n424, A3 => n507, ZN => n509);
   U163 : XOR2_X1 port map( A => B(13), B => A(13), Z => n512);
   U164 : XOR2_X1 port map( A => n513, B => n515, Z => SUM(12));
   U165 : XOR2_X1 port map( A => B(12), B => A(12), Z => n515);
   U166 : XOR2_X1 port map( A => n519, B => n521, Z => SUM(10));
   U167 : XOR2_X1 port map( A => B(10), B => A(10), Z => n521);
   U168 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : OR2_X1 port map( A1 => A(31), A2 => n395, ZN => n438);
   U2 : AOI21_X1 port map( B1 => n498, B2 => n499, A => n413, ZN => n495);
   U3 : NAND2_X1 port map( A1 => n409, A2 => n487, ZN => n486);
   U4 : INV_X1 port map( A => A(23), ZN => n405);
   U5 : INV_X1 port map( A => A(28), ZN => n397);
   U6 : INV_X1 port map( A => A(11), ZN => n423);
   U7 : NAND2_X1 port map( A1 => A(16), A2 => n500, ZN => n498);
   U8 : INV_X1 port map( A => A(7), ZN => n429);
   U9 : INV_X1 port map( A => A(14), ZN => n417);
   U10 : INV_X1 port map( A => n439, ZN => n395);
   U11 : INV_X1 port map( A => n482, ZN => n408);
   U12 : INV_X1 port map( A => n470, ZN => n403);
   U13 : XNOR2_X1 port map( A => A(18), B => B(18), ZN => n494);
   U14 : XNOR2_X1 port map( A => B(37), B => A(37), ZN => n451);
   U15 : AOI22_X1 port map( A1 => carry_36_port, A2 => n453, B1 => A(36), B2 =>
                           B(36), ZN => n452);
   U16 : XNOR2_X1 port map( A => A(15), B => B(15), ZN => n504);
   U17 : OAI221_X1 port map( B1 => n508, B2 => n424, C1 => n507, C2 => n506, A 
                           => n509, ZN => SUM(14));
   U18 : XNOR2_X1 port map( A => n507, B => A(14), ZN => n508);
   U19 : XNOR2_X1 port map( A => n476, B => n478, ZN => SUM(23));
   U20 : XNOR2_X1 port map( A => B(23), B => n405, ZN => n478);
   U21 : OAI22_X1 port map( A1 => n502, A2 => n415, B1 => n503, B2 => n422, ZN 
                           => n500);
   U22 : AND2_X1 port map( A1 => n502, A2 => n415, ZN => n503);
   U23 : INV_X1 port map( A => A(15), ZN => n415);
   U24 : INV_X1 port map( A => B(15), ZN => n422);
   U25 : AOI22_X1 port map( A1 => n479, A2 => A(22), B1 => n480, B2 => B(22), 
                           ZN => n476);
   U26 : OR2_X1 port map( A1 => n479, A2 => A(22), ZN => n480);
   U27 : OAI22_X1 port map( A1 => n492, A2 => n411, B1 => n493, B2 => n416, ZN 
                           => n489);
   U28 : AND2_X1 port map( A1 => n492, A2 => n411, ZN => n493);
   U29 : INV_X1 port map( A => A(18), ZN => n411);
   U30 : INV_X1 port map( A => B(18), ZN => n416);
   U31 : AOI22_X1 port map( A1 => n442, A2 => A(8), B1 => n523, B2 => B(8), ZN 
                           => n440);
   U32 : OR2_X1 port map( A1 => A(8), A2 => n442, ZN => n523);
   U33 : AOI21_X1 port map( B1 => n420, B2 => A(13), A => n419, ZN => n507);
   U34 : INV_X1 port map( A => n510, ZN => n419);
   U35 : OAI21_X1 port map( B1 => n420, B2 => A(13), A => B(13), ZN => n510);
   U36 : INV_X1 port map( A => n511, ZN => n420);
   U37 : OAI21_X1 port map( B1 => B(4), B2 => A(4), A => n434, ZN => n448);
   U38 : INV_X1 port map( A => n527, ZN => n434);
   U39 : AOI21_X1 port map( B1 => A(4), B2 => B(4), A => carry_4_port, ZN => 
                           n527);
   U40 : AOI21_X1 port map( B1 => n405, B2 => n476, A => n477, ZN => n473);
   U41 : AOI21_X1 port map( B1 => n406, B2 => A(23), A => B(23), ZN => n477);
   U42 : INV_X1 port map( A => n476, ZN => n406);
   U43 : XNOR2_X1 port map( A => B(17), B => n497, ZN => SUM(17));
   U44 : NAND2_X1 port map( A1 => n496, A2 => n412, ZN => n497);
   U45 : INV_X1 port map( A => n495, ZN => n412);
   U46 : AOI22_X1 port map( A1 => n458, A2 => A(29), B1 => n459, B2 => B(29), 
                           ZN => n456);
   U47 : OR2_X1 port map( A1 => A(29), A2 => n458, ZN => n459);
   U48 : AOI22_X1 port map( A1 => n396, A2 => A(30), B1 => n455, B2 => B(30), 
                           ZN => n439);
   U49 : OR2_X1 port map( A1 => A(30), A2 => n396, ZN => n455);
   U50 : INV_X1 port map( A => n456, ZN => n396);
   U51 : OAI21_X1 port map( B1 => A(6), B2 => n446, A => n431, ZN => n444);
   U52 : INV_X1 port map( A => n525, ZN => n431);
   U53 : AOI21_X1 port map( B1 => n446, B2 => A(6), A => B(6), ZN => n525);
   U54 : OAI21_X1 port map( B1 => A(27), B2 => n400, A => n399, ZN => n461);
   U55 : INV_X1 port map( A => n464, ZN => n399);
   U56 : AOI21_X1 port map( B1 => n400, B2 => A(27), A => B(27), ZN => n464);
   U57 : INV_X1 port map( A => n465, ZN => n400);
   U58 : OAI21_X1 port map( B1 => A(10), B2 => n519, A => n426, ZN => n516);
   U59 : INV_X1 port map( A => n520, ZN => n426);
   U60 : AOI21_X1 port map( B1 => n519, B2 => A(10), A => B(10), ZN => n520);
   U61 : AOI21_X1 port map( B1 => n402, B2 => n470, A => n471, ZN => n467);
   U62 : INV_X1 port map( A => A(25), ZN => n402);
   U63 : AOI21_X1 port map( B1 => n403, B2 => A(25), A => B(25), ZN => n471);
   U64 : OAI21_X1 port map( B1 => B(17), B2 => n495, A => n496, ZN => n492);
   U65 : OAI21_X1 port map( B1 => A(19), B2 => n489, A => n410, ZN => n487);
   U66 : INV_X1 port map( A => n490, ZN => n410);
   U67 : AOI21_X1 port map( B1 => n489, B2 => A(19), A => B(19), ZN => n490);
   U68 : XNOR2_X1 port map( A => n440, B => n441, ZN => SUM(9));
   U69 : XNOR2_X1 port map( A => n516, B => n518, ZN => SUM(11));
   U70 : XNOR2_X1 port map( A => B(11), B => n423, ZN => n518);
   U71 : XNOR2_X1 port map( A => n511, B => n512, ZN => SUM(13));
   U72 : XNOR2_X1 port map( A => n473, B => n475, ZN => SUM(24));
   U73 : XNOR2_X1 port map( A => A(24), B => B(24), ZN => n475);
   U74 : OAI21_X1 port map( B1 => n448, B2 => n432, A => n526, ZN => n446);
   U75 : INV_X1 port map( A => A(5), ZN => n432);
   U76 : OAI21_X1 port map( B1 => n433, B2 => A(5), A => B(5), ZN => n526);
   U77 : INV_X1 port map( A => n448, ZN => n433);
   U78 : OAI21_X1 port map( B1 => n440, B2 => n427, A => n522, ZN => n519);
   U79 : INV_X1 port map( A => A(9), ZN => n427);
   U80 : OAI21_X1 port map( B1 => A(9), B2 => n428, A => B(9), ZN => n522);
   U81 : INV_X1 port map( A => n440, ZN => n428);
   U82 : OAI21_X1 port map( B1 => n516, B2 => n423, A => n517, ZN => n513);
   U83 : OAI21_X1 port map( B1 => n425, B2 => A(11), A => B(11), ZN => n517);
   U84 : INV_X1 port map( A => n516, ZN => n425);
   U85 : XNOR2_X1 port map( A => B(20), B => n488, ZN => SUM(20));
   U86 : OAI21_X1 port map( B1 => n487, B2 => n409, A => n486, ZN => n488);
   U87 : AOI21_X1 port map( B1 => n407, B2 => n482, A => n483, ZN => n479);
   U88 : INV_X1 port map( A => A(21), ZN => n407);
   U89 : AOI21_X1 port map( B1 => n408, B2 => A(21), A => B(21), ZN => n483);
   U90 : AOI21_X1 port map( B1 => n467, B2 => A(26), A => n401, ZN => n465);
   U91 : INV_X1 port map( A => n468, ZN => n401);
   U92 : OAI21_X1 port map( B1 => n467, B2 => A(26), A => B(26), ZN => n468);
   U93 : AOI21_X1 port map( B1 => n473, B2 => A(24), A => n404, ZN => n470);
   U94 : INV_X1 port map( A => n474, ZN => n404);
   U95 : OAI21_X1 port map( B1 => n473, B2 => A(24), A => B(24), ZN => n474);
   U96 : OAI21_X1 port map( B1 => n444, B2 => n429, A => n524, ZN => n442);
   U97 : OAI21_X1 port map( B1 => n430, B2 => A(7), A => B(7), ZN => n524);
   U98 : INV_X1 port map( A => n444, ZN => n430);
   U99 : OAI21_X1 port map( B1 => n461, B2 => n397, A => n462, ZN => n458);
   U100 : OAI21_X1 port map( B1 => n398, B2 => A(28), A => B(28), ZN => n462);
   U101 : INV_X1 port map( A => n461, ZN => n398);
   U102 : OAI21_X1 port map( B1 => n505, B2 => n418, A => n506, ZN => n502);
   U103 : INV_X1 port map( A => n507, ZN => n418);
   U104 : NOR2_X1 port map( A1 => n417, A2 => n424, ZN => n505);
   U105 : OAI21_X1 port map( B1 => A(12), B2 => n513, A => n421, ZN => n511);
   U106 : INV_X1 port map( A => n514, ZN => n421);
   U107 : AOI21_X1 port map( B1 => n513, B2 => A(12), A => B(12), ZN => n514);
   U108 : XNOR2_X1 port map( A => n444, B => n445, ZN => SUM(7));
   U109 : XNOR2_X1 port map( A => B(7), B => n429, ZN => n445);
   U110 : XNOR2_X1 port map( A => n456, B => n457, ZN => SUM(30));
   U111 : OAI21_X1 port map( B1 => A(16), B2 => n500, A => B(16), ZN => n499);
   U112 : INV_X1 port map( A => n435, ZN => n393);
   U113 : AOI22_X1 port map( A1 => B(34), A2 => A(34), B1 => n436, B2 => 
                           carry_34_port, ZN => n435);
   U114 : INV_X1 port map( A => A(20), ZN => n409);
   U115 : XNOR2_X1 port map( A => n465, B => n466, ZN => SUM(27));
   U116 : XNOR2_X1 port map( A => n461, B => n463, ZN => SUM(28));
   U117 : XNOR2_X1 port map( A => B(28), B => n397, ZN => n463);
   U118 : INV_X1 port map( A => n437, ZN => n394);
   U119 : AOI22_X1 port map( A1 => n395, A2 => A(31), B1 => n438, B2 => B(31), 
                           ZN => n437);
   U120 : NAND2_X1 port map( A1 => n417, A2 => n424, ZN => n506);
   U121 : NAND2_X1 port map( A1 => n485, A2 => n486, ZN => n482);
   U122 : OAI21_X1 port map( B1 => n487, B2 => n409, A => n414, ZN => n485);
   U123 : INV_X1 port map( A => B(20), ZN => n414);
   U124 : XNOR2_X1 port map( A => n408, B => n484, ZN => SUM(21));
   U125 : XNOR2_X1 port map( A => A(21), B => B(21), ZN => n484);
   U126 : XNOR2_X1 port map( A => n439, B => n454, ZN => SUM(31));
   U127 : INV_X1 port map( A => A(17), ZN => n413);
   U128 : INV_X1 port map( A => B(14), ZN => n424);
   U129 : XNOR2_X1 port map( A => n448, B => n449, ZN => SUM(5));
   U130 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT36_DW01_add_0 is

   port( A, B : in std_logic_vector (35 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (35 downto 0);  CO : out std_logic);

end RCA_NBIT36_DW01_add_0;

architecture SYN_rpl of RCA_NBIT36_DW01_add_0 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_33_port, carry_2_port, n1, n446, n447, n448, n449, n450, n451, 
      n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, 
      n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, 
      n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, 
      n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, 
      n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, 
      n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, 
      n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, 
      n536, n537, n538, n539, n403, n404, n405, n406, n407, n408, n409, n410, 
      n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, 
      n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, 
      n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n_1064 
      : std_logic;

begin
   
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => n403, CO => n_1064, S 
                           => SUM(35));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => n405, CO => 
                           carry_33_port, S => SUM(32));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n1, CO => carry_2_port, S
                           => SUM(1));
   U140 : XOR2_X1 port map( A => n453, B => n454, Z => SUM(8));
   U141 : XOR2_X1 port map( A => B(8), B => A(8), Z => n454);
   U142 : XOR2_X1 port map( A => n456, B => n457, Z => SUM(6));
   U143 : XOR2_X1 port map( A => B(6), B => A(6), Z => n457);
   U144 : XOR2_X1 port map( A => n459, B => n460, Z => SUM(4));
   U145 : XOR2_X1 port map( A => B(4), B => A(4), Z => n460);
   U146 : XOR2_X1 port map( A => A(34), B => B(34), Z => n450);
   U147 : XOR2_X1 port map( A => carry_33_port, B => n463, Z => SUM(33));
   U148 : XOR2_X1 port map( A => A(33), B => B(33), Z => n463);
   U149 : XOR2_X1 port map( A => n447, B => n448, Z => SUM(31));
   U150 : XOR2_X1 port map( A => A(31), B => B(31), Z => n448);
   U151 : XOR2_X1 port map( A => B(30), B => A(30), Z => n466);
   U152 : XOR2_X1 port map( A => A(2), B => n469, Z => SUM(2));
   U153 : XOR2_X1 port map( A => carry_2_port, B => B(2), Z => n469);
   U154 : XOR2_X1 port map( A => B(29), B => A(29), Z => n470);
   U155 : XOR2_X1 port map( A => B(28), B => A(28), Z => n473);
   U156 : XOR2_X1 port map( A => n474, B => n476, Z => SUM(27));
   U157 : XOR2_X1 port map( A => B(27), B => A(27), Z => n476);
   U158 : XOR2_X1 port map( A => n480, B => n482, Z => SUM(25));
   U159 : XOR2_X1 port map( A => B(25), B => A(25), Z => n482);
   U160 : XOR2_X1 port map( A => n486, B => n488, Z => SUM(23));
   U161 : XOR2_X1 port map( A => B(23), B => A(23), Z => n488);
   U162 : XOR2_X1 port map( A => n419, B => B(20), Z => n497);
   U163 : XOR2_X1 port map( A => n422, B => B(18), Z => n503);
   U164 : XOR2_X1 port map( A => n425, B => B(16), Z => n509);
   U165 : XOR2_X1 port map( A => n428, B => B(14), Z => n515);
   U166 : XOR2_X1 port map( A => n517, B => n518, Z => SUM(13));
   U167 : XOR2_X1 port map( A => B(13), B => A(13), Z => n518);
   U168 : XOR2_X1 port map( A => B(12), B => A(12), Z => n521);
   U169 : XOR2_X1 port map( A => B(11), B => A(11), Z => n524);
   U170 : XOR2_X1 port map( A => n525, B => n529, Z => SUM(10));
   U171 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U1 : XNOR2_X1 port map( A => n451, B => n450, ZN => SUM(34));
   U2 : INV_X1 port map( A => n527, ZN => n435);
   U3 : INV_X1 port map( A => n513, ZN => n429);
   U4 : INV_X1 port map( A => n535, ZN => n441);
   U5 : INV_X1 port map( A => n532, ZN => n438);
   U6 : INV_X1 port map( A => n477, ZN => n411);
   U7 : INV_X1 port map( A => n489, ZN => n417);
   U8 : INV_X1 port map( A => n507, ZN => n426);
   U9 : INV_X1 port map( A => n501, ZN => n423);
   U10 : INV_X1 port map( A => n495, ZN => n420);
   U11 : INV_X1 port map( A => n451, ZN => n404);
   U12 : XNOR2_X1 port map( A => B(10), B => n433, ZN => n529);
   U13 : OAI22_X1 port map( A1 => n522, A2 => B(11), B1 => A(11), B2 => n432, 
                           ZN => n519);
   U14 : AND2_X1 port map( A1 => n432, A2 => A(11), ZN => n522);
   U15 : INV_X1 port map( A => n523, ZN => n432);
   U16 : AOI22_X1 port map( A1 => n408, A2 => A(29), B1 => n467, B2 => B(29), 
                           ZN => n464);
   U17 : OR2_X1 port map( A1 => A(29), A2 => n408, ZN => n467);
   U18 : INV_X1 port map( A => n468, ZN => n408);
   U19 : OAI22_X1 port map( A1 => A(10), A2 => n525, B1 => B(10), B2 => n526, 
                           ZN => n523);
   U20 : AOI211_X1 port map( C1 => n527, C2 => n434, A => n433, B => n528, ZN 
                           => n526);
   U21 : AOI21_X1 port map( B1 => A(9), B2 => n435, A => B(9), ZN => n528);
   U22 : AOI21_X1 port map( B1 => n486, B2 => A(23), A => n415, ZN => n483);
   U23 : INV_X1 port map( A => n487, ZN => n415);
   U24 : OAI21_X1 port map( B1 => A(23), B2 => n486, A => B(23), ZN => n487);
   U25 : OAI22_X1 port map( A1 => n516, A2 => B(13), B1 => A(13), B2 => n517, 
                           ZN => n513);
   U26 : AND2_X1 port map( A1 => n517, A2 => A(13), ZN => n516);
   U27 : AOI21_X1 port map( B1 => A(2), B2 => B(2), A => n445, ZN => n461);
   U28 : INV_X1 port map( A => n539, ZN => n445);
   U29 : OAI21_X1 port map( B1 => A(2), B2 => B(2), A => carry_2_port, ZN => 
                           n539);
   U30 : OAI21_X1 port map( B1 => A(8), B2 => n453, A => n436, ZN => n527);
   U31 : INV_X1 port map( A => n531, ZN => n436);
   U32 : AOI21_X1 port map( B1 => n453, B2 => A(8), A => B(8), ZN => n531);
   U33 : AOI21_X1 port map( B1 => n428, B2 => n513, A => n514, ZN => n510);
   U34 : AOI21_X1 port map( B1 => n429, B2 => A(14), A => B(14), ZN => n514);
   U35 : AOI21_X1 port map( B1 => n425, B2 => n507, A => n508, ZN => n504);
   U36 : AOI21_X1 port map( B1 => n426, B2 => A(16), A => B(16), ZN => n508);
   U37 : AOI21_X1 port map( B1 => n422, B2 => n501, A => n502, ZN => n498);
   U38 : AOI21_X1 port map( B1 => n423, B2 => A(18), A => B(18), ZN => n502);
   U39 : AOI21_X1 port map( B1 => n419, B2 => n495, A => n496, ZN => n492);
   U40 : AOI21_X1 port map( B1 => n420, B2 => A(20), A => B(20), ZN => n496);
   U41 : AOI22_X1 port map( A1 => n474, A2 => A(27), B1 => n475, B2 => B(27), 
                           ZN => n472);
   U42 : OR2_X1 port map( A1 => A(27), A2 => n474, ZN => n475);
   U43 : AOI22_X1 port map( A1 => n409, A2 => A(28), B1 => n471, B2 => B(28), 
                           ZN => n468);
   U44 : OR2_X1 port map( A1 => A(28), A2 => n409, ZN => n471);
   U45 : INV_X1 port map( A => n472, ZN => n409);
   U46 : XNOR2_X1 port map( A => n483, B => n485, ZN => SUM(24));
   U47 : XNOR2_X1 port map( A => B(24), B => n413, ZN => n485);
   U48 : XNOR2_X1 port map( A => n492, B => n494, ZN => SUM(21));
   U49 : XNOR2_X1 port map( A => A(21), B => B(21), ZN => n494);
   U50 : AOI22_X1 port map( A1 => n463, A2 => carry_33_port, B1 => A(33), B2 =>
                           B(33), ZN => n451);
   U51 : AOI21_X1 port map( B1 => n510, B2 => A(15), A => n427, ZN => n507);
   U52 : INV_X1 port map( A => n511, ZN => n427);
   U53 : OAI21_X1 port map( B1 => n510, B2 => A(15), A => B(15), ZN => n511);
   U54 : AOI21_X1 port map( B1 => n504, B2 => A(17), A => n424, ZN => n501);
   U55 : INV_X1 port map( A => n505, ZN => n424);
   U56 : OAI21_X1 port map( B1 => n504, B2 => A(17), A => B(17), ZN => n505);
   U57 : AOI21_X1 port map( B1 => n498, B2 => A(19), A => n421, ZN => n495);
   U58 : INV_X1 port map( A => n499, ZN => n421);
   U59 : OAI21_X1 port map( B1 => n498, B2 => A(19), A => B(19), ZN => n499);
   U60 : AOI21_X1 port map( B1 => n492, B2 => A(21), A => n418, ZN => n489);
   U61 : INV_X1 port map( A => n493, ZN => n418);
   U62 : OAI21_X1 port map( B1 => n492, B2 => A(21), A => B(21), ZN => n493);
   U63 : AOI21_X1 port map( B1 => n443, B2 => n461, A => n538, ZN => n459);
   U64 : AOI21_X1 port map( B1 => n444, B2 => A(3), A => B(3), ZN => n538);
   U65 : INV_X1 port map( A => n461, ZN => n444);
   U66 : AOI21_X1 port map( B1 => n413, B2 => n483, A => n484, ZN => n480);
   U67 : AOI21_X1 port map( B1 => n414, B2 => A(24), A => B(24), ZN => n484);
   U68 : INV_X1 port map( A => n483, ZN => n414);
   U69 : XNOR2_X1 port map( A => n429, B => n515, ZN => SUM(14));
   U70 : XNOR2_X1 port map( A => n411, B => n479, ZN => SUM(26));
   U71 : XNOR2_X1 port map( A => A(26), B => B(26), ZN => n479);
   U72 : XNOR2_X1 port map( A => n519, B => n521, ZN => SUM(12));
   U73 : OAI21_X1 port map( B1 => A(4), B2 => n459, A => n442, ZN => n535);
   U74 : INV_X1 port map( A => n537, ZN => n442);
   U75 : AOI21_X1 port map( B1 => n459, B2 => A(4), A => B(4), ZN => n537);
   U76 : OAI21_X1 port map( B1 => A(6), B2 => n456, A => n439, ZN => n532);
   U77 : INV_X1 port map( A => n534, ZN => n439);
   U78 : AOI21_X1 port map( B1 => n456, B2 => A(6), A => B(6), ZN => n534);
   U79 : OAI21_X1 port map( B1 => A(25), B2 => n480, A => n412, ZN => n477);
   U80 : INV_X1 port map( A => n481, ZN => n412);
   U81 : AOI21_X1 port map( B1 => n480, B2 => A(25), A => B(25), ZN => n481);
   U82 : XNOR2_X1 port map( A => n498, B => n500, ZN => SUM(19));
   U83 : XNOR2_X1 port map( A => A(19), B => B(19), ZN => n500);
   U84 : XNOR2_X1 port map( A => n441, B => n458, ZN => SUM(5));
   U85 : XNOR2_X1 port map( A => A(5), B => B(5), ZN => n458);
   U86 : XNOR2_X1 port map( A => n435, B => n452, ZN => SUM(9));
   U87 : XNOR2_X1 port map( A => B(9), B => A(9), ZN => n452);
   U88 : OAI21_X1 port map( B1 => n535, B2 => n440, A => n536, ZN => n456);
   U89 : INV_X1 port map( A => A(5), ZN => n440);
   U90 : OAI21_X1 port map( B1 => n441, B2 => A(5), A => B(5), ZN => n536);
   U91 : OAI21_X1 port map( B1 => n532, B2 => n437, A => n533, ZN => n453);
   U92 : INV_X1 port map( A => A(7), ZN => n437);
   U93 : OAI21_X1 port map( B1 => n438, B2 => A(7), A => B(7), ZN => n533);
   U94 : XNOR2_X1 port map( A => n509, B => n426, ZN => SUM(16));
   U95 : OAI21_X1 port map( B1 => n489, B2 => n416, A => n490, ZN => n486);
   U96 : INV_X1 port map( A => A(22), ZN => n416);
   U97 : OAI21_X1 port map( B1 => A(22), B2 => n417, A => B(22), ZN => n490);
   U98 : XNOR2_X1 port map( A => n464, B => n466, ZN => SUM(30));
   U99 : XNOR2_X1 port map( A => n468, B => n470, ZN => SUM(29));
   U100 : XNOR2_X1 port map( A => n491, B => n417, ZN => SUM(22));
   U101 : XNOR2_X1 port map( A => A(22), B => B(22), ZN => n491);
   U102 : OAI21_X1 port map( B1 => n519, B2 => n430, A => n520, ZN => n517);
   U103 : INV_X1 port map( A => A(12), ZN => n430);
   U104 : OAI21_X1 port map( B1 => n431, B2 => A(12), A => B(12), ZN => n520);
   U105 : INV_X1 port map( A => n519, ZN => n431);
   U106 : OAI21_X1 port map( B1 => n477, B2 => n410, A => n478, ZN => n474);
   U107 : INV_X1 port map( A => A(26), ZN => n410);
   U108 : OAI21_X1 port map( B1 => n411, B2 => A(26), A => B(26), ZN => n478);
   U109 : XNOR2_X1 port map( A => B(3), B => n443, ZN => n462);
   U110 : XNOR2_X1 port map( A => n510, B => n512, ZN => SUM(15));
   U111 : XNOR2_X1 port map( A => A(15), B => B(15), ZN => n512);
   U112 : AOI22_X1 port map( A1 => B(31), A2 => A(31), B1 => n447, B2 => n448, 
                           ZN => n446);
   U113 : XNOR2_X1 port map( A => n503, B => n423, ZN => SUM(18));
   U114 : XNOR2_X1 port map( A => n523, B => n524, ZN => SUM(11));
   U115 : XNOR2_X1 port map( A => n472, B => n473, ZN => SUM(28));
   U116 : XNOR2_X1 port map( A => n438, B => n455, ZN => SUM(7));
   U117 : XNOR2_X1 port map( A => A(7), B => B(7), ZN => n455);
   U118 : OAI21_X1 port map( B1 => n527, B2 => n434, A => n530, ZN => n525);
   U119 : OAI21_X1 port map( B1 => n435, B2 => A(9), A => B(9), ZN => n530);
   U120 : OAI21_X1 port map( B1 => n464, B2 => n406, A => n465, ZN => n447);
   U121 : INV_X1 port map( A => A(30), ZN => n406);
   U122 : OAI21_X1 port map( B1 => A(30), B2 => n407, A => B(30), ZN => n465);
   U123 : INV_X1 port map( A => n464, ZN => n407);
   U124 : INV_X1 port map( A => A(9), ZN => n434);
   U125 : INV_X1 port map( A => A(3), ZN => n443);
   U126 : INV_X1 port map( A => A(24), ZN => n413);
   U127 : INV_X1 port map( A => A(10), ZN => n433);
   U128 : INV_X1 port map( A => n446, ZN => n405);
   U129 : INV_X1 port map( A => A(14), ZN => n428);
   U130 : INV_X1 port map( A => A(16), ZN => n425);
   U131 : INV_X1 port map( A => A(18), ZN => n422);
   U132 : INV_X1 port map( A => A(20), ZN => n419);
   U133 : XNOR2_X1 port map( A => n497, B => n420, ZN => SUM(20));
   U134 : XNOR2_X1 port map( A => n504, B => n506, ZN => SUM(17));
   U135 : XNOR2_X1 port map( A => A(17), B => B(17), ZN => n506);
   U136 : INV_X1 port map( A => n449, ZN => n403);
   U137 : AOI22_X1 port map( A1 => B(34), A2 => A(34), B1 => n404, B2 => n450, 
                           ZN => n449);
   U138 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => n1);
   U139 : XNOR2_X1 port map( A => n461, B => n462, ZN => SUM(3));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT64 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64;

architecture SYN_DIRECT of RCA_NBIT64 is

   component RCA_NBIT64_DW01_add_0
      port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (63 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1065 : std_logic;

begin
   
   Co <= '0';
   n2 <= '0';
   add_95 : RCA_NBIT64_DW01_add_0 port map( A(63) => A(63), A(62) => A(62), 
                           A(61) => A(61), A(60) => A(60), A(59) => A(59), 
                           A(58) => A(58), A(57) => A(57), A(56) => A(56), 
                           A(55) => A(55), A(54) => A(54), A(53) => A(53), 
                           A(52) => A(52), A(51) => A(51), A(50) => A(50), 
                           A(49) => A(49), A(48) => A(48), A(47) => A(47), 
                           A(46) => A(46), A(45) => A(45), A(44) => A(44), 
                           A(43) => A(43), A(42) => A(42), A(41) => A(41), 
                           A(40) => A(40), A(39) => A(39), A(38) => A(38), 
                           A(37) => A(37), A(36) => A(36), A(35) => A(35), 
                           A(34) => A(34), A(33) => A(33), A(32) => A(32), 
                           A(31) => A(31), A(30) => A(30), A(29) => A(29), 
                           A(28) => A(28), A(27) => A(27), A(26) => A(26), 
                           A(25) => A(25), A(24) => A(24), A(23) => A(23), 
                           A(22) => A(22), A(21) => A(21), A(20) => A(20), 
                           A(19) => A(19), A(18) => A(18), A(17) => A(17), 
                           A(16) => A(16), A(15) => A(15), A(14) => A(14), 
                           A(13) => A(13), A(12) => A(12), A(11) => A(11), 
                           A(10) => A(10), A(9) => A(9), A(8) => A(8), A(7) => 
                           A(7), A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3)
                           => A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(63) => B(63), B(62) => B(62), B(61) => B(61), 
                           B(60) => B(60), B(59) => B(59), B(58) => B(58), 
                           B(57) => B(57), B(56) => B(56), B(55) => B(55), 
                           B(54) => B(54), B(53) => B(53), B(52) => B(52), 
                           B(51) => B(51), B(50) => B(50), B(49) => B(49), 
                           B(48) => B(48), B(47) => B(47), B(46) => B(46), 
                           B(45) => B(45), B(44) => B(44), B(43) => B(43), 
                           B(42) => B(42), B(41) => B(41), B(40) => B(40), 
                           B(39) => B(39), B(38) => B(38), B(37) => B(37), 
                           B(36) => B(36), B(35) => B(35), B(34) => B(34), 
                           B(33) => B(33), B(32) => B(32), B(31) => B(31), 
                           B(30) => B(30), B(29) => B(29), B(28) => B(28), 
                           B(27) => B(27), B(26) => B(26), B(25) => B(25), 
                           B(24) => B(24), B(23) => B(23), B(22) => B(22), 
                           B(21) => B(21), B(20) => B(20), B(19) => B(19), 
                           B(18) => B(18), B(17) => B(17), B(16) => B(16), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => B(0), CI => n2, SUM(63) 
                           => S(63), SUM(62) => S(62), SUM(61) => S(61), 
                           SUM(60) => S(60), SUM(59) => S(59), SUM(58) => S(58)
                           , SUM(57) => S(57), SUM(56) => S(56), SUM(55) => 
                           S(55), SUM(54) => S(54), SUM(53) => S(53), SUM(52) 
                           => S(52), SUM(51) => S(51), SUM(50) => S(50), 
                           SUM(49) => S(49), SUM(48) => S(48), SUM(47) => S(47)
                           , SUM(46) => S(46), SUM(45) => S(45), SUM(44) => 
                           S(44), SUM(43) => S(43), SUM(42) => S(42), SUM(41) 
                           => S(41), SUM(40) => S(40), SUM(39) => S(39), 
                           SUM(38) => S(38), SUM(37) => S(37), SUM(36) => S(36)
                           , SUM(35) => S(35), SUM(34) => S(34), SUM(33) => 
                           S(33), SUM(32) => S(32), SUM(31) => S(31), SUM(30) 
                           => S(30), SUM(29) => S(29), SUM(28) => S(28), 
                           SUM(27) => S(27), SUM(26) => S(26), SUM(25) => S(25)
                           , SUM(24) => S(24), SUM(23) => S(23), SUM(22) => 
                           S(22), SUM(21) => S(21), SUM(20) => S(20), SUM(19) 
                           => S(19), SUM(18) => S(18), SUM(17) => S(17), 
                           SUM(16) => S(16), SUM(15) => S(15), SUM(14) => S(14)
                           , SUM(13) => S(13), SUM(12) => S(12), SUM(11) => 
                           S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) => 
                           S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5)
                           , SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1065);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT62 is

   port( A, B : in std_logic_vector (61 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (61 downto 0);  Co : out std_logic);

end RCA_NBIT62;

architecture SYN_DIRECT of RCA_NBIT62 is

   component RCA_NBIT62_DW01_add_0
      port( A, B : in std_logic_vector (61 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (61 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1066 : std_logic;

begin
   
   Co <= '0';
   n2 <= '0';
   add_95 : RCA_NBIT62_DW01_add_0 port map( A(61) => A(61), A(60) => A(60), 
                           A(59) => A(59), A(58) => A(58), A(57) => A(57), 
                           A(56) => A(56), A(55) => A(55), A(54) => A(54), 
                           A(53) => A(53), A(52) => A(52), A(51) => A(51), 
                           A(50) => A(50), A(49) => A(49), A(48) => A(48), 
                           A(47) => A(47), A(46) => A(46), A(45) => A(45), 
                           A(44) => A(44), A(43) => A(43), A(42) => A(42), 
                           A(41) => A(41), A(40) => A(40), A(39) => A(39), 
                           A(38) => A(38), A(37) => A(37), A(36) => A(36), 
                           A(35) => A(35), A(34) => A(34), A(33) => A(33), 
                           A(32) => A(32), A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(61) => B(61), B(60) => B(60), 
                           B(59) => B(59), B(58) => B(58), B(57) => B(57), 
                           B(56) => B(56), B(55) => B(55), B(54) => B(54), 
                           B(53) => B(53), B(52) => B(52), B(51) => B(51), 
                           B(50) => B(50), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => n2, SUM(61) => S(61), 
                           SUM(60) => S(60), SUM(59) => S(59), SUM(58) => S(58)
                           , SUM(57) => S(57), SUM(56) => S(56), SUM(55) => 
                           S(55), SUM(54) => S(54), SUM(53) => S(53), SUM(52) 
                           => S(52), SUM(51) => S(51), SUM(50) => S(50), 
                           SUM(49) => S(49), SUM(48) => S(48), SUM(47) => S(47)
                           , SUM(46) => S(46), SUM(45) => S(45), SUM(44) => 
                           S(44), SUM(43) => S(43), SUM(42) => S(42), SUM(41) 
                           => S(41), SUM(40) => S(40), SUM(39) => S(39), 
                           SUM(38) => S(38), SUM(37) => S(37), SUM(36) => S(36)
                           , SUM(35) => S(35), SUM(34) => S(34), SUM(33) => 
                           S(33), SUM(32) => S(32), SUM(31) => S(31), SUM(30) 
                           => S(30), SUM(29) => S(29), SUM(28) => S(28), 
                           SUM(27) => S(27), SUM(26) => S(26), SUM(25) => S(25)
                           , SUM(24) => S(24), SUM(23) => S(23), SUM(22) => 
                           S(22), SUM(21) => S(21), SUM(20) => S(20), SUM(19) 
                           => S(19), SUM(18) => S(18), SUM(17) => S(17), 
                           SUM(16) => S(16), SUM(15) => S(15), SUM(14) => S(14)
                           , SUM(13) => S(13), SUM(12) => S(12), SUM(11) => 
                           S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) => 
                           S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5)
                           , SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1066);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT60 is

   port( A, B : in std_logic_vector (59 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (59 downto 0);  Co : out std_logic);

end RCA_NBIT60;

architecture SYN_DIRECT of RCA_NBIT60 is

   component RCA_NBIT60_DW01_add_0
      port( A, B : in std_logic_vector (59 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (59 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1067 : std_logic;

begin
   
   Co <= '0';
   n2 <= '0';
   add_95 : RCA_NBIT60_DW01_add_0 port map( A(59) => A(59), A(58) => A(58), 
                           A(57) => A(57), A(56) => A(56), A(55) => A(55), 
                           A(54) => A(54), A(53) => A(53), A(52) => A(52), 
                           A(51) => A(51), A(50) => A(50), A(49) => A(49), 
                           A(48) => A(48), A(47) => A(47), A(46) => A(46), 
                           A(45) => A(45), A(44) => A(44), A(43) => A(43), 
                           A(42) => A(42), A(41) => A(41), A(40) => A(40), 
                           A(39) => A(39), A(38) => A(38), A(37) => A(37), 
                           A(36) => A(36), A(35) => A(35), A(34) => A(34), 
                           A(33) => A(33), A(32) => A(32), A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(59) => B(59), 
                           B(58) => B(58), B(57) => B(57), B(56) => B(56), 
                           B(55) => B(55), B(54) => B(54), B(53) => B(53), 
                           B(52) => B(52), B(51) => B(51), B(50) => B(50), 
                           B(49) => B(49), B(48) => B(48), B(47) => B(47), 
                           B(46) => B(46), B(45) => B(45), B(44) => B(44), 
                           B(43) => B(43), B(42) => B(42), B(41) => B(41), 
                           B(40) => B(40), B(39) => B(39), B(38) => B(38), 
                           B(37) => B(37), B(36) => B(36), B(35) => B(35), 
                           B(34) => B(34), B(33) => B(33), B(32) => B(32), 
                           B(31) => B(31), B(30) => B(30), B(29) => B(29), 
                           B(28) => B(28), B(27) => B(27), B(26) => B(26), 
                           B(25) => B(25), B(24) => B(24), B(23) => B(23), 
                           B(22) => B(22), B(21) => B(21), B(20) => B(20), 
                           B(19) => B(19), B(18) => B(18), B(17) => B(17), 
                           B(16) => B(16), B(15) => B(15), B(14) => B(14), 
                           B(13) => B(13), B(12) => B(12), B(11) => B(11), 
                           B(10) => B(10), B(9) => B(9), B(8) => B(8), B(7) => 
                           B(7), B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3)
                           => B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), 
                           CI => n2, SUM(59) => S(59), SUM(58) => S(58), 
                           SUM(57) => S(57), SUM(56) => S(56), SUM(55) => S(55)
                           , SUM(54) => S(54), SUM(53) => S(53), SUM(52) => 
                           S(52), SUM(51) => S(51), SUM(50) => S(50), SUM(49) 
                           => S(49), SUM(48) => S(48), SUM(47) => S(47), 
                           SUM(46) => S(46), SUM(45) => S(45), SUM(44) => S(44)
                           , SUM(43) => S(43), SUM(42) => S(42), SUM(41) => 
                           S(41), SUM(40) => S(40), SUM(39) => S(39), SUM(38) 
                           => S(38), SUM(37) => S(37), SUM(36) => S(36), 
                           SUM(35) => S(35), SUM(34) => S(34), SUM(33) => S(33)
                           , SUM(32) => S(32), SUM(31) => S(31), SUM(30) => 
                           S(30), SUM(29) => S(29), SUM(28) => S(28), SUM(27) 
                           => S(27), SUM(26) => S(26), SUM(25) => S(25), 
                           SUM(24) => S(24), SUM(23) => S(23), SUM(22) => S(22)
                           , SUM(21) => S(21), SUM(20) => S(20), SUM(19) => 
                           S(19), SUM(18) => S(18), SUM(17) => S(17), SUM(16) 
                           => S(16), SUM(15) => S(15), SUM(14) => S(14), 
                           SUM(13) => S(13), SUM(12) => S(12), SUM(11) => S(11)
                           , SUM(10) => S(10), SUM(9) => S(9), SUM(8) => S(8), 
                           SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5), 
                           SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1067);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT58 is

   port( A, B : in std_logic_vector (57 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (57 downto 0);  Co : out std_logic);

end RCA_NBIT58;

architecture SYN_DIRECT of RCA_NBIT58 is

   component RCA_NBIT58_DW01_add_0
      port( A, B : in std_logic_vector (57 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (57 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1068 : std_logic;

begin
   
   Co <= '0';
   n2 <= '0';
   add_95 : RCA_NBIT58_DW01_add_0 port map( A(57) => A(57), A(56) => A(56), 
                           A(55) => A(55), A(54) => A(54), A(53) => A(53), 
                           A(52) => A(52), A(51) => A(51), A(50) => A(50), 
                           A(49) => A(49), A(48) => A(48), A(47) => A(47), 
                           A(46) => A(46), A(45) => A(45), A(44) => A(44), 
                           A(43) => A(43), A(42) => A(42), A(41) => A(41), 
                           A(40) => A(40), A(39) => A(39), A(38) => A(38), 
                           A(37) => A(37), A(36) => A(36), A(35) => A(35), 
                           A(34) => A(34), A(33) => A(33), A(32) => A(32), 
                           A(31) => A(31), A(30) => A(30), A(29) => A(29), 
                           A(28) => A(28), A(27) => A(27), A(26) => A(26), 
                           A(25) => A(25), A(24) => A(24), A(23) => A(23), 
                           A(22) => A(22), A(21) => A(21), A(20) => A(20), 
                           A(19) => A(19), A(18) => A(18), A(17) => A(17), 
                           A(16) => A(16), A(15) => A(15), A(14) => A(14), 
                           A(13) => A(13), A(12) => A(12), A(11) => A(11), 
                           A(10) => A(10), A(9) => A(9), A(8) => A(8), A(7) => 
                           A(7), A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3)
                           => A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(57) => B(57), B(56) => B(56), B(55) => B(55), 
                           B(54) => B(54), B(53) => B(53), B(52) => B(52), 
                           B(51) => B(51), B(50) => B(50), B(49) => B(49), 
                           B(48) => B(48), B(47) => B(47), B(46) => B(46), 
                           B(45) => B(45), B(44) => B(44), B(43) => B(43), 
                           B(42) => B(42), B(41) => B(41), B(40) => B(40), 
                           B(39) => B(39), B(38) => B(38), B(37) => B(37), 
                           B(36) => B(36), B(35) => B(35), B(34) => B(34), 
                           B(33) => B(33), B(32) => B(32), B(31) => B(31), 
                           B(30) => B(30), B(29) => B(29), B(28) => B(28), 
                           B(27) => B(27), B(26) => B(26), B(25) => B(25), 
                           B(24) => B(24), B(23) => B(23), B(22) => B(22), 
                           B(21) => B(21), B(20) => B(20), B(19) => B(19), 
                           B(18) => B(18), B(17) => B(17), B(16) => B(16), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => B(0), CI => n2, SUM(57) 
                           => S(57), SUM(56) => S(56), SUM(55) => S(55), 
                           SUM(54) => S(54), SUM(53) => S(53), SUM(52) => S(52)
                           , SUM(51) => S(51), SUM(50) => S(50), SUM(49) => 
                           S(49), SUM(48) => S(48), SUM(47) => S(47), SUM(46) 
                           => S(46), SUM(45) => S(45), SUM(44) => S(44), 
                           SUM(43) => S(43), SUM(42) => S(42), SUM(41) => S(41)
                           , SUM(40) => S(40), SUM(39) => S(39), SUM(38) => 
                           S(38), SUM(37) => S(37), SUM(36) => S(36), SUM(35) 
                           => S(35), SUM(34) => S(34), SUM(33) => S(33), 
                           SUM(32) => S(32), SUM(31) => S(31), SUM(30) => S(30)
                           , SUM(29) => S(29), SUM(28) => S(28), SUM(27) => 
                           S(27), SUM(26) => S(26), SUM(25) => S(25), SUM(24) 
                           => S(24), SUM(23) => S(23), SUM(22) => S(22), 
                           SUM(21) => S(21), SUM(20) => S(20), SUM(19) => S(19)
                           , SUM(18) => S(18), SUM(17) => S(17), SUM(16) => 
                           S(16), SUM(15) => S(15), SUM(14) => S(14), SUM(13) 
                           => S(13), SUM(12) => S(12), SUM(11) => S(11), 
                           SUM(10) => S(10), SUM(9) => S(9), SUM(8) => S(8), 
                           SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5), 
                           SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1068);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT56 is

   port( A, B : in std_logic_vector (55 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (55 downto 0);  Co : out std_logic);

end RCA_NBIT56;

architecture SYN_DIRECT of RCA_NBIT56 is

   component RCA_NBIT56_DW01_add_0
      port( A, B : in std_logic_vector (55 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (55 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1069 : std_logic;

begin
   
   Co <= '0';
   n2 <= '0';
   add_95 : RCA_NBIT56_DW01_add_0 port map( A(55) => A(55), A(54) => A(54), 
                           A(53) => A(53), A(52) => A(52), A(51) => A(51), 
                           A(50) => A(50), A(49) => A(49), A(48) => A(48), 
                           A(47) => A(47), A(46) => A(46), A(45) => A(45), 
                           A(44) => A(44), A(43) => A(43), A(42) => A(42), 
                           A(41) => A(41), A(40) => A(40), A(39) => A(39), 
                           A(38) => A(38), A(37) => A(37), A(36) => A(36), 
                           A(35) => A(35), A(34) => A(34), A(33) => A(33), 
                           A(32) => A(32), A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(55) => B(55), B(54) => B(54), 
                           B(53) => B(53), B(52) => B(52), B(51) => B(51), 
                           B(50) => B(50), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => n2, SUM(55) => S(55), 
                           SUM(54) => S(54), SUM(53) => S(53), SUM(52) => S(52)
                           , SUM(51) => S(51), SUM(50) => S(50), SUM(49) => 
                           S(49), SUM(48) => S(48), SUM(47) => S(47), SUM(46) 
                           => S(46), SUM(45) => S(45), SUM(44) => S(44), 
                           SUM(43) => S(43), SUM(42) => S(42), SUM(41) => S(41)
                           , SUM(40) => S(40), SUM(39) => S(39), SUM(38) => 
                           S(38), SUM(37) => S(37), SUM(36) => S(36), SUM(35) 
                           => S(35), SUM(34) => S(34), SUM(33) => S(33), 
                           SUM(32) => S(32), SUM(31) => S(31), SUM(30) => S(30)
                           , SUM(29) => S(29), SUM(28) => S(28), SUM(27) => 
                           S(27), SUM(26) => S(26), SUM(25) => S(25), SUM(24) 
                           => S(24), SUM(23) => S(23), SUM(22) => S(22), 
                           SUM(21) => S(21), SUM(20) => S(20), SUM(19) => S(19)
                           , SUM(18) => S(18), SUM(17) => S(17), SUM(16) => 
                           S(16), SUM(15) => S(15), SUM(14) => S(14), SUM(13) 
                           => S(13), SUM(12) => S(12), SUM(11) => S(11), 
                           SUM(10) => S(10), SUM(9) => S(9), SUM(8) => S(8), 
                           SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5), 
                           SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1069);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT54 is

   port( A, B : in std_logic_vector (53 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (53 downto 0);  Co : out std_logic);

end RCA_NBIT54;

architecture SYN_DIRECT of RCA_NBIT54 is

   component RCA_NBIT54_DW01_add_0
      port( A, B : in std_logic_vector (53 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (53 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1070 : std_logic;

begin
   
   Co <= '0';
   n2 <= '0';
   add_95 : RCA_NBIT54_DW01_add_0 port map( A(53) => A(53), A(52) => A(52), 
                           A(51) => A(51), A(50) => A(50), A(49) => A(49), 
                           A(48) => A(48), A(47) => A(47), A(46) => A(46), 
                           A(45) => A(45), A(44) => A(44), A(43) => A(43), 
                           A(42) => A(42), A(41) => A(41), A(40) => A(40), 
                           A(39) => A(39), A(38) => A(38), A(37) => A(37), 
                           A(36) => A(36), A(35) => A(35), A(34) => A(34), 
                           A(33) => A(33), A(32) => A(32), A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(53) => B(53), 
                           B(52) => B(52), B(51) => B(51), B(50) => B(50), 
                           B(49) => B(49), B(48) => B(48), B(47) => B(47), 
                           B(46) => B(46), B(45) => B(45), B(44) => B(44), 
                           B(43) => B(43), B(42) => B(42), B(41) => B(41), 
                           B(40) => B(40), B(39) => B(39), B(38) => B(38), 
                           B(37) => B(37), B(36) => B(36), B(35) => B(35), 
                           B(34) => B(34), B(33) => B(33), B(32) => B(32), 
                           B(31) => B(31), B(30) => B(30), B(29) => B(29), 
                           B(28) => B(28), B(27) => B(27), B(26) => B(26), 
                           B(25) => B(25), B(24) => B(24), B(23) => B(23), 
                           B(22) => B(22), B(21) => B(21), B(20) => B(20), 
                           B(19) => B(19), B(18) => B(18), B(17) => B(17), 
                           B(16) => B(16), B(15) => B(15), B(14) => B(14), 
                           B(13) => B(13), B(12) => B(12), B(11) => B(11), 
                           B(10) => B(10), B(9) => B(9), B(8) => B(8), B(7) => 
                           B(7), B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3)
                           => B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), 
                           CI => n2, SUM(53) => S(53), SUM(52) => S(52), 
                           SUM(51) => S(51), SUM(50) => S(50), SUM(49) => S(49)
                           , SUM(48) => S(48), SUM(47) => S(47), SUM(46) => 
                           S(46), SUM(45) => S(45), SUM(44) => S(44), SUM(43) 
                           => S(43), SUM(42) => S(42), SUM(41) => S(41), 
                           SUM(40) => S(40), SUM(39) => S(39), SUM(38) => S(38)
                           , SUM(37) => S(37), SUM(36) => S(36), SUM(35) => 
                           S(35), SUM(34) => S(34), SUM(33) => S(33), SUM(32) 
                           => S(32), SUM(31) => S(31), SUM(30) => S(30), 
                           SUM(29) => S(29), SUM(28) => S(28), SUM(27) => S(27)
                           , SUM(26) => S(26), SUM(25) => S(25), SUM(24) => 
                           S(24), SUM(23) => S(23), SUM(22) => S(22), SUM(21) 
                           => S(21), SUM(20) => S(20), SUM(19) => S(19), 
                           SUM(18) => S(18), SUM(17) => S(17), SUM(16) => S(16)
                           , SUM(15) => S(15), SUM(14) => S(14), SUM(13) => 
                           S(13), SUM(12) => S(12), SUM(11) => S(11), SUM(10) 
                           => S(10), SUM(9) => S(9), SUM(8) => S(8), SUM(7) => 
                           S(7), SUM(6) => S(6), SUM(5) => S(5), SUM(4) => S(4)
                           , SUM(3) => S(3), SUM(2) => S(2), SUM(1) => S(1), 
                           SUM(0) => S(0), CO => n_1070);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT52 is

   port( A, B : in std_logic_vector (51 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (51 downto 0);  Co : out std_logic);

end RCA_NBIT52;

architecture SYN_DIRECT of RCA_NBIT52 is

   component RCA_NBIT52_DW01_add_0
      port( A, B : in std_logic_vector (51 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (51 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1071 : std_logic;

begin
   
   Co <= '0';
   n2 <= '0';
   add_95 : RCA_NBIT52_DW01_add_0 port map( A(51) => A(51), A(50) => A(50), 
                           A(49) => A(49), A(48) => A(48), A(47) => A(47), 
                           A(46) => A(46), A(45) => A(45), A(44) => A(44), 
                           A(43) => A(43), A(42) => A(42), A(41) => A(41), 
                           A(40) => A(40), A(39) => A(39), A(38) => A(38), 
                           A(37) => A(37), A(36) => A(36), A(35) => A(35), 
                           A(34) => A(34), A(33) => A(33), A(32) => A(32), 
                           A(31) => A(31), A(30) => A(30), A(29) => A(29), 
                           A(28) => A(28), A(27) => A(27), A(26) => A(26), 
                           A(25) => A(25), A(24) => A(24), A(23) => A(23), 
                           A(22) => A(22), A(21) => A(21), A(20) => A(20), 
                           A(19) => A(19), A(18) => A(18), A(17) => A(17), 
                           A(16) => A(16), A(15) => A(15), A(14) => A(14), 
                           A(13) => A(13), A(12) => A(12), A(11) => A(11), 
                           A(10) => A(10), A(9) => A(9), A(8) => A(8), A(7) => 
                           A(7), A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3)
                           => A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(51) => B(51), B(50) => B(50), B(49) => B(49), 
                           B(48) => B(48), B(47) => B(47), B(46) => B(46), 
                           B(45) => B(45), B(44) => B(44), B(43) => B(43), 
                           B(42) => B(42), B(41) => B(41), B(40) => B(40), 
                           B(39) => B(39), B(38) => B(38), B(37) => B(37), 
                           B(36) => B(36), B(35) => B(35), B(34) => B(34), 
                           B(33) => B(33), B(32) => B(32), B(31) => B(31), 
                           B(30) => B(30), B(29) => B(29), B(28) => B(28), 
                           B(27) => B(27), B(26) => B(26), B(25) => B(25), 
                           B(24) => B(24), B(23) => B(23), B(22) => B(22), 
                           B(21) => B(21), B(20) => B(20), B(19) => B(19), 
                           B(18) => B(18), B(17) => B(17), B(16) => B(16), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => B(0), CI => n2, SUM(51) 
                           => S(51), SUM(50) => S(50), SUM(49) => S(49), 
                           SUM(48) => S(48), SUM(47) => S(47), SUM(46) => S(46)
                           , SUM(45) => S(45), SUM(44) => S(44), SUM(43) => 
                           S(43), SUM(42) => S(42), SUM(41) => S(41), SUM(40) 
                           => S(40), SUM(39) => S(39), SUM(38) => S(38), 
                           SUM(37) => S(37), SUM(36) => S(36), SUM(35) => S(35)
                           , SUM(34) => S(34), SUM(33) => S(33), SUM(32) => 
                           S(32), SUM(31) => S(31), SUM(30) => S(30), SUM(29) 
                           => S(29), SUM(28) => S(28), SUM(27) => S(27), 
                           SUM(26) => S(26), SUM(25) => S(25), SUM(24) => S(24)
                           , SUM(23) => S(23), SUM(22) => S(22), SUM(21) => 
                           S(21), SUM(20) => S(20), SUM(19) => S(19), SUM(18) 
                           => S(18), SUM(17) => S(17), SUM(16) => S(16), 
                           SUM(15) => S(15), SUM(14) => S(14), SUM(13) => S(13)
                           , SUM(12) => S(12), SUM(11) => S(11), SUM(10) => 
                           S(10), SUM(9) => S(9), SUM(8) => S(8), SUM(7) => 
                           S(7), SUM(6) => S(6), SUM(5) => S(5), SUM(4) => S(4)
                           , SUM(3) => S(3), SUM(2) => S(2), SUM(1) => S(1), 
                           SUM(0) => S(0), CO => n_1071);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT50 is

   port( A, B : in std_logic_vector (49 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (49 downto 0);  Co : out std_logic);

end RCA_NBIT50;

architecture SYN_DIRECT of RCA_NBIT50 is

   component RCA_NBIT50_DW01_add_0
      port( A, B : in std_logic_vector (49 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (49 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1072 : std_logic;

begin
   
   Co <= '0';
   n2 <= '0';
   add_95 : RCA_NBIT50_DW01_add_0 port map( A(49) => A(49), A(48) => A(48), 
                           A(47) => A(47), A(46) => A(46), A(45) => A(45), 
                           A(44) => A(44), A(43) => A(43), A(42) => A(42), 
                           A(41) => A(41), A(40) => A(40), A(39) => A(39), 
                           A(38) => A(38), A(37) => A(37), A(36) => A(36), 
                           A(35) => A(35), A(34) => A(34), A(33) => A(33), 
                           A(32) => A(32), A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => n2, SUM(49) => S(49), 
                           SUM(48) => S(48), SUM(47) => S(47), SUM(46) => S(46)
                           , SUM(45) => S(45), SUM(44) => S(44), SUM(43) => 
                           S(43), SUM(42) => S(42), SUM(41) => S(41), SUM(40) 
                           => S(40), SUM(39) => S(39), SUM(38) => S(38), 
                           SUM(37) => S(37), SUM(36) => S(36), SUM(35) => S(35)
                           , SUM(34) => S(34), SUM(33) => S(33), SUM(32) => 
                           S(32), SUM(31) => S(31), SUM(30) => S(30), SUM(29) 
                           => S(29), SUM(28) => S(28), SUM(27) => S(27), 
                           SUM(26) => S(26), SUM(25) => S(25), SUM(24) => S(24)
                           , SUM(23) => S(23), SUM(22) => S(22), SUM(21) => 
                           S(21), SUM(20) => S(20), SUM(19) => S(19), SUM(18) 
                           => S(18), SUM(17) => S(17), SUM(16) => S(16), 
                           SUM(15) => S(15), SUM(14) => S(14), SUM(13) => S(13)
                           , SUM(12) => S(12), SUM(11) => S(11), SUM(10) => 
                           S(10), SUM(9) => S(9), SUM(8) => S(8), SUM(7) => 
                           S(7), SUM(6) => S(6), SUM(5) => S(5), SUM(4) => S(4)
                           , SUM(3) => S(3), SUM(2) => S(2), SUM(1) => S(1), 
                           SUM(0) => S(0), CO => n_1072);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT48 is

   port( A, B : in std_logic_vector (47 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (47 downto 0);  Co : out std_logic);

end RCA_NBIT48;

architecture SYN_DIRECT of RCA_NBIT48 is

   component RCA_NBIT48_DW01_add_0
      port( A, B : in std_logic_vector (47 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (47 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1073 : std_logic;

begin
   
   Co <= '0';
   n2 <= '0';
   add_95 : RCA_NBIT48_DW01_add_0 port map( A(47) => A(47), A(46) => A(46), 
                           A(45) => A(45), A(44) => A(44), A(43) => A(43), 
                           A(42) => A(42), A(41) => A(41), A(40) => A(40), 
                           A(39) => A(39), A(38) => A(38), A(37) => A(37), 
                           A(36) => A(36), A(35) => A(35), A(34) => A(34), 
                           A(33) => A(33), A(32) => A(32), A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(47) => B(47), 
                           B(46) => B(46), B(45) => B(45), B(44) => B(44), 
                           B(43) => B(43), B(42) => B(42), B(41) => B(41), 
                           B(40) => B(40), B(39) => B(39), B(38) => B(38), 
                           B(37) => B(37), B(36) => B(36), B(35) => B(35), 
                           B(34) => B(34), B(33) => B(33), B(32) => B(32), 
                           B(31) => B(31), B(30) => B(30), B(29) => B(29), 
                           B(28) => B(28), B(27) => B(27), B(26) => B(26), 
                           B(25) => B(25), B(24) => B(24), B(23) => B(23), 
                           B(22) => B(22), B(21) => B(21), B(20) => B(20), 
                           B(19) => B(19), B(18) => B(18), B(17) => B(17), 
                           B(16) => B(16), B(15) => B(15), B(14) => B(14), 
                           B(13) => B(13), B(12) => B(12), B(11) => B(11), 
                           B(10) => B(10), B(9) => B(9), B(8) => B(8), B(7) => 
                           B(7), B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3)
                           => B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), 
                           CI => n2, SUM(47) => S(47), SUM(46) => S(46), 
                           SUM(45) => S(45), SUM(44) => S(44), SUM(43) => S(43)
                           , SUM(42) => S(42), SUM(41) => S(41), SUM(40) => 
                           S(40), SUM(39) => S(39), SUM(38) => S(38), SUM(37) 
                           => S(37), SUM(36) => S(36), SUM(35) => S(35), 
                           SUM(34) => S(34), SUM(33) => S(33), SUM(32) => S(32)
                           , SUM(31) => S(31), SUM(30) => S(30), SUM(29) => 
                           S(29), SUM(28) => S(28), SUM(27) => S(27), SUM(26) 
                           => S(26), SUM(25) => S(25), SUM(24) => S(24), 
                           SUM(23) => S(23), SUM(22) => S(22), SUM(21) => S(21)
                           , SUM(20) => S(20), SUM(19) => S(19), SUM(18) => 
                           S(18), SUM(17) => S(17), SUM(16) => S(16), SUM(15) 
                           => S(15), SUM(14) => S(14), SUM(13) => S(13), 
                           SUM(12) => S(12), SUM(11) => S(11), SUM(10) => S(10)
                           , SUM(9) => S(9), SUM(8) => S(8), SUM(7) => S(7), 
                           SUM(6) => S(6), SUM(5) => S(5), SUM(4) => S(4), 
                           SUM(3) => S(3), SUM(2) => S(2), SUM(1) => S(1), 
                           SUM(0) => S(0), CO => n_1073);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT46 is

   port( A, B : in std_logic_vector (45 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (45 downto 0);  Co : out std_logic);

end RCA_NBIT46;

architecture SYN_DIRECT of RCA_NBIT46 is

   component RCA_NBIT46_DW01_add_0
      port( A, B : in std_logic_vector (45 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (45 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1074 : std_logic;

begin
   
   Co <= '0';
   n2 <= '0';
   add_95 : RCA_NBIT46_DW01_add_0 port map( A(45) => A(45), A(44) => A(44), 
                           A(43) => A(43), A(42) => A(42), A(41) => A(41), 
                           A(40) => A(40), A(39) => A(39), A(38) => A(38), 
                           A(37) => A(37), A(36) => A(36), A(35) => A(35), 
                           A(34) => A(34), A(33) => A(33), A(32) => A(32), 
                           A(31) => A(31), A(30) => A(30), A(29) => A(29), 
                           A(28) => A(28), A(27) => A(27), A(26) => A(26), 
                           A(25) => A(25), A(24) => A(24), A(23) => A(23), 
                           A(22) => A(22), A(21) => A(21), A(20) => A(20), 
                           A(19) => A(19), A(18) => A(18), A(17) => A(17), 
                           A(16) => A(16), A(15) => A(15), A(14) => A(14), 
                           A(13) => A(13), A(12) => A(12), A(11) => A(11), 
                           A(10) => A(10), A(9) => A(9), A(8) => A(8), A(7) => 
                           A(7), A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3)
                           => A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(45) => B(45), B(44) => B(44), B(43) => B(43), 
                           B(42) => B(42), B(41) => B(41), B(40) => B(40), 
                           B(39) => B(39), B(38) => B(38), B(37) => B(37), 
                           B(36) => B(36), B(35) => B(35), B(34) => B(34), 
                           B(33) => B(33), B(32) => B(32), B(31) => B(31), 
                           B(30) => B(30), B(29) => B(29), B(28) => B(28), 
                           B(27) => B(27), B(26) => B(26), B(25) => B(25), 
                           B(24) => B(24), B(23) => B(23), B(22) => B(22), 
                           B(21) => B(21), B(20) => B(20), B(19) => B(19), 
                           B(18) => B(18), B(17) => B(17), B(16) => B(16), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => B(0), CI => n2, SUM(45) 
                           => S(45), SUM(44) => S(44), SUM(43) => S(43), 
                           SUM(42) => S(42), SUM(41) => S(41), SUM(40) => S(40)
                           , SUM(39) => S(39), SUM(38) => S(38), SUM(37) => 
                           S(37), SUM(36) => S(36), SUM(35) => S(35), SUM(34) 
                           => S(34), SUM(33) => S(33), SUM(32) => S(32), 
                           SUM(31) => S(31), SUM(30) => S(30), SUM(29) => S(29)
                           , SUM(28) => S(28), SUM(27) => S(27), SUM(26) => 
                           S(26), SUM(25) => S(25), SUM(24) => S(24), SUM(23) 
                           => S(23), SUM(22) => S(22), SUM(21) => S(21), 
                           SUM(20) => S(20), SUM(19) => S(19), SUM(18) => S(18)
                           , SUM(17) => S(17), SUM(16) => S(16), SUM(15) => 
                           S(15), SUM(14) => S(14), SUM(13) => S(13), SUM(12) 
                           => S(12), SUM(11) => S(11), SUM(10) => S(10), SUM(9)
                           => S(9), SUM(8) => S(8), SUM(7) => S(7), SUM(6) => 
                           S(6), SUM(5) => S(5), SUM(4) => S(4), SUM(3) => S(3)
                           , SUM(2) => S(2), SUM(1) => S(1), SUM(0) => S(0), CO
                           => n_1074);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT44 is

   port( A, B : in std_logic_vector (43 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (43 downto 0);  Co : out std_logic);

end RCA_NBIT44;

architecture SYN_DIRECT of RCA_NBIT44 is

   component RCA_NBIT44_DW01_add_0
      port( A, B : in std_logic_vector (43 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (43 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1075 : std_logic;

begin
   
   Co <= '0';
   n2 <= '0';
   add_95 : RCA_NBIT44_DW01_add_0 port map( A(43) => A(43), A(42) => A(42), 
                           A(41) => A(41), A(40) => A(40), A(39) => A(39), 
                           A(38) => A(38), A(37) => A(37), A(36) => A(36), 
                           A(35) => A(35), A(34) => A(34), A(33) => A(33), 
                           A(32) => A(32), A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => n2, SUM(43) => S(43), 
                           SUM(42) => S(42), SUM(41) => S(41), SUM(40) => S(40)
                           , SUM(39) => S(39), SUM(38) => S(38), SUM(37) => 
                           S(37), SUM(36) => S(36), SUM(35) => S(35), SUM(34) 
                           => S(34), SUM(33) => S(33), SUM(32) => S(32), 
                           SUM(31) => S(31), SUM(30) => S(30), SUM(29) => S(29)
                           , SUM(28) => S(28), SUM(27) => S(27), SUM(26) => 
                           S(26), SUM(25) => S(25), SUM(24) => S(24), SUM(23) 
                           => S(23), SUM(22) => S(22), SUM(21) => S(21), 
                           SUM(20) => S(20), SUM(19) => S(19), SUM(18) => S(18)
                           , SUM(17) => S(17), SUM(16) => S(16), SUM(15) => 
                           S(15), SUM(14) => S(14), SUM(13) => S(13), SUM(12) 
                           => S(12), SUM(11) => S(11), SUM(10) => S(10), SUM(9)
                           => S(9), SUM(8) => S(8), SUM(7) => S(7), SUM(6) => 
                           S(6), SUM(5) => S(5), SUM(4) => S(4), SUM(3) => S(3)
                           , SUM(2) => S(2), SUM(1) => S(1), SUM(0) => S(0), CO
                           => n_1075);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT42 is

   port( A, B : in std_logic_vector (41 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (41 downto 0);  Co : out std_logic);

end RCA_NBIT42;

architecture SYN_DIRECT of RCA_NBIT42 is

   component RCA_NBIT42_DW01_add_0
      port( A, B : in std_logic_vector (41 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (41 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1076 : std_logic;

begin
   
   Co <= '0';
   n2 <= '0';
   add_95 : RCA_NBIT42_DW01_add_0 port map( A(41) => A(41), A(40) => A(40), 
                           A(39) => A(39), A(38) => A(38), A(37) => A(37), 
                           A(36) => A(36), A(35) => A(35), A(34) => A(34), 
                           A(33) => A(33), A(32) => A(32), A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(41) => B(41), 
                           B(40) => B(40), B(39) => B(39), B(38) => B(38), 
                           B(37) => B(37), B(36) => B(36), B(35) => B(35), 
                           B(34) => B(34), B(33) => B(33), B(32) => B(32), 
                           B(31) => B(31), B(30) => B(30), B(29) => B(29), 
                           B(28) => B(28), B(27) => B(27), B(26) => B(26), 
                           B(25) => B(25), B(24) => B(24), B(23) => B(23), 
                           B(22) => B(22), B(21) => B(21), B(20) => B(20), 
                           B(19) => B(19), B(18) => B(18), B(17) => B(17), 
                           B(16) => B(16), B(15) => B(15), B(14) => B(14), 
                           B(13) => B(13), B(12) => B(12), B(11) => B(11), 
                           B(10) => B(10), B(9) => B(9), B(8) => B(8), B(7) => 
                           B(7), B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3)
                           => B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), 
                           CI => n2, SUM(41) => S(41), SUM(40) => S(40), 
                           SUM(39) => S(39), SUM(38) => S(38), SUM(37) => S(37)
                           , SUM(36) => S(36), SUM(35) => S(35), SUM(34) => 
                           S(34), SUM(33) => S(33), SUM(32) => S(32), SUM(31) 
                           => S(31), SUM(30) => S(30), SUM(29) => S(29), 
                           SUM(28) => S(28), SUM(27) => S(27), SUM(26) => S(26)
                           , SUM(25) => S(25), SUM(24) => S(24), SUM(23) => 
                           S(23), SUM(22) => S(22), SUM(21) => S(21), SUM(20) 
                           => S(20), SUM(19) => S(19), SUM(18) => S(18), 
                           SUM(17) => S(17), SUM(16) => S(16), SUM(15) => S(15)
                           , SUM(14) => S(14), SUM(13) => S(13), SUM(12) => 
                           S(12), SUM(11) => S(11), SUM(10) => S(10), SUM(9) =>
                           S(9), SUM(8) => S(8), SUM(7) => S(7), SUM(6) => S(6)
                           , SUM(5) => S(5), SUM(4) => S(4), SUM(3) => S(3), 
                           SUM(2) => S(2), SUM(1) => S(1), SUM(0) => S(0), CO 
                           => n_1076);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT40 is

   port( A, B : in std_logic_vector (39 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (39 downto 0);  Co : out std_logic);

end RCA_NBIT40;

architecture SYN_DIRECT of RCA_NBIT40 is

   component RCA_NBIT40_DW01_add_0
      port( A, B : in std_logic_vector (39 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (39 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1077 : std_logic;

begin
   
   Co <= '0';
   n2 <= '0';
   add_95 : RCA_NBIT40_DW01_add_0 port map( A(39) => A(39), A(38) => A(38), 
                           A(37) => A(37), A(36) => A(36), A(35) => A(35), 
                           A(34) => A(34), A(33) => A(33), A(32) => A(32), 
                           A(31) => A(31), A(30) => A(30), A(29) => A(29), 
                           A(28) => A(28), A(27) => A(27), A(26) => A(26), 
                           A(25) => A(25), A(24) => A(24), A(23) => A(23), 
                           A(22) => A(22), A(21) => A(21), A(20) => A(20), 
                           A(19) => A(19), A(18) => A(18), A(17) => A(17), 
                           A(16) => A(16), A(15) => A(15), A(14) => A(14), 
                           A(13) => A(13), A(12) => A(12), A(11) => A(11), 
                           A(10) => A(10), A(9) => A(9), A(8) => A(8), A(7) => 
                           A(7), A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3)
                           => A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(39) => B(39), B(38) => B(38), B(37) => B(37), 
                           B(36) => B(36), B(35) => B(35), B(34) => B(34), 
                           B(33) => B(33), B(32) => B(32), B(31) => B(31), 
                           B(30) => B(30), B(29) => B(29), B(28) => B(28), 
                           B(27) => B(27), B(26) => B(26), B(25) => B(25), 
                           B(24) => B(24), B(23) => B(23), B(22) => B(22), 
                           B(21) => B(21), B(20) => B(20), B(19) => B(19), 
                           B(18) => B(18), B(17) => B(17), B(16) => B(16), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => B(0), CI => n2, SUM(39) 
                           => S(39), SUM(38) => S(38), SUM(37) => S(37), 
                           SUM(36) => S(36), SUM(35) => S(35), SUM(34) => S(34)
                           , SUM(33) => S(33), SUM(32) => S(32), SUM(31) => 
                           S(31), SUM(30) => S(30), SUM(29) => S(29), SUM(28) 
                           => S(28), SUM(27) => S(27), SUM(26) => S(26), 
                           SUM(25) => S(25), SUM(24) => S(24), SUM(23) => S(23)
                           , SUM(22) => S(22), SUM(21) => S(21), SUM(20) => 
                           S(20), SUM(19) => S(19), SUM(18) => S(18), SUM(17) 
                           => S(17), SUM(16) => S(16), SUM(15) => S(15), 
                           SUM(14) => S(14), SUM(13) => S(13), SUM(12) => S(12)
                           , SUM(11) => S(11), SUM(10) => S(10), SUM(9) => S(9)
                           , SUM(8) => S(8), SUM(7) => S(7), SUM(6) => S(6), 
                           SUM(5) => S(5), SUM(4) => S(4), SUM(3) => S(3), 
                           SUM(2) => S(2), SUM(1) => S(1), SUM(0) => S(0), CO 
                           => n_1077);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT38 is

   port( A, B : in std_logic_vector (37 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (37 downto 0);  Co : out std_logic);

end RCA_NBIT38;

architecture SYN_DIRECT of RCA_NBIT38 is

   component RCA_NBIT38_DW01_add_0
      port( A, B : in std_logic_vector (37 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (37 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1078 : std_logic;

begin
   
   Co <= '0';
   n2 <= '0';
   add_95 : RCA_NBIT38_DW01_add_0 port map( A(37) => A(37), A(36) => A(36), 
                           A(35) => A(35), A(34) => A(34), A(33) => A(33), 
                           A(32) => A(32), A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => n2, SUM(37) => S(37), 
                           SUM(36) => S(36), SUM(35) => S(35), SUM(34) => S(34)
                           , SUM(33) => S(33), SUM(32) => S(32), SUM(31) => 
                           S(31), SUM(30) => S(30), SUM(29) => S(29), SUM(28) 
                           => S(28), SUM(27) => S(27), SUM(26) => S(26), 
                           SUM(25) => S(25), SUM(24) => S(24), SUM(23) => S(23)
                           , SUM(22) => S(22), SUM(21) => S(21), SUM(20) => 
                           S(20), SUM(19) => S(19), SUM(18) => S(18), SUM(17) 
                           => S(17), SUM(16) => S(16), SUM(15) => S(15), 
                           SUM(14) => S(14), SUM(13) => S(13), SUM(12) => S(12)
                           , SUM(11) => S(11), SUM(10) => S(10), SUM(9) => S(9)
                           , SUM(8) => S(8), SUM(7) => S(7), SUM(6) => S(6), 
                           SUM(5) => S(5), SUM(4) => S(4), SUM(3) => S(3), 
                           SUM(2) => S(2), SUM(1) => S(1), SUM(0) => S(0), CO 
                           => n_1078);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity RCA_NBIT36 is

   port( A, B : in std_logic_vector (35 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (35 downto 0);  Co : out std_logic);

end RCA_NBIT36;

architecture SYN_DIRECT of RCA_NBIT36 is

   component RCA_NBIT36_DW01_add_0
      port( A, B : in std_logic_vector (35 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (35 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1079 : std_logic;

begin
   
   Co <= '0';
   n2 <= '0';
   add_95 : RCA_NBIT36_DW01_add_0 port map( A(35) => A(35), A(34) => A(34), 
                           A(33) => A(33), A(32) => A(32), A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(35) => B(35), 
                           B(34) => B(34), B(33) => B(33), B(32) => B(32), 
                           B(31) => B(31), B(30) => B(30), B(29) => B(29), 
                           B(28) => B(28), B(27) => B(27), B(26) => B(26), 
                           B(25) => B(25), B(24) => B(24), B(23) => B(23), 
                           B(22) => B(22), B(21) => B(21), B(20) => B(20), 
                           B(19) => B(19), B(18) => B(18), B(17) => B(17), 
                           B(16) => B(16), B(15) => B(15), B(14) => B(14), 
                           B(13) => B(13), B(12) => B(12), B(11) => B(11), 
                           B(10) => B(10), B(9) => B(9), B(8) => B(8), B(7) => 
                           B(7), B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3)
                           => B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), 
                           CI => n2, SUM(35) => S(35), SUM(34) => S(34), 
                           SUM(33) => S(33), SUM(32) => S(32), SUM(31) => S(31)
                           , SUM(30) => S(30), SUM(29) => S(29), SUM(28) => 
                           S(28), SUM(27) => S(27), SUM(26) => S(26), SUM(25) 
                           => S(25), SUM(24) => S(24), SUM(23) => S(23), 
                           SUM(22) => S(22), SUM(21) => S(21), SUM(20) => S(20)
                           , SUM(19) => S(19), SUM(18) => S(18), SUM(17) => 
                           S(17), SUM(16) => S(16), SUM(15) => S(15), SUM(14) 
                           => S(14), SUM(13) => S(13), SUM(12) => S(12), 
                           SUM(11) => S(11), SUM(10) => S(10), SUM(9) => S(9), 
                           SUM(8) => S(8), SUM(7) => S(7), SUM(6) => S(6), 
                           SUM(5) => S(5), SUM(4) => S(4), SUM(3) => S(3), 
                           SUM(2) => S(2), SUM(1) => S(1), SUM(0) => S(0), CO 
                           => n_1079);

end SYN_DIRECT;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT64_i30 is

   port( A_s, A_ns, B : in std_logic_vector (63 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (63 downto 0));

end BOOTHENC_NBIT64_i30;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT64_i30 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, O_63_port, O_62_port, O_61_port, O_60_port, O_59_port,
      O_58_port, O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, 
      O_52_port, O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, 
      O_46_port, O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, 
      O_40_port, O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, 
      O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, 
      O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, 
      O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, 
      O_16_port, O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, 
      O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, 
      O_3_port, O_2_port, O_1_port, n890, n891, n892, n893, n894, n895, n896, 
      n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, 
      n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, 
      n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, 
      n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, 
      n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, 
      n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, 
      n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, 
      n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, 
      n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, 
      n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, 
      n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, 
      n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, 
      n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, 
      n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, 
      n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, 
      n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, 
      n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, 
      n1084 : std_logic;

begin
   O <= ( O_63_port, O_62_port, O_61_port, O_60_port, O_59_port, O_58_port, 
      O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, O_52_port, 
      O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, O_46_port, 
      O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, O_40_port, 
      O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, 
      O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, 
      O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, 
      O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, O_16_port, 
      O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, O_10_port, 
      O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, O_3_port, 
      O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(61), A_s(60), A_s(59), A_s(58), A_s(57), A_s(56), A_s(55), 
      A_s(54), A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), 
      A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), 
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   A_nso <= ( A_ns(61), A_ns(60), A_ns(59), A_ns(58), A_ns(57), A_ns(56), 
      A_ns(55), A_ns(54), A_ns(53), A_ns(52), A_ns(51), A_ns(50), A_ns(49), 
      A_ns(48), A_ns(47), A_ns(46), A_ns(45), A_ns(44), A_ns(43), A_ns(42), 
      A_ns(41), A_ns(40), A_ns(39), A_ns(38), A_ns(37), A_ns(36), A_ns(35), 
      A_ns(34), A_ns(33), A_ns(32), A_ns(31), A_ns(30), A_ns(29), A_ns(28), 
      A_ns(27), A_ns(26), A_ns(25), A_ns(24), A_ns(23), A_ns(22), A_ns(21), 
      A_ns(20), A_ns(19), A_ns(18), A_ns(17), A_ns(16), A_ns(15), A_ns(14), 
      A_ns(13), A_ns(12), A_ns(11), A_ns(10), A_ns(9), A_ns(8), A_ns(7), 
      A_ns(6), A_ns(5), A_ns(4), A_ns(3), A_ns(2), A_ns(1), A_ns(0), 
      X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : AND3_X1 port map( A1 => B(30), A2 => n1084, A3 => B(29), ZN => n890);
   U3 : INV_X4 port map( A => n890, ZN => n891);
   U4 : INV_X4 port map( A => n1051, ZN => n897);
   U5 : INV_X4 port map( A => n1052, ZN => n896);
   U6 : OR3_X4 port map( A1 => B(29), A2 => B(30), A3 => n1084, ZN => n892);
   U7 : OAI221_X1 port map( B1 => n892, B2 => n893, C1 => n891, C2 => n894, A 
                           => n895, ZN => O_9_port);
   U8 : AOI22_X1 port map( A1 => A_ns(8), A2 => n896, B1 => A_s(8), B2 => n897,
                           ZN => n895);
   U9 : INV_X1 port map( A => A_s(7), ZN => n894);
   U10 : INV_X1 port map( A => A_ns(7), ZN => n893);
   U11 : OAI221_X1 port map( B1 => n892, B2 => n898, C1 => n891, C2 => n899, A 
                           => n900, ZN => O_8_port);
   U12 : AOI22_X1 port map( A1 => A_ns(7), A2 => n896, B1 => A_s(7), B2 => n897
                           , ZN => n900);
   U13 : INV_X1 port map( A => A_s(6), ZN => n899);
   U14 : INV_X1 port map( A => A_ns(6), ZN => n898);
   U15 : OAI221_X1 port map( B1 => n892, B2 => n901, C1 => n891, C2 => n902, A 
                           => n903, ZN => O_7_port);
   U16 : AOI22_X1 port map( A1 => A_ns(6), A2 => n896, B1 => A_s(6), B2 => n897
                           , ZN => n903);
   U17 : INV_X1 port map( A => A_s(5), ZN => n902);
   U18 : INV_X1 port map( A => A_ns(5), ZN => n901);
   U19 : OAI221_X1 port map( B1 => n892, B2 => n904, C1 => n891, C2 => n905, A 
                           => n906, ZN => O_6_port);
   U20 : AOI22_X1 port map( A1 => A_ns(5), A2 => n896, B1 => A_s(5), B2 => n897
                           , ZN => n906);
   U21 : INV_X1 port map( A => A_s(4), ZN => n905);
   U22 : INV_X1 port map( A => A_ns(4), ZN => n904);
   U23 : OAI221_X1 port map( B1 => n892, B2 => n907, C1 => n891, C2 => n908, A 
                           => n909, ZN => O_63_port);
   U24 : AOI22_X1 port map( A1 => A_ns(62), A2 => n896, B1 => A_s(62), B2 => 
                           n897, ZN => n909);
   U25 : INV_X1 port map( A => A_s(61), ZN => n908);
   U26 : INV_X1 port map( A => A_ns(61), ZN => n907);
   U27 : OAI221_X1 port map( B1 => n892, B2 => n910, C1 => n891, C2 => n911, A 
                           => n912, ZN => O_62_port);
   U28 : AOI22_X1 port map( A1 => A_ns(61), A2 => n896, B1 => A_s(61), B2 => 
                           n897, ZN => n912);
   U29 : INV_X1 port map( A => A_s(60), ZN => n911);
   U30 : INV_X1 port map( A => A_ns(60), ZN => n910);
   U31 : OAI221_X1 port map( B1 => n892, B2 => n913, C1 => n891, C2 => n914, A 
                           => n915, ZN => O_61_port);
   U32 : AOI22_X1 port map( A1 => A_ns(60), A2 => n896, B1 => A_s(60), B2 => 
                           n897, ZN => n915);
   U33 : INV_X1 port map( A => A_s(59), ZN => n914);
   U34 : INV_X1 port map( A => A_ns(59), ZN => n913);
   U35 : OAI221_X1 port map( B1 => n892, B2 => n916, C1 => n891, C2 => n917, A 
                           => n918, ZN => O_60_port);
   U36 : AOI22_X1 port map( A1 => A_ns(59), A2 => n896, B1 => A_s(59), B2 => 
                           n897, ZN => n918);
   U37 : INV_X1 port map( A => A_s(58), ZN => n917);
   U38 : INV_X1 port map( A => A_ns(58), ZN => n916);
   U39 : OAI221_X1 port map( B1 => n892, B2 => n919, C1 => n891, C2 => n920, A 
                           => n921, ZN => O_5_port);
   U40 : AOI22_X1 port map( A1 => A_ns(4), A2 => n896, B1 => A_s(4), B2 => n897
                           , ZN => n921);
   U41 : INV_X1 port map( A => A_s(3), ZN => n920);
   U42 : INV_X1 port map( A => A_ns(3), ZN => n919);
   U43 : OAI221_X1 port map( B1 => n892, B2 => n922, C1 => n891, C2 => n923, A 
                           => n924, ZN => O_59_port);
   U44 : AOI22_X1 port map( A1 => A_ns(58), A2 => n896, B1 => A_s(58), B2 => 
                           n897, ZN => n924);
   U45 : INV_X1 port map( A => A_s(57), ZN => n923);
   U46 : INV_X1 port map( A => A_ns(57), ZN => n922);
   U47 : OAI221_X1 port map( B1 => n892, B2 => n925, C1 => n891, C2 => n926, A 
                           => n927, ZN => O_58_port);
   U48 : AOI22_X1 port map( A1 => A_ns(57), A2 => n896, B1 => A_s(57), B2 => 
                           n897, ZN => n927);
   U49 : INV_X1 port map( A => A_s(56), ZN => n926);
   U50 : INV_X1 port map( A => A_ns(56), ZN => n925);
   U51 : OAI221_X1 port map( B1 => n892, B2 => n928, C1 => n891, C2 => n929, A 
                           => n930, ZN => O_57_port);
   U52 : AOI22_X1 port map( A1 => A_ns(56), A2 => n896, B1 => A_s(56), B2 => 
                           n897, ZN => n930);
   U53 : INV_X1 port map( A => A_s(55), ZN => n929);
   U54 : INV_X1 port map( A => A_ns(55), ZN => n928);
   U55 : OAI221_X1 port map( B1 => n892, B2 => n931, C1 => n891, C2 => n932, A 
                           => n933, ZN => O_56_port);
   U56 : AOI22_X1 port map( A1 => A_ns(55), A2 => n896, B1 => A_s(55), B2 => 
                           n897, ZN => n933);
   U57 : INV_X1 port map( A => A_s(54), ZN => n932);
   U58 : INV_X1 port map( A => A_ns(54), ZN => n931);
   U59 : OAI221_X1 port map( B1 => n892, B2 => n934, C1 => n891, C2 => n935, A 
                           => n936, ZN => O_55_port);
   U60 : AOI22_X1 port map( A1 => A_ns(54), A2 => n896, B1 => A_s(54), B2 => 
                           n897, ZN => n936);
   U61 : INV_X1 port map( A => A_s(53), ZN => n935);
   U62 : INV_X1 port map( A => A_ns(53), ZN => n934);
   U63 : OAI221_X1 port map( B1 => n892, B2 => n937, C1 => n891, C2 => n938, A 
                           => n939, ZN => O_54_port);
   U64 : AOI22_X1 port map( A1 => A_ns(53), A2 => n896, B1 => A_s(53), B2 => 
                           n897, ZN => n939);
   U65 : INV_X1 port map( A => A_s(52), ZN => n938);
   U66 : INV_X1 port map( A => A_ns(52), ZN => n937);
   U67 : OAI221_X1 port map( B1 => n892, B2 => n940, C1 => n891, C2 => n941, A 
                           => n942, ZN => O_53_port);
   U68 : AOI22_X1 port map( A1 => A_ns(52), A2 => n896, B1 => A_s(52), B2 => 
                           n897, ZN => n942);
   U69 : INV_X1 port map( A => A_s(51), ZN => n941);
   U70 : INV_X1 port map( A => A_ns(51), ZN => n940);
   U71 : OAI221_X1 port map( B1 => n892, B2 => n943, C1 => n891, C2 => n944, A 
                           => n945, ZN => O_52_port);
   U72 : AOI22_X1 port map( A1 => A_ns(51), A2 => n896, B1 => A_s(51), B2 => 
                           n897, ZN => n945);
   U73 : INV_X1 port map( A => A_s(50), ZN => n944);
   U74 : INV_X1 port map( A => A_ns(50), ZN => n943);
   U75 : OAI221_X1 port map( B1 => n892, B2 => n946, C1 => n891, C2 => n947, A 
                           => n948, ZN => O_51_port);
   U76 : AOI22_X1 port map( A1 => A_ns(50), A2 => n896, B1 => A_s(50), B2 => 
                           n897, ZN => n948);
   U77 : INV_X1 port map( A => A_s(49), ZN => n947);
   U78 : INV_X1 port map( A => A_ns(49), ZN => n946);
   U79 : OAI221_X1 port map( B1 => n892, B2 => n949, C1 => n891, C2 => n950, A 
                           => n951, ZN => O_50_port);
   U80 : AOI22_X1 port map( A1 => A_ns(49), A2 => n896, B1 => A_s(49), B2 => 
                           n897, ZN => n951);
   U81 : INV_X1 port map( A => A_s(48), ZN => n950);
   U82 : INV_X1 port map( A => A_ns(48), ZN => n949);
   U83 : OAI221_X1 port map( B1 => n892, B2 => n952, C1 => n891, C2 => n953, A 
                           => n954, ZN => O_4_port);
   U84 : AOI22_X1 port map( A1 => A_ns(3), A2 => n896, B1 => A_s(3), B2 => n897
                           , ZN => n954);
   U85 : INV_X1 port map( A => A_s(2), ZN => n953);
   U86 : INV_X1 port map( A => A_ns(2), ZN => n952);
   U87 : OAI221_X1 port map( B1 => n892, B2 => n955, C1 => n891, C2 => n956, A 
                           => n957, ZN => O_49_port);
   U88 : AOI22_X1 port map( A1 => A_ns(48), A2 => n896, B1 => A_s(48), B2 => 
                           n897, ZN => n957);
   U89 : INV_X1 port map( A => A_s(47), ZN => n956);
   U90 : INV_X1 port map( A => A_ns(47), ZN => n955);
   U91 : OAI221_X1 port map( B1 => n892, B2 => n958, C1 => n891, C2 => n959, A 
                           => n960, ZN => O_48_port);
   U92 : AOI22_X1 port map( A1 => A_ns(47), A2 => n896, B1 => A_s(47), B2 => 
                           n897, ZN => n960);
   U93 : INV_X1 port map( A => A_s(46), ZN => n959);
   U94 : INV_X1 port map( A => A_ns(46), ZN => n958);
   U95 : OAI221_X1 port map( B1 => n892, B2 => n961, C1 => n891, C2 => n962, A 
                           => n963, ZN => O_47_port);
   U96 : AOI22_X1 port map( A1 => A_ns(46), A2 => n896, B1 => A_s(46), B2 => 
                           n897, ZN => n963);
   U97 : INV_X1 port map( A => A_s(45), ZN => n962);
   U98 : INV_X1 port map( A => A_ns(45), ZN => n961);
   U99 : OAI221_X1 port map( B1 => n892, B2 => n964, C1 => n891, C2 => n965, A 
                           => n966, ZN => O_46_port);
   U100 : AOI22_X1 port map( A1 => A_ns(45), A2 => n896, B1 => A_s(45), B2 => 
                           n897, ZN => n966);
   U101 : INV_X1 port map( A => A_s(44), ZN => n965);
   U102 : INV_X1 port map( A => A_ns(44), ZN => n964);
   U103 : OAI221_X1 port map( B1 => n892, B2 => n967, C1 => n891, C2 => n968, A
                           => n969, ZN => O_45_port);
   U104 : AOI22_X1 port map( A1 => A_ns(44), A2 => n896, B1 => A_s(44), B2 => 
                           n897, ZN => n969);
   U105 : INV_X1 port map( A => A_s(43), ZN => n968);
   U106 : INV_X1 port map( A => A_ns(43), ZN => n967);
   U107 : OAI221_X1 port map( B1 => n892, B2 => n970, C1 => n891, C2 => n971, A
                           => n972, ZN => O_44_port);
   U108 : AOI22_X1 port map( A1 => A_ns(43), A2 => n896, B1 => A_s(43), B2 => 
                           n897, ZN => n972);
   U109 : INV_X1 port map( A => A_s(42), ZN => n971);
   U110 : INV_X1 port map( A => A_ns(42), ZN => n970);
   U111 : OAI221_X1 port map( B1 => n892, B2 => n973, C1 => n891, C2 => n974, A
                           => n975, ZN => O_43_port);
   U112 : AOI22_X1 port map( A1 => A_ns(42), A2 => n896, B1 => A_s(42), B2 => 
                           n897, ZN => n975);
   U113 : INV_X1 port map( A => A_s(41), ZN => n974);
   U114 : INV_X1 port map( A => A_ns(41), ZN => n973);
   U115 : OAI221_X1 port map( B1 => n892, B2 => n976, C1 => n891, C2 => n977, A
                           => n978, ZN => O_42_port);
   U116 : AOI22_X1 port map( A1 => A_ns(41), A2 => n896, B1 => A_s(41), B2 => 
                           n897, ZN => n978);
   U117 : INV_X1 port map( A => A_s(40), ZN => n977);
   U118 : INV_X1 port map( A => A_ns(40), ZN => n976);
   U119 : OAI221_X1 port map( B1 => n892, B2 => n979, C1 => n891, C2 => n980, A
                           => n981, ZN => O_41_port);
   U120 : AOI22_X1 port map( A1 => A_ns(40), A2 => n896, B1 => A_s(40), B2 => 
                           n897, ZN => n981);
   U121 : INV_X1 port map( A => A_s(39), ZN => n980);
   U122 : INV_X1 port map( A => A_ns(39), ZN => n979);
   U123 : OAI221_X1 port map( B1 => n892, B2 => n982, C1 => n891, C2 => n983, A
                           => n984, ZN => O_40_port);
   U124 : AOI22_X1 port map( A1 => A_ns(39), A2 => n896, B1 => A_s(39), B2 => 
                           n897, ZN => n984);
   U125 : INV_X1 port map( A => A_s(38), ZN => n983);
   U126 : INV_X1 port map( A => A_ns(38), ZN => n982);
   U127 : OAI221_X1 port map( B1 => n892, B2 => n985, C1 => n891, C2 => n986, A
                           => n987, ZN => O_3_port);
   U128 : AOI22_X1 port map( A1 => A_ns(2), A2 => n896, B1 => A_s(2), B2 => 
                           n897, ZN => n987);
   U129 : INV_X1 port map( A => A_s(1), ZN => n986);
   U130 : INV_X1 port map( A => A_ns(1), ZN => n985);
   U131 : OAI221_X1 port map( B1 => n892, B2 => n988, C1 => n891, C2 => n989, A
                           => n990, ZN => O_39_port);
   U132 : AOI22_X1 port map( A1 => A_ns(38), A2 => n896, B1 => A_s(38), B2 => 
                           n897, ZN => n990);
   U133 : INV_X1 port map( A => A_s(37), ZN => n989);
   U134 : INV_X1 port map( A => A_ns(37), ZN => n988);
   U135 : OAI221_X1 port map( B1 => n892, B2 => n991, C1 => n891, C2 => n992, A
                           => n993, ZN => O_38_port);
   U136 : AOI22_X1 port map( A1 => A_ns(37), A2 => n896, B1 => A_s(37), B2 => 
                           n897, ZN => n993);
   U137 : INV_X1 port map( A => A_s(36), ZN => n992);
   U138 : INV_X1 port map( A => A_ns(36), ZN => n991);
   U139 : OAI221_X1 port map( B1 => n892, B2 => n994, C1 => n891, C2 => n995, A
                           => n996, ZN => O_37_port);
   U140 : AOI22_X1 port map( A1 => A_ns(36), A2 => n896, B1 => A_s(36), B2 => 
                           n897, ZN => n996);
   U141 : INV_X1 port map( A => A_s(35), ZN => n995);
   U142 : INV_X1 port map( A => A_ns(35), ZN => n994);
   U143 : OAI221_X1 port map( B1 => n892, B2 => n997, C1 => n891, C2 => n998, A
                           => n999, ZN => O_36_port);
   U144 : AOI22_X1 port map( A1 => A_ns(35), A2 => n896, B1 => A_s(35), B2 => 
                           n897, ZN => n999);
   U145 : INV_X1 port map( A => A_s(34), ZN => n998);
   U146 : INV_X1 port map( A => A_ns(34), ZN => n997);
   U147 : OAI221_X1 port map( B1 => n892, B2 => n1000, C1 => n891, C2 => n1001,
                           A => n1002, ZN => O_35_port);
   U148 : AOI22_X1 port map( A1 => A_ns(34), A2 => n896, B1 => A_s(34), B2 => 
                           n897, ZN => n1002);
   U149 : INV_X1 port map( A => A_s(33), ZN => n1001);
   U150 : INV_X1 port map( A => A_ns(33), ZN => n1000);
   U151 : OAI221_X1 port map( B1 => n892, B2 => n1003, C1 => n891, C2 => n1004,
                           A => n1005, ZN => O_34_port);
   U152 : AOI22_X1 port map( A1 => A_ns(33), A2 => n896, B1 => A_s(33), B2 => 
                           n897, ZN => n1005);
   U153 : INV_X1 port map( A => A_s(32), ZN => n1004);
   U154 : INV_X1 port map( A => A_ns(32), ZN => n1003);
   U155 : OAI221_X1 port map( B1 => n892, B2 => n1006, C1 => n891, C2 => n1007,
                           A => n1008, ZN => O_33_port);
   U156 : AOI22_X1 port map( A1 => A_ns(32), A2 => n896, B1 => A_s(32), B2 => 
                           n897, ZN => n1008);
   U157 : INV_X1 port map( A => A_s(31), ZN => n1007);
   U158 : INV_X1 port map( A => A_ns(31), ZN => n1006);
   U159 : OAI221_X1 port map( B1 => n892, B2 => n1009, C1 => n891, C2 => n1010,
                           A => n1011, ZN => O_32_port);
   U160 : AOI22_X1 port map( A1 => A_ns(31), A2 => n896, B1 => A_s(31), B2 => 
                           n897, ZN => n1011);
   U161 : INV_X1 port map( A => A_s(30), ZN => n1010);
   U162 : INV_X1 port map( A => A_ns(30), ZN => n1009);
   U163 : OAI221_X1 port map( B1 => n892, B2 => n1012, C1 => n891, C2 => n1013,
                           A => n1014, ZN => O_31_port);
   U164 : AOI22_X1 port map( A1 => A_ns(30), A2 => n896, B1 => A_s(30), B2 => 
                           n897, ZN => n1014);
   U165 : INV_X1 port map( A => A_s(29), ZN => n1013);
   U166 : INV_X1 port map( A => A_ns(29), ZN => n1012);
   U167 : OAI221_X1 port map( B1 => n892, B2 => n1015, C1 => n891, C2 => n1016,
                           A => n1017, ZN => O_30_port);
   U168 : AOI22_X1 port map( A1 => A_ns(29), A2 => n896, B1 => A_s(29), B2 => 
                           n897, ZN => n1017);
   U169 : INV_X1 port map( A => A_s(28), ZN => n1016);
   U170 : INV_X1 port map( A => A_ns(28), ZN => n1015);
   U171 : OAI221_X1 port map( B1 => n892, B2 => n1018, C1 => n891, C2 => n1019,
                           A => n1020, ZN => O_2_port);
   U172 : AOI22_X1 port map( A1 => A_ns(1), A2 => n896, B1 => A_s(1), B2 => 
                           n897, ZN => n1020);
   U173 : OAI221_X1 port map( B1 => n892, B2 => n1021, C1 => n891, C2 => n1022,
                           A => n1023, ZN => O_29_port);
   U174 : AOI22_X1 port map( A1 => A_ns(28), A2 => n896, B1 => A_s(28), B2 => 
                           n897, ZN => n1023);
   U175 : INV_X1 port map( A => A_s(27), ZN => n1022);
   U176 : INV_X1 port map( A => A_ns(27), ZN => n1021);
   U177 : OAI221_X1 port map( B1 => n892, B2 => n1024, C1 => n891, C2 => n1025,
                           A => n1026, ZN => O_28_port);
   U178 : AOI22_X1 port map( A1 => A_ns(27), A2 => n896, B1 => A_s(27), B2 => 
                           n897, ZN => n1026);
   U179 : INV_X1 port map( A => A_s(26), ZN => n1025);
   U180 : INV_X1 port map( A => A_ns(26), ZN => n1024);
   U181 : OAI221_X1 port map( B1 => n892, B2 => n1027, C1 => n891, C2 => n1028,
                           A => n1029, ZN => O_27_port);
   U182 : AOI22_X1 port map( A1 => A_ns(26), A2 => n896, B1 => A_s(26), B2 => 
                           n897, ZN => n1029);
   U183 : INV_X1 port map( A => A_s(25), ZN => n1028);
   U184 : INV_X1 port map( A => A_ns(25), ZN => n1027);
   U185 : OAI221_X1 port map( B1 => n892, B2 => n1030, C1 => n891, C2 => n1031,
                           A => n1032, ZN => O_26_port);
   U186 : AOI22_X1 port map( A1 => A_ns(25), A2 => n896, B1 => A_s(25), B2 => 
                           n897, ZN => n1032);
   U187 : INV_X1 port map( A => A_s(24), ZN => n1031);
   U188 : INV_X1 port map( A => A_ns(24), ZN => n1030);
   U189 : OAI221_X1 port map( B1 => n892, B2 => n1033, C1 => n891, C2 => n1034,
                           A => n1035, ZN => O_25_port);
   U190 : AOI22_X1 port map( A1 => A_ns(24), A2 => n896, B1 => A_s(24), B2 => 
                           n897, ZN => n1035);
   U191 : INV_X1 port map( A => A_s(23), ZN => n1034);
   U192 : INV_X1 port map( A => A_ns(23), ZN => n1033);
   U193 : OAI221_X1 port map( B1 => n892, B2 => n1036, C1 => n891, C2 => n1037,
                           A => n1038, ZN => O_24_port);
   U194 : AOI22_X1 port map( A1 => A_ns(23), A2 => n896, B1 => A_s(23), B2 => 
                           n897, ZN => n1038);
   U195 : INV_X1 port map( A => A_s(22), ZN => n1037);
   U196 : INV_X1 port map( A => A_ns(22), ZN => n1036);
   U197 : OAI221_X1 port map( B1 => n892, B2 => n1039, C1 => n891, C2 => n1040,
                           A => n1041, ZN => O_23_port);
   U198 : AOI22_X1 port map( A1 => A_ns(22), A2 => n896, B1 => A_s(22), B2 => 
                           n897, ZN => n1041);
   U199 : INV_X1 port map( A => A_s(21), ZN => n1040);
   U200 : INV_X1 port map( A => A_ns(21), ZN => n1039);
   U201 : OAI221_X1 port map( B1 => n892, B2 => n1042, C1 => n891, C2 => n1043,
                           A => n1044, ZN => O_22_port);
   U202 : AOI22_X1 port map( A1 => A_ns(21), A2 => n896, B1 => A_s(21), B2 => 
                           n897, ZN => n1044);
   U203 : INV_X1 port map( A => A_s(20), ZN => n1043);
   U204 : INV_X1 port map( A => A_ns(20), ZN => n1042);
   U205 : OAI221_X1 port map( B1 => n892, B2 => n1045, C1 => n891, C2 => n1046,
                           A => n1047, ZN => O_21_port);
   U206 : AOI22_X1 port map( A1 => A_ns(20), A2 => n896, B1 => A_s(20), B2 => 
                           n897, ZN => n1047);
   U207 : INV_X1 port map( A => A_s(19), ZN => n1046);
   U208 : INV_X1 port map( A => A_ns(19), ZN => n1045);
   U209 : OAI221_X1 port map( B1 => n892, B2 => n1048, C1 => n891, C2 => n1049,
                           A => n1050, ZN => O_20_port);
   U210 : AOI22_X1 port map( A1 => A_ns(19), A2 => n896, B1 => A_s(19), B2 => 
                           n897, ZN => n1050);
   U211 : INV_X1 port map( A => A_s(18), ZN => n1049);
   U212 : INV_X1 port map( A => A_ns(18), ZN => n1048);
   U213 : OAI22_X1 port map( A1 => n1051, A2 => n1019, B1 => n1052, B2 => n1018
                           , ZN => O_1_port);
   U214 : INV_X1 port map( A => A_ns(0), ZN => n1018);
   U215 : INV_X1 port map( A => A_s(0), ZN => n1019);
   U216 : OAI221_X1 port map( B1 => n892, B2 => n1053, C1 => n891, C2 => n1054,
                           A => n1055, ZN => O_19_port);
   U217 : AOI22_X1 port map( A1 => A_ns(18), A2 => n896, B1 => A_s(18), B2 => 
                           n897, ZN => n1055);
   U218 : INV_X1 port map( A => A_s(17), ZN => n1054);
   U219 : INV_X1 port map( A => A_ns(17), ZN => n1053);
   U220 : OAI221_X1 port map( B1 => n892, B2 => n1056, C1 => n891, C2 => n1057,
                           A => n1058, ZN => O_18_port);
   U221 : AOI22_X1 port map( A1 => A_ns(17), A2 => n896, B1 => A_s(17), B2 => 
                           n897, ZN => n1058);
   U222 : INV_X1 port map( A => A_s(16), ZN => n1057);
   U223 : INV_X1 port map( A => A_ns(16), ZN => n1056);
   U224 : OAI221_X1 port map( B1 => n892, B2 => n1059, C1 => n891, C2 => n1060,
                           A => n1061, ZN => O_17_port);
   U225 : AOI22_X1 port map( A1 => A_ns(16), A2 => n896, B1 => A_s(16), B2 => 
                           n897, ZN => n1061);
   U226 : INV_X1 port map( A => A_s(15), ZN => n1060);
   U227 : INV_X1 port map( A => A_ns(15), ZN => n1059);
   U228 : OAI221_X1 port map( B1 => n892, B2 => n1062, C1 => n891, C2 => n1063,
                           A => n1064, ZN => O_16_port);
   U229 : AOI22_X1 port map( A1 => A_ns(15), A2 => n896, B1 => A_s(15), B2 => 
                           n897, ZN => n1064);
   U230 : INV_X1 port map( A => A_s(14), ZN => n1063);
   U231 : INV_X1 port map( A => A_ns(14), ZN => n1062);
   U232 : OAI221_X1 port map( B1 => n892, B2 => n1065, C1 => n891, C2 => n1066,
                           A => n1067, ZN => O_15_port);
   U233 : AOI22_X1 port map( A1 => A_ns(14), A2 => n896, B1 => A_s(14), B2 => 
                           n897, ZN => n1067);
   U234 : INV_X1 port map( A => A_s(13), ZN => n1066);
   U235 : INV_X1 port map( A => A_ns(13), ZN => n1065);
   U236 : OAI221_X1 port map( B1 => n892, B2 => n1068, C1 => n891, C2 => n1069,
                           A => n1070, ZN => O_14_port);
   U237 : AOI22_X1 port map( A1 => A_ns(13), A2 => n896, B1 => A_s(13), B2 => 
                           n897, ZN => n1070);
   U238 : INV_X1 port map( A => A_s(12), ZN => n1069);
   U239 : INV_X1 port map( A => A_ns(12), ZN => n1068);
   U240 : OAI221_X1 port map( B1 => n892, B2 => n1071, C1 => n891, C2 => n1072,
                           A => n1073, ZN => O_13_port);
   U241 : AOI22_X1 port map( A1 => A_ns(12), A2 => n896, B1 => A_s(12), B2 => 
                           n897, ZN => n1073);
   U242 : INV_X1 port map( A => A_s(11), ZN => n1072);
   U243 : INV_X1 port map( A => A_ns(11), ZN => n1071);
   U244 : OAI221_X1 port map( B1 => n892, B2 => n1074, C1 => n891, C2 => n1075,
                           A => n1076, ZN => O_12_port);
   U245 : AOI22_X1 port map( A1 => A_ns(11), A2 => n896, B1 => A_s(11), B2 => 
                           n897, ZN => n1076);
   U246 : INV_X1 port map( A => A_s(10), ZN => n1075);
   U247 : INV_X1 port map( A => A_ns(10), ZN => n1074);
   U248 : OAI221_X1 port map( B1 => n892, B2 => n1077, C1 => n891, C2 => n1078,
                           A => n1079, ZN => O_11_port);
   U249 : AOI22_X1 port map( A1 => A_ns(10), A2 => n896, B1 => A_s(10), B2 => 
                           n897, ZN => n1079);
   U250 : INV_X1 port map( A => A_s(9), ZN => n1078);
   U251 : INV_X1 port map( A => A_ns(9), ZN => n1077);
   U252 : OAI221_X1 port map( B1 => n1080, B2 => n892, C1 => n1081, C2 => n891,
                           A => n1082, ZN => O_10_port);
   U253 : AOI22_X1 port map( A1 => A_ns(9), A2 => n896, B1 => A_s(9), B2 => 
                           n897, ZN => n1082);
   U254 : NAND2_X1 port map( A1 => n1083, A2 => n1051, ZN => n1052);
   U255 : NAND2_X1 port map( A1 => n1083, A2 => n1084, ZN => n1051);
   U256 : XOR2_X1 port map( A => B(29), B => B(30), Z => n1083);
   U257 : INV_X1 port map( A => A_s(8), ZN => n1081);
   U258 : INV_X1 port map( A => B(31), ZN => n1084);
   U259 : INV_X1 port map( A => A_ns(8), ZN => n1080);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT62_i28 is

   port( A_s, A_ns, B : in std_logic_vector (61 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (61 downto 0));

end BOOTHENC_NBIT62_i28;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT62_i28 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, O_61_port, O_60_port, O_59_port, O_58_port, O_57_port,
      O_56_port, O_55_port, O_54_port, O_53_port, O_52_port, O_51_port, 
      O_50_port, O_49_port, O_48_port, O_47_port, O_46_port, O_45_port, 
      O_44_port, O_43_port, O_42_port, O_41_port, O_40_port, O_39_port, 
      O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, O_33_port, 
      O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, O_27_port, 
      O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, O_21_port, 
      O_20_port, O_19_port, O_18_port, O_17_port, O_16_port, O_15_port, 
      O_14_port, O_13_port, O_12_port, O_11_port, O_10_port, O_9_port, O_8_port
      , O_7_port, O_6_port, O_5_port, O_4_port, O_3_port, O_2_port, O_1_port, 
      n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, 
      n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, 
      n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, 
      n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, 
      n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, 
      n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, 
      n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, 
      n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, 
      n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, 
      n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, 
      n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
      n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, 
      n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, 
      n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, 
      n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, 
      n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, 
      n1052, n1053, n1054, n1055, n1056, n1057, n1058 : std_logic;

begin
   O <= ( O_61_port, O_60_port, O_59_port, O_58_port, O_57_port, O_56_port, 
      O_55_port, O_54_port, O_53_port, O_52_port, O_51_port, O_50_port, 
      O_49_port, O_48_port, O_47_port, O_46_port, O_45_port, O_44_port, 
      O_43_port, O_42_port, O_41_port, O_40_port, O_39_port, O_38_port, 
      O_37_port, O_36_port, O_35_port, O_34_port, O_33_port, O_32_port, 
      O_31_port, O_30_port, O_29_port, O_28_port, O_27_port, O_26_port, 
      O_25_port, O_24_port, O_23_port, O_22_port, O_21_port, O_20_port, 
      O_19_port, O_18_port, O_17_port, O_16_port, O_15_port, O_14_port, 
      O_13_port, O_12_port, O_11_port, O_10_port, O_9_port, O_8_port, O_7_port,
      O_6_port, O_5_port, O_4_port, O_3_port, O_2_port, O_1_port, X_Logic0_port
      );
   A_so <= ( A_s(59), A_s(58), A_s(57), A_s(56), A_s(55), A_s(54), A_s(53), 
      A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), A_s(46), A_s(45), 
      A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), A_s(38), A_s(37), 
      A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), A_s(30), A_s(29), 
      A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), A_s(22), A_s(21), 
      A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), A_s(14), A_s(13), 
      A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), A_s(6), A_s(5), A_s(4)
      , A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, X_Logic0_port );
   A_nso <= ( A_ns(59), A_ns(58), A_ns(57), A_ns(56), A_ns(55), A_ns(54), 
      A_ns(53), A_ns(52), A_ns(51), A_ns(50), A_ns(49), A_ns(48), A_ns(47), 
      A_ns(46), A_ns(45), A_ns(44), A_ns(43), A_ns(42), A_ns(41), A_ns(40), 
      A_ns(39), A_ns(38), A_ns(37), A_ns(36), A_ns(35), A_ns(34), A_ns(33), 
      A_ns(32), A_ns(31), A_ns(30), A_ns(29), A_ns(28), A_ns(27), A_ns(26), 
      A_ns(25), A_ns(24), A_ns(23), A_ns(22), A_ns(21), A_ns(20), A_ns(19), 
      A_ns(18), A_ns(17), A_ns(16), A_ns(15), A_ns(14), A_ns(13), A_ns(12), 
      A_ns(11), A_ns(10), A_ns(9), A_ns(8), A_ns(7), A_ns(6), A_ns(5), A_ns(4),
      A_ns(3), A_ns(2), A_ns(1), A_ns(0), X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : AND3_X1 port map( A1 => B(28), A2 => n1058, A3 => B(27), ZN => n870);
   U3 : INV_X4 port map( A => n870, ZN => n871);
   U4 : INV_X4 port map( A => n1025, ZN => n877);
   U5 : INV_X4 port map( A => n1026, ZN => n876);
   U6 : OR3_X4 port map( A1 => B(27), A2 => B(28), A3 => n1058, ZN => n872);
   U7 : OAI221_X1 port map( B1 => n872, B2 => n873, C1 => n871, C2 => n874, A 
                           => n875, ZN => O_9_port);
   U8 : AOI22_X1 port map( A1 => A_ns(8), A2 => n876, B1 => A_s(8), B2 => n877,
                           ZN => n875);
   U9 : INV_X1 port map( A => A_s(7), ZN => n874);
   U10 : INV_X1 port map( A => A_ns(7), ZN => n873);
   U11 : OAI221_X1 port map( B1 => n872, B2 => n878, C1 => n871, C2 => n879, A 
                           => n880, ZN => O_8_port);
   U12 : AOI22_X1 port map( A1 => A_ns(7), A2 => n876, B1 => A_s(7), B2 => n877
                           , ZN => n880);
   U13 : INV_X1 port map( A => A_s(6), ZN => n879);
   U14 : INV_X1 port map( A => A_ns(6), ZN => n878);
   U15 : OAI221_X1 port map( B1 => n872, B2 => n881, C1 => n871, C2 => n882, A 
                           => n883, ZN => O_7_port);
   U16 : AOI22_X1 port map( A1 => A_ns(6), A2 => n876, B1 => A_s(6), B2 => n877
                           , ZN => n883);
   U17 : INV_X1 port map( A => A_s(5), ZN => n882);
   U18 : INV_X1 port map( A => A_ns(5), ZN => n881);
   U19 : OAI221_X1 port map( B1 => n872, B2 => n884, C1 => n871, C2 => n885, A 
                           => n886, ZN => O_6_port);
   U20 : AOI22_X1 port map( A1 => A_ns(5), A2 => n876, B1 => A_s(5), B2 => n877
                           , ZN => n886);
   U21 : INV_X1 port map( A => A_s(4), ZN => n885);
   U22 : INV_X1 port map( A => A_ns(4), ZN => n884);
   U23 : OAI221_X1 port map( B1 => n872, B2 => n887, C1 => n871, C2 => n888, A 
                           => n889, ZN => O_61_port);
   U24 : AOI22_X1 port map( A1 => A_ns(60), A2 => n876, B1 => A_s(60), B2 => 
                           n877, ZN => n889);
   U25 : INV_X1 port map( A => A_s(59), ZN => n888);
   U26 : INV_X1 port map( A => A_ns(59), ZN => n887);
   U27 : OAI221_X1 port map( B1 => n872, B2 => n890, C1 => n871, C2 => n891, A 
                           => n892, ZN => O_60_port);
   U28 : AOI22_X1 port map( A1 => A_ns(59), A2 => n876, B1 => A_s(59), B2 => 
                           n877, ZN => n892);
   U29 : INV_X1 port map( A => A_s(58), ZN => n891);
   U30 : INV_X1 port map( A => A_ns(58), ZN => n890);
   U31 : OAI221_X1 port map( B1 => n872, B2 => n893, C1 => n871, C2 => n894, A 
                           => n895, ZN => O_5_port);
   U32 : AOI22_X1 port map( A1 => A_ns(4), A2 => n876, B1 => A_s(4), B2 => n877
                           , ZN => n895);
   U33 : INV_X1 port map( A => A_s(3), ZN => n894);
   U34 : INV_X1 port map( A => A_ns(3), ZN => n893);
   U35 : OAI221_X1 port map( B1 => n872, B2 => n896, C1 => n871, C2 => n897, A 
                           => n898, ZN => O_59_port);
   U36 : AOI22_X1 port map( A1 => A_ns(58), A2 => n876, B1 => A_s(58), B2 => 
                           n877, ZN => n898);
   U37 : INV_X1 port map( A => A_s(57), ZN => n897);
   U38 : INV_X1 port map( A => A_ns(57), ZN => n896);
   U39 : OAI221_X1 port map( B1 => n872, B2 => n899, C1 => n871, C2 => n900, A 
                           => n901, ZN => O_58_port);
   U40 : AOI22_X1 port map( A1 => A_ns(57), A2 => n876, B1 => A_s(57), B2 => 
                           n877, ZN => n901);
   U41 : INV_X1 port map( A => A_s(56), ZN => n900);
   U42 : INV_X1 port map( A => A_ns(56), ZN => n899);
   U43 : OAI221_X1 port map( B1 => n872, B2 => n902, C1 => n871, C2 => n903, A 
                           => n904, ZN => O_57_port);
   U44 : AOI22_X1 port map( A1 => A_ns(56), A2 => n876, B1 => A_s(56), B2 => 
                           n877, ZN => n904);
   U45 : INV_X1 port map( A => A_s(55), ZN => n903);
   U46 : INV_X1 port map( A => A_ns(55), ZN => n902);
   U47 : OAI221_X1 port map( B1 => n872, B2 => n905, C1 => n871, C2 => n906, A 
                           => n907, ZN => O_56_port);
   U48 : AOI22_X1 port map( A1 => A_ns(55), A2 => n876, B1 => A_s(55), B2 => 
                           n877, ZN => n907);
   U49 : INV_X1 port map( A => A_s(54), ZN => n906);
   U50 : INV_X1 port map( A => A_ns(54), ZN => n905);
   U51 : OAI221_X1 port map( B1 => n872, B2 => n908, C1 => n871, C2 => n909, A 
                           => n910, ZN => O_55_port);
   U52 : AOI22_X1 port map( A1 => A_ns(54), A2 => n876, B1 => A_s(54), B2 => 
                           n877, ZN => n910);
   U53 : INV_X1 port map( A => A_s(53), ZN => n909);
   U54 : INV_X1 port map( A => A_ns(53), ZN => n908);
   U55 : OAI221_X1 port map( B1 => n872, B2 => n911, C1 => n871, C2 => n912, A 
                           => n913, ZN => O_54_port);
   U56 : AOI22_X1 port map( A1 => A_ns(53), A2 => n876, B1 => A_s(53), B2 => 
                           n877, ZN => n913);
   U57 : INV_X1 port map( A => A_s(52), ZN => n912);
   U58 : INV_X1 port map( A => A_ns(52), ZN => n911);
   U59 : OAI221_X1 port map( B1 => n872, B2 => n914, C1 => n871, C2 => n915, A 
                           => n916, ZN => O_53_port);
   U60 : AOI22_X1 port map( A1 => A_ns(52), A2 => n876, B1 => A_s(52), B2 => 
                           n877, ZN => n916);
   U61 : INV_X1 port map( A => A_s(51), ZN => n915);
   U62 : INV_X1 port map( A => A_ns(51), ZN => n914);
   U63 : OAI221_X1 port map( B1 => n872, B2 => n917, C1 => n871, C2 => n918, A 
                           => n919, ZN => O_52_port);
   U64 : AOI22_X1 port map( A1 => A_ns(51), A2 => n876, B1 => A_s(51), B2 => 
                           n877, ZN => n919);
   U65 : INV_X1 port map( A => A_s(50), ZN => n918);
   U66 : INV_X1 port map( A => A_ns(50), ZN => n917);
   U67 : OAI221_X1 port map( B1 => n872, B2 => n920, C1 => n871, C2 => n921, A 
                           => n922, ZN => O_51_port);
   U68 : AOI22_X1 port map( A1 => A_ns(50), A2 => n876, B1 => A_s(50), B2 => 
                           n877, ZN => n922);
   U69 : INV_X1 port map( A => A_s(49), ZN => n921);
   U70 : INV_X1 port map( A => A_ns(49), ZN => n920);
   U71 : OAI221_X1 port map( B1 => n872, B2 => n923, C1 => n871, C2 => n924, A 
                           => n925, ZN => O_50_port);
   U72 : AOI22_X1 port map( A1 => A_ns(49), A2 => n876, B1 => A_s(49), B2 => 
                           n877, ZN => n925);
   U73 : INV_X1 port map( A => A_s(48), ZN => n924);
   U74 : INV_X1 port map( A => A_ns(48), ZN => n923);
   U75 : OAI221_X1 port map( B1 => n872, B2 => n926, C1 => n871, C2 => n927, A 
                           => n928, ZN => O_4_port);
   U76 : AOI22_X1 port map( A1 => A_ns(3), A2 => n876, B1 => A_s(3), B2 => n877
                           , ZN => n928);
   U77 : INV_X1 port map( A => A_s(2), ZN => n927);
   U78 : INV_X1 port map( A => A_ns(2), ZN => n926);
   U79 : OAI221_X1 port map( B1 => n872, B2 => n929, C1 => n871, C2 => n930, A 
                           => n931, ZN => O_49_port);
   U80 : AOI22_X1 port map( A1 => A_ns(48), A2 => n876, B1 => A_s(48), B2 => 
                           n877, ZN => n931);
   U81 : INV_X1 port map( A => A_s(47), ZN => n930);
   U82 : INV_X1 port map( A => A_ns(47), ZN => n929);
   U83 : OAI221_X1 port map( B1 => n872, B2 => n932, C1 => n871, C2 => n933, A 
                           => n934, ZN => O_48_port);
   U84 : AOI22_X1 port map( A1 => A_ns(47), A2 => n876, B1 => A_s(47), B2 => 
                           n877, ZN => n934);
   U85 : INV_X1 port map( A => A_s(46), ZN => n933);
   U86 : INV_X1 port map( A => A_ns(46), ZN => n932);
   U87 : OAI221_X1 port map( B1 => n872, B2 => n935, C1 => n871, C2 => n936, A 
                           => n937, ZN => O_47_port);
   U88 : AOI22_X1 port map( A1 => A_ns(46), A2 => n876, B1 => A_s(46), B2 => 
                           n877, ZN => n937);
   U89 : INV_X1 port map( A => A_s(45), ZN => n936);
   U90 : INV_X1 port map( A => A_ns(45), ZN => n935);
   U91 : OAI221_X1 port map( B1 => n872, B2 => n938, C1 => n871, C2 => n939, A 
                           => n940, ZN => O_46_port);
   U92 : AOI22_X1 port map( A1 => A_ns(45), A2 => n876, B1 => A_s(45), B2 => 
                           n877, ZN => n940);
   U93 : INV_X1 port map( A => A_s(44), ZN => n939);
   U94 : INV_X1 port map( A => A_ns(44), ZN => n938);
   U95 : OAI221_X1 port map( B1 => n872, B2 => n941, C1 => n871, C2 => n942, A 
                           => n943, ZN => O_45_port);
   U96 : AOI22_X1 port map( A1 => A_ns(44), A2 => n876, B1 => A_s(44), B2 => 
                           n877, ZN => n943);
   U97 : INV_X1 port map( A => A_s(43), ZN => n942);
   U98 : INV_X1 port map( A => A_ns(43), ZN => n941);
   U99 : OAI221_X1 port map( B1 => n872, B2 => n944, C1 => n871, C2 => n945, A 
                           => n946, ZN => O_44_port);
   U100 : AOI22_X1 port map( A1 => A_ns(43), A2 => n876, B1 => A_s(43), B2 => 
                           n877, ZN => n946);
   U101 : INV_X1 port map( A => A_s(42), ZN => n945);
   U102 : INV_X1 port map( A => A_ns(42), ZN => n944);
   U103 : OAI221_X1 port map( B1 => n872, B2 => n947, C1 => n871, C2 => n948, A
                           => n949, ZN => O_43_port);
   U104 : AOI22_X1 port map( A1 => A_ns(42), A2 => n876, B1 => A_s(42), B2 => 
                           n877, ZN => n949);
   U105 : INV_X1 port map( A => A_s(41), ZN => n948);
   U106 : INV_X1 port map( A => A_ns(41), ZN => n947);
   U107 : OAI221_X1 port map( B1 => n872, B2 => n950, C1 => n871, C2 => n951, A
                           => n952, ZN => O_42_port);
   U108 : AOI22_X1 port map( A1 => A_ns(41), A2 => n876, B1 => A_s(41), B2 => 
                           n877, ZN => n952);
   U109 : INV_X1 port map( A => A_s(40), ZN => n951);
   U110 : INV_X1 port map( A => A_ns(40), ZN => n950);
   U111 : OAI221_X1 port map( B1 => n872, B2 => n953, C1 => n871, C2 => n954, A
                           => n955, ZN => O_41_port);
   U112 : AOI22_X1 port map( A1 => A_ns(40), A2 => n876, B1 => A_s(40), B2 => 
                           n877, ZN => n955);
   U113 : INV_X1 port map( A => A_s(39), ZN => n954);
   U114 : INV_X1 port map( A => A_ns(39), ZN => n953);
   U115 : OAI221_X1 port map( B1 => n872, B2 => n956, C1 => n871, C2 => n957, A
                           => n958, ZN => O_40_port);
   U116 : AOI22_X1 port map( A1 => A_ns(39), A2 => n876, B1 => A_s(39), B2 => 
                           n877, ZN => n958);
   U117 : INV_X1 port map( A => A_s(38), ZN => n957);
   U118 : INV_X1 port map( A => A_ns(38), ZN => n956);
   U119 : OAI221_X1 port map( B1 => n872, B2 => n959, C1 => n871, C2 => n960, A
                           => n961, ZN => O_3_port);
   U120 : AOI22_X1 port map( A1 => A_ns(2), A2 => n876, B1 => A_s(2), B2 => 
                           n877, ZN => n961);
   U121 : INV_X1 port map( A => A_s(1), ZN => n960);
   U122 : INV_X1 port map( A => A_ns(1), ZN => n959);
   U123 : OAI221_X1 port map( B1 => n872, B2 => n962, C1 => n871, C2 => n963, A
                           => n964, ZN => O_39_port);
   U124 : AOI22_X1 port map( A1 => A_ns(38), A2 => n876, B1 => A_s(38), B2 => 
                           n877, ZN => n964);
   U125 : INV_X1 port map( A => A_s(37), ZN => n963);
   U126 : INV_X1 port map( A => A_ns(37), ZN => n962);
   U127 : OAI221_X1 port map( B1 => n872, B2 => n965, C1 => n871, C2 => n966, A
                           => n967, ZN => O_38_port);
   U128 : AOI22_X1 port map( A1 => A_ns(37), A2 => n876, B1 => A_s(37), B2 => 
                           n877, ZN => n967);
   U129 : INV_X1 port map( A => A_s(36), ZN => n966);
   U130 : INV_X1 port map( A => A_ns(36), ZN => n965);
   U131 : OAI221_X1 port map( B1 => n872, B2 => n968, C1 => n871, C2 => n969, A
                           => n970, ZN => O_37_port);
   U132 : AOI22_X1 port map( A1 => A_ns(36), A2 => n876, B1 => A_s(36), B2 => 
                           n877, ZN => n970);
   U133 : INV_X1 port map( A => A_s(35), ZN => n969);
   U134 : INV_X1 port map( A => A_ns(35), ZN => n968);
   U135 : OAI221_X1 port map( B1 => n872, B2 => n971, C1 => n871, C2 => n972, A
                           => n973, ZN => O_36_port);
   U136 : AOI22_X1 port map( A1 => A_ns(35), A2 => n876, B1 => A_s(35), B2 => 
                           n877, ZN => n973);
   U137 : INV_X1 port map( A => A_s(34), ZN => n972);
   U138 : INV_X1 port map( A => A_ns(34), ZN => n971);
   U139 : OAI221_X1 port map( B1 => n872, B2 => n974, C1 => n871, C2 => n975, A
                           => n976, ZN => O_35_port);
   U140 : AOI22_X1 port map( A1 => A_ns(34), A2 => n876, B1 => A_s(34), B2 => 
                           n877, ZN => n976);
   U141 : INV_X1 port map( A => A_s(33), ZN => n975);
   U142 : INV_X1 port map( A => A_ns(33), ZN => n974);
   U143 : OAI221_X1 port map( B1 => n872, B2 => n977, C1 => n871, C2 => n978, A
                           => n979, ZN => O_34_port);
   U144 : AOI22_X1 port map( A1 => A_ns(33), A2 => n876, B1 => A_s(33), B2 => 
                           n877, ZN => n979);
   U145 : INV_X1 port map( A => A_s(32), ZN => n978);
   U146 : INV_X1 port map( A => A_ns(32), ZN => n977);
   U147 : OAI221_X1 port map( B1 => n872, B2 => n980, C1 => n871, C2 => n981, A
                           => n982, ZN => O_33_port);
   U148 : AOI22_X1 port map( A1 => A_ns(32), A2 => n876, B1 => A_s(32), B2 => 
                           n877, ZN => n982);
   U149 : INV_X1 port map( A => A_s(31), ZN => n981);
   U150 : INV_X1 port map( A => A_ns(31), ZN => n980);
   U151 : OAI221_X1 port map( B1 => n872, B2 => n983, C1 => n871, C2 => n984, A
                           => n985, ZN => O_32_port);
   U152 : AOI22_X1 port map( A1 => A_ns(31), A2 => n876, B1 => A_s(31), B2 => 
                           n877, ZN => n985);
   U153 : INV_X1 port map( A => A_s(30), ZN => n984);
   U154 : INV_X1 port map( A => A_ns(30), ZN => n983);
   U155 : OAI221_X1 port map( B1 => n872, B2 => n986, C1 => n871, C2 => n987, A
                           => n988, ZN => O_31_port);
   U156 : AOI22_X1 port map( A1 => A_ns(30), A2 => n876, B1 => A_s(30), B2 => 
                           n877, ZN => n988);
   U157 : INV_X1 port map( A => A_s(29), ZN => n987);
   U158 : INV_X1 port map( A => A_ns(29), ZN => n986);
   U159 : OAI221_X1 port map( B1 => n872, B2 => n989, C1 => n871, C2 => n990, A
                           => n991, ZN => O_30_port);
   U160 : AOI22_X1 port map( A1 => A_ns(29), A2 => n876, B1 => A_s(29), B2 => 
                           n877, ZN => n991);
   U161 : INV_X1 port map( A => A_s(28), ZN => n990);
   U162 : INV_X1 port map( A => A_ns(28), ZN => n989);
   U163 : OAI221_X1 port map( B1 => n872, B2 => n992, C1 => n871, C2 => n993, A
                           => n994, ZN => O_2_port);
   U164 : AOI22_X1 port map( A1 => A_ns(1), A2 => n876, B1 => A_s(1), B2 => 
                           n877, ZN => n994);
   U165 : OAI221_X1 port map( B1 => n872, B2 => n995, C1 => n871, C2 => n996, A
                           => n997, ZN => O_29_port);
   U166 : AOI22_X1 port map( A1 => A_ns(28), A2 => n876, B1 => A_s(28), B2 => 
                           n877, ZN => n997);
   U167 : INV_X1 port map( A => A_s(27), ZN => n996);
   U168 : INV_X1 port map( A => A_ns(27), ZN => n995);
   U169 : OAI221_X1 port map( B1 => n872, B2 => n998, C1 => n871, C2 => n999, A
                           => n1000, ZN => O_28_port);
   U170 : AOI22_X1 port map( A1 => A_ns(27), A2 => n876, B1 => A_s(27), B2 => 
                           n877, ZN => n1000);
   U171 : INV_X1 port map( A => A_s(26), ZN => n999);
   U172 : INV_X1 port map( A => A_ns(26), ZN => n998);
   U173 : OAI221_X1 port map( B1 => n872, B2 => n1001, C1 => n871, C2 => n1002,
                           A => n1003, ZN => O_27_port);
   U174 : AOI22_X1 port map( A1 => A_ns(26), A2 => n876, B1 => A_s(26), B2 => 
                           n877, ZN => n1003);
   U175 : INV_X1 port map( A => A_s(25), ZN => n1002);
   U176 : INV_X1 port map( A => A_ns(25), ZN => n1001);
   U177 : OAI221_X1 port map( B1 => n872, B2 => n1004, C1 => n871, C2 => n1005,
                           A => n1006, ZN => O_26_port);
   U178 : AOI22_X1 port map( A1 => A_ns(25), A2 => n876, B1 => A_s(25), B2 => 
                           n877, ZN => n1006);
   U179 : INV_X1 port map( A => A_s(24), ZN => n1005);
   U180 : INV_X1 port map( A => A_ns(24), ZN => n1004);
   U181 : OAI221_X1 port map( B1 => n872, B2 => n1007, C1 => n871, C2 => n1008,
                           A => n1009, ZN => O_25_port);
   U182 : AOI22_X1 port map( A1 => A_ns(24), A2 => n876, B1 => A_s(24), B2 => 
                           n877, ZN => n1009);
   U183 : INV_X1 port map( A => A_s(23), ZN => n1008);
   U184 : INV_X1 port map( A => A_ns(23), ZN => n1007);
   U185 : OAI221_X1 port map( B1 => n872, B2 => n1010, C1 => n871, C2 => n1011,
                           A => n1012, ZN => O_24_port);
   U186 : AOI22_X1 port map( A1 => A_ns(23), A2 => n876, B1 => A_s(23), B2 => 
                           n877, ZN => n1012);
   U187 : INV_X1 port map( A => A_s(22), ZN => n1011);
   U188 : INV_X1 port map( A => A_ns(22), ZN => n1010);
   U189 : OAI221_X1 port map( B1 => n872, B2 => n1013, C1 => n871, C2 => n1014,
                           A => n1015, ZN => O_23_port);
   U190 : AOI22_X1 port map( A1 => A_ns(22), A2 => n876, B1 => A_s(22), B2 => 
                           n877, ZN => n1015);
   U191 : INV_X1 port map( A => A_s(21), ZN => n1014);
   U192 : INV_X1 port map( A => A_ns(21), ZN => n1013);
   U193 : OAI221_X1 port map( B1 => n872, B2 => n1016, C1 => n871, C2 => n1017,
                           A => n1018, ZN => O_22_port);
   U194 : AOI22_X1 port map( A1 => A_ns(21), A2 => n876, B1 => A_s(21), B2 => 
                           n877, ZN => n1018);
   U195 : INV_X1 port map( A => A_s(20), ZN => n1017);
   U196 : INV_X1 port map( A => A_ns(20), ZN => n1016);
   U197 : OAI221_X1 port map( B1 => n872, B2 => n1019, C1 => n871, C2 => n1020,
                           A => n1021, ZN => O_21_port);
   U198 : AOI22_X1 port map( A1 => A_ns(20), A2 => n876, B1 => A_s(20), B2 => 
                           n877, ZN => n1021);
   U199 : INV_X1 port map( A => A_s(19), ZN => n1020);
   U200 : INV_X1 port map( A => A_ns(19), ZN => n1019);
   U201 : OAI221_X1 port map( B1 => n872, B2 => n1022, C1 => n871, C2 => n1023,
                           A => n1024, ZN => O_20_port);
   U202 : AOI22_X1 port map( A1 => A_ns(19), A2 => n876, B1 => A_s(19), B2 => 
                           n877, ZN => n1024);
   U203 : INV_X1 port map( A => A_s(18), ZN => n1023);
   U204 : INV_X1 port map( A => A_ns(18), ZN => n1022);
   U205 : OAI22_X1 port map( A1 => n1025, A2 => n993, B1 => n1026, B2 => n992, 
                           ZN => O_1_port);
   U206 : INV_X1 port map( A => A_ns(0), ZN => n992);
   U207 : INV_X1 port map( A => A_s(0), ZN => n993);
   U208 : OAI221_X1 port map( B1 => n872, B2 => n1027, C1 => n871, C2 => n1028,
                           A => n1029, ZN => O_19_port);
   U209 : AOI22_X1 port map( A1 => A_ns(18), A2 => n876, B1 => A_s(18), B2 => 
                           n877, ZN => n1029);
   U210 : INV_X1 port map( A => A_s(17), ZN => n1028);
   U211 : INV_X1 port map( A => A_ns(17), ZN => n1027);
   U212 : OAI221_X1 port map( B1 => n872, B2 => n1030, C1 => n871, C2 => n1031,
                           A => n1032, ZN => O_18_port);
   U213 : AOI22_X1 port map( A1 => A_ns(17), A2 => n876, B1 => A_s(17), B2 => 
                           n877, ZN => n1032);
   U214 : INV_X1 port map( A => A_s(16), ZN => n1031);
   U215 : INV_X1 port map( A => A_ns(16), ZN => n1030);
   U216 : OAI221_X1 port map( B1 => n872, B2 => n1033, C1 => n871, C2 => n1034,
                           A => n1035, ZN => O_17_port);
   U217 : AOI22_X1 port map( A1 => A_ns(16), A2 => n876, B1 => A_s(16), B2 => 
                           n877, ZN => n1035);
   U218 : INV_X1 port map( A => A_s(15), ZN => n1034);
   U219 : INV_X1 port map( A => A_ns(15), ZN => n1033);
   U220 : OAI221_X1 port map( B1 => n872, B2 => n1036, C1 => n871, C2 => n1037,
                           A => n1038, ZN => O_16_port);
   U221 : AOI22_X1 port map( A1 => A_ns(15), A2 => n876, B1 => A_s(15), B2 => 
                           n877, ZN => n1038);
   U222 : INV_X1 port map( A => A_s(14), ZN => n1037);
   U223 : INV_X1 port map( A => A_ns(14), ZN => n1036);
   U224 : OAI221_X1 port map( B1 => n872, B2 => n1039, C1 => n871, C2 => n1040,
                           A => n1041, ZN => O_15_port);
   U225 : AOI22_X1 port map( A1 => A_ns(14), A2 => n876, B1 => A_s(14), B2 => 
                           n877, ZN => n1041);
   U226 : INV_X1 port map( A => A_s(13), ZN => n1040);
   U227 : INV_X1 port map( A => A_ns(13), ZN => n1039);
   U228 : OAI221_X1 port map( B1 => n872, B2 => n1042, C1 => n871, C2 => n1043,
                           A => n1044, ZN => O_14_port);
   U229 : AOI22_X1 port map( A1 => A_ns(13), A2 => n876, B1 => A_s(13), B2 => 
                           n877, ZN => n1044);
   U230 : INV_X1 port map( A => A_s(12), ZN => n1043);
   U231 : INV_X1 port map( A => A_ns(12), ZN => n1042);
   U232 : OAI221_X1 port map( B1 => n872, B2 => n1045, C1 => n871, C2 => n1046,
                           A => n1047, ZN => O_13_port);
   U233 : AOI22_X1 port map( A1 => A_ns(12), A2 => n876, B1 => A_s(12), B2 => 
                           n877, ZN => n1047);
   U234 : INV_X1 port map( A => A_s(11), ZN => n1046);
   U235 : INV_X1 port map( A => A_ns(11), ZN => n1045);
   U236 : OAI221_X1 port map( B1 => n872, B2 => n1048, C1 => n871, C2 => n1049,
                           A => n1050, ZN => O_12_port);
   U237 : AOI22_X1 port map( A1 => A_ns(11), A2 => n876, B1 => A_s(11), B2 => 
                           n877, ZN => n1050);
   U238 : INV_X1 port map( A => A_s(10), ZN => n1049);
   U239 : INV_X1 port map( A => A_ns(10), ZN => n1048);
   U240 : OAI221_X1 port map( B1 => n872, B2 => n1051, C1 => n871, C2 => n1052,
                           A => n1053, ZN => O_11_port);
   U241 : AOI22_X1 port map( A1 => A_ns(10), A2 => n876, B1 => A_s(10), B2 => 
                           n877, ZN => n1053);
   U242 : INV_X1 port map( A => A_s(9), ZN => n1052);
   U243 : INV_X1 port map( A => A_ns(9), ZN => n1051);
   U244 : OAI221_X1 port map( B1 => n1054, B2 => n872, C1 => n1055, C2 => n871,
                           A => n1056, ZN => O_10_port);
   U245 : AOI22_X1 port map( A1 => A_ns(9), A2 => n876, B1 => A_s(9), B2 => 
                           n877, ZN => n1056);
   U246 : NAND2_X1 port map( A1 => n1057, A2 => n1025, ZN => n1026);
   U247 : NAND2_X1 port map( A1 => n1057, A2 => n1058, ZN => n1025);
   U248 : XOR2_X1 port map( A => B(27), B => B(28), Z => n1057);
   U249 : INV_X1 port map( A => A_s(8), ZN => n1055);
   U250 : INV_X1 port map( A => B(29), ZN => n1058);
   U251 : INV_X1 port map( A => A_ns(8), ZN => n1054);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT60_i26 is

   port( A_s, A_ns, B : in std_logic_vector (59 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (59 downto 0));

end BOOTHENC_NBIT60_i26;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT60_i26 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, O_59_port, O_58_port, O_57_port, O_56_port, O_55_port,
      O_54_port, O_53_port, O_52_port, O_51_port, O_50_port, O_49_port, 
      O_48_port, O_47_port, O_46_port, O_45_port, O_44_port, O_43_port, 
      O_42_port, O_41_port, O_40_port, O_39_port, O_38_port, O_37_port, 
      O_36_port, O_35_port, O_34_port, O_33_port, O_32_port, O_31_port, 
      O_30_port, O_29_port, O_28_port, O_27_port, O_26_port, O_25_port, 
      O_24_port, O_23_port, O_22_port, O_21_port, O_20_port, O_19_port, 
      O_18_port, O_17_port, O_16_port, O_15_port, O_14_port, O_13_port, 
      O_12_port, O_11_port, O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, 
      O_5_port, O_4_port, O_3_port, O_2_port, O_1_port, n844, n845, n846, n847,
      n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, 
      n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, 
      n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, 
      n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, 
      n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, 
      n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, 
      n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, 
      n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, 
      n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, 
      n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, 
      n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, 
      n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, 
      n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, 
      n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, 
      n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, 
      n1023, n1024, n1025, n1026 : std_logic;

begin
   O <= ( O_59_port, O_58_port, O_57_port, O_56_port, O_55_port, O_54_port, 
      O_53_port, O_52_port, O_51_port, O_50_port, O_49_port, O_48_port, 
      O_47_port, O_46_port, O_45_port, O_44_port, O_43_port, O_42_port, 
      O_41_port, O_40_port, O_39_port, O_38_port, O_37_port, O_36_port, 
      O_35_port, O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, 
      O_29_port, O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, 
      O_23_port, O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, 
      O_17_port, O_16_port, O_15_port, O_14_port, O_13_port, O_12_port, 
      O_11_port, O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, 
      O_4_port, O_3_port, O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(57), A_s(56), A_s(55), A_s(54), A_s(53), A_s(52), A_s(51), 
      A_s(50), A_s(49), A_s(48), A_s(47), A_s(46), A_s(45), A_s(44), A_s(43), 
      A_s(42), A_s(41), A_s(40), A_s(39), A_s(38), A_s(37), A_s(36), A_s(35), 
      A_s(34), A_s(33), A_s(32), A_s(31), A_s(30), A_s(29), A_s(28), A_s(27), 
      A_s(26), A_s(25), A_s(24), A_s(23), A_s(22), A_s(21), A_s(20), A_s(19), 
      A_s(18), A_s(17), A_s(16), A_s(15), A_s(14), A_s(13), A_s(12), A_s(11), 
      A_s(10), A_s(9), A_s(8), A_s(7), A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), 
      A_s(1), A_s(0), X_Logic0_port, X_Logic0_port );
   A_nso <= ( A_ns(57), A_ns(56), A_ns(55), A_ns(54), A_ns(53), A_ns(52), 
      A_ns(51), A_ns(50), A_ns(49), A_ns(48), A_ns(47), A_ns(46), A_ns(45), 
      A_ns(44), A_ns(43), A_ns(42), A_ns(41), A_ns(40), A_ns(39), A_ns(38), 
      A_ns(37), A_ns(36), A_ns(35), A_ns(34), A_ns(33), A_ns(32), A_ns(31), 
      A_ns(30), A_ns(29), A_ns(28), A_ns(27), A_ns(26), A_ns(25), A_ns(24), 
      A_ns(23), A_ns(22), A_ns(21), A_ns(20), A_ns(19), A_ns(18), A_ns(17), 
      A_ns(16), A_ns(15), A_ns(14), A_ns(13), A_ns(12), A_ns(11), A_ns(10), 
      A_ns(9), A_ns(8), A_ns(7), A_ns(6), A_ns(5), A_ns(4), A_ns(3), A_ns(2), 
      A_ns(1), A_ns(0), X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : AND3_X1 port map( A1 => B(26), A2 => n1026, A3 => B(25), ZN => n844);
   U3 : INV_X4 port map( A => n844, ZN => n845);
   U4 : INV_X4 port map( A => n993, ZN => n851);
   U5 : INV_X4 port map( A => n994, ZN => n850);
   U6 : OR3_X4 port map( A1 => B(25), A2 => B(26), A3 => n1026, ZN => n846);
   U7 : OAI221_X1 port map( B1 => n846, B2 => n847, C1 => n845, C2 => n848, A 
                           => n849, ZN => O_9_port);
   U8 : AOI22_X1 port map( A1 => A_ns(8), A2 => n850, B1 => A_s(8), B2 => n851,
                           ZN => n849);
   U9 : INV_X1 port map( A => A_s(7), ZN => n848);
   U10 : INV_X1 port map( A => A_ns(7), ZN => n847);
   U11 : OAI221_X1 port map( B1 => n846, B2 => n852, C1 => n845, C2 => n853, A 
                           => n854, ZN => O_8_port);
   U12 : AOI22_X1 port map( A1 => A_ns(7), A2 => n850, B1 => A_s(7), B2 => n851
                           , ZN => n854);
   U13 : INV_X1 port map( A => A_s(6), ZN => n853);
   U14 : INV_X1 port map( A => A_ns(6), ZN => n852);
   U15 : OAI221_X1 port map( B1 => n846, B2 => n855, C1 => n845, C2 => n856, A 
                           => n857, ZN => O_7_port);
   U16 : AOI22_X1 port map( A1 => A_ns(6), A2 => n850, B1 => A_s(6), B2 => n851
                           , ZN => n857);
   U17 : INV_X1 port map( A => A_s(5), ZN => n856);
   U18 : INV_X1 port map( A => A_ns(5), ZN => n855);
   U19 : OAI221_X1 port map( B1 => n846, B2 => n858, C1 => n845, C2 => n859, A 
                           => n860, ZN => O_6_port);
   U20 : AOI22_X1 port map( A1 => A_ns(5), A2 => n850, B1 => A_s(5), B2 => n851
                           , ZN => n860);
   U21 : INV_X1 port map( A => A_s(4), ZN => n859);
   U22 : INV_X1 port map( A => A_ns(4), ZN => n858);
   U23 : OAI221_X1 port map( B1 => n846, B2 => n861, C1 => n845, C2 => n862, A 
                           => n863, ZN => O_5_port);
   U24 : AOI22_X1 port map( A1 => A_ns(4), A2 => n850, B1 => A_s(4), B2 => n851
                           , ZN => n863);
   U25 : INV_X1 port map( A => A_s(3), ZN => n862);
   U26 : INV_X1 port map( A => A_ns(3), ZN => n861);
   U27 : OAI221_X1 port map( B1 => n846, B2 => n864, C1 => n845, C2 => n865, A 
                           => n866, ZN => O_59_port);
   U28 : AOI22_X1 port map( A1 => A_ns(58), A2 => n850, B1 => A_s(58), B2 => 
                           n851, ZN => n866);
   U29 : INV_X1 port map( A => A_s(57), ZN => n865);
   U30 : INV_X1 port map( A => A_ns(57), ZN => n864);
   U31 : OAI221_X1 port map( B1 => n846, B2 => n867, C1 => n845, C2 => n868, A 
                           => n869, ZN => O_58_port);
   U32 : AOI22_X1 port map( A1 => A_ns(57), A2 => n850, B1 => A_s(57), B2 => 
                           n851, ZN => n869);
   U33 : INV_X1 port map( A => A_s(56), ZN => n868);
   U34 : INV_X1 port map( A => A_ns(56), ZN => n867);
   U35 : OAI221_X1 port map( B1 => n846, B2 => n870, C1 => n845, C2 => n871, A 
                           => n872, ZN => O_57_port);
   U36 : AOI22_X1 port map( A1 => A_ns(56), A2 => n850, B1 => A_s(56), B2 => 
                           n851, ZN => n872);
   U37 : INV_X1 port map( A => A_s(55), ZN => n871);
   U38 : INV_X1 port map( A => A_ns(55), ZN => n870);
   U39 : OAI221_X1 port map( B1 => n846, B2 => n873, C1 => n845, C2 => n874, A 
                           => n875, ZN => O_56_port);
   U40 : AOI22_X1 port map( A1 => A_ns(55), A2 => n850, B1 => A_s(55), B2 => 
                           n851, ZN => n875);
   U41 : INV_X1 port map( A => A_s(54), ZN => n874);
   U42 : INV_X1 port map( A => A_ns(54), ZN => n873);
   U43 : OAI221_X1 port map( B1 => n846, B2 => n876, C1 => n845, C2 => n877, A 
                           => n878, ZN => O_55_port);
   U44 : AOI22_X1 port map( A1 => A_ns(54), A2 => n850, B1 => A_s(54), B2 => 
                           n851, ZN => n878);
   U45 : INV_X1 port map( A => A_s(53), ZN => n877);
   U46 : INV_X1 port map( A => A_ns(53), ZN => n876);
   U47 : OAI221_X1 port map( B1 => n846, B2 => n879, C1 => n845, C2 => n880, A 
                           => n881, ZN => O_54_port);
   U48 : AOI22_X1 port map( A1 => A_ns(53), A2 => n850, B1 => A_s(53), B2 => 
                           n851, ZN => n881);
   U49 : INV_X1 port map( A => A_s(52), ZN => n880);
   U50 : INV_X1 port map( A => A_ns(52), ZN => n879);
   U51 : OAI221_X1 port map( B1 => n846, B2 => n882, C1 => n845, C2 => n883, A 
                           => n884, ZN => O_53_port);
   U52 : AOI22_X1 port map( A1 => A_ns(52), A2 => n850, B1 => A_s(52), B2 => 
                           n851, ZN => n884);
   U53 : INV_X1 port map( A => A_s(51), ZN => n883);
   U54 : INV_X1 port map( A => A_ns(51), ZN => n882);
   U55 : OAI221_X1 port map( B1 => n846, B2 => n885, C1 => n845, C2 => n886, A 
                           => n887, ZN => O_52_port);
   U56 : AOI22_X1 port map( A1 => A_ns(51), A2 => n850, B1 => A_s(51), B2 => 
                           n851, ZN => n887);
   U57 : INV_X1 port map( A => A_s(50), ZN => n886);
   U58 : INV_X1 port map( A => A_ns(50), ZN => n885);
   U59 : OAI221_X1 port map( B1 => n846, B2 => n888, C1 => n845, C2 => n889, A 
                           => n890, ZN => O_51_port);
   U60 : AOI22_X1 port map( A1 => A_ns(50), A2 => n850, B1 => A_s(50), B2 => 
                           n851, ZN => n890);
   U61 : INV_X1 port map( A => A_s(49), ZN => n889);
   U62 : INV_X1 port map( A => A_ns(49), ZN => n888);
   U63 : OAI221_X1 port map( B1 => n846, B2 => n891, C1 => n845, C2 => n892, A 
                           => n893, ZN => O_50_port);
   U64 : AOI22_X1 port map( A1 => A_ns(49), A2 => n850, B1 => A_s(49), B2 => 
                           n851, ZN => n893);
   U65 : INV_X1 port map( A => A_s(48), ZN => n892);
   U66 : INV_X1 port map( A => A_ns(48), ZN => n891);
   U67 : OAI221_X1 port map( B1 => n846, B2 => n894, C1 => n845, C2 => n895, A 
                           => n896, ZN => O_4_port);
   U68 : AOI22_X1 port map( A1 => A_ns(3), A2 => n850, B1 => A_s(3), B2 => n851
                           , ZN => n896);
   U69 : INV_X1 port map( A => A_s(2), ZN => n895);
   U70 : INV_X1 port map( A => A_ns(2), ZN => n894);
   U71 : OAI221_X1 port map( B1 => n846, B2 => n897, C1 => n845, C2 => n898, A 
                           => n899, ZN => O_49_port);
   U72 : AOI22_X1 port map( A1 => A_ns(48), A2 => n850, B1 => A_s(48), B2 => 
                           n851, ZN => n899);
   U73 : INV_X1 port map( A => A_s(47), ZN => n898);
   U74 : INV_X1 port map( A => A_ns(47), ZN => n897);
   U75 : OAI221_X1 port map( B1 => n846, B2 => n900, C1 => n845, C2 => n901, A 
                           => n902, ZN => O_48_port);
   U76 : AOI22_X1 port map( A1 => A_ns(47), A2 => n850, B1 => A_s(47), B2 => 
                           n851, ZN => n902);
   U77 : INV_X1 port map( A => A_s(46), ZN => n901);
   U78 : INV_X1 port map( A => A_ns(46), ZN => n900);
   U79 : OAI221_X1 port map( B1 => n846, B2 => n903, C1 => n845, C2 => n904, A 
                           => n905, ZN => O_47_port);
   U80 : AOI22_X1 port map( A1 => A_ns(46), A2 => n850, B1 => A_s(46), B2 => 
                           n851, ZN => n905);
   U81 : INV_X1 port map( A => A_s(45), ZN => n904);
   U82 : INV_X1 port map( A => A_ns(45), ZN => n903);
   U83 : OAI221_X1 port map( B1 => n846, B2 => n906, C1 => n845, C2 => n907, A 
                           => n908, ZN => O_46_port);
   U84 : AOI22_X1 port map( A1 => A_ns(45), A2 => n850, B1 => A_s(45), B2 => 
                           n851, ZN => n908);
   U85 : INV_X1 port map( A => A_s(44), ZN => n907);
   U86 : INV_X1 port map( A => A_ns(44), ZN => n906);
   U87 : OAI221_X1 port map( B1 => n846, B2 => n909, C1 => n845, C2 => n910, A 
                           => n911, ZN => O_45_port);
   U88 : AOI22_X1 port map( A1 => A_ns(44), A2 => n850, B1 => A_s(44), B2 => 
                           n851, ZN => n911);
   U89 : INV_X1 port map( A => A_s(43), ZN => n910);
   U90 : INV_X1 port map( A => A_ns(43), ZN => n909);
   U91 : OAI221_X1 port map( B1 => n846, B2 => n912, C1 => n845, C2 => n913, A 
                           => n914, ZN => O_44_port);
   U92 : AOI22_X1 port map( A1 => A_ns(43), A2 => n850, B1 => A_s(43), B2 => 
                           n851, ZN => n914);
   U93 : INV_X1 port map( A => A_s(42), ZN => n913);
   U94 : INV_X1 port map( A => A_ns(42), ZN => n912);
   U95 : OAI221_X1 port map( B1 => n846, B2 => n915, C1 => n845, C2 => n916, A 
                           => n917, ZN => O_43_port);
   U96 : AOI22_X1 port map( A1 => A_ns(42), A2 => n850, B1 => A_s(42), B2 => 
                           n851, ZN => n917);
   U97 : INV_X1 port map( A => A_s(41), ZN => n916);
   U98 : INV_X1 port map( A => A_ns(41), ZN => n915);
   U99 : OAI221_X1 port map( B1 => n846, B2 => n918, C1 => n845, C2 => n919, A 
                           => n920, ZN => O_42_port);
   U100 : AOI22_X1 port map( A1 => A_ns(41), A2 => n850, B1 => A_s(41), B2 => 
                           n851, ZN => n920);
   U101 : INV_X1 port map( A => A_s(40), ZN => n919);
   U102 : INV_X1 port map( A => A_ns(40), ZN => n918);
   U103 : OAI221_X1 port map( B1 => n846, B2 => n921, C1 => n845, C2 => n922, A
                           => n923, ZN => O_41_port);
   U104 : AOI22_X1 port map( A1 => A_ns(40), A2 => n850, B1 => A_s(40), B2 => 
                           n851, ZN => n923);
   U105 : INV_X1 port map( A => A_s(39), ZN => n922);
   U106 : INV_X1 port map( A => A_ns(39), ZN => n921);
   U107 : OAI221_X1 port map( B1 => n846, B2 => n924, C1 => n845, C2 => n925, A
                           => n926, ZN => O_40_port);
   U108 : AOI22_X1 port map( A1 => A_ns(39), A2 => n850, B1 => A_s(39), B2 => 
                           n851, ZN => n926);
   U109 : INV_X1 port map( A => A_s(38), ZN => n925);
   U110 : INV_X1 port map( A => A_ns(38), ZN => n924);
   U111 : OAI221_X1 port map( B1 => n846, B2 => n927, C1 => n845, C2 => n928, A
                           => n929, ZN => O_3_port);
   U112 : AOI22_X1 port map( A1 => A_ns(2), A2 => n850, B1 => A_s(2), B2 => 
                           n851, ZN => n929);
   U113 : INV_X1 port map( A => A_s(1), ZN => n928);
   U114 : INV_X1 port map( A => A_ns(1), ZN => n927);
   U115 : OAI221_X1 port map( B1 => n846, B2 => n930, C1 => n845, C2 => n931, A
                           => n932, ZN => O_39_port);
   U116 : AOI22_X1 port map( A1 => A_ns(38), A2 => n850, B1 => A_s(38), B2 => 
                           n851, ZN => n932);
   U117 : INV_X1 port map( A => A_s(37), ZN => n931);
   U118 : INV_X1 port map( A => A_ns(37), ZN => n930);
   U119 : OAI221_X1 port map( B1 => n846, B2 => n933, C1 => n845, C2 => n934, A
                           => n935, ZN => O_38_port);
   U120 : AOI22_X1 port map( A1 => A_ns(37), A2 => n850, B1 => A_s(37), B2 => 
                           n851, ZN => n935);
   U121 : INV_X1 port map( A => A_s(36), ZN => n934);
   U122 : INV_X1 port map( A => A_ns(36), ZN => n933);
   U123 : OAI221_X1 port map( B1 => n846, B2 => n936, C1 => n845, C2 => n937, A
                           => n938, ZN => O_37_port);
   U124 : AOI22_X1 port map( A1 => A_ns(36), A2 => n850, B1 => A_s(36), B2 => 
                           n851, ZN => n938);
   U125 : INV_X1 port map( A => A_s(35), ZN => n937);
   U126 : INV_X1 port map( A => A_ns(35), ZN => n936);
   U127 : OAI221_X1 port map( B1 => n846, B2 => n939, C1 => n845, C2 => n940, A
                           => n941, ZN => O_36_port);
   U128 : AOI22_X1 port map( A1 => A_ns(35), A2 => n850, B1 => A_s(35), B2 => 
                           n851, ZN => n941);
   U129 : INV_X1 port map( A => A_s(34), ZN => n940);
   U130 : INV_X1 port map( A => A_ns(34), ZN => n939);
   U131 : OAI221_X1 port map( B1 => n846, B2 => n942, C1 => n845, C2 => n943, A
                           => n944, ZN => O_35_port);
   U132 : AOI22_X1 port map( A1 => A_ns(34), A2 => n850, B1 => A_s(34), B2 => 
                           n851, ZN => n944);
   U133 : INV_X1 port map( A => A_s(33), ZN => n943);
   U134 : INV_X1 port map( A => A_ns(33), ZN => n942);
   U135 : OAI221_X1 port map( B1 => n846, B2 => n945, C1 => n845, C2 => n946, A
                           => n947, ZN => O_34_port);
   U136 : AOI22_X1 port map( A1 => A_ns(33), A2 => n850, B1 => A_s(33), B2 => 
                           n851, ZN => n947);
   U137 : INV_X1 port map( A => A_s(32), ZN => n946);
   U138 : INV_X1 port map( A => A_ns(32), ZN => n945);
   U139 : OAI221_X1 port map( B1 => n846, B2 => n948, C1 => n845, C2 => n949, A
                           => n950, ZN => O_33_port);
   U140 : AOI22_X1 port map( A1 => A_ns(32), A2 => n850, B1 => A_s(32), B2 => 
                           n851, ZN => n950);
   U141 : INV_X1 port map( A => A_s(31), ZN => n949);
   U142 : INV_X1 port map( A => A_ns(31), ZN => n948);
   U143 : OAI221_X1 port map( B1 => n846, B2 => n951, C1 => n845, C2 => n952, A
                           => n953, ZN => O_32_port);
   U144 : AOI22_X1 port map( A1 => A_ns(31), A2 => n850, B1 => A_s(31), B2 => 
                           n851, ZN => n953);
   U145 : INV_X1 port map( A => A_s(30), ZN => n952);
   U146 : INV_X1 port map( A => A_ns(30), ZN => n951);
   U147 : OAI221_X1 port map( B1 => n846, B2 => n954, C1 => n845, C2 => n955, A
                           => n956, ZN => O_31_port);
   U148 : AOI22_X1 port map( A1 => A_ns(30), A2 => n850, B1 => A_s(30), B2 => 
                           n851, ZN => n956);
   U149 : INV_X1 port map( A => A_s(29), ZN => n955);
   U150 : INV_X1 port map( A => A_ns(29), ZN => n954);
   U151 : OAI221_X1 port map( B1 => n846, B2 => n957, C1 => n845, C2 => n958, A
                           => n959, ZN => O_30_port);
   U152 : AOI22_X1 port map( A1 => A_ns(29), A2 => n850, B1 => A_s(29), B2 => 
                           n851, ZN => n959);
   U153 : INV_X1 port map( A => A_s(28), ZN => n958);
   U154 : INV_X1 port map( A => A_ns(28), ZN => n957);
   U155 : OAI221_X1 port map( B1 => n846, B2 => n960, C1 => n845, C2 => n961, A
                           => n962, ZN => O_2_port);
   U156 : AOI22_X1 port map( A1 => A_ns(1), A2 => n850, B1 => A_s(1), B2 => 
                           n851, ZN => n962);
   U157 : OAI221_X1 port map( B1 => n846, B2 => n963, C1 => n845, C2 => n964, A
                           => n965, ZN => O_29_port);
   U158 : AOI22_X1 port map( A1 => A_ns(28), A2 => n850, B1 => A_s(28), B2 => 
                           n851, ZN => n965);
   U159 : INV_X1 port map( A => A_s(27), ZN => n964);
   U160 : INV_X1 port map( A => A_ns(27), ZN => n963);
   U161 : OAI221_X1 port map( B1 => n846, B2 => n966, C1 => n845, C2 => n967, A
                           => n968, ZN => O_28_port);
   U162 : AOI22_X1 port map( A1 => A_ns(27), A2 => n850, B1 => A_s(27), B2 => 
                           n851, ZN => n968);
   U163 : INV_X1 port map( A => A_s(26), ZN => n967);
   U164 : INV_X1 port map( A => A_ns(26), ZN => n966);
   U165 : OAI221_X1 port map( B1 => n846, B2 => n969, C1 => n845, C2 => n970, A
                           => n971, ZN => O_27_port);
   U166 : AOI22_X1 port map( A1 => A_ns(26), A2 => n850, B1 => A_s(26), B2 => 
                           n851, ZN => n971);
   U167 : INV_X1 port map( A => A_s(25), ZN => n970);
   U168 : INV_X1 port map( A => A_ns(25), ZN => n969);
   U169 : OAI221_X1 port map( B1 => n846, B2 => n972, C1 => n845, C2 => n973, A
                           => n974, ZN => O_26_port);
   U170 : AOI22_X1 port map( A1 => A_ns(25), A2 => n850, B1 => A_s(25), B2 => 
                           n851, ZN => n974);
   U171 : INV_X1 port map( A => A_s(24), ZN => n973);
   U172 : INV_X1 port map( A => A_ns(24), ZN => n972);
   U173 : OAI221_X1 port map( B1 => n846, B2 => n975, C1 => n845, C2 => n976, A
                           => n977, ZN => O_25_port);
   U174 : AOI22_X1 port map( A1 => A_ns(24), A2 => n850, B1 => A_s(24), B2 => 
                           n851, ZN => n977);
   U175 : INV_X1 port map( A => A_s(23), ZN => n976);
   U176 : INV_X1 port map( A => A_ns(23), ZN => n975);
   U177 : OAI221_X1 port map( B1 => n846, B2 => n978, C1 => n845, C2 => n979, A
                           => n980, ZN => O_24_port);
   U178 : AOI22_X1 port map( A1 => A_ns(23), A2 => n850, B1 => A_s(23), B2 => 
                           n851, ZN => n980);
   U179 : INV_X1 port map( A => A_s(22), ZN => n979);
   U180 : INV_X1 port map( A => A_ns(22), ZN => n978);
   U181 : OAI221_X1 port map( B1 => n846, B2 => n981, C1 => n845, C2 => n982, A
                           => n983, ZN => O_23_port);
   U182 : AOI22_X1 port map( A1 => A_ns(22), A2 => n850, B1 => A_s(22), B2 => 
                           n851, ZN => n983);
   U183 : INV_X1 port map( A => A_s(21), ZN => n982);
   U184 : INV_X1 port map( A => A_ns(21), ZN => n981);
   U185 : OAI221_X1 port map( B1 => n846, B2 => n984, C1 => n845, C2 => n985, A
                           => n986, ZN => O_22_port);
   U186 : AOI22_X1 port map( A1 => A_ns(21), A2 => n850, B1 => A_s(21), B2 => 
                           n851, ZN => n986);
   U187 : INV_X1 port map( A => A_s(20), ZN => n985);
   U188 : INV_X1 port map( A => A_ns(20), ZN => n984);
   U189 : OAI221_X1 port map( B1 => n846, B2 => n987, C1 => n845, C2 => n988, A
                           => n989, ZN => O_21_port);
   U190 : AOI22_X1 port map( A1 => A_ns(20), A2 => n850, B1 => A_s(20), B2 => 
                           n851, ZN => n989);
   U191 : INV_X1 port map( A => A_s(19), ZN => n988);
   U192 : INV_X1 port map( A => A_ns(19), ZN => n987);
   U193 : OAI221_X1 port map( B1 => n846, B2 => n990, C1 => n845, C2 => n991, A
                           => n992, ZN => O_20_port);
   U194 : AOI22_X1 port map( A1 => A_ns(19), A2 => n850, B1 => A_s(19), B2 => 
                           n851, ZN => n992);
   U195 : INV_X1 port map( A => A_s(18), ZN => n991);
   U196 : INV_X1 port map( A => A_ns(18), ZN => n990);
   U197 : OAI22_X1 port map( A1 => n993, A2 => n961, B1 => n994, B2 => n960, ZN
                           => O_1_port);
   U198 : INV_X1 port map( A => A_ns(0), ZN => n960);
   U199 : INV_X1 port map( A => A_s(0), ZN => n961);
   U200 : OAI221_X1 port map( B1 => n846, B2 => n995, C1 => n845, C2 => n996, A
                           => n997, ZN => O_19_port);
   U201 : AOI22_X1 port map( A1 => A_ns(18), A2 => n850, B1 => A_s(18), B2 => 
                           n851, ZN => n997);
   U202 : INV_X1 port map( A => A_s(17), ZN => n996);
   U203 : INV_X1 port map( A => A_ns(17), ZN => n995);
   U204 : OAI221_X1 port map( B1 => n846, B2 => n998, C1 => n845, C2 => n999, A
                           => n1000, ZN => O_18_port);
   U205 : AOI22_X1 port map( A1 => A_ns(17), A2 => n850, B1 => A_s(17), B2 => 
                           n851, ZN => n1000);
   U206 : INV_X1 port map( A => A_s(16), ZN => n999);
   U207 : INV_X1 port map( A => A_ns(16), ZN => n998);
   U208 : OAI221_X1 port map( B1 => n846, B2 => n1001, C1 => n845, C2 => n1002,
                           A => n1003, ZN => O_17_port);
   U209 : AOI22_X1 port map( A1 => A_ns(16), A2 => n850, B1 => A_s(16), B2 => 
                           n851, ZN => n1003);
   U210 : INV_X1 port map( A => A_s(15), ZN => n1002);
   U211 : INV_X1 port map( A => A_ns(15), ZN => n1001);
   U212 : OAI221_X1 port map( B1 => n846, B2 => n1004, C1 => n845, C2 => n1005,
                           A => n1006, ZN => O_16_port);
   U213 : AOI22_X1 port map( A1 => A_ns(15), A2 => n850, B1 => A_s(15), B2 => 
                           n851, ZN => n1006);
   U214 : INV_X1 port map( A => A_s(14), ZN => n1005);
   U215 : INV_X1 port map( A => A_ns(14), ZN => n1004);
   U216 : OAI221_X1 port map( B1 => n846, B2 => n1007, C1 => n845, C2 => n1008,
                           A => n1009, ZN => O_15_port);
   U217 : AOI22_X1 port map( A1 => A_ns(14), A2 => n850, B1 => A_s(14), B2 => 
                           n851, ZN => n1009);
   U218 : INV_X1 port map( A => A_s(13), ZN => n1008);
   U219 : INV_X1 port map( A => A_ns(13), ZN => n1007);
   U220 : OAI221_X1 port map( B1 => n846, B2 => n1010, C1 => n845, C2 => n1011,
                           A => n1012, ZN => O_14_port);
   U221 : AOI22_X1 port map( A1 => A_ns(13), A2 => n850, B1 => A_s(13), B2 => 
                           n851, ZN => n1012);
   U222 : INV_X1 port map( A => A_s(12), ZN => n1011);
   U223 : INV_X1 port map( A => A_ns(12), ZN => n1010);
   U224 : OAI221_X1 port map( B1 => n846, B2 => n1013, C1 => n845, C2 => n1014,
                           A => n1015, ZN => O_13_port);
   U225 : AOI22_X1 port map( A1 => A_ns(12), A2 => n850, B1 => A_s(12), B2 => 
                           n851, ZN => n1015);
   U226 : INV_X1 port map( A => A_s(11), ZN => n1014);
   U227 : INV_X1 port map( A => A_ns(11), ZN => n1013);
   U228 : OAI221_X1 port map( B1 => n846, B2 => n1016, C1 => n845, C2 => n1017,
                           A => n1018, ZN => O_12_port);
   U229 : AOI22_X1 port map( A1 => A_ns(11), A2 => n850, B1 => A_s(11), B2 => 
                           n851, ZN => n1018);
   U230 : INV_X1 port map( A => A_s(10), ZN => n1017);
   U231 : INV_X1 port map( A => A_ns(10), ZN => n1016);
   U232 : OAI221_X1 port map( B1 => n846, B2 => n1019, C1 => n845, C2 => n1020,
                           A => n1021, ZN => O_11_port);
   U233 : AOI22_X1 port map( A1 => A_ns(10), A2 => n850, B1 => A_s(10), B2 => 
                           n851, ZN => n1021);
   U234 : INV_X1 port map( A => A_s(9), ZN => n1020);
   U235 : INV_X1 port map( A => A_ns(9), ZN => n1019);
   U236 : OAI221_X1 port map( B1 => n1022, B2 => n846, C1 => n1023, C2 => n845,
                           A => n1024, ZN => O_10_port);
   U237 : AOI22_X1 port map( A1 => A_ns(9), A2 => n850, B1 => A_s(9), B2 => 
                           n851, ZN => n1024);
   U238 : NAND2_X1 port map( A1 => n1025, A2 => n993, ZN => n994);
   U239 : NAND2_X1 port map( A1 => n1025, A2 => n1026, ZN => n993);
   U240 : XOR2_X1 port map( A => B(25), B => B(26), Z => n1025);
   U241 : INV_X1 port map( A => A_s(8), ZN => n1023);
   U242 : INV_X1 port map( A => B(27), ZN => n1026);
   U243 : INV_X1 port map( A => A_ns(8), ZN => n1022);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT58_i24 is

   port( A_s, A_ns, B : in std_logic_vector (57 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (57 downto 0));

end BOOTHENC_NBIT58_i24;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT58_i24 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, O_57_port, O_56_port, O_55_port, O_54_port, O_53_port,
      O_52_port, O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, 
      O_46_port, O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, 
      O_40_port, O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, 
      O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, 
      O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, 
      O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, 
      O_16_port, O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, 
      O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, 
      O_3_port, O_2_port, O_1_port, n827, n828, n829, n830, n831, n832, n833, 
      n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, 
      n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, 
      n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, 
      n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, 
      n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, 
      n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, 
      n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, 
      n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, 
      n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, 
      n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, 
      n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, 
      n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, 
      n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, 
      n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
      n1002, n1003 : std_logic;

begin
   O <= ( O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, O_52_port, 
      O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, O_46_port, 
      O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, O_40_port, 
      O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, 
      O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, 
      O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, 
      O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, O_16_port, 
      O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, O_10_port, 
      O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, O_3_port, 
      O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(55), A_s(54), A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), 
      A_s(48), A_s(47), A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), 
      A_s(40), A_s(39), A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), 
      A_s(32), A_s(31), A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), 
      A_s(24), A_s(23), A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), 
      A_s(16), A_s(15), A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), 
      A_s(8), A_s(7), A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), 
      X_Logic0_port, X_Logic0_port );
   A_nso <= ( A_ns(55), A_ns(54), A_ns(53), A_ns(52), A_ns(51), A_ns(50), 
      A_ns(49), A_ns(48), A_ns(47), A_ns(46), A_ns(45), A_ns(44), A_ns(43), 
      A_ns(42), A_ns(41), A_ns(40), A_ns(39), A_ns(38), A_ns(37), A_ns(36), 
      A_ns(35), A_ns(34), A_ns(33), A_ns(32), A_ns(31), A_ns(30), A_ns(29), 
      A_ns(28), A_ns(27), A_ns(26), A_ns(25), A_ns(24), A_ns(23), A_ns(22), 
      A_ns(21), A_ns(20), A_ns(19), A_ns(18), A_ns(17), A_ns(16), A_ns(15), 
      A_ns(14), A_ns(13), A_ns(12), A_ns(11), A_ns(10), A_ns(9), A_ns(8), 
      A_ns(7), A_ns(6), A_ns(5), A_ns(4), A_ns(3), A_ns(2), A_ns(1), A_ns(0), 
      X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : AND3_X1 port map( A1 => B(24), A2 => n1003, A3 => B(23), ZN => n827);
   U3 : INV_X4 port map( A => n827, ZN => n828);
   U4 : INV_X4 port map( A => n970, ZN => n834);
   U5 : INV_X4 port map( A => n971, ZN => n833);
   U6 : OR3_X4 port map( A1 => B(23), A2 => B(24), A3 => n1003, ZN => n829);
   U7 : OAI221_X1 port map( B1 => n829, B2 => n830, C1 => n828, C2 => n831, A 
                           => n832, ZN => O_9_port);
   U8 : AOI22_X1 port map( A1 => A_ns(8), A2 => n833, B1 => A_s(8), B2 => n834,
                           ZN => n832);
   U9 : INV_X1 port map( A => A_s(7), ZN => n831);
   U10 : INV_X1 port map( A => A_ns(7), ZN => n830);
   U11 : OAI221_X1 port map( B1 => n829, B2 => n835, C1 => n828, C2 => n836, A 
                           => n837, ZN => O_8_port);
   U12 : AOI22_X1 port map( A1 => A_ns(7), A2 => n833, B1 => A_s(7), B2 => n834
                           , ZN => n837);
   U13 : INV_X1 port map( A => A_s(6), ZN => n836);
   U14 : INV_X1 port map( A => A_ns(6), ZN => n835);
   U15 : OAI221_X1 port map( B1 => n829, B2 => n838, C1 => n828, C2 => n839, A 
                           => n840, ZN => O_7_port);
   U16 : AOI22_X1 port map( A1 => A_ns(6), A2 => n833, B1 => A_s(6), B2 => n834
                           , ZN => n840);
   U17 : INV_X1 port map( A => A_s(5), ZN => n839);
   U18 : INV_X1 port map( A => A_ns(5), ZN => n838);
   U19 : OAI221_X1 port map( B1 => n829, B2 => n841, C1 => n828, C2 => n842, A 
                           => n843, ZN => O_6_port);
   U20 : AOI22_X1 port map( A1 => A_ns(5), A2 => n833, B1 => A_s(5), B2 => n834
                           , ZN => n843);
   U21 : INV_X1 port map( A => A_s(4), ZN => n842);
   U22 : INV_X1 port map( A => A_ns(4), ZN => n841);
   U23 : OAI221_X1 port map( B1 => n829, B2 => n844, C1 => n828, C2 => n845, A 
                           => n846, ZN => O_5_port);
   U24 : AOI22_X1 port map( A1 => A_ns(4), A2 => n833, B1 => A_s(4), B2 => n834
                           , ZN => n846);
   U25 : INV_X1 port map( A => A_s(3), ZN => n845);
   U26 : INV_X1 port map( A => A_ns(3), ZN => n844);
   U27 : OAI221_X1 port map( B1 => n829, B2 => n847, C1 => n828, C2 => n848, A 
                           => n849, ZN => O_57_port);
   U28 : AOI22_X1 port map( A1 => A_ns(56), A2 => n833, B1 => A_s(56), B2 => 
                           n834, ZN => n849);
   U29 : INV_X1 port map( A => A_s(55), ZN => n848);
   U30 : INV_X1 port map( A => A_ns(55), ZN => n847);
   U31 : OAI221_X1 port map( B1 => n829, B2 => n850, C1 => n828, C2 => n851, A 
                           => n852, ZN => O_56_port);
   U32 : AOI22_X1 port map( A1 => A_ns(55), A2 => n833, B1 => A_s(55), B2 => 
                           n834, ZN => n852);
   U33 : INV_X1 port map( A => A_s(54), ZN => n851);
   U34 : INV_X1 port map( A => A_ns(54), ZN => n850);
   U35 : OAI221_X1 port map( B1 => n829, B2 => n853, C1 => n828, C2 => n854, A 
                           => n855, ZN => O_55_port);
   U36 : AOI22_X1 port map( A1 => A_ns(54), A2 => n833, B1 => A_s(54), B2 => 
                           n834, ZN => n855);
   U37 : INV_X1 port map( A => A_s(53), ZN => n854);
   U38 : INV_X1 port map( A => A_ns(53), ZN => n853);
   U39 : OAI221_X1 port map( B1 => n829, B2 => n856, C1 => n828, C2 => n857, A 
                           => n858, ZN => O_54_port);
   U40 : AOI22_X1 port map( A1 => A_ns(53), A2 => n833, B1 => A_s(53), B2 => 
                           n834, ZN => n858);
   U41 : INV_X1 port map( A => A_s(52), ZN => n857);
   U42 : INV_X1 port map( A => A_ns(52), ZN => n856);
   U43 : OAI221_X1 port map( B1 => n829, B2 => n859, C1 => n828, C2 => n860, A 
                           => n861, ZN => O_53_port);
   U44 : AOI22_X1 port map( A1 => A_ns(52), A2 => n833, B1 => A_s(52), B2 => 
                           n834, ZN => n861);
   U45 : INV_X1 port map( A => A_s(51), ZN => n860);
   U46 : INV_X1 port map( A => A_ns(51), ZN => n859);
   U47 : OAI221_X1 port map( B1 => n829, B2 => n862, C1 => n828, C2 => n863, A 
                           => n864, ZN => O_52_port);
   U48 : AOI22_X1 port map( A1 => A_ns(51), A2 => n833, B1 => A_s(51), B2 => 
                           n834, ZN => n864);
   U49 : INV_X1 port map( A => A_s(50), ZN => n863);
   U50 : INV_X1 port map( A => A_ns(50), ZN => n862);
   U51 : OAI221_X1 port map( B1 => n829, B2 => n865, C1 => n828, C2 => n866, A 
                           => n867, ZN => O_51_port);
   U52 : AOI22_X1 port map( A1 => A_ns(50), A2 => n833, B1 => A_s(50), B2 => 
                           n834, ZN => n867);
   U53 : INV_X1 port map( A => A_s(49), ZN => n866);
   U54 : INV_X1 port map( A => A_ns(49), ZN => n865);
   U55 : OAI221_X1 port map( B1 => n829, B2 => n868, C1 => n828, C2 => n869, A 
                           => n870, ZN => O_50_port);
   U56 : AOI22_X1 port map( A1 => A_ns(49), A2 => n833, B1 => A_s(49), B2 => 
                           n834, ZN => n870);
   U57 : INV_X1 port map( A => A_s(48), ZN => n869);
   U58 : INV_X1 port map( A => A_ns(48), ZN => n868);
   U59 : OAI221_X1 port map( B1 => n829, B2 => n871, C1 => n828, C2 => n872, A 
                           => n873, ZN => O_4_port);
   U60 : AOI22_X1 port map( A1 => A_ns(3), A2 => n833, B1 => A_s(3), B2 => n834
                           , ZN => n873);
   U61 : INV_X1 port map( A => A_s(2), ZN => n872);
   U62 : INV_X1 port map( A => A_ns(2), ZN => n871);
   U63 : OAI221_X1 port map( B1 => n829, B2 => n874, C1 => n828, C2 => n875, A 
                           => n876, ZN => O_49_port);
   U64 : AOI22_X1 port map( A1 => A_ns(48), A2 => n833, B1 => A_s(48), B2 => 
                           n834, ZN => n876);
   U65 : INV_X1 port map( A => A_s(47), ZN => n875);
   U66 : INV_X1 port map( A => A_ns(47), ZN => n874);
   U67 : OAI221_X1 port map( B1 => n829, B2 => n877, C1 => n828, C2 => n878, A 
                           => n879, ZN => O_48_port);
   U68 : AOI22_X1 port map( A1 => A_ns(47), A2 => n833, B1 => A_s(47), B2 => 
                           n834, ZN => n879);
   U69 : INV_X1 port map( A => A_s(46), ZN => n878);
   U70 : INV_X1 port map( A => A_ns(46), ZN => n877);
   U71 : OAI221_X1 port map( B1 => n829, B2 => n880, C1 => n828, C2 => n881, A 
                           => n882, ZN => O_47_port);
   U72 : AOI22_X1 port map( A1 => A_ns(46), A2 => n833, B1 => A_s(46), B2 => 
                           n834, ZN => n882);
   U73 : INV_X1 port map( A => A_s(45), ZN => n881);
   U74 : INV_X1 port map( A => A_ns(45), ZN => n880);
   U75 : OAI221_X1 port map( B1 => n829, B2 => n883, C1 => n828, C2 => n884, A 
                           => n885, ZN => O_46_port);
   U76 : AOI22_X1 port map( A1 => A_ns(45), A2 => n833, B1 => A_s(45), B2 => 
                           n834, ZN => n885);
   U77 : INV_X1 port map( A => A_s(44), ZN => n884);
   U78 : INV_X1 port map( A => A_ns(44), ZN => n883);
   U79 : OAI221_X1 port map( B1 => n829, B2 => n886, C1 => n828, C2 => n887, A 
                           => n888, ZN => O_45_port);
   U80 : AOI22_X1 port map( A1 => A_ns(44), A2 => n833, B1 => A_s(44), B2 => 
                           n834, ZN => n888);
   U81 : INV_X1 port map( A => A_s(43), ZN => n887);
   U82 : INV_X1 port map( A => A_ns(43), ZN => n886);
   U83 : OAI221_X1 port map( B1 => n829, B2 => n889, C1 => n828, C2 => n890, A 
                           => n891, ZN => O_44_port);
   U84 : AOI22_X1 port map( A1 => A_ns(43), A2 => n833, B1 => A_s(43), B2 => 
                           n834, ZN => n891);
   U85 : INV_X1 port map( A => A_s(42), ZN => n890);
   U86 : INV_X1 port map( A => A_ns(42), ZN => n889);
   U87 : OAI221_X1 port map( B1 => n829, B2 => n892, C1 => n828, C2 => n893, A 
                           => n894, ZN => O_43_port);
   U88 : AOI22_X1 port map( A1 => A_ns(42), A2 => n833, B1 => A_s(42), B2 => 
                           n834, ZN => n894);
   U89 : INV_X1 port map( A => A_s(41), ZN => n893);
   U90 : INV_X1 port map( A => A_ns(41), ZN => n892);
   U91 : OAI221_X1 port map( B1 => n829, B2 => n895, C1 => n828, C2 => n896, A 
                           => n897, ZN => O_42_port);
   U92 : AOI22_X1 port map( A1 => A_ns(41), A2 => n833, B1 => A_s(41), B2 => 
                           n834, ZN => n897);
   U93 : INV_X1 port map( A => A_s(40), ZN => n896);
   U94 : INV_X1 port map( A => A_ns(40), ZN => n895);
   U95 : OAI221_X1 port map( B1 => n829, B2 => n898, C1 => n828, C2 => n899, A 
                           => n900, ZN => O_41_port);
   U96 : AOI22_X1 port map( A1 => A_ns(40), A2 => n833, B1 => A_s(40), B2 => 
                           n834, ZN => n900);
   U97 : INV_X1 port map( A => A_s(39), ZN => n899);
   U98 : INV_X1 port map( A => A_ns(39), ZN => n898);
   U99 : OAI221_X1 port map( B1 => n829, B2 => n901, C1 => n828, C2 => n902, A 
                           => n903, ZN => O_40_port);
   U100 : AOI22_X1 port map( A1 => A_ns(39), A2 => n833, B1 => A_s(39), B2 => 
                           n834, ZN => n903);
   U101 : INV_X1 port map( A => A_s(38), ZN => n902);
   U102 : INV_X1 port map( A => A_ns(38), ZN => n901);
   U103 : OAI221_X1 port map( B1 => n829, B2 => n904, C1 => n828, C2 => n905, A
                           => n906, ZN => O_3_port);
   U104 : AOI22_X1 port map( A1 => A_ns(2), A2 => n833, B1 => A_s(2), B2 => 
                           n834, ZN => n906);
   U105 : INV_X1 port map( A => A_s(1), ZN => n905);
   U106 : INV_X1 port map( A => A_ns(1), ZN => n904);
   U107 : OAI221_X1 port map( B1 => n829, B2 => n907, C1 => n828, C2 => n908, A
                           => n909, ZN => O_39_port);
   U108 : AOI22_X1 port map( A1 => A_ns(38), A2 => n833, B1 => A_s(38), B2 => 
                           n834, ZN => n909);
   U109 : INV_X1 port map( A => A_s(37), ZN => n908);
   U110 : INV_X1 port map( A => A_ns(37), ZN => n907);
   U111 : OAI221_X1 port map( B1 => n829, B2 => n910, C1 => n828, C2 => n911, A
                           => n912, ZN => O_38_port);
   U112 : AOI22_X1 port map( A1 => A_ns(37), A2 => n833, B1 => A_s(37), B2 => 
                           n834, ZN => n912);
   U113 : INV_X1 port map( A => A_s(36), ZN => n911);
   U114 : INV_X1 port map( A => A_ns(36), ZN => n910);
   U115 : OAI221_X1 port map( B1 => n829, B2 => n913, C1 => n828, C2 => n914, A
                           => n915, ZN => O_37_port);
   U116 : AOI22_X1 port map( A1 => A_ns(36), A2 => n833, B1 => A_s(36), B2 => 
                           n834, ZN => n915);
   U117 : INV_X1 port map( A => A_s(35), ZN => n914);
   U118 : INV_X1 port map( A => A_ns(35), ZN => n913);
   U119 : OAI221_X1 port map( B1 => n829, B2 => n916, C1 => n828, C2 => n917, A
                           => n918, ZN => O_36_port);
   U120 : AOI22_X1 port map( A1 => A_ns(35), A2 => n833, B1 => A_s(35), B2 => 
                           n834, ZN => n918);
   U121 : INV_X1 port map( A => A_s(34), ZN => n917);
   U122 : INV_X1 port map( A => A_ns(34), ZN => n916);
   U123 : OAI221_X1 port map( B1 => n829, B2 => n919, C1 => n828, C2 => n920, A
                           => n921, ZN => O_35_port);
   U124 : AOI22_X1 port map( A1 => A_ns(34), A2 => n833, B1 => A_s(34), B2 => 
                           n834, ZN => n921);
   U125 : INV_X1 port map( A => A_s(33), ZN => n920);
   U126 : INV_X1 port map( A => A_ns(33), ZN => n919);
   U127 : OAI221_X1 port map( B1 => n829, B2 => n922, C1 => n828, C2 => n923, A
                           => n924, ZN => O_34_port);
   U128 : AOI22_X1 port map( A1 => A_ns(33), A2 => n833, B1 => A_s(33), B2 => 
                           n834, ZN => n924);
   U129 : INV_X1 port map( A => A_s(32), ZN => n923);
   U130 : INV_X1 port map( A => A_ns(32), ZN => n922);
   U131 : OAI221_X1 port map( B1 => n829, B2 => n925, C1 => n828, C2 => n926, A
                           => n927, ZN => O_33_port);
   U132 : AOI22_X1 port map( A1 => A_ns(32), A2 => n833, B1 => A_s(32), B2 => 
                           n834, ZN => n927);
   U133 : INV_X1 port map( A => A_s(31), ZN => n926);
   U134 : INV_X1 port map( A => A_ns(31), ZN => n925);
   U135 : OAI221_X1 port map( B1 => n829, B2 => n928, C1 => n828, C2 => n929, A
                           => n930, ZN => O_32_port);
   U136 : AOI22_X1 port map( A1 => A_ns(31), A2 => n833, B1 => A_s(31), B2 => 
                           n834, ZN => n930);
   U137 : INV_X1 port map( A => A_s(30), ZN => n929);
   U138 : INV_X1 port map( A => A_ns(30), ZN => n928);
   U139 : OAI221_X1 port map( B1 => n829, B2 => n931, C1 => n828, C2 => n932, A
                           => n933, ZN => O_31_port);
   U140 : AOI22_X1 port map( A1 => A_ns(30), A2 => n833, B1 => A_s(30), B2 => 
                           n834, ZN => n933);
   U141 : INV_X1 port map( A => A_s(29), ZN => n932);
   U142 : INV_X1 port map( A => A_ns(29), ZN => n931);
   U143 : OAI221_X1 port map( B1 => n829, B2 => n934, C1 => n828, C2 => n935, A
                           => n936, ZN => O_30_port);
   U144 : AOI22_X1 port map( A1 => A_ns(29), A2 => n833, B1 => A_s(29), B2 => 
                           n834, ZN => n936);
   U145 : INV_X1 port map( A => A_s(28), ZN => n935);
   U146 : INV_X1 port map( A => A_ns(28), ZN => n934);
   U147 : OAI221_X1 port map( B1 => n829, B2 => n937, C1 => n828, C2 => n938, A
                           => n939, ZN => O_2_port);
   U148 : AOI22_X1 port map( A1 => A_ns(1), A2 => n833, B1 => A_s(1), B2 => 
                           n834, ZN => n939);
   U149 : OAI221_X1 port map( B1 => n829, B2 => n940, C1 => n828, C2 => n941, A
                           => n942, ZN => O_29_port);
   U150 : AOI22_X1 port map( A1 => A_ns(28), A2 => n833, B1 => A_s(28), B2 => 
                           n834, ZN => n942);
   U151 : INV_X1 port map( A => A_s(27), ZN => n941);
   U152 : INV_X1 port map( A => A_ns(27), ZN => n940);
   U153 : OAI221_X1 port map( B1 => n829, B2 => n943, C1 => n828, C2 => n944, A
                           => n945, ZN => O_28_port);
   U154 : AOI22_X1 port map( A1 => A_ns(27), A2 => n833, B1 => A_s(27), B2 => 
                           n834, ZN => n945);
   U155 : INV_X1 port map( A => A_s(26), ZN => n944);
   U156 : INV_X1 port map( A => A_ns(26), ZN => n943);
   U157 : OAI221_X1 port map( B1 => n829, B2 => n946, C1 => n828, C2 => n947, A
                           => n948, ZN => O_27_port);
   U158 : AOI22_X1 port map( A1 => A_ns(26), A2 => n833, B1 => A_s(26), B2 => 
                           n834, ZN => n948);
   U159 : INV_X1 port map( A => A_s(25), ZN => n947);
   U160 : INV_X1 port map( A => A_ns(25), ZN => n946);
   U161 : OAI221_X1 port map( B1 => n829, B2 => n949, C1 => n828, C2 => n950, A
                           => n951, ZN => O_26_port);
   U162 : AOI22_X1 port map( A1 => A_ns(25), A2 => n833, B1 => A_s(25), B2 => 
                           n834, ZN => n951);
   U163 : INV_X1 port map( A => A_s(24), ZN => n950);
   U164 : INV_X1 port map( A => A_ns(24), ZN => n949);
   U165 : OAI221_X1 port map( B1 => n829, B2 => n952, C1 => n828, C2 => n953, A
                           => n954, ZN => O_25_port);
   U166 : AOI22_X1 port map( A1 => A_ns(24), A2 => n833, B1 => A_s(24), B2 => 
                           n834, ZN => n954);
   U167 : INV_X1 port map( A => A_s(23), ZN => n953);
   U168 : INV_X1 port map( A => A_ns(23), ZN => n952);
   U169 : OAI221_X1 port map( B1 => n829, B2 => n955, C1 => n828, C2 => n956, A
                           => n957, ZN => O_24_port);
   U170 : AOI22_X1 port map( A1 => A_ns(23), A2 => n833, B1 => A_s(23), B2 => 
                           n834, ZN => n957);
   U171 : INV_X1 port map( A => A_s(22), ZN => n956);
   U172 : INV_X1 port map( A => A_ns(22), ZN => n955);
   U173 : OAI221_X1 port map( B1 => n829, B2 => n958, C1 => n828, C2 => n959, A
                           => n960, ZN => O_23_port);
   U174 : AOI22_X1 port map( A1 => A_ns(22), A2 => n833, B1 => A_s(22), B2 => 
                           n834, ZN => n960);
   U175 : INV_X1 port map( A => A_s(21), ZN => n959);
   U176 : INV_X1 port map( A => A_ns(21), ZN => n958);
   U177 : OAI221_X1 port map( B1 => n829, B2 => n961, C1 => n828, C2 => n962, A
                           => n963, ZN => O_22_port);
   U178 : AOI22_X1 port map( A1 => A_ns(21), A2 => n833, B1 => A_s(21), B2 => 
                           n834, ZN => n963);
   U179 : INV_X1 port map( A => A_s(20), ZN => n962);
   U180 : INV_X1 port map( A => A_ns(20), ZN => n961);
   U181 : OAI221_X1 port map( B1 => n829, B2 => n964, C1 => n828, C2 => n965, A
                           => n966, ZN => O_21_port);
   U182 : AOI22_X1 port map( A1 => A_ns(20), A2 => n833, B1 => A_s(20), B2 => 
                           n834, ZN => n966);
   U183 : INV_X1 port map( A => A_s(19), ZN => n965);
   U184 : INV_X1 port map( A => A_ns(19), ZN => n964);
   U185 : OAI221_X1 port map( B1 => n829, B2 => n967, C1 => n828, C2 => n968, A
                           => n969, ZN => O_20_port);
   U186 : AOI22_X1 port map( A1 => A_ns(19), A2 => n833, B1 => A_s(19), B2 => 
                           n834, ZN => n969);
   U187 : INV_X1 port map( A => A_s(18), ZN => n968);
   U188 : INV_X1 port map( A => A_ns(18), ZN => n967);
   U189 : OAI22_X1 port map( A1 => n970, A2 => n938, B1 => n971, B2 => n937, ZN
                           => O_1_port);
   U190 : INV_X1 port map( A => A_ns(0), ZN => n937);
   U191 : INV_X1 port map( A => A_s(0), ZN => n938);
   U192 : OAI221_X1 port map( B1 => n829, B2 => n972, C1 => n828, C2 => n973, A
                           => n974, ZN => O_19_port);
   U193 : AOI22_X1 port map( A1 => A_ns(18), A2 => n833, B1 => A_s(18), B2 => 
                           n834, ZN => n974);
   U194 : INV_X1 port map( A => A_s(17), ZN => n973);
   U195 : INV_X1 port map( A => A_ns(17), ZN => n972);
   U196 : OAI221_X1 port map( B1 => n829, B2 => n975, C1 => n828, C2 => n976, A
                           => n977, ZN => O_18_port);
   U197 : AOI22_X1 port map( A1 => A_ns(17), A2 => n833, B1 => A_s(17), B2 => 
                           n834, ZN => n977);
   U198 : INV_X1 port map( A => A_s(16), ZN => n976);
   U199 : INV_X1 port map( A => A_ns(16), ZN => n975);
   U200 : OAI221_X1 port map( B1 => n829, B2 => n978, C1 => n828, C2 => n979, A
                           => n980, ZN => O_17_port);
   U201 : AOI22_X1 port map( A1 => A_ns(16), A2 => n833, B1 => A_s(16), B2 => 
                           n834, ZN => n980);
   U202 : INV_X1 port map( A => A_s(15), ZN => n979);
   U203 : INV_X1 port map( A => A_ns(15), ZN => n978);
   U204 : OAI221_X1 port map( B1 => n829, B2 => n981, C1 => n828, C2 => n982, A
                           => n983, ZN => O_16_port);
   U205 : AOI22_X1 port map( A1 => A_ns(15), A2 => n833, B1 => A_s(15), B2 => 
                           n834, ZN => n983);
   U206 : INV_X1 port map( A => A_s(14), ZN => n982);
   U207 : INV_X1 port map( A => A_ns(14), ZN => n981);
   U208 : OAI221_X1 port map( B1 => n829, B2 => n984, C1 => n828, C2 => n985, A
                           => n986, ZN => O_15_port);
   U209 : AOI22_X1 port map( A1 => A_ns(14), A2 => n833, B1 => A_s(14), B2 => 
                           n834, ZN => n986);
   U210 : INV_X1 port map( A => A_s(13), ZN => n985);
   U211 : INV_X1 port map( A => A_ns(13), ZN => n984);
   U212 : OAI221_X1 port map( B1 => n829, B2 => n987, C1 => n828, C2 => n988, A
                           => n989, ZN => O_14_port);
   U213 : AOI22_X1 port map( A1 => A_ns(13), A2 => n833, B1 => A_s(13), B2 => 
                           n834, ZN => n989);
   U214 : INV_X1 port map( A => A_s(12), ZN => n988);
   U215 : INV_X1 port map( A => A_ns(12), ZN => n987);
   U216 : OAI221_X1 port map( B1 => n829, B2 => n990, C1 => n828, C2 => n991, A
                           => n992, ZN => O_13_port);
   U217 : AOI22_X1 port map( A1 => A_ns(12), A2 => n833, B1 => A_s(12), B2 => 
                           n834, ZN => n992);
   U218 : INV_X1 port map( A => A_s(11), ZN => n991);
   U219 : INV_X1 port map( A => A_ns(11), ZN => n990);
   U220 : OAI221_X1 port map( B1 => n829, B2 => n993, C1 => n828, C2 => n994, A
                           => n995, ZN => O_12_port);
   U221 : AOI22_X1 port map( A1 => A_ns(11), A2 => n833, B1 => A_s(11), B2 => 
                           n834, ZN => n995);
   U222 : INV_X1 port map( A => A_s(10), ZN => n994);
   U223 : INV_X1 port map( A => A_ns(10), ZN => n993);
   U224 : OAI221_X1 port map( B1 => n829, B2 => n996, C1 => n828, C2 => n997, A
                           => n998, ZN => O_11_port);
   U225 : AOI22_X1 port map( A1 => A_ns(10), A2 => n833, B1 => A_s(10), B2 => 
                           n834, ZN => n998);
   U226 : INV_X1 port map( A => A_s(9), ZN => n997);
   U227 : INV_X1 port map( A => A_ns(9), ZN => n996);
   U228 : OAI221_X1 port map( B1 => n999, B2 => n829, C1 => n1000, C2 => n828, 
                           A => n1001, ZN => O_10_port);
   U229 : AOI22_X1 port map( A1 => A_ns(9), A2 => n833, B1 => A_s(9), B2 => 
                           n834, ZN => n1001);
   U230 : NAND2_X1 port map( A1 => n1002, A2 => n970, ZN => n971);
   U231 : NAND2_X1 port map( A1 => n1002, A2 => n1003, ZN => n970);
   U232 : XOR2_X1 port map( A => B(23), B => B(24), Z => n1002);
   U233 : INV_X1 port map( A => A_s(8), ZN => n1000);
   U234 : INV_X1 port map( A => B(25), ZN => n1003);
   U235 : INV_X1 port map( A => A_ns(8), ZN => n999);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT56_i22 is

   port( A_s, A_ns, B : in std_logic_vector (55 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (55 downto 0));

end BOOTHENC_NBIT56_i22;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT56_i22 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, O_55_port, O_54_port, O_53_port, O_52_port, O_51_port,
      O_50_port, O_49_port, O_48_port, O_47_port, O_46_port, O_45_port, 
      O_44_port, O_43_port, O_42_port, O_41_port, O_40_port, O_39_port, 
      O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, O_33_port, 
      O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, O_27_port, 
      O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, O_21_port, 
      O_20_port, O_19_port, O_18_port, O_17_port, O_16_port, O_15_port, 
      O_14_port, O_13_port, O_12_port, O_11_port, O_9_port, O_8_port, O_7_port,
      O_6_port, O_5_port, O_4_port, O_3_port, O_2_port, O_10_port, n782, n783, 
      n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, 
      n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, 
      n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, 
      n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, 
      n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, 
      n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, 
      n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, 
      n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, 
      n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, 
      n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, 
      n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, 
      n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, 
      n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, 
      n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, 
      n952, O_1_port : std_logic;

begin
   O <= ( O_55_port, O_54_port, O_53_port, O_52_port, O_51_port, O_50_port, 
      O_49_port, O_48_port, O_47_port, O_46_port, O_45_port, O_44_port, 
      O_43_port, O_42_port, O_41_port, O_40_port, O_39_port, O_38_port, 
      O_37_port, O_36_port, O_35_port, O_34_port, O_33_port, O_32_port, 
      O_31_port, O_30_port, O_29_port, O_28_port, O_27_port, O_26_port, 
      O_25_port, O_24_port, O_23_port, O_22_port, O_21_port, O_20_port, 
      O_19_port, O_18_port, O_17_port, O_16_port, O_15_port, O_14_port, 
      O_13_port, O_12_port, O_11_port, O_10_port, O_9_port, O_8_port, O_7_port,
      O_6_port, O_5_port, O_4_port, O_3_port, O_2_port, O_1_port, X_Logic0_port
      );
   A_so <= ( A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), 
      A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), 
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   A_nso <= ( A_ns(53), A_ns(52), A_ns(51), A_ns(50), A_ns(49), A_ns(48), 
      A_ns(47), A_ns(46), A_ns(45), A_ns(44), A_ns(43), A_ns(42), A_ns(41), 
      A_ns(40), A_ns(39), A_ns(38), A_ns(37), A_ns(36), A_ns(35), A_ns(34), 
      A_ns(33), A_ns(32), A_ns(31), A_ns(30), A_ns(29), A_ns(28), A_ns(27), 
      A_ns(26), A_ns(25), A_ns(24), A_ns(23), A_ns(22), A_ns(21), A_ns(20), 
      A_ns(19), A_ns(18), A_ns(17), A_ns(16), A_ns(15), A_ns(14), A_ns(13), 
      A_ns(12), A_ns(11), A_ns(10), A_ns(9), A_ns(8), A_ns(7), A_ns(6), A_ns(5)
      , A_ns(4), A_ns(3), A_ns(2), A_ns(1), A_ns(0), X_Logic0_port, 
      X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : AND3_X1 port map( A1 => B(22), A2 => n952, A3 => B(21), ZN => n782);
   U3 : INV_X4 port map( A => n782, ZN => n783);
   U4 : INV_X4 port map( A => n784, ZN => n793);
   U5 : INV_X4 port map( A => n786, ZN => n792);
   U6 : OR3_X4 port map( A1 => B(21), A2 => B(22), A3 => n952, ZN => n788);
   U7 : OAI22_X1 port map( A1 => n784, A2 => n785, B1 => n786, B2 => n787, ZN 
                           => O_1_port);
   U8 : OAI221_X1 port map( B1 => n788, B2 => n789, C1 => n783, C2 => n790, A 
                           => n791, ZN => O_9_port);
   U9 : AOI22_X1 port map( A1 => A_ns(8), A2 => n792, B1 => A_s(8), B2 => n793,
                           ZN => n791);
   U10 : INV_X1 port map( A => A_s(7), ZN => n790);
   U11 : INV_X1 port map( A => A_ns(7), ZN => n789);
   U12 : OAI221_X1 port map( B1 => n788, B2 => n794, C1 => n783, C2 => n795, A 
                           => n796, ZN => O_8_port);
   U13 : AOI22_X1 port map( A1 => A_ns(7), A2 => n792, B1 => A_s(7), B2 => n793
                           , ZN => n796);
   U14 : INV_X1 port map( A => A_s(6), ZN => n795);
   U15 : INV_X1 port map( A => A_ns(6), ZN => n794);
   U16 : OAI221_X1 port map( B1 => n788, B2 => n797, C1 => n783, C2 => n798, A 
                           => n799, ZN => O_7_port);
   U17 : AOI22_X1 port map( A1 => A_ns(6), A2 => n792, B1 => A_s(6), B2 => n793
                           , ZN => n799);
   U18 : INV_X1 port map( A => A_s(5), ZN => n798);
   U19 : INV_X1 port map( A => A_ns(5), ZN => n797);
   U20 : OAI221_X1 port map( B1 => n788, B2 => n800, C1 => n783, C2 => n801, A 
                           => n802, ZN => O_6_port);
   U21 : AOI22_X1 port map( A1 => A_ns(5), A2 => n792, B1 => A_s(5), B2 => n793
                           , ZN => n802);
   U22 : INV_X1 port map( A => A_s(4), ZN => n801);
   U23 : INV_X1 port map( A => A_ns(4), ZN => n800);
   U24 : OAI221_X1 port map( B1 => n788, B2 => n803, C1 => n783, C2 => n804, A 
                           => n805, ZN => O_5_port);
   U25 : AOI22_X1 port map( A1 => A_ns(4), A2 => n792, B1 => A_s(4), B2 => n793
                           , ZN => n805);
   U26 : INV_X1 port map( A => A_s(3), ZN => n804);
   U27 : INV_X1 port map( A => A_ns(3), ZN => n803);
   U28 : OAI221_X1 port map( B1 => n788, B2 => n806, C1 => n783, C2 => n807, A 
                           => n808, ZN => O_55_port);
   U29 : AOI22_X1 port map( A1 => A_ns(54), A2 => n792, B1 => A_s(54), B2 => 
                           n793, ZN => n808);
   U30 : INV_X1 port map( A => A_s(53), ZN => n807);
   U31 : INV_X1 port map( A => A_ns(53), ZN => n806);
   U32 : OAI221_X1 port map( B1 => n788, B2 => n809, C1 => n783, C2 => n810, A 
                           => n811, ZN => O_54_port);
   U33 : AOI22_X1 port map( A1 => A_ns(53), A2 => n792, B1 => A_s(53), B2 => 
                           n793, ZN => n811);
   U34 : INV_X1 port map( A => A_s(52), ZN => n810);
   U35 : INV_X1 port map( A => A_ns(52), ZN => n809);
   U36 : OAI221_X1 port map( B1 => n788, B2 => n812, C1 => n783, C2 => n813, A 
                           => n814, ZN => O_53_port);
   U37 : AOI22_X1 port map( A1 => A_ns(52), A2 => n792, B1 => A_s(52), B2 => 
                           n793, ZN => n814);
   U38 : INV_X1 port map( A => A_s(51), ZN => n813);
   U39 : INV_X1 port map( A => A_ns(51), ZN => n812);
   U40 : OAI221_X1 port map( B1 => n788, B2 => n815, C1 => n783, C2 => n816, A 
                           => n817, ZN => O_52_port);
   U41 : AOI22_X1 port map( A1 => A_ns(51), A2 => n792, B1 => A_s(51), B2 => 
                           n793, ZN => n817);
   U42 : INV_X1 port map( A => A_s(50), ZN => n816);
   U43 : INV_X1 port map( A => A_ns(50), ZN => n815);
   U44 : OAI221_X1 port map( B1 => n788, B2 => n818, C1 => n783, C2 => n819, A 
                           => n820, ZN => O_51_port);
   U45 : AOI22_X1 port map( A1 => A_ns(50), A2 => n792, B1 => A_s(50), B2 => 
                           n793, ZN => n820);
   U46 : INV_X1 port map( A => A_s(49), ZN => n819);
   U47 : INV_X1 port map( A => A_ns(49), ZN => n818);
   U48 : OAI221_X1 port map( B1 => n788, B2 => n821, C1 => n783, C2 => n822, A 
                           => n823, ZN => O_50_port);
   U49 : AOI22_X1 port map( A1 => A_ns(49), A2 => n792, B1 => A_s(49), B2 => 
                           n793, ZN => n823);
   U50 : INV_X1 port map( A => A_s(48), ZN => n822);
   U51 : INV_X1 port map( A => A_ns(48), ZN => n821);
   U52 : OAI221_X1 port map( B1 => n788, B2 => n824, C1 => n783, C2 => n825, A 
                           => n826, ZN => O_4_port);
   U53 : AOI22_X1 port map( A1 => A_ns(3), A2 => n792, B1 => A_s(3), B2 => n793
                           , ZN => n826);
   U54 : INV_X1 port map( A => A_s(2), ZN => n825);
   U55 : INV_X1 port map( A => A_ns(2), ZN => n824);
   U56 : OAI221_X1 port map( B1 => n788, B2 => n827, C1 => n783, C2 => n828, A 
                           => n829, ZN => O_49_port);
   U57 : AOI22_X1 port map( A1 => A_ns(48), A2 => n792, B1 => A_s(48), B2 => 
                           n793, ZN => n829);
   U58 : INV_X1 port map( A => A_s(47), ZN => n828);
   U59 : INV_X1 port map( A => A_ns(47), ZN => n827);
   U60 : OAI221_X1 port map( B1 => n788, B2 => n830, C1 => n783, C2 => n831, A 
                           => n832, ZN => O_48_port);
   U61 : AOI22_X1 port map( A1 => A_ns(47), A2 => n792, B1 => A_s(47), B2 => 
                           n793, ZN => n832);
   U62 : INV_X1 port map( A => A_s(46), ZN => n831);
   U63 : INV_X1 port map( A => A_ns(46), ZN => n830);
   U64 : OAI221_X1 port map( B1 => n788, B2 => n833, C1 => n783, C2 => n834, A 
                           => n835, ZN => O_47_port);
   U65 : AOI22_X1 port map( A1 => A_ns(46), A2 => n792, B1 => A_s(46), B2 => 
                           n793, ZN => n835);
   U66 : INV_X1 port map( A => A_s(45), ZN => n834);
   U67 : INV_X1 port map( A => A_ns(45), ZN => n833);
   U68 : OAI221_X1 port map( B1 => n788, B2 => n836, C1 => n783, C2 => n837, A 
                           => n838, ZN => O_46_port);
   U69 : AOI22_X1 port map( A1 => A_ns(45), A2 => n792, B1 => A_s(45), B2 => 
                           n793, ZN => n838);
   U70 : INV_X1 port map( A => A_s(44), ZN => n837);
   U71 : INV_X1 port map( A => A_ns(44), ZN => n836);
   U72 : OAI221_X1 port map( B1 => n788, B2 => n839, C1 => n783, C2 => n840, A 
                           => n841, ZN => O_45_port);
   U73 : AOI22_X1 port map( A1 => A_ns(44), A2 => n792, B1 => A_s(44), B2 => 
                           n793, ZN => n841);
   U74 : INV_X1 port map( A => A_s(43), ZN => n840);
   U75 : INV_X1 port map( A => A_ns(43), ZN => n839);
   U76 : OAI221_X1 port map( B1 => n788, B2 => n842, C1 => n783, C2 => n843, A 
                           => n844, ZN => O_44_port);
   U77 : AOI22_X1 port map( A1 => A_ns(43), A2 => n792, B1 => A_s(43), B2 => 
                           n793, ZN => n844);
   U78 : INV_X1 port map( A => A_s(42), ZN => n843);
   U79 : INV_X1 port map( A => A_ns(42), ZN => n842);
   U80 : OAI221_X1 port map( B1 => n788, B2 => n845, C1 => n783, C2 => n846, A 
                           => n847, ZN => O_43_port);
   U81 : AOI22_X1 port map( A1 => A_ns(42), A2 => n792, B1 => A_s(42), B2 => 
                           n793, ZN => n847);
   U82 : INV_X1 port map( A => A_s(41), ZN => n846);
   U83 : INV_X1 port map( A => A_ns(41), ZN => n845);
   U84 : OAI221_X1 port map( B1 => n788, B2 => n848, C1 => n783, C2 => n849, A 
                           => n850, ZN => O_42_port);
   U85 : AOI22_X1 port map( A1 => A_ns(41), A2 => n792, B1 => A_s(41), B2 => 
                           n793, ZN => n850);
   U86 : INV_X1 port map( A => A_s(40), ZN => n849);
   U87 : INV_X1 port map( A => A_ns(40), ZN => n848);
   U88 : OAI221_X1 port map( B1 => n788, B2 => n851, C1 => n783, C2 => n852, A 
                           => n853, ZN => O_41_port);
   U89 : AOI22_X1 port map( A1 => A_ns(40), A2 => n792, B1 => A_s(40), B2 => 
                           n793, ZN => n853);
   U90 : INV_X1 port map( A => A_s(39), ZN => n852);
   U91 : INV_X1 port map( A => A_ns(39), ZN => n851);
   U92 : OAI221_X1 port map( B1 => n788, B2 => n854, C1 => n783, C2 => n855, A 
                           => n856, ZN => O_40_port);
   U93 : AOI22_X1 port map( A1 => A_ns(39), A2 => n792, B1 => A_s(39), B2 => 
                           n793, ZN => n856);
   U94 : INV_X1 port map( A => A_s(38), ZN => n855);
   U95 : INV_X1 port map( A => A_ns(38), ZN => n854);
   U96 : OAI221_X1 port map( B1 => n788, B2 => n857, C1 => n783, C2 => n858, A 
                           => n859, ZN => O_3_port);
   U97 : AOI22_X1 port map( A1 => A_ns(2), A2 => n792, B1 => A_s(2), B2 => n793
                           , ZN => n859);
   U98 : INV_X1 port map( A => A_s(1), ZN => n858);
   U99 : INV_X1 port map( A => A_ns(1), ZN => n857);
   U100 : OAI221_X1 port map( B1 => n788, B2 => n860, C1 => n783, C2 => n861, A
                           => n862, ZN => O_39_port);
   U101 : AOI22_X1 port map( A1 => A_ns(38), A2 => n792, B1 => A_s(38), B2 => 
                           n793, ZN => n862);
   U102 : INV_X1 port map( A => A_s(37), ZN => n861);
   U103 : INV_X1 port map( A => A_ns(37), ZN => n860);
   U104 : OAI221_X1 port map( B1 => n788, B2 => n863, C1 => n783, C2 => n864, A
                           => n865, ZN => O_38_port);
   U105 : AOI22_X1 port map( A1 => A_ns(37), A2 => n792, B1 => A_s(37), B2 => 
                           n793, ZN => n865);
   U106 : INV_X1 port map( A => A_s(36), ZN => n864);
   U107 : INV_X1 port map( A => A_ns(36), ZN => n863);
   U108 : OAI221_X1 port map( B1 => n788, B2 => n866, C1 => n783, C2 => n867, A
                           => n868, ZN => O_37_port);
   U109 : AOI22_X1 port map( A1 => A_ns(36), A2 => n792, B1 => A_s(36), B2 => 
                           n793, ZN => n868);
   U110 : INV_X1 port map( A => A_s(35), ZN => n867);
   U111 : INV_X1 port map( A => A_ns(35), ZN => n866);
   U112 : OAI221_X1 port map( B1 => n788, B2 => n869, C1 => n783, C2 => n870, A
                           => n871, ZN => O_36_port);
   U113 : AOI22_X1 port map( A1 => A_ns(35), A2 => n792, B1 => A_s(35), B2 => 
                           n793, ZN => n871);
   U114 : INV_X1 port map( A => A_s(34), ZN => n870);
   U115 : INV_X1 port map( A => A_ns(34), ZN => n869);
   U116 : OAI221_X1 port map( B1 => n788, B2 => n872, C1 => n783, C2 => n873, A
                           => n874, ZN => O_35_port);
   U117 : AOI22_X1 port map( A1 => A_ns(34), A2 => n792, B1 => A_s(34), B2 => 
                           n793, ZN => n874);
   U118 : INV_X1 port map( A => A_s(33), ZN => n873);
   U119 : INV_X1 port map( A => A_ns(33), ZN => n872);
   U120 : OAI221_X1 port map( B1 => n788, B2 => n875, C1 => n783, C2 => n876, A
                           => n877, ZN => O_34_port);
   U121 : AOI22_X1 port map( A1 => A_ns(33), A2 => n792, B1 => A_s(33), B2 => 
                           n793, ZN => n877);
   U122 : INV_X1 port map( A => A_s(32), ZN => n876);
   U123 : INV_X1 port map( A => A_ns(32), ZN => n875);
   U124 : OAI221_X1 port map( B1 => n788, B2 => n878, C1 => n783, C2 => n879, A
                           => n880, ZN => O_33_port);
   U125 : AOI22_X1 port map( A1 => A_ns(32), A2 => n792, B1 => A_s(32), B2 => 
                           n793, ZN => n880);
   U126 : INV_X1 port map( A => A_s(31), ZN => n879);
   U127 : INV_X1 port map( A => A_ns(31), ZN => n878);
   U128 : OAI221_X1 port map( B1 => n788, B2 => n881, C1 => n783, C2 => n882, A
                           => n883, ZN => O_32_port);
   U129 : AOI22_X1 port map( A1 => A_ns(31), A2 => n792, B1 => A_s(31), B2 => 
                           n793, ZN => n883);
   U130 : INV_X1 port map( A => A_s(30), ZN => n882);
   U131 : INV_X1 port map( A => A_ns(30), ZN => n881);
   U132 : OAI221_X1 port map( B1 => n788, B2 => n884, C1 => n783, C2 => n885, A
                           => n886, ZN => O_31_port);
   U133 : AOI22_X1 port map( A1 => A_ns(30), A2 => n792, B1 => A_s(30), B2 => 
                           n793, ZN => n886);
   U134 : INV_X1 port map( A => A_s(29), ZN => n885);
   U135 : INV_X1 port map( A => A_ns(29), ZN => n884);
   U136 : OAI221_X1 port map( B1 => n788, B2 => n887, C1 => n783, C2 => n888, A
                           => n889, ZN => O_30_port);
   U137 : AOI22_X1 port map( A1 => A_ns(29), A2 => n792, B1 => A_s(29), B2 => 
                           n793, ZN => n889);
   U138 : INV_X1 port map( A => A_s(28), ZN => n888);
   U139 : INV_X1 port map( A => A_ns(28), ZN => n887);
   U140 : OAI221_X1 port map( B1 => n787, B2 => n788, C1 => n785, C2 => n783, A
                           => n890, ZN => O_2_port);
   U141 : AOI22_X1 port map( A1 => A_ns(1), A2 => n792, B1 => A_s(1), B2 => 
                           n793, ZN => n890);
   U142 : INV_X1 port map( A => A_s(0), ZN => n785);
   U143 : INV_X1 port map( A => A_ns(0), ZN => n787);
   U144 : OAI221_X1 port map( B1 => n788, B2 => n891, C1 => n783, C2 => n892, A
                           => n893, ZN => O_29_port);
   U145 : AOI22_X1 port map( A1 => A_ns(28), A2 => n792, B1 => A_s(28), B2 => 
                           n793, ZN => n893);
   U146 : INV_X1 port map( A => A_s(27), ZN => n892);
   U147 : INV_X1 port map( A => A_ns(27), ZN => n891);
   U148 : OAI221_X1 port map( B1 => n788, B2 => n894, C1 => n783, C2 => n895, A
                           => n896, ZN => O_28_port);
   U149 : AOI22_X1 port map( A1 => A_ns(27), A2 => n792, B1 => A_s(27), B2 => 
                           n793, ZN => n896);
   U150 : INV_X1 port map( A => A_s(26), ZN => n895);
   U151 : INV_X1 port map( A => A_ns(26), ZN => n894);
   U152 : OAI221_X1 port map( B1 => n788, B2 => n897, C1 => n783, C2 => n898, A
                           => n899, ZN => O_27_port);
   U153 : AOI22_X1 port map( A1 => A_ns(26), A2 => n792, B1 => A_s(26), B2 => 
                           n793, ZN => n899);
   U154 : INV_X1 port map( A => A_s(25), ZN => n898);
   U155 : INV_X1 port map( A => A_ns(25), ZN => n897);
   U156 : OAI221_X1 port map( B1 => n788, B2 => n900, C1 => n783, C2 => n901, A
                           => n902, ZN => O_26_port);
   U157 : AOI22_X1 port map( A1 => A_ns(25), A2 => n792, B1 => A_s(25), B2 => 
                           n793, ZN => n902);
   U158 : INV_X1 port map( A => A_s(24), ZN => n901);
   U159 : INV_X1 port map( A => A_ns(24), ZN => n900);
   U160 : OAI221_X1 port map( B1 => n788, B2 => n903, C1 => n783, C2 => n904, A
                           => n905, ZN => O_25_port);
   U161 : AOI22_X1 port map( A1 => A_ns(24), A2 => n792, B1 => A_s(24), B2 => 
                           n793, ZN => n905);
   U162 : INV_X1 port map( A => A_s(23), ZN => n904);
   U163 : INV_X1 port map( A => A_ns(23), ZN => n903);
   U164 : OAI221_X1 port map( B1 => n788, B2 => n906, C1 => n783, C2 => n907, A
                           => n908, ZN => O_24_port);
   U165 : AOI22_X1 port map( A1 => A_ns(23), A2 => n792, B1 => A_s(23), B2 => 
                           n793, ZN => n908);
   U166 : INV_X1 port map( A => A_s(22), ZN => n907);
   U167 : INV_X1 port map( A => A_ns(22), ZN => n906);
   U168 : OAI221_X1 port map( B1 => n788, B2 => n909, C1 => n783, C2 => n910, A
                           => n911, ZN => O_23_port);
   U169 : AOI22_X1 port map( A1 => A_ns(22), A2 => n792, B1 => A_s(22), B2 => 
                           n793, ZN => n911);
   U170 : INV_X1 port map( A => A_s(21), ZN => n910);
   U171 : INV_X1 port map( A => A_ns(21), ZN => n909);
   U172 : OAI221_X1 port map( B1 => n788, B2 => n912, C1 => n783, C2 => n913, A
                           => n914, ZN => O_22_port);
   U173 : AOI22_X1 port map( A1 => A_ns(21), A2 => n792, B1 => A_s(21), B2 => 
                           n793, ZN => n914);
   U174 : INV_X1 port map( A => A_s(20), ZN => n913);
   U175 : INV_X1 port map( A => A_ns(20), ZN => n912);
   U176 : OAI221_X1 port map( B1 => n788, B2 => n915, C1 => n783, C2 => n916, A
                           => n917, ZN => O_21_port);
   U177 : AOI22_X1 port map( A1 => A_ns(20), A2 => n792, B1 => A_s(20), B2 => 
                           n793, ZN => n917);
   U178 : INV_X1 port map( A => A_s(19), ZN => n916);
   U179 : INV_X1 port map( A => A_ns(19), ZN => n915);
   U180 : OAI221_X1 port map( B1 => n788, B2 => n918, C1 => n783, C2 => n919, A
                           => n920, ZN => O_20_port);
   U181 : AOI22_X1 port map( A1 => A_ns(19), A2 => n792, B1 => A_s(19), B2 => 
                           n793, ZN => n920);
   U182 : INV_X1 port map( A => A_s(18), ZN => n919);
   U183 : INV_X1 port map( A => A_ns(18), ZN => n918);
   U184 : OAI221_X1 port map( B1 => n788, B2 => n921, C1 => n783, C2 => n922, A
                           => n923, ZN => O_19_port);
   U185 : AOI22_X1 port map( A1 => A_ns(18), A2 => n792, B1 => A_s(18), B2 => 
                           n793, ZN => n923);
   U186 : INV_X1 port map( A => A_s(17), ZN => n922);
   U187 : INV_X1 port map( A => A_ns(17), ZN => n921);
   U188 : OAI221_X1 port map( B1 => n788, B2 => n924, C1 => n783, C2 => n925, A
                           => n926, ZN => O_18_port);
   U189 : AOI22_X1 port map( A1 => A_ns(17), A2 => n792, B1 => A_s(17), B2 => 
                           n793, ZN => n926);
   U190 : INV_X1 port map( A => A_s(16), ZN => n925);
   U191 : INV_X1 port map( A => A_ns(16), ZN => n924);
   U192 : OAI221_X1 port map( B1 => n788, B2 => n927, C1 => n783, C2 => n928, A
                           => n929, ZN => O_17_port);
   U193 : AOI22_X1 port map( A1 => A_ns(16), A2 => n792, B1 => A_s(16), B2 => 
                           n793, ZN => n929);
   U194 : INV_X1 port map( A => A_s(15), ZN => n928);
   U195 : INV_X1 port map( A => A_ns(15), ZN => n927);
   U196 : OAI221_X1 port map( B1 => n788, B2 => n930, C1 => n783, C2 => n931, A
                           => n932, ZN => O_16_port);
   U197 : AOI22_X1 port map( A1 => A_ns(15), A2 => n792, B1 => A_s(15), B2 => 
                           n793, ZN => n932);
   U198 : INV_X1 port map( A => A_s(14), ZN => n931);
   U199 : INV_X1 port map( A => A_ns(14), ZN => n930);
   U200 : OAI221_X1 port map( B1 => n788, B2 => n933, C1 => n783, C2 => n934, A
                           => n935, ZN => O_15_port);
   U201 : AOI22_X1 port map( A1 => A_ns(14), A2 => n792, B1 => A_s(14), B2 => 
                           n793, ZN => n935);
   U202 : INV_X1 port map( A => A_s(13), ZN => n934);
   U203 : INV_X1 port map( A => A_ns(13), ZN => n933);
   U204 : OAI221_X1 port map( B1 => n788, B2 => n936, C1 => n783, C2 => n937, A
                           => n938, ZN => O_14_port);
   U205 : AOI22_X1 port map( A1 => A_ns(13), A2 => n792, B1 => A_s(13), B2 => 
                           n793, ZN => n938);
   U206 : INV_X1 port map( A => A_s(12), ZN => n937);
   U207 : INV_X1 port map( A => A_ns(12), ZN => n936);
   U208 : OAI221_X1 port map( B1 => n788, B2 => n939, C1 => n783, C2 => n940, A
                           => n941, ZN => O_13_port);
   U209 : AOI22_X1 port map( A1 => A_ns(12), A2 => n792, B1 => A_s(12), B2 => 
                           n793, ZN => n941);
   U210 : INV_X1 port map( A => A_s(11), ZN => n940);
   U211 : INV_X1 port map( A => A_ns(11), ZN => n939);
   U212 : OAI221_X1 port map( B1 => n788, B2 => n942, C1 => n783, C2 => n943, A
                           => n944, ZN => O_12_port);
   U213 : AOI22_X1 port map( A1 => A_ns(11), A2 => n792, B1 => A_s(11), B2 => 
                           n793, ZN => n944);
   U214 : INV_X1 port map( A => A_s(10), ZN => n943);
   U215 : INV_X1 port map( A => A_ns(10), ZN => n942);
   U216 : OAI221_X1 port map( B1 => n788, B2 => n945, C1 => n783, C2 => n946, A
                           => n947, ZN => O_11_port);
   U217 : AOI22_X1 port map( A1 => A_ns(10), A2 => n792, B1 => A_s(10), B2 => 
                           n793, ZN => n947);
   U218 : INV_X1 port map( A => A_s(9), ZN => n946);
   U219 : INV_X1 port map( A => A_ns(9), ZN => n945);
   U220 : OAI221_X1 port map( B1 => n948, B2 => n788, C1 => n949, C2 => n783, A
                           => n950, ZN => O_10_port);
   U221 : AOI22_X1 port map( A1 => A_ns(9), A2 => n792, B1 => A_s(9), B2 => 
                           n793, ZN => n950);
   U222 : NAND2_X1 port map( A1 => n951, A2 => n784, ZN => n786);
   U223 : NAND2_X1 port map( A1 => n951, A2 => n952, ZN => n784);
   U224 : XOR2_X1 port map( A => B(21), B => B(22), Z => n951);
   U225 : INV_X1 port map( A => A_s(8), ZN => n949);
   U226 : INV_X1 port map( A => B(23), ZN => n952);
   U227 : INV_X1 port map( A => A_ns(8), ZN => n948);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT54_i20 is

   port( A_s, A_ns, B : in std_logic_vector (53 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (53 downto 0));

end BOOTHENC_NBIT54_i20;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT54_i20 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, O_53_port, O_52_port, O_51_port, O_50_port, O_49_port,
      O_48_port, O_47_port, O_46_port, O_45_port, O_44_port, O_43_port, 
      O_42_port, O_41_port, O_40_port, O_39_port, O_38_port, O_37_port, 
      O_36_port, O_35_port, O_34_port, O_33_port, O_32_port, O_31_port, 
      O_30_port, O_29_port, O_28_port, O_27_port, O_26_port, O_25_port, 
      O_24_port, O_23_port, O_22_port, O_21_port, O_20_port, O_19_port, 
      O_18_port, O_17_port, O_16_port, O_15_port, O_14_port, O_13_port, 
      O_12_port, O_11_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, 
      O_4_port, O_3_port, O_2_port, O_10_port, n759, n760, n761, n762, n763, 
      n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, 
      n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, 
      n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, 
      n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, 
      n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, 
      n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, 
      n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, 
      n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, 
      n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, 
      n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, 
      n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, 
      n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, 
      n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, 
      n920, n921, n922, n923, n924, O_1_port : std_logic;

begin
   O <= ( O_53_port, O_52_port, O_51_port, O_50_port, O_49_port, O_48_port, 
      O_47_port, O_46_port, O_45_port, O_44_port, O_43_port, O_42_port, 
      O_41_port, O_40_port, O_39_port, O_38_port, O_37_port, O_36_port, 
      O_35_port, O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, 
      O_29_port, O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, 
      O_23_port, O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, 
      O_17_port, O_16_port, O_15_port, O_14_port, O_13_port, O_12_port, 
      O_11_port, O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, 
      O_4_port, O_3_port, O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), A_s(46), A_s(45), 
      A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), A_s(38), A_s(37), 
      A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), A_s(30), A_s(29), 
      A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), A_s(22), A_s(21), 
      A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), A_s(14), A_s(13), 
      A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), A_s(6), A_s(5), A_s(4)
      , A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, X_Logic0_port );
   A_nso <= ( A_ns(51), A_ns(50), A_ns(49), A_ns(48), A_ns(47), A_ns(46), 
      A_ns(45), A_ns(44), A_ns(43), A_ns(42), A_ns(41), A_ns(40), A_ns(39), 
      A_ns(38), A_ns(37), A_ns(36), A_ns(35), A_ns(34), A_ns(33), A_ns(32), 
      A_ns(31), A_ns(30), A_ns(29), A_ns(28), A_ns(27), A_ns(26), A_ns(25), 
      A_ns(24), A_ns(23), A_ns(22), A_ns(21), A_ns(20), A_ns(19), A_ns(18), 
      A_ns(17), A_ns(16), A_ns(15), A_ns(14), A_ns(13), A_ns(12), A_ns(11), 
      A_ns(10), A_ns(9), A_ns(8), A_ns(7), A_ns(6), A_ns(5), A_ns(4), A_ns(3), 
      A_ns(2), A_ns(1), A_ns(0), X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : AND3_X1 port map( A1 => B(20), A2 => n924, A3 => B(19), ZN => n759);
   U3 : INV_X1 port map( A => n759, ZN => n760);
   U4 : INV_X1 port map( A => n759, ZN => n761);
   U5 : INV_X4 port map( A => n762, ZN => n771);
   U6 : INV_X4 port map( A => n764, ZN => n770);
   U7 : OR3_X4 port map( A1 => B(19), A2 => B(20), A3 => n924, ZN => n766);
   U8 : OAI22_X1 port map( A1 => n762, A2 => n763, B1 => n764, B2 => n765, ZN 
                           => O_1_port);
   U9 : OAI221_X1 port map( B1 => n766, B2 => n767, C1 => n761, C2 => n768, A 
                           => n769, ZN => O_9_port);
   U10 : AOI22_X1 port map( A1 => A_ns(8), A2 => n770, B1 => A_s(8), B2 => n771
                           , ZN => n769);
   U11 : INV_X1 port map( A => A_s(7), ZN => n768);
   U12 : INV_X1 port map( A => A_ns(7), ZN => n767);
   U13 : OAI221_X1 port map( B1 => n766, B2 => n772, C1 => n760, C2 => n773, A 
                           => n774, ZN => O_8_port);
   U14 : AOI22_X1 port map( A1 => A_ns(7), A2 => n770, B1 => A_s(7), B2 => n771
                           , ZN => n774);
   U15 : INV_X1 port map( A => A_s(6), ZN => n773);
   U16 : INV_X1 port map( A => A_ns(6), ZN => n772);
   U17 : OAI221_X1 port map( B1 => n766, B2 => n775, C1 => n761, C2 => n776, A 
                           => n777, ZN => O_7_port);
   U18 : AOI22_X1 port map( A1 => A_ns(6), A2 => n770, B1 => A_s(6), B2 => n771
                           , ZN => n777);
   U19 : INV_X1 port map( A => A_s(5), ZN => n776);
   U20 : INV_X1 port map( A => A_ns(5), ZN => n775);
   U21 : OAI221_X1 port map( B1 => n766, B2 => n778, C1 => n760, C2 => n779, A 
                           => n780, ZN => O_6_port);
   U22 : AOI22_X1 port map( A1 => A_ns(5), A2 => n770, B1 => A_s(5), B2 => n771
                           , ZN => n780);
   U23 : INV_X1 port map( A => A_s(4), ZN => n779);
   U24 : INV_X1 port map( A => A_ns(4), ZN => n778);
   U25 : OAI221_X1 port map( B1 => n766, B2 => n781, C1 => n761, C2 => n782, A 
                           => n783, ZN => O_5_port);
   U26 : AOI22_X1 port map( A1 => A_ns(4), A2 => n770, B1 => A_s(4), B2 => n771
                           , ZN => n783);
   U27 : INV_X1 port map( A => A_s(3), ZN => n782);
   U28 : INV_X1 port map( A => A_ns(3), ZN => n781);
   U29 : OAI221_X1 port map( B1 => n766, B2 => n784, C1 => n760, C2 => n785, A 
                           => n786, ZN => O_53_port);
   U30 : AOI22_X1 port map( A1 => A_ns(52), A2 => n770, B1 => A_s(52), B2 => 
                           n771, ZN => n786);
   U31 : INV_X1 port map( A => A_s(51), ZN => n785);
   U32 : INV_X1 port map( A => A_ns(51), ZN => n784);
   U33 : OAI221_X1 port map( B1 => n766, B2 => n787, C1 => n761, C2 => n788, A 
                           => n789, ZN => O_52_port);
   U34 : AOI22_X1 port map( A1 => A_ns(51), A2 => n770, B1 => A_s(51), B2 => 
                           n771, ZN => n789);
   U35 : INV_X1 port map( A => A_s(50), ZN => n788);
   U36 : INV_X1 port map( A => A_ns(50), ZN => n787);
   U37 : OAI221_X1 port map( B1 => n766, B2 => n790, C1 => n760, C2 => n791, A 
                           => n792, ZN => O_51_port);
   U38 : AOI22_X1 port map( A1 => A_ns(50), A2 => n770, B1 => A_s(50), B2 => 
                           n771, ZN => n792);
   U39 : INV_X1 port map( A => A_s(49), ZN => n791);
   U40 : INV_X1 port map( A => A_ns(49), ZN => n790);
   U41 : OAI221_X1 port map( B1 => n766, B2 => n793, C1 => n761, C2 => n794, A 
                           => n795, ZN => O_50_port);
   U42 : AOI22_X1 port map( A1 => A_ns(49), A2 => n770, B1 => A_s(49), B2 => 
                           n771, ZN => n795);
   U43 : INV_X1 port map( A => A_s(48), ZN => n794);
   U44 : INV_X1 port map( A => A_ns(48), ZN => n793);
   U45 : OAI221_X1 port map( B1 => n766, B2 => n796, C1 => n760, C2 => n797, A 
                           => n798, ZN => O_4_port);
   U46 : AOI22_X1 port map( A1 => A_ns(3), A2 => n770, B1 => A_s(3), B2 => n771
                           , ZN => n798);
   U47 : INV_X1 port map( A => A_s(2), ZN => n797);
   U48 : INV_X1 port map( A => A_ns(2), ZN => n796);
   U49 : OAI221_X1 port map( B1 => n766, B2 => n799, C1 => n761, C2 => n800, A 
                           => n801, ZN => O_49_port);
   U50 : AOI22_X1 port map( A1 => A_ns(48), A2 => n770, B1 => A_s(48), B2 => 
                           n771, ZN => n801);
   U51 : INV_X1 port map( A => A_s(47), ZN => n800);
   U52 : INV_X1 port map( A => A_ns(47), ZN => n799);
   U53 : OAI221_X1 port map( B1 => n766, B2 => n802, C1 => n760, C2 => n803, A 
                           => n804, ZN => O_48_port);
   U54 : AOI22_X1 port map( A1 => A_ns(47), A2 => n770, B1 => A_s(47), B2 => 
                           n771, ZN => n804);
   U55 : INV_X1 port map( A => A_s(46), ZN => n803);
   U56 : INV_X1 port map( A => A_ns(46), ZN => n802);
   U57 : OAI221_X1 port map( B1 => n766, B2 => n805, C1 => n761, C2 => n806, A 
                           => n807, ZN => O_47_port);
   U58 : AOI22_X1 port map( A1 => A_ns(46), A2 => n770, B1 => A_s(46), B2 => 
                           n771, ZN => n807);
   U59 : INV_X1 port map( A => A_s(45), ZN => n806);
   U60 : INV_X1 port map( A => A_ns(45), ZN => n805);
   U61 : OAI221_X1 port map( B1 => n766, B2 => n808, C1 => n760, C2 => n809, A 
                           => n810, ZN => O_46_port);
   U62 : AOI22_X1 port map( A1 => A_ns(45), A2 => n770, B1 => A_s(45), B2 => 
                           n771, ZN => n810);
   U63 : INV_X1 port map( A => A_s(44), ZN => n809);
   U64 : INV_X1 port map( A => A_ns(44), ZN => n808);
   U65 : OAI221_X1 port map( B1 => n766, B2 => n811, C1 => n761, C2 => n812, A 
                           => n813, ZN => O_45_port);
   U66 : AOI22_X1 port map( A1 => A_ns(44), A2 => n770, B1 => A_s(44), B2 => 
                           n771, ZN => n813);
   U67 : INV_X1 port map( A => A_s(43), ZN => n812);
   U68 : INV_X1 port map( A => A_ns(43), ZN => n811);
   U69 : OAI221_X1 port map( B1 => n766, B2 => n814, C1 => n760, C2 => n815, A 
                           => n816, ZN => O_44_port);
   U70 : AOI22_X1 port map( A1 => A_ns(43), A2 => n770, B1 => A_s(43), B2 => 
                           n771, ZN => n816);
   U71 : INV_X1 port map( A => A_s(42), ZN => n815);
   U72 : INV_X1 port map( A => A_ns(42), ZN => n814);
   U73 : OAI221_X1 port map( B1 => n766, B2 => n817, C1 => n761, C2 => n818, A 
                           => n819, ZN => O_43_port);
   U74 : AOI22_X1 port map( A1 => A_ns(42), A2 => n770, B1 => A_s(42), B2 => 
                           n771, ZN => n819);
   U75 : INV_X1 port map( A => A_s(41), ZN => n818);
   U76 : INV_X1 port map( A => A_ns(41), ZN => n817);
   U77 : OAI221_X1 port map( B1 => n766, B2 => n820, C1 => n760, C2 => n821, A 
                           => n822, ZN => O_42_port);
   U78 : AOI22_X1 port map( A1 => A_ns(41), A2 => n770, B1 => A_s(41), B2 => 
                           n771, ZN => n822);
   U79 : INV_X1 port map( A => A_s(40), ZN => n821);
   U80 : INV_X1 port map( A => A_ns(40), ZN => n820);
   U81 : OAI221_X1 port map( B1 => n766, B2 => n823, C1 => n761, C2 => n824, A 
                           => n825, ZN => O_41_port);
   U82 : AOI22_X1 port map( A1 => A_ns(40), A2 => n770, B1 => A_s(40), B2 => 
                           n771, ZN => n825);
   U83 : INV_X1 port map( A => A_s(39), ZN => n824);
   U84 : INV_X1 port map( A => A_ns(39), ZN => n823);
   U85 : OAI221_X1 port map( B1 => n766, B2 => n826, C1 => n760, C2 => n827, A 
                           => n828, ZN => O_40_port);
   U86 : AOI22_X1 port map( A1 => A_ns(39), A2 => n770, B1 => A_s(39), B2 => 
                           n771, ZN => n828);
   U87 : INV_X1 port map( A => A_s(38), ZN => n827);
   U88 : INV_X1 port map( A => A_ns(38), ZN => n826);
   U89 : OAI221_X1 port map( B1 => n766, B2 => n829, C1 => n761, C2 => n830, A 
                           => n831, ZN => O_3_port);
   U90 : AOI22_X1 port map( A1 => A_ns(2), A2 => n770, B1 => A_s(2), B2 => n771
                           , ZN => n831);
   U91 : INV_X1 port map( A => A_s(1), ZN => n830);
   U92 : INV_X1 port map( A => A_ns(1), ZN => n829);
   U93 : OAI221_X1 port map( B1 => n766, B2 => n832, C1 => n760, C2 => n833, A 
                           => n834, ZN => O_39_port);
   U94 : AOI22_X1 port map( A1 => A_ns(38), A2 => n770, B1 => A_s(38), B2 => 
                           n771, ZN => n834);
   U95 : INV_X1 port map( A => A_s(37), ZN => n833);
   U96 : INV_X1 port map( A => A_ns(37), ZN => n832);
   U97 : OAI221_X1 port map( B1 => n766, B2 => n835, C1 => n761, C2 => n836, A 
                           => n837, ZN => O_38_port);
   U98 : AOI22_X1 port map( A1 => A_ns(37), A2 => n770, B1 => A_s(37), B2 => 
                           n771, ZN => n837);
   U99 : INV_X1 port map( A => A_s(36), ZN => n836);
   U100 : INV_X1 port map( A => A_ns(36), ZN => n835);
   U101 : OAI221_X1 port map( B1 => n766, B2 => n838, C1 => n760, C2 => n839, A
                           => n840, ZN => O_37_port);
   U102 : AOI22_X1 port map( A1 => A_ns(36), A2 => n770, B1 => A_s(36), B2 => 
                           n771, ZN => n840);
   U103 : INV_X1 port map( A => A_s(35), ZN => n839);
   U104 : INV_X1 port map( A => A_ns(35), ZN => n838);
   U105 : OAI221_X1 port map( B1 => n766, B2 => n841, C1 => n761, C2 => n842, A
                           => n843, ZN => O_36_port);
   U106 : AOI22_X1 port map( A1 => A_ns(35), A2 => n770, B1 => A_s(35), B2 => 
                           n771, ZN => n843);
   U107 : INV_X1 port map( A => A_s(34), ZN => n842);
   U108 : INV_X1 port map( A => A_ns(34), ZN => n841);
   U109 : OAI221_X1 port map( B1 => n766, B2 => n844, C1 => n760, C2 => n845, A
                           => n846, ZN => O_35_port);
   U110 : AOI22_X1 port map( A1 => A_ns(34), A2 => n770, B1 => A_s(34), B2 => 
                           n771, ZN => n846);
   U111 : INV_X1 port map( A => A_s(33), ZN => n845);
   U112 : INV_X1 port map( A => A_ns(33), ZN => n844);
   U113 : OAI221_X1 port map( B1 => n766, B2 => n847, C1 => n761, C2 => n848, A
                           => n849, ZN => O_34_port);
   U114 : AOI22_X1 port map( A1 => A_ns(33), A2 => n770, B1 => A_s(33), B2 => 
                           n771, ZN => n849);
   U115 : INV_X1 port map( A => A_s(32), ZN => n848);
   U116 : INV_X1 port map( A => A_ns(32), ZN => n847);
   U117 : OAI221_X1 port map( B1 => n766, B2 => n850, C1 => n760, C2 => n851, A
                           => n852, ZN => O_33_port);
   U118 : AOI22_X1 port map( A1 => A_ns(32), A2 => n770, B1 => A_s(32), B2 => 
                           n771, ZN => n852);
   U119 : INV_X1 port map( A => A_s(31), ZN => n851);
   U120 : INV_X1 port map( A => A_ns(31), ZN => n850);
   U121 : OAI221_X1 port map( B1 => n766, B2 => n853, C1 => n761, C2 => n854, A
                           => n855, ZN => O_32_port);
   U122 : AOI22_X1 port map( A1 => A_ns(31), A2 => n770, B1 => A_s(31), B2 => 
                           n771, ZN => n855);
   U123 : INV_X1 port map( A => A_s(30), ZN => n854);
   U124 : INV_X1 port map( A => A_ns(30), ZN => n853);
   U125 : OAI221_X1 port map( B1 => n766, B2 => n856, C1 => n760, C2 => n857, A
                           => n858, ZN => O_31_port);
   U126 : AOI22_X1 port map( A1 => A_ns(30), A2 => n770, B1 => A_s(30), B2 => 
                           n771, ZN => n858);
   U127 : INV_X1 port map( A => A_s(29), ZN => n857);
   U128 : INV_X1 port map( A => A_ns(29), ZN => n856);
   U129 : OAI221_X1 port map( B1 => n766, B2 => n859, C1 => n761, C2 => n860, A
                           => n861, ZN => O_30_port);
   U130 : AOI22_X1 port map( A1 => A_ns(29), A2 => n770, B1 => A_s(29), B2 => 
                           n771, ZN => n861);
   U131 : INV_X1 port map( A => A_s(28), ZN => n860);
   U132 : INV_X1 port map( A => A_ns(28), ZN => n859);
   U133 : OAI221_X1 port map( B1 => n765, B2 => n766, C1 => n763, C2 => n761, A
                           => n862, ZN => O_2_port);
   U134 : AOI22_X1 port map( A1 => A_ns(1), A2 => n770, B1 => A_s(1), B2 => 
                           n771, ZN => n862);
   U135 : INV_X1 port map( A => A_s(0), ZN => n763);
   U136 : INV_X1 port map( A => A_ns(0), ZN => n765);
   U137 : OAI221_X1 port map( B1 => n766, B2 => n863, C1 => n760, C2 => n864, A
                           => n865, ZN => O_29_port);
   U138 : AOI22_X1 port map( A1 => A_ns(28), A2 => n770, B1 => A_s(28), B2 => 
                           n771, ZN => n865);
   U139 : INV_X1 port map( A => A_s(27), ZN => n864);
   U140 : INV_X1 port map( A => A_ns(27), ZN => n863);
   U141 : OAI221_X1 port map( B1 => n766, B2 => n866, C1 => n761, C2 => n867, A
                           => n868, ZN => O_28_port);
   U142 : AOI22_X1 port map( A1 => A_ns(27), A2 => n770, B1 => A_s(27), B2 => 
                           n771, ZN => n868);
   U143 : INV_X1 port map( A => A_s(26), ZN => n867);
   U144 : INV_X1 port map( A => A_ns(26), ZN => n866);
   U145 : OAI221_X1 port map( B1 => n766, B2 => n869, C1 => n760, C2 => n870, A
                           => n871, ZN => O_27_port);
   U146 : AOI22_X1 port map( A1 => A_ns(26), A2 => n770, B1 => A_s(26), B2 => 
                           n771, ZN => n871);
   U147 : INV_X1 port map( A => A_s(25), ZN => n870);
   U148 : INV_X1 port map( A => A_ns(25), ZN => n869);
   U149 : OAI221_X1 port map( B1 => n766, B2 => n872, C1 => n761, C2 => n873, A
                           => n874, ZN => O_26_port);
   U150 : AOI22_X1 port map( A1 => A_ns(25), A2 => n770, B1 => A_s(25), B2 => 
                           n771, ZN => n874);
   U151 : INV_X1 port map( A => A_s(24), ZN => n873);
   U152 : INV_X1 port map( A => A_ns(24), ZN => n872);
   U153 : OAI221_X1 port map( B1 => n766, B2 => n875, C1 => n760, C2 => n876, A
                           => n877, ZN => O_25_port);
   U154 : AOI22_X1 port map( A1 => A_ns(24), A2 => n770, B1 => A_s(24), B2 => 
                           n771, ZN => n877);
   U155 : INV_X1 port map( A => A_s(23), ZN => n876);
   U156 : INV_X1 port map( A => A_ns(23), ZN => n875);
   U157 : OAI221_X1 port map( B1 => n766, B2 => n878, C1 => n761, C2 => n879, A
                           => n880, ZN => O_24_port);
   U158 : AOI22_X1 port map( A1 => A_ns(23), A2 => n770, B1 => A_s(23), B2 => 
                           n771, ZN => n880);
   U159 : INV_X1 port map( A => A_s(22), ZN => n879);
   U160 : INV_X1 port map( A => A_ns(22), ZN => n878);
   U161 : OAI221_X1 port map( B1 => n766, B2 => n881, C1 => n760, C2 => n882, A
                           => n883, ZN => O_23_port);
   U162 : AOI22_X1 port map( A1 => A_ns(22), A2 => n770, B1 => A_s(22), B2 => 
                           n771, ZN => n883);
   U163 : INV_X1 port map( A => A_s(21), ZN => n882);
   U164 : INV_X1 port map( A => A_ns(21), ZN => n881);
   U165 : OAI221_X1 port map( B1 => n766, B2 => n884, C1 => n761, C2 => n885, A
                           => n886, ZN => O_22_port);
   U166 : AOI22_X1 port map( A1 => A_ns(21), A2 => n770, B1 => A_s(21), B2 => 
                           n771, ZN => n886);
   U167 : INV_X1 port map( A => A_s(20), ZN => n885);
   U168 : INV_X1 port map( A => A_ns(20), ZN => n884);
   U169 : OAI221_X1 port map( B1 => n766, B2 => n887, C1 => n760, C2 => n888, A
                           => n889, ZN => O_21_port);
   U170 : AOI22_X1 port map( A1 => A_ns(20), A2 => n770, B1 => A_s(20), B2 => 
                           n771, ZN => n889);
   U171 : INV_X1 port map( A => A_s(19), ZN => n888);
   U172 : INV_X1 port map( A => A_ns(19), ZN => n887);
   U173 : OAI221_X1 port map( B1 => n766, B2 => n890, C1 => n761, C2 => n891, A
                           => n892, ZN => O_20_port);
   U174 : AOI22_X1 port map( A1 => A_ns(19), A2 => n770, B1 => A_s(19), B2 => 
                           n771, ZN => n892);
   U175 : INV_X1 port map( A => A_s(18), ZN => n891);
   U176 : INV_X1 port map( A => A_ns(18), ZN => n890);
   U177 : OAI221_X1 port map( B1 => n766, B2 => n893, C1 => n760, C2 => n894, A
                           => n895, ZN => O_19_port);
   U178 : AOI22_X1 port map( A1 => A_ns(18), A2 => n770, B1 => A_s(18), B2 => 
                           n771, ZN => n895);
   U179 : INV_X1 port map( A => A_s(17), ZN => n894);
   U180 : INV_X1 port map( A => A_ns(17), ZN => n893);
   U181 : OAI221_X1 port map( B1 => n766, B2 => n896, C1 => n761, C2 => n897, A
                           => n898, ZN => O_18_port);
   U182 : AOI22_X1 port map( A1 => A_ns(17), A2 => n770, B1 => A_s(17), B2 => 
                           n771, ZN => n898);
   U183 : INV_X1 port map( A => A_s(16), ZN => n897);
   U184 : INV_X1 port map( A => A_ns(16), ZN => n896);
   U185 : OAI221_X1 port map( B1 => n766, B2 => n899, C1 => n760, C2 => n900, A
                           => n901, ZN => O_17_port);
   U186 : AOI22_X1 port map( A1 => A_ns(16), A2 => n770, B1 => A_s(16), B2 => 
                           n771, ZN => n901);
   U187 : INV_X1 port map( A => A_s(15), ZN => n900);
   U188 : INV_X1 port map( A => A_ns(15), ZN => n899);
   U189 : OAI221_X1 port map( B1 => n766, B2 => n902, C1 => n761, C2 => n903, A
                           => n904, ZN => O_16_port);
   U190 : AOI22_X1 port map( A1 => A_ns(15), A2 => n770, B1 => A_s(15), B2 => 
                           n771, ZN => n904);
   U191 : INV_X1 port map( A => A_s(14), ZN => n903);
   U192 : INV_X1 port map( A => A_ns(14), ZN => n902);
   U193 : OAI221_X1 port map( B1 => n766, B2 => n905, C1 => n760, C2 => n906, A
                           => n907, ZN => O_15_port);
   U194 : AOI22_X1 port map( A1 => A_ns(14), A2 => n770, B1 => A_s(14), B2 => 
                           n771, ZN => n907);
   U195 : INV_X1 port map( A => A_s(13), ZN => n906);
   U196 : INV_X1 port map( A => A_ns(13), ZN => n905);
   U197 : OAI221_X1 port map( B1 => n766, B2 => n908, C1 => n761, C2 => n909, A
                           => n910, ZN => O_14_port);
   U198 : AOI22_X1 port map( A1 => A_ns(13), A2 => n770, B1 => A_s(13), B2 => 
                           n771, ZN => n910);
   U199 : INV_X1 port map( A => A_s(12), ZN => n909);
   U200 : INV_X1 port map( A => A_ns(12), ZN => n908);
   U201 : OAI221_X1 port map( B1 => n766, B2 => n911, C1 => n760, C2 => n912, A
                           => n913, ZN => O_13_port);
   U202 : AOI22_X1 port map( A1 => A_ns(12), A2 => n770, B1 => A_s(12), B2 => 
                           n771, ZN => n913);
   U203 : INV_X1 port map( A => A_s(11), ZN => n912);
   U204 : INV_X1 port map( A => A_ns(11), ZN => n911);
   U205 : OAI221_X1 port map( B1 => n766, B2 => n914, C1 => n761, C2 => n915, A
                           => n916, ZN => O_12_port);
   U206 : AOI22_X1 port map( A1 => A_ns(11), A2 => n770, B1 => A_s(11), B2 => 
                           n771, ZN => n916);
   U207 : INV_X1 port map( A => A_s(10), ZN => n915);
   U208 : INV_X1 port map( A => A_ns(10), ZN => n914);
   U209 : OAI221_X1 port map( B1 => n766, B2 => n917, C1 => n760, C2 => n918, A
                           => n919, ZN => O_11_port);
   U210 : AOI22_X1 port map( A1 => A_ns(10), A2 => n770, B1 => A_s(10), B2 => 
                           n771, ZN => n919);
   U211 : INV_X1 port map( A => A_s(9), ZN => n918);
   U212 : INV_X1 port map( A => A_ns(9), ZN => n917);
   U213 : OAI221_X1 port map( B1 => n920, B2 => n766, C1 => n921, C2 => n760, A
                           => n922, ZN => O_10_port);
   U214 : AOI22_X1 port map( A1 => A_ns(9), A2 => n770, B1 => A_s(9), B2 => 
                           n771, ZN => n922);
   U215 : NAND2_X1 port map( A1 => n923, A2 => n762, ZN => n764);
   U216 : NAND2_X1 port map( A1 => n923, A2 => n924, ZN => n762);
   U217 : XOR2_X1 port map( A => B(19), B => B(20), Z => n923);
   U218 : INV_X1 port map( A => A_s(8), ZN => n921);
   U219 : INV_X1 port map( A => B(21), ZN => n924);
   U220 : INV_X1 port map( A => A_ns(8), ZN => n920);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT52_i18 is

   port( A_s, A_ns, B : in std_logic_vector (51 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (51 downto 0));

end BOOTHENC_NBIT52_i18;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT52_i18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, O_49_port, O_50_port, O_51_port, O_48_port, O_47_port,
      O_46_port, O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, 
      O_40_port, O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, 
      O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, 
      O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, 
      O_22_port, O_21_port, O_20_port, O_19_port, O_2_port, O_3_port, O_4_port,
      O_5_port, O_6_port, O_7_port, O_8_port, O_9_port, O_10_port, O_11_port, 
      O_12_port, O_13_port, O_14_port, O_15_port, O_16_port, O_17_port, 
      O_18_port, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, 
      n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, 
      n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, 
      n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, 
      n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, 
      n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, 
      n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, 
      n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, 
      n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, 
      n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, 
      n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, 
      n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, 
      n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, 
      n943, n944, n945, n946, n947, O_1_port : std_logic;

begin
   O <= ( O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, O_46_port, 
      O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, O_40_port, 
      O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, 
      O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, 
      O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, 
      O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, O_16_port, 
      O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, O_10_port, 
      O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, O_3_port, 
      O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(49), A_s(48), A_s(47), A_s(46), A_s(45), A_s(44), A_s(43), 
      A_s(42), A_s(41), A_s(40), A_s(39), A_s(38), A_s(37), A_s(36), A_s(35), 
      A_s(34), A_s(33), A_s(32), A_s(31), A_s(30), A_s(29), A_s(28), A_s(27), 
      A_s(26), A_s(25), A_s(24), A_s(23), A_s(22), A_s(21), A_s(20), A_s(19), 
      A_s(18), A_s(17), A_s(16), A_s(15), A_s(14), A_s(13), A_s(12), A_s(11), 
      A_s(10), A_s(9), A_s(8), A_s(7), A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), 
      A_s(1), A_s(0), X_Logic0_port, X_Logic0_port );
   A_nso <= ( A_ns(49), A_ns(48), A_ns(47), A_ns(46), A_ns(45), A_ns(44), 
      A_ns(43), A_ns(42), A_ns(41), A_ns(40), A_ns(39), A_ns(38), A_ns(37), 
      A_ns(36), A_ns(35), A_ns(34), A_ns(33), A_ns(32), A_ns(31), A_ns(30), 
      A_ns(29), A_ns(28), A_ns(27), A_ns(26), A_ns(25), A_ns(24), A_ns(23), 
      A_ns(22), A_ns(21), A_ns(20), A_ns(19), A_ns(18), A_ns(17), A_ns(16), 
      A_ns(15), A_ns(14), A_ns(13), A_ns(12), A_ns(11), A_ns(10), A_ns(9), 
      A_ns(8), A_ns(7), A_ns(6), A_ns(5), A_ns(4), A_ns(3), A_ns(2), A_ns(1), 
      A_ns(0), X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : AND3_X1 port map( A1 => B(18), A2 => n947, A3 => B(17), ZN => n789);
   U3 : INV_X2 port map( A => n789, ZN => n790);
   U4 : OR3_X4 port map( A1 => B(17), A2 => B(18), A3 => n947, ZN => n795);
   U5 : INV_X4 port map( A => n793, ZN => n799);
   U6 : INV_X2 port map( A => n791, ZN => n800);
   U7 : OAI22_X1 port map( A1 => n791, A2 => n792, B1 => n793, B2 => n794, ZN 
                           => O_1_port);
   U8 : OAI221_X1 port map( B1 => n795, B2 => n796, C1 => n790, C2 => n797, A 
                           => n798, ZN => O_9_port);
   U9 : AOI22_X1 port map( A1 => A_ns(8), A2 => n799, B1 => A_s(8), B2 => n800,
                           ZN => n798);
   U10 : INV_X1 port map( A => A_s(7), ZN => n797);
   U11 : INV_X1 port map( A => A_ns(7), ZN => n796);
   U12 : OAI221_X1 port map( B1 => n795, B2 => n801, C1 => n790, C2 => n802, A 
                           => n803, ZN => O_8_port);
   U13 : AOI22_X1 port map( A1 => A_ns(7), A2 => n799, B1 => A_s(7), B2 => n800
                           , ZN => n803);
   U14 : INV_X1 port map( A => A_s(6), ZN => n802);
   U15 : INV_X1 port map( A => A_ns(6), ZN => n801);
   U16 : OAI221_X1 port map( B1 => n795, B2 => n804, C1 => n790, C2 => n805, A 
                           => n806, ZN => O_7_port);
   U17 : AOI22_X1 port map( A1 => A_ns(6), A2 => n799, B1 => A_s(6), B2 => n800
                           , ZN => n806);
   U18 : INV_X1 port map( A => A_s(5), ZN => n805);
   U19 : INV_X1 port map( A => A_ns(5), ZN => n804);
   U20 : OAI221_X1 port map( B1 => n795, B2 => n807, C1 => n790, C2 => n808, A 
                           => n809, ZN => O_6_port);
   U21 : AOI22_X1 port map( A1 => A_ns(5), A2 => n799, B1 => A_s(5), B2 => n800
                           , ZN => n809);
   U22 : INV_X1 port map( A => A_s(4), ZN => n808);
   U23 : INV_X1 port map( A => A_ns(4), ZN => n807);
   U24 : OAI221_X1 port map( B1 => n795, B2 => n810, C1 => n790, C2 => n811, A 
                           => n812, ZN => O_5_port);
   U25 : AOI22_X1 port map( A1 => A_ns(4), A2 => n799, B1 => A_s(4), B2 => n800
                           , ZN => n812);
   U26 : INV_X1 port map( A => A_s(3), ZN => n811);
   U27 : INV_X1 port map( A => A_ns(3), ZN => n810);
   U28 : OAI221_X1 port map( B1 => n795, B2 => n813, C1 => n790, C2 => n814, A 
                           => n815, ZN => O_51_port);
   U29 : AOI22_X1 port map( A1 => A_ns(50), A2 => n799, B1 => A_s(50), B2 => 
                           n800, ZN => n815);
   U30 : INV_X1 port map( A => A_s(49), ZN => n814);
   U31 : INV_X1 port map( A => A_ns(49), ZN => n813);
   U32 : OAI221_X1 port map( B1 => n795, B2 => n816, C1 => n790, C2 => n817, A 
                           => n818, ZN => O_50_port);
   U33 : AOI22_X1 port map( A1 => A_ns(49), A2 => n799, B1 => A_s(49), B2 => 
                           n800, ZN => n818);
   U34 : INV_X1 port map( A => A_s(48), ZN => n817);
   U35 : INV_X1 port map( A => A_ns(48), ZN => n816);
   U36 : OAI221_X1 port map( B1 => n795, B2 => n819, C1 => n790, C2 => n820, A 
                           => n821, ZN => O_4_port);
   U37 : AOI22_X1 port map( A1 => A_ns(3), A2 => n799, B1 => A_s(3), B2 => n800
                           , ZN => n821);
   U38 : INV_X1 port map( A => A_s(2), ZN => n820);
   U39 : INV_X1 port map( A => A_ns(2), ZN => n819);
   U40 : OAI221_X1 port map( B1 => n795, B2 => n822, C1 => n790, C2 => n823, A 
                           => n824, ZN => O_49_port);
   U41 : AOI22_X1 port map( A1 => A_ns(48), A2 => n799, B1 => A_s(48), B2 => 
                           n800, ZN => n824);
   U42 : INV_X1 port map( A => A_s(47), ZN => n823);
   U43 : INV_X1 port map( A => A_ns(47), ZN => n822);
   U44 : OAI221_X1 port map( B1 => n795, B2 => n825, C1 => n790, C2 => n826, A 
                           => n827, ZN => O_48_port);
   U45 : AOI22_X1 port map( A1 => A_ns(47), A2 => n799, B1 => A_s(47), B2 => 
                           n800, ZN => n827);
   U46 : INV_X1 port map( A => A_s(46), ZN => n826);
   U47 : INV_X1 port map( A => A_ns(46), ZN => n825);
   U48 : OAI221_X1 port map( B1 => n795, B2 => n828, C1 => n790, C2 => n829, A 
                           => n830, ZN => O_47_port);
   U49 : AOI22_X1 port map( A1 => A_ns(46), A2 => n799, B1 => A_s(46), B2 => 
                           n800, ZN => n830);
   U50 : INV_X1 port map( A => A_s(45), ZN => n829);
   U51 : INV_X1 port map( A => A_ns(45), ZN => n828);
   U52 : OAI221_X1 port map( B1 => n795, B2 => n831, C1 => n790, C2 => n832, A 
                           => n833, ZN => O_46_port);
   U53 : AOI22_X1 port map( A1 => A_ns(45), A2 => n799, B1 => A_s(45), B2 => 
                           n800, ZN => n833);
   U54 : INV_X1 port map( A => A_s(44), ZN => n832);
   U55 : INV_X1 port map( A => A_ns(44), ZN => n831);
   U56 : OAI221_X1 port map( B1 => n795, B2 => n834, C1 => n790, C2 => n835, A 
                           => n836, ZN => O_45_port);
   U57 : AOI22_X1 port map( A1 => A_ns(44), A2 => n799, B1 => A_s(44), B2 => 
                           n800, ZN => n836);
   U58 : INV_X1 port map( A => A_s(43), ZN => n835);
   U59 : INV_X1 port map( A => A_ns(43), ZN => n834);
   U60 : OAI221_X1 port map( B1 => n795, B2 => n837, C1 => n790, C2 => n838, A 
                           => n839, ZN => O_44_port);
   U61 : AOI22_X1 port map( A1 => A_ns(43), A2 => n799, B1 => A_s(43), B2 => 
                           n800, ZN => n839);
   U62 : INV_X1 port map( A => A_s(42), ZN => n838);
   U63 : INV_X1 port map( A => A_ns(42), ZN => n837);
   U64 : OAI221_X1 port map( B1 => n795, B2 => n840, C1 => n790, C2 => n841, A 
                           => n842, ZN => O_43_port);
   U65 : AOI22_X1 port map( A1 => A_ns(42), A2 => n799, B1 => A_s(42), B2 => 
                           n800, ZN => n842);
   U66 : INV_X1 port map( A => A_s(41), ZN => n841);
   U67 : INV_X1 port map( A => A_ns(41), ZN => n840);
   U68 : OAI221_X1 port map( B1 => n795, B2 => n843, C1 => n790, C2 => n844, A 
                           => n845, ZN => O_42_port);
   U69 : AOI22_X1 port map( A1 => A_ns(41), A2 => n799, B1 => A_s(41), B2 => 
                           n800, ZN => n845);
   U70 : INV_X1 port map( A => A_s(40), ZN => n844);
   U71 : INV_X1 port map( A => A_ns(40), ZN => n843);
   U72 : OAI221_X1 port map( B1 => n795, B2 => n846, C1 => n790, C2 => n847, A 
                           => n848, ZN => O_41_port);
   U73 : AOI22_X1 port map( A1 => A_ns(40), A2 => n799, B1 => A_s(40), B2 => 
                           n800, ZN => n848);
   U74 : INV_X1 port map( A => A_s(39), ZN => n847);
   U75 : INV_X1 port map( A => A_ns(39), ZN => n846);
   U76 : OAI221_X1 port map( B1 => n795, B2 => n849, C1 => n790, C2 => n850, A 
                           => n851, ZN => O_40_port);
   U77 : AOI22_X1 port map( A1 => A_ns(39), A2 => n799, B1 => A_s(39), B2 => 
                           n800, ZN => n851);
   U78 : INV_X1 port map( A => A_s(38), ZN => n850);
   U79 : INV_X1 port map( A => A_ns(38), ZN => n849);
   U80 : OAI221_X1 port map( B1 => n795, B2 => n852, C1 => n790, C2 => n853, A 
                           => n854, ZN => O_3_port);
   U81 : AOI22_X1 port map( A1 => A_ns(2), A2 => n799, B1 => A_s(2), B2 => n800
                           , ZN => n854);
   U82 : INV_X1 port map( A => A_s(1), ZN => n853);
   U83 : INV_X1 port map( A => A_ns(1), ZN => n852);
   U84 : OAI221_X1 port map( B1 => n795, B2 => n855, C1 => n790, C2 => n856, A 
                           => n857, ZN => O_39_port);
   U85 : AOI22_X1 port map( A1 => A_ns(38), A2 => n799, B1 => A_s(38), B2 => 
                           n800, ZN => n857);
   U86 : INV_X1 port map( A => A_s(37), ZN => n856);
   U87 : INV_X1 port map( A => A_ns(37), ZN => n855);
   U88 : OAI221_X1 port map( B1 => n795, B2 => n858, C1 => n790, C2 => n859, A 
                           => n860, ZN => O_38_port);
   U89 : AOI22_X1 port map( A1 => A_ns(37), A2 => n799, B1 => A_s(37), B2 => 
                           n800, ZN => n860);
   U90 : INV_X1 port map( A => A_s(36), ZN => n859);
   U91 : INV_X1 port map( A => A_ns(36), ZN => n858);
   U92 : OAI221_X1 port map( B1 => n795, B2 => n861, C1 => n790, C2 => n862, A 
                           => n863, ZN => O_37_port);
   U93 : AOI22_X1 port map( A1 => A_ns(36), A2 => n799, B1 => A_s(36), B2 => 
                           n800, ZN => n863);
   U94 : INV_X1 port map( A => A_s(35), ZN => n862);
   U95 : INV_X1 port map( A => A_ns(35), ZN => n861);
   U96 : OAI221_X1 port map( B1 => n795, B2 => n864, C1 => n790, C2 => n865, A 
                           => n866, ZN => O_36_port);
   U97 : AOI22_X1 port map( A1 => A_ns(35), A2 => n799, B1 => A_s(35), B2 => 
                           n800, ZN => n866);
   U98 : INV_X1 port map( A => A_s(34), ZN => n865);
   U99 : INV_X1 port map( A => A_ns(34), ZN => n864);
   U100 : OAI221_X1 port map( B1 => n795, B2 => n867, C1 => n790, C2 => n868, A
                           => n869, ZN => O_35_port);
   U101 : AOI22_X1 port map( A1 => A_ns(34), A2 => n799, B1 => A_s(34), B2 => 
                           n800, ZN => n869);
   U102 : INV_X1 port map( A => A_s(33), ZN => n868);
   U103 : INV_X1 port map( A => A_ns(33), ZN => n867);
   U104 : OAI221_X1 port map( B1 => n795, B2 => n870, C1 => n790, C2 => n871, A
                           => n872, ZN => O_34_port);
   U105 : AOI22_X1 port map( A1 => A_ns(33), A2 => n799, B1 => A_s(33), B2 => 
                           n800, ZN => n872);
   U106 : INV_X1 port map( A => A_s(32), ZN => n871);
   U107 : INV_X1 port map( A => A_ns(32), ZN => n870);
   U108 : OAI221_X1 port map( B1 => n795, B2 => n873, C1 => n790, C2 => n874, A
                           => n875, ZN => O_33_port);
   U109 : AOI22_X1 port map( A1 => A_ns(32), A2 => n799, B1 => A_s(32), B2 => 
                           n800, ZN => n875);
   U110 : INV_X1 port map( A => A_s(31), ZN => n874);
   U111 : INV_X1 port map( A => A_ns(31), ZN => n873);
   U112 : OAI221_X1 port map( B1 => n795, B2 => n876, C1 => n790, C2 => n877, A
                           => n878, ZN => O_32_port);
   U113 : AOI22_X1 port map( A1 => A_ns(31), A2 => n799, B1 => A_s(31), B2 => 
                           n800, ZN => n878);
   U114 : INV_X1 port map( A => A_s(30), ZN => n877);
   U115 : INV_X1 port map( A => A_ns(30), ZN => n876);
   U116 : OAI221_X1 port map( B1 => n795, B2 => n879, C1 => n790, C2 => n880, A
                           => n881, ZN => O_31_port);
   U117 : AOI22_X1 port map( A1 => A_ns(30), A2 => n799, B1 => A_s(30), B2 => 
                           n800, ZN => n881);
   U118 : INV_X1 port map( A => A_s(29), ZN => n880);
   U119 : INV_X1 port map( A => A_ns(29), ZN => n879);
   U120 : OAI221_X1 port map( B1 => n795, B2 => n882, C1 => n790, C2 => n883, A
                           => n884, ZN => O_30_port);
   U121 : AOI22_X1 port map( A1 => A_ns(29), A2 => n799, B1 => A_s(29), B2 => 
                           n800, ZN => n884);
   U122 : INV_X1 port map( A => A_s(28), ZN => n883);
   U123 : INV_X1 port map( A => A_ns(28), ZN => n882);
   U124 : OAI221_X1 port map( B1 => n794, B2 => n795, C1 => n792, C2 => n790, A
                           => n885, ZN => O_2_port);
   U125 : AOI22_X1 port map( A1 => A_ns(1), A2 => n799, B1 => A_s(1), B2 => 
                           n800, ZN => n885);
   U126 : INV_X1 port map( A => A_s(0), ZN => n792);
   U127 : INV_X1 port map( A => A_ns(0), ZN => n794);
   U128 : OAI221_X1 port map( B1 => n795, B2 => n886, C1 => n790, C2 => n887, A
                           => n888, ZN => O_29_port);
   U129 : AOI22_X1 port map( A1 => A_ns(28), A2 => n799, B1 => A_s(28), B2 => 
                           n800, ZN => n888);
   U130 : INV_X1 port map( A => A_s(27), ZN => n887);
   U131 : INV_X1 port map( A => A_ns(27), ZN => n886);
   U132 : OAI221_X1 port map( B1 => n795, B2 => n889, C1 => n790, C2 => n890, A
                           => n891, ZN => O_28_port);
   U133 : AOI22_X1 port map( A1 => A_ns(27), A2 => n799, B1 => A_s(27), B2 => 
                           n800, ZN => n891);
   U134 : INV_X1 port map( A => A_s(26), ZN => n890);
   U135 : INV_X1 port map( A => A_ns(26), ZN => n889);
   U136 : OAI221_X1 port map( B1 => n795, B2 => n892, C1 => n790, C2 => n893, A
                           => n894, ZN => O_27_port);
   U137 : AOI22_X1 port map( A1 => A_ns(26), A2 => n799, B1 => A_s(26), B2 => 
                           n800, ZN => n894);
   U138 : INV_X1 port map( A => A_s(25), ZN => n893);
   U139 : INV_X1 port map( A => A_ns(25), ZN => n892);
   U140 : OAI221_X1 port map( B1 => n795, B2 => n895, C1 => n790, C2 => n896, A
                           => n897, ZN => O_26_port);
   U141 : AOI22_X1 port map( A1 => A_ns(25), A2 => n799, B1 => A_s(25), B2 => 
                           n800, ZN => n897);
   U142 : INV_X1 port map( A => A_s(24), ZN => n896);
   U143 : INV_X1 port map( A => A_ns(24), ZN => n895);
   U144 : OAI221_X1 port map( B1 => n795, B2 => n898, C1 => n790, C2 => n899, A
                           => n900, ZN => O_25_port);
   U145 : AOI22_X1 port map( A1 => A_ns(24), A2 => n799, B1 => A_s(24), B2 => 
                           n800, ZN => n900);
   U146 : INV_X1 port map( A => A_s(23), ZN => n899);
   U147 : INV_X1 port map( A => A_ns(23), ZN => n898);
   U148 : OAI221_X1 port map( B1 => n795, B2 => n901, C1 => n790, C2 => n902, A
                           => n903, ZN => O_24_port);
   U149 : AOI22_X1 port map( A1 => A_ns(23), A2 => n799, B1 => A_s(23), B2 => 
                           n800, ZN => n903);
   U150 : INV_X1 port map( A => A_s(22), ZN => n902);
   U151 : INV_X1 port map( A => A_ns(22), ZN => n901);
   U152 : OAI221_X1 port map( B1 => n795, B2 => n904, C1 => n790, C2 => n905, A
                           => n906, ZN => O_23_port);
   U153 : AOI22_X1 port map( A1 => A_ns(22), A2 => n799, B1 => A_s(22), B2 => 
                           n800, ZN => n906);
   U154 : INV_X1 port map( A => A_s(21), ZN => n905);
   U155 : INV_X1 port map( A => A_ns(21), ZN => n904);
   U156 : OAI221_X1 port map( B1 => n795, B2 => n907, C1 => n790, C2 => n908, A
                           => n909, ZN => O_22_port);
   U157 : AOI22_X1 port map( A1 => A_ns(21), A2 => n799, B1 => A_s(21), B2 => 
                           n800, ZN => n909);
   U158 : INV_X1 port map( A => A_s(20), ZN => n908);
   U159 : INV_X1 port map( A => A_ns(20), ZN => n907);
   U160 : OAI221_X1 port map( B1 => n795, B2 => n910, C1 => n790, C2 => n911, A
                           => n912, ZN => O_21_port);
   U161 : AOI22_X1 port map( A1 => A_ns(20), A2 => n799, B1 => A_s(20), B2 => 
                           n800, ZN => n912);
   U162 : INV_X1 port map( A => A_s(19), ZN => n911);
   U163 : INV_X1 port map( A => A_ns(19), ZN => n910);
   U164 : OAI221_X1 port map( B1 => n795, B2 => n913, C1 => n790, C2 => n914, A
                           => n915, ZN => O_20_port);
   U165 : AOI22_X1 port map( A1 => A_ns(19), A2 => n799, B1 => A_s(19), B2 => 
                           n800, ZN => n915);
   U166 : INV_X1 port map( A => A_s(18), ZN => n914);
   U167 : INV_X1 port map( A => A_ns(18), ZN => n913);
   U168 : OAI221_X1 port map( B1 => n795, B2 => n916, C1 => n790, C2 => n917, A
                           => n918, ZN => O_19_port);
   U169 : AOI22_X1 port map( A1 => A_ns(18), A2 => n799, B1 => A_s(18), B2 => 
                           n800, ZN => n918);
   U170 : INV_X1 port map( A => A_s(17), ZN => n917);
   U171 : INV_X1 port map( A => A_ns(17), ZN => n916);
   U172 : OAI221_X1 port map( B1 => n795, B2 => n919, C1 => n790, C2 => n920, A
                           => n921, ZN => O_18_port);
   U173 : AOI22_X1 port map( A1 => A_ns(17), A2 => n799, B1 => A_s(17), B2 => 
                           n800, ZN => n921);
   U174 : INV_X1 port map( A => A_s(16), ZN => n920);
   U175 : INV_X1 port map( A => A_ns(16), ZN => n919);
   U176 : OAI221_X1 port map( B1 => n795, B2 => n922, C1 => n790, C2 => n923, A
                           => n924, ZN => O_17_port);
   U177 : AOI22_X1 port map( A1 => A_ns(16), A2 => n799, B1 => A_s(16), B2 => 
                           n800, ZN => n924);
   U178 : INV_X1 port map( A => A_s(15), ZN => n923);
   U179 : INV_X1 port map( A => A_ns(15), ZN => n922);
   U180 : OAI221_X1 port map( B1 => n795, B2 => n925, C1 => n790, C2 => n926, A
                           => n927, ZN => O_16_port);
   U181 : AOI22_X1 port map( A1 => A_ns(15), A2 => n799, B1 => A_s(15), B2 => 
                           n800, ZN => n927);
   U182 : INV_X1 port map( A => A_s(14), ZN => n926);
   U183 : INV_X1 port map( A => A_ns(14), ZN => n925);
   U184 : OAI221_X1 port map( B1 => n795, B2 => n928, C1 => n790, C2 => n929, A
                           => n930, ZN => O_15_port);
   U185 : AOI22_X1 port map( A1 => A_ns(14), A2 => n799, B1 => A_s(14), B2 => 
                           n800, ZN => n930);
   U186 : INV_X1 port map( A => A_s(13), ZN => n929);
   U187 : INV_X1 port map( A => A_ns(13), ZN => n928);
   U188 : OAI221_X1 port map( B1 => n795, B2 => n931, C1 => n790, C2 => n932, A
                           => n933, ZN => O_14_port);
   U189 : AOI22_X1 port map( A1 => A_ns(13), A2 => n799, B1 => A_s(13), B2 => 
                           n800, ZN => n933);
   U190 : INV_X1 port map( A => A_s(12), ZN => n932);
   U191 : INV_X1 port map( A => A_ns(12), ZN => n931);
   U192 : OAI221_X1 port map( B1 => n795, B2 => n934, C1 => n790, C2 => n935, A
                           => n936, ZN => O_13_port);
   U193 : AOI22_X1 port map( A1 => A_ns(12), A2 => n799, B1 => A_s(12), B2 => 
                           n800, ZN => n936);
   U194 : INV_X1 port map( A => A_s(11), ZN => n935);
   U195 : INV_X1 port map( A => A_ns(11), ZN => n934);
   U196 : OAI221_X1 port map( B1 => n795, B2 => n937, C1 => n790, C2 => n938, A
                           => n939, ZN => O_12_port);
   U197 : AOI22_X1 port map( A1 => A_ns(11), A2 => n799, B1 => A_s(11), B2 => 
                           n800, ZN => n939);
   U198 : INV_X1 port map( A => A_s(10), ZN => n938);
   U199 : INV_X1 port map( A => A_ns(10), ZN => n937);
   U200 : OAI221_X1 port map( B1 => n795, B2 => n940, C1 => n790, C2 => n941, A
                           => n942, ZN => O_11_port);
   U201 : AOI22_X1 port map( A1 => A_ns(10), A2 => n799, B1 => A_s(10), B2 => 
                           n800, ZN => n942);
   U202 : INV_X1 port map( A => A_s(9), ZN => n941);
   U203 : INV_X1 port map( A => A_ns(9), ZN => n940);
   U204 : OAI221_X1 port map( B1 => n943, B2 => n795, C1 => n944, C2 => n790, A
                           => n945, ZN => O_10_port);
   U205 : AOI22_X1 port map( A1 => A_ns(9), A2 => n799, B1 => A_s(9), B2 => 
                           n800, ZN => n945);
   U206 : NAND2_X1 port map( A1 => n946, A2 => n791, ZN => n793);
   U207 : NAND2_X1 port map( A1 => n946, A2 => n947, ZN => n791);
   U208 : XOR2_X1 port map( A => B(17), B => B(18), Z => n946);
   U209 : INV_X1 port map( A => A_s(8), ZN => n944);
   U210 : INV_X1 port map( A => B(19), ZN => n947);
   U211 : INV_X1 port map( A => A_ns(8), ZN => n943);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT50_i16 is

   port( A_s, A_ns, B : in std_logic_vector (49 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (49 downto 0));

end BOOTHENC_NBIT50_i16;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT50_i16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, O_47_port, O_48_port, O_49_port, O_46_port, O_45_port,
      O_44_port, O_43_port, O_42_port, O_41_port, O_40_port, O_39_port, 
      O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, O_33_port, 
      O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, O_27_port, 
      O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, O_21_port, 
      O_20_port, O_19_port, O_18_port, O_17_port, O_2_port, O_3_port, O_4_port,
      O_5_port, O_6_port, O_7_port, O_8_port, O_9_port, O_10_port, O_11_port, 
      O_12_port, O_13_port, O_14_port, O_15_port, O_16_port, n805, n806, n807, 
      n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, 
      n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, 
      n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, 
      n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, 
      n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, 
      n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, 
      n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, 
      n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, 
      n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, 
      n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, 
      n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, 
      n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, 
      n952, n953, n954, n955, n956, O_1_port : std_logic;

begin
   O <= ( O_49_port, O_48_port, O_47_port, O_46_port, O_45_port, O_44_port, 
      O_43_port, O_42_port, O_41_port, O_40_port, O_39_port, O_38_port, 
      O_37_port, O_36_port, O_35_port, O_34_port, O_33_port, O_32_port, 
      O_31_port, O_30_port, O_29_port, O_28_port, O_27_port, O_26_port, 
      O_25_port, O_24_port, O_23_port, O_22_port, O_21_port, O_20_port, 
      O_19_port, O_18_port, O_17_port, O_16_port, O_15_port, O_14_port, 
      O_13_port, O_12_port, O_11_port, O_10_port, O_9_port, O_8_port, O_7_port,
      O_6_port, O_5_port, O_4_port, O_3_port, O_2_port, O_1_port, X_Logic0_port
      );
   A_so <= ( A_s(47), A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), 
      A_s(40), A_s(39), A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), 
      A_s(32), A_s(31), A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), 
      A_s(24), A_s(23), A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), 
      A_s(16), A_s(15), A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), 
      A_s(8), A_s(7), A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), 
      X_Logic0_port, X_Logic0_port );
   A_nso <= ( A_ns(47), A_ns(46), A_ns(45), A_ns(44), A_ns(43), A_ns(42), 
      A_ns(41), A_ns(40), A_ns(39), A_ns(38), A_ns(37), A_ns(36), A_ns(35), 
      A_ns(34), A_ns(33), A_ns(32), A_ns(31), A_ns(30), A_ns(29), A_ns(28), 
      A_ns(27), A_ns(26), A_ns(25), A_ns(24), A_ns(23), A_ns(22), A_ns(21), 
      A_ns(20), A_ns(19), A_ns(18), A_ns(17), A_ns(16), A_ns(15), A_ns(14), 
      A_ns(13), A_ns(12), A_ns(11), A_ns(10), A_ns(9), A_ns(8), A_ns(7), 
      A_ns(6), A_ns(5), A_ns(4), A_ns(3), A_ns(2), A_ns(1), A_ns(0), 
      X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : NAND3_X2 port map( A1 => B(16), A2 => n956, A3 => B(15), ZN => n811);
   U3 : INV_X2 port map( A => n805, ZN => n815);
   U4 : OR3_X2 port map( A1 => B(15), A2 => B(16), A3 => n956, ZN => n809);
   U5 : INV_X2 port map( A => n807, ZN => n814);
   U6 : OAI22_X1 port map( A1 => n805, A2 => n806, B1 => n807, B2 => n808, ZN 
                           => O_1_port);
   U7 : OAI221_X1 port map( B1 => n809, B2 => n810, C1 => n811, C2 => n812, A 
                           => n813, ZN => O_9_port);
   U8 : AOI22_X1 port map( A1 => A_ns(8), A2 => n814, B1 => A_s(8), B2 => n815,
                           ZN => n813);
   U9 : INV_X1 port map( A => A_s(7), ZN => n812);
   U10 : INV_X1 port map( A => A_ns(7), ZN => n810);
   U11 : OAI221_X1 port map( B1 => n809, B2 => n816, C1 => n811, C2 => n817, A 
                           => n818, ZN => O_8_port);
   U12 : AOI22_X1 port map( A1 => A_ns(7), A2 => n814, B1 => A_s(7), B2 => n815
                           , ZN => n818);
   U13 : INV_X1 port map( A => A_s(6), ZN => n817);
   U14 : INV_X1 port map( A => A_ns(6), ZN => n816);
   U15 : OAI221_X1 port map( B1 => n809, B2 => n819, C1 => n811, C2 => n820, A 
                           => n821, ZN => O_7_port);
   U16 : AOI22_X1 port map( A1 => A_ns(6), A2 => n814, B1 => A_s(6), B2 => n815
                           , ZN => n821);
   U17 : INV_X1 port map( A => A_s(5), ZN => n820);
   U18 : INV_X1 port map( A => A_ns(5), ZN => n819);
   U19 : OAI221_X1 port map( B1 => n809, B2 => n822, C1 => n811, C2 => n823, A 
                           => n824, ZN => O_6_port);
   U20 : AOI22_X1 port map( A1 => A_ns(5), A2 => n814, B1 => A_s(5), B2 => n815
                           , ZN => n824);
   U21 : INV_X1 port map( A => A_s(4), ZN => n823);
   U22 : INV_X1 port map( A => A_ns(4), ZN => n822);
   U23 : OAI221_X1 port map( B1 => n809, B2 => n825, C1 => n811, C2 => n826, A 
                           => n827, ZN => O_5_port);
   U24 : AOI22_X1 port map( A1 => A_ns(4), A2 => n814, B1 => A_s(4), B2 => n815
                           , ZN => n827);
   U25 : INV_X1 port map( A => A_s(3), ZN => n826);
   U26 : INV_X1 port map( A => A_ns(3), ZN => n825);
   U27 : OAI221_X1 port map( B1 => n809, B2 => n828, C1 => n811, C2 => n829, A 
                           => n830, ZN => O_4_port);
   U28 : AOI22_X1 port map( A1 => A_ns(3), A2 => n814, B1 => A_s(3), B2 => n815
                           , ZN => n830);
   U29 : INV_X1 port map( A => A_s(2), ZN => n829);
   U30 : INV_X1 port map( A => A_ns(2), ZN => n828);
   U31 : OAI221_X1 port map( B1 => n809, B2 => n831, C1 => n811, C2 => n832, A 
                           => n833, ZN => O_49_port);
   U32 : AOI22_X1 port map( A1 => A_ns(48), A2 => n814, B1 => A_s(48), B2 => 
                           n815, ZN => n833);
   U33 : INV_X1 port map( A => A_s(47), ZN => n832);
   U34 : INV_X1 port map( A => A_ns(47), ZN => n831);
   U35 : OAI221_X1 port map( B1 => n809, B2 => n834, C1 => n811, C2 => n835, A 
                           => n836, ZN => O_48_port);
   U36 : AOI22_X1 port map( A1 => A_ns(47), A2 => n814, B1 => A_s(47), B2 => 
                           n815, ZN => n836);
   U37 : INV_X1 port map( A => A_s(46), ZN => n835);
   U38 : INV_X1 port map( A => A_ns(46), ZN => n834);
   U39 : OAI221_X1 port map( B1 => n809, B2 => n837, C1 => n811, C2 => n838, A 
                           => n839, ZN => O_47_port);
   U40 : AOI22_X1 port map( A1 => A_ns(46), A2 => n814, B1 => A_s(46), B2 => 
                           n815, ZN => n839);
   U41 : INV_X1 port map( A => A_s(45), ZN => n838);
   U42 : INV_X1 port map( A => A_ns(45), ZN => n837);
   U43 : OAI221_X1 port map( B1 => n809, B2 => n840, C1 => n811, C2 => n841, A 
                           => n842, ZN => O_46_port);
   U44 : AOI22_X1 port map( A1 => A_ns(45), A2 => n814, B1 => A_s(45), B2 => 
                           n815, ZN => n842);
   U45 : INV_X1 port map( A => A_s(44), ZN => n841);
   U46 : INV_X1 port map( A => A_ns(44), ZN => n840);
   U47 : OAI221_X1 port map( B1 => n809, B2 => n843, C1 => n811, C2 => n844, A 
                           => n845, ZN => O_45_port);
   U48 : AOI22_X1 port map( A1 => A_ns(44), A2 => n814, B1 => A_s(44), B2 => 
                           n815, ZN => n845);
   U49 : INV_X1 port map( A => A_s(43), ZN => n844);
   U50 : INV_X1 port map( A => A_ns(43), ZN => n843);
   U51 : OAI221_X1 port map( B1 => n809, B2 => n846, C1 => n811, C2 => n847, A 
                           => n848, ZN => O_44_port);
   U52 : AOI22_X1 port map( A1 => A_ns(43), A2 => n814, B1 => A_s(43), B2 => 
                           n815, ZN => n848);
   U53 : INV_X1 port map( A => A_s(42), ZN => n847);
   U54 : INV_X1 port map( A => A_ns(42), ZN => n846);
   U55 : OAI221_X1 port map( B1 => n809, B2 => n849, C1 => n811, C2 => n850, A 
                           => n851, ZN => O_43_port);
   U56 : AOI22_X1 port map( A1 => A_ns(42), A2 => n814, B1 => A_s(42), B2 => 
                           n815, ZN => n851);
   U57 : INV_X1 port map( A => A_s(41), ZN => n850);
   U58 : INV_X1 port map( A => A_ns(41), ZN => n849);
   U59 : OAI221_X1 port map( B1 => n809, B2 => n852, C1 => n811, C2 => n853, A 
                           => n854, ZN => O_42_port);
   U60 : AOI22_X1 port map( A1 => A_ns(41), A2 => n814, B1 => A_s(41), B2 => 
                           n815, ZN => n854);
   U61 : INV_X1 port map( A => A_s(40), ZN => n853);
   U62 : INV_X1 port map( A => A_ns(40), ZN => n852);
   U63 : OAI221_X1 port map( B1 => n809, B2 => n855, C1 => n811, C2 => n856, A 
                           => n857, ZN => O_41_port);
   U64 : AOI22_X1 port map( A1 => A_ns(40), A2 => n814, B1 => A_s(40), B2 => 
                           n815, ZN => n857);
   U65 : INV_X1 port map( A => A_s(39), ZN => n856);
   U66 : INV_X1 port map( A => A_ns(39), ZN => n855);
   U67 : OAI221_X1 port map( B1 => n809, B2 => n858, C1 => n811, C2 => n859, A 
                           => n860, ZN => O_40_port);
   U68 : AOI22_X1 port map( A1 => A_ns(39), A2 => n814, B1 => A_s(39), B2 => 
                           n815, ZN => n860);
   U69 : INV_X1 port map( A => A_s(38), ZN => n859);
   U70 : INV_X1 port map( A => A_ns(38), ZN => n858);
   U71 : OAI221_X1 port map( B1 => n809, B2 => n861, C1 => n811, C2 => n862, A 
                           => n863, ZN => O_3_port);
   U72 : AOI22_X1 port map( A1 => A_ns(2), A2 => n814, B1 => A_s(2), B2 => n815
                           , ZN => n863);
   U73 : INV_X1 port map( A => A_s(1), ZN => n862);
   U74 : INV_X1 port map( A => A_ns(1), ZN => n861);
   U75 : OAI221_X1 port map( B1 => n809, B2 => n864, C1 => n811, C2 => n865, A 
                           => n866, ZN => O_39_port);
   U76 : AOI22_X1 port map( A1 => A_ns(38), A2 => n814, B1 => A_s(38), B2 => 
                           n815, ZN => n866);
   U77 : INV_X1 port map( A => A_s(37), ZN => n865);
   U78 : INV_X1 port map( A => A_ns(37), ZN => n864);
   U79 : OAI221_X1 port map( B1 => n809, B2 => n867, C1 => n811, C2 => n868, A 
                           => n869, ZN => O_38_port);
   U80 : AOI22_X1 port map( A1 => A_ns(37), A2 => n814, B1 => A_s(37), B2 => 
                           n815, ZN => n869);
   U81 : INV_X1 port map( A => A_s(36), ZN => n868);
   U82 : INV_X1 port map( A => A_ns(36), ZN => n867);
   U83 : OAI221_X1 port map( B1 => n809, B2 => n870, C1 => n811, C2 => n871, A 
                           => n872, ZN => O_37_port);
   U84 : AOI22_X1 port map( A1 => A_ns(36), A2 => n814, B1 => A_s(36), B2 => 
                           n815, ZN => n872);
   U85 : INV_X1 port map( A => A_s(35), ZN => n871);
   U86 : INV_X1 port map( A => A_ns(35), ZN => n870);
   U87 : OAI221_X1 port map( B1 => n809, B2 => n873, C1 => n811, C2 => n874, A 
                           => n875, ZN => O_36_port);
   U88 : AOI22_X1 port map( A1 => A_ns(35), A2 => n814, B1 => A_s(35), B2 => 
                           n815, ZN => n875);
   U89 : INV_X1 port map( A => A_s(34), ZN => n874);
   U90 : INV_X1 port map( A => A_ns(34), ZN => n873);
   U91 : OAI221_X1 port map( B1 => n809, B2 => n876, C1 => n811, C2 => n877, A 
                           => n878, ZN => O_35_port);
   U92 : AOI22_X1 port map( A1 => A_ns(34), A2 => n814, B1 => A_s(34), B2 => 
                           n815, ZN => n878);
   U93 : INV_X1 port map( A => A_s(33), ZN => n877);
   U94 : INV_X1 port map( A => A_ns(33), ZN => n876);
   U95 : OAI221_X1 port map( B1 => n809, B2 => n879, C1 => n811, C2 => n880, A 
                           => n881, ZN => O_34_port);
   U96 : AOI22_X1 port map( A1 => A_ns(33), A2 => n814, B1 => A_s(33), B2 => 
                           n815, ZN => n881);
   U97 : INV_X1 port map( A => A_s(32), ZN => n880);
   U98 : INV_X1 port map( A => A_ns(32), ZN => n879);
   U99 : OAI221_X1 port map( B1 => n809, B2 => n882, C1 => n811, C2 => n883, A 
                           => n884, ZN => O_33_port);
   U100 : AOI22_X1 port map( A1 => A_ns(32), A2 => n814, B1 => A_s(32), B2 => 
                           n815, ZN => n884);
   U101 : INV_X1 port map( A => A_s(31), ZN => n883);
   U102 : INV_X1 port map( A => A_ns(31), ZN => n882);
   U103 : OAI221_X1 port map( B1 => n809, B2 => n885, C1 => n811, C2 => n886, A
                           => n887, ZN => O_32_port);
   U104 : AOI22_X1 port map( A1 => A_ns(31), A2 => n814, B1 => A_s(31), B2 => 
                           n815, ZN => n887);
   U105 : INV_X1 port map( A => A_s(30), ZN => n886);
   U106 : INV_X1 port map( A => A_ns(30), ZN => n885);
   U107 : OAI221_X1 port map( B1 => n809, B2 => n888, C1 => n811, C2 => n889, A
                           => n890, ZN => O_31_port);
   U108 : AOI22_X1 port map( A1 => A_ns(30), A2 => n814, B1 => A_s(30), B2 => 
                           n815, ZN => n890);
   U109 : INV_X1 port map( A => A_s(29), ZN => n889);
   U110 : INV_X1 port map( A => A_ns(29), ZN => n888);
   U111 : OAI221_X1 port map( B1 => n809, B2 => n891, C1 => n811, C2 => n892, A
                           => n893, ZN => O_30_port);
   U112 : AOI22_X1 port map( A1 => A_ns(29), A2 => n814, B1 => A_s(29), B2 => 
                           n815, ZN => n893);
   U113 : INV_X1 port map( A => A_s(28), ZN => n892);
   U114 : INV_X1 port map( A => A_ns(28), ZN => n891);
   U115 : OAI221_X1 port map( B1 => n808, B2 => n809, C1 => n806, C2 => n811, A
                           => n894, ZN => O_2_port);
   U116 : AOI22_X1 port map( A1 => A_ns(1), A2 => n814, B1 => A_s(1), B2 => 
                           n815, ZN => n894);
   U117 : INV_X1 port map( A => A_s(0), ZN => n806);
   U118 : INV_X1 port map( A => A_ns(0), ZN => n808);
   U119 : OAI221_X1 port map( B1 => n809, B2 => n895, C1 => n811, C2 => n896, A
                           => n897, ZN => O_29_port);
   U120 : AOI22_X1 port map( A1 => A_ns(28), A2 => n814, B1 => A_s(28), B2 => 
                           n815, ZN => n897);
   U121 : INV_X1 port map( A => A_s(27), ZN => n896);
   U122 : INV_X1 port map( A => A_ns(27), ZN => n895);
   U123 : OAI221_X1 port map( B1 => n809, B2 => n898, C1 => n811, C2 => n899, A
                           => n900, ZN => O_28_port);
   U124 : AOI22_X1 port map( A1 => A_ns(27), A2 => n814, B1 => A_s(27), B2 => 
                           n815, ZN => n900);
   U125 : INV_X1 port map( A => A_s(26), ZN => n899);
   U126 : INV_X1 port map( A => A_ns(26), ZN => n898);
   U127 : OAI221_X1 port map( B1 => n809, B2 => n901, C1 => n811, C2 => n902, A
                           => n903, ZN => O_27_port);
   U128 : AOI22_X1 port map( A1 => A_ns(26), A2 => n814, B1 => A_s(26), B2 => 
                           n815, ZN => n903);
   U129 : INV_X1 port map( A => A_s(25), ZN => n902);
   U130 : INV_X1 port map( A => A_ns(25), ZN => n901);
   U131 : OAI221_X1 port map( B1 => n809, B2 => n904, C1 => n811, C2 => n905, A
                           => n906, ZN => O_26_port);
   U132 : AOI22_X1 port map( A1 => A_ns(25), A2 => n814, B1 => A_s(25), B2 => 
                           n815, ZN => n906);
   U133 : INV_X1 port map( A => A_s(24), ZN => n905);
   U134 : INV_X1 port map( A => A_ns(24), ZN => n904);
   U135 : OAI221_X1 port map( B1 => n809, B2 => n907, C1 => n811, C2 => n908, A
                           => n909, ZN => O_25_port);
   U136 : AOI22_X1 port map( A1 => A_ns(24), A2 => n814, B1 => A_s(24), B2 => 
                           n815, ZN => n909);
   U137 : INV_X1 port map( A => A_s(23), ZN => n908);
   U138 : INV_X1 port map( A => A_ns(23), ZN => n907);
   U139 : OAI221_X1 port map( B1 => n809, B2 => n910, C1 => n811, C2 => n911, A
                           => n912, ZN => O_24_port);
   U140 : AOI22_X1 port map( A1 => A_ns(23), A2 => n814, B1 => A_s(23), B2 => 
                           n815, ZN => n912);
   U141 : INV_X1 port map( A => A_s(22), ZN => n911);
   U142 : INV_X1 port map( A => A_ns(22), ZN => n910);
   U143 : OAI221_X1 port map( B1 => n809, B2 => n913, C1 => n811, C2 => n914, A
                           => n915, ZN => O_23_port);
   U144 : AOI22_X1 port map( A1 => A_ns(22), A2 => n814, B1 => A_s(22), B2 => 
                           n815, ZN => n915);
   U145 : INV_X1 port map( A => A_s(21), ZN => n914);
   U146 : INV_X1 port map( A => A_ns(21), ZN => n913);
   U147 : OAI221_X1 port map( B1 => n809, B2 => n916, C1 => n811, C2 => n917, A
                           => n918, ZN => O_22_port);
   U148 : AOI22_X1 port map( A1 => A_ns(21), A2 => n814, B1 => A_s(21), B2 => 
                           n815, ZN => n918);
   U149 : INV_X1 port map( A => A_s(20), ZN => n917);
   U150 : INV_X1 port map( A => A_ns(20), ZN => n916);
   U151 : OAI221_X1 port map( B1 => n809, B2 => n919, C1 => n811, C2 => n920, A
                           => n921, ZN => O_21_port);
   U152 : AOI22_X1 port map( A1 => A_ns(20), A2 => n814, B1 => A_s(20), B2 => 
                           n815, ZN => n921);
   U153 : INV_X1 port map( A => A_s(19), ZN => n920);
   U154 : INV_X1 port map( A => A_ns(19), ZN => n919);
   U155 : OAI221_X1 port map( B1 => n809, B2 => n922, C1 => n811, C2 => n923, A
                           => n924, ZN => O_20_port);
   U156 : AOI22_X1 port map( A1 => A_ns(19), A2 => n814, B1 => A_s(19), B2 => 
                           n815, ZN => n924);
   U157 : INV_X1 port map( A => A_s(18), ZN => n923);
   U158 : INV_X1 port map( A => A_ns(18), ZN => n922);
   U159 : OAI221_X1 port map( B1 => n809, B2 => n925, C1 => n811, C2 => n926, A
                           => n927, ZN => O_19_port);
   U160 : AOI22_X1 port map( A1 => A_ns(18), A2 => n814, B1 => A_s(18), B2 => 
                           n815, ZN => n927);
   U161 : INV_X1 port map( A => A_s(17), ZN => n926);
   U162 : INV_X1 port map( A => A_ns(17), ZN => n925);
   U163 : OAI221_X1 port map( B1 => n809, B2 => n928, C1 => n811, C2 => n929, A
                           => n930, ZN => O_18_port);
   U164 : AOI22_X1 port map( A1 => A_ns(17), A2 => n814, B1 => A_s(17), B2 => 
                           n815, ZN => n930);
   U165 : INV_X1 port map( A => A_s(16), ZN => n929);
   U166 : INV_X1 port map( A => A_ns(16), ZN => n928);
   U167 : OAI221_X1 port map( B1 => n809, B2 => n931, C1 => n811, C2 => n932, A
                           => n933, ZN => O_17_port);
   U168 : AOI22_X1 port map( A1 => A_ns(16), A2 => n814, B1 => A_s(16), B2 => 
                           n815, ZN => n933);
   U169 : INV_X1 port map( A => A_s(15), ZN => n932);
   U170 : INV_X1 port map( A => A_ns(15), ZN => n931);
   U171 : OAI221_X1 port map( B1 => n809, B2 => n934, C1 => n811, C2 => n935, A
                           => n936, ZN => O_16_port);
   U172 : AOI22_X1 port map( A1 => A_ns(15), A2 => n814, B1 => A_s(15), B2 => 
                           n815, ZN => n936);
   U173 : INV_X1 port map( A => A_s(14), ZN => n935);
   U174 : INV_X1 port map( A => A_ns(14), ZN => n934);
   U175 : OAI221_X1 port map( B1 => n809, B2 => n937, C1 => n811, C2 => n938, A
                           => n939, ZN => O_15_port);
   U176 : AOI22_X1 port map( A1 => A_ns(14), A2 => n814, B1 => A_s(14), B2 => 
                           n815, ZN => n939);
   U177 : INV_X1 port map( A => A_s(13), ZN => n938);
   U178 : INV_X1 port map( A => A_ns(13), ZN => n937);
   U179 : OAI221_X1 port map( B1 => n809, B2 => n940, C1 => n811, C2 => n941, A
                           => n942, ZN => O_14_port);
   U180 : AOI22_X1 port map( A1 => A_ns(13), A2 => n814, B1 => A_s(13), B2 => 
                           n815, ZN => n942);
   U181 : INV_X1 port map( A => A_s(12), ZN => n941);
   U182 : INV_X1 port map( A => A_ns(12), ZN => n940);
   U183 : OAI221_X1 port map( B1 => n809, B2 => n943, C1 => n811, C2 => n944, A
                           => n945, ZN => O_13_port);
   U184 : AOI22_X1 port map( A1 => A_ns(12), A2 => n814, B1 => A_s(12), B2 => 
                           n815, ZN => n945);
   U185 : INV_X1 port map( A => A_s(11), ZN => n944);
   U186 : INV_X1 port map( A => A_ns(11), ZN => n943);
   U187 : OAI221_X1 port map( B1 => n809, B2 => n946, C1 => n811, C2 => n947, A
                           => n948, ZN => O_12_port);
   U188 : AOI22_X1 port map( A1 => A_ns(11), A2 => n814, B1 => A_s(11), B2 => 
                           n815, ZN => n948);
   U189 : INV_X1 port map( A => A_s(10), ZN => n947);
   U190 : INV_X1 port map( A => A_ns(10), ZN => n946);
   U191 : OAI221_X1 port map( B1 => n809, B2 => n949, C1 => n811, C2 => n950, A
                           => n951, ZN => O_11_port);
   U192 : AOI22_X1 port map( A1 => A_ns(10), A2 => n814, B1 => A_s(10), B2 => 
                           n815, ZN => n951);
   U193 : INV_X1 port map( A => A_s(9), ZN => n950);
   U194 : INV_X1 port map( A => A_ns(9), ZN => n949);
   U195 : OAI221_X1 port map( B1 => n952, B2 => n809, C1 => n953, C2 => n811, A
                           => n954, ZN => O_10_port);
   U196 : AOI22_X1 port map( A1 => A_ns(9), A2 => n814, B1 => A_s(9), B2 => 
                           n815, ZN => n954);
   U197 : NAND2_X1 port map( A1 => n955, A2 => n805, ZN => n807);
   U198 : NAND2_X1 port map( A1 => n955, A2 => n956, ZN => n805);
   U199 : XOR2_X1 port map( A => B(15), B => B(16), Z => n955);
   U200 : INV_X1 port map( A => A_s(8), ZN => n953);
   U201 : INV_X1 port map( A => B(17), ZN => n956);
   U202 : INV_X1 port map( A => A_ns(8), ZN => n952);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT48_i14 is

   port( A_s, A_ns, B : in std_logic_vector (47 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (47 downto 0));

end BOOTHENC_NBIT48_i14;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT48_i14 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, n813, n814, n815, n816, n817, n818, n819, n820, n821, 
      n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, 
      n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, 
      n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, 
      n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, 
      n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, 
      n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, 
      n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, 
      n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, 
      n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, 
      n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, 
      n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, O_45_port, 
      O_46_port, O_47_port, O_44_port, O_43_port, O_42_port, O_41_port, 
      O_40_port, O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, 
      O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, 
      O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, 
      O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, 
      O_16_port, O_15_port, O_1_port, O_2_port, O_3_port, O_4_port, O_5_port, 
      O_6_port, O_7_port, O_8_port, O_9_port, O_10_port, O_11_port, O_12_port, 
      O_13_port, O_14_port : std_logic;

begin
   O <= ( O_47_port, O_46_port, O_45_port, O_44_port, O_43_port, O_42_port, 
      O_41_port, O_40_port, O_39_port, O_38_port, O_37_port, O_36_port, 
      O_35_port, O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, 
      O_29_port, O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, 
      O_23_port, O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, 
      O_17_port, O_16_port, O_15_port, O_14_port, O_13_port, O_12_port, 
      O_11_port, O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, 
      O_4_port, O_3_port, O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), 
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   A_nso <= ( A_ns(45), A_ns(44), A_ns(43), A_ns(42), A_ns(41), A_ns(40), 
      A_ns(39), A_ns(38), A_ns(37), A_ns(36), A_ns(35), A_ns(34), A_ns(33), 
      A_ns(32), A_ns(31), A_ns(30), A_ns(29), A_ns(28), A_ns(27), A_ns(26), 
      A_ns(25), A_ns(24), A_ns(23), A_ns(22), A_ns(21), A_ns(20), A_ns(19), 
      A_ns(18), A_ns(17), A_ns(16), A_ns(15), A_ns(14), A_ns(13), A_ns(12), 
      A_ns(11), A_ns(10), A_ns(9), A_ns(8), A_ns(7), A_ns(6), A_ns(5), A_ns(4),
      A_ns(3), A_ns(2), A_ns(1), A_ns(0), X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : OR3_X1 port map( A1 => B(13), A2 => B(14), A3 => n950, ZN => n813);
   U3 : INV_X2 port map( A => n813, ZN => n814);
   U4 : NAND2_X2 port map( A1 => n951, A2 => n817, ZN => n815);
   U5 : INV_X2 port map( A => n824, ZN => n820);
   U6 : NAND2_X2 port map( A1 => n951, A2 => n950, ZN => n817);
   U7 : OAI221_X1 port map( B1 => n815, B2 => n816, C1 => n817, C2 => n818, A 
                           => n819, ZN => O_45_port);
   U8 : AOI22_X1 port map( A1 => A_ns(43), A2 => n814, B1 => A_s(43), B2 => 
                           n820, ZN => n819);
   U9 : INV_X1 port map( A => A_s(44), ZN => n818);
   U10 : INV_X1 port map( A => A_ns(44), ZN => n816);
   U11 : OAI221_X1 port map( B1 => n815, B2 => n821, C1 => n817, C2 => n822, A 
                           => n823, ZN => O_46_port);
   U12 : AOI22_X1 port map( A1 => A_ns(44), A2 => n814, B1 => A_s(44), B2 => 
                           n820, ZN => n823);
   U13 : OAI221_X1 port map( B1 => n813, B2 => n821, C1 => n824, C2 => n822, A 
                           => n825, ZN => O_47_port);
   U14 : AOI22_X1 port map( A1 => A_ns(46), A2 => n826, B1 => A_s(46), B2 => 
                           n827, ZN => n825);
   U15 : INV_X1 port map( A => A_s(45), ZN => n822);
   U16 : INV_X1 port map( A => A_ns(45), ZN => n821);
   U17 : OAI221_X1 port map( B1 => n813, B2 => n828, C1 => n824, C2 => n829, A 
                           => n830, ZN => O_44_port);
   U18 : AOI22_X1 port map( A1 => n826, A2 => A_ns(43), B1 => n827, B2 => 
                           A_s(43), ZN => n830);
   U19 : OAI221_X1 port map( B1 => n815, B2 => n828, C1 => n817, C2 => n829, A 
                           => n831, ZN => O_43_port);
   U20 : AOI22_X1 port map( A1 => A_ns(41), A2 => n814, B1 => A_s(41), B2 => 
                           n820, ZN => n831);
   U21 : INV_X1 port map( A => A_s(42), ZN => n829);
   U22 : INV_X1 port map( A => A_ns(42), ZN => n828);
   U23 : OAI221_X1 port map( B1 => n815, B2 => n832, C1 => n817, C2 => n833, A 
                           => n834, ZN => O_42_port);
   U24 : AOI22_X1 port map( A1 => A_ns(40), A2 => n814, B1 => A_s(40), B2 => 
                           n820, ZN => n834);
   U25 : INV_X1 port map( A => A_s(41), ZN => n833);
   U26 : INV_X1 port map( A => A_ns(41), ZN => n832);
   U27 : OAI221_X1 port map( B1 => n815, B2 => n835, C1 => n817, C2 => n836, A 
                           => n837, ZN => O_41_port);
   U28 : AOI22_X1 port map( A1 => A_ns(39), A2 => n814, B1 => A_s(39), B2 => 
                           n820, ZN => n837);
   U29 : INV_X1 port map( A => A_s(40), ZN => n836);
   U30 : INV_X1 port map( A => A_ns(40), ZN => n835);
   U31 : OAI221_X1 port map( B1 => n815, B2 => n838, C1 => n817, C2 => n839, A 
                           => n840, ZN => O_40_port);
   U32 : AOI22_X1 port map( A1 => A_ns(38), A2 => n814, B1 => A_s(38), B2 => 
                           n820, ZN => n840);
   U33 : INV_X1 port map( A => A_s(39), ZN => n839);
   U34 : INV_X1 port map( A => A_ns(39), ZN => n838);
   U35 : OAI221_X1 port map( B1 => n815, B2 => n841, C1 => n817, C2 => n842, A 
                           => n843, ZN => O_39_port);
   U36 : AOI22_X1 port map( A1 => A_ns(37), A2 => n814, B1 => A_s(37), B2 => 
                           n820, ZN => n843);
   U37 : INV_X1 port map( A => A_s(38), ZN => n842);
   U38 : INV_X1 port map( A => A_ns(38), ZN => n841);
   U39 : OAI221_X1 port map( B1 => n815, B2 => n844, C1 => n817, C2 => n845, A 
                           => n846, ZN => O_38_port);
   U40 : AOI22_X1 port map( A1 => A_ns(36), A2 => n814, B1 => A_s(36), B2 => 
                           n820, ZN => n846);
   U41 : INV_X1 port map( A => A_s(37), ZN => n845);
   U42 : INV_X1 port map( A => A_ns(37), ZN => n844);
   U43 : OAI221_X1 port map( B1 => n815, B2 => n847, C1 => n817, C2 => n848, A 
                           => n849, ZN => O_37_port);
   U44 : AOI22_X1 port map( A1 => A_ns(35), A2 => n814, B1 => A_s(35), B2 => 
                           n820, ZN => n849);
   U45 : INV_X1 port map( A => A_s(36), ZN => n848);
   U46 : INV_X1 port map( A => A_ns(36), ZN => n847);
   U47 : OAI221_X1 port map( B1 => n815, B2 => n850, C1 => n817, C2 => n851, A 
                           => n852, ZN => O_36_port);
   U48 : AOI22_X1 port map( A1 => A_ns(34), A2 => n814, B1 => A_s(34), B2 => 
                           n820, ZN => n852);
   U49 : INV_X1 port map( A => A_s(35), ZN => n851);
   U50 : INV_X1 port map( A => A_ns(35), ZN => n850);
   U51 : OAI221_X1 port map( B1 => n815, B2 => n853, C1 => n817, C2 => n854, A 
                           => n855, ZN => O_35_port);
   U52 : AOI22_X1 port map( A1 => A_ns(33), A2 => n814, B1 => A_s(33), B2 => 
                           n820, ZN => n855);
   U53 : INV_X1 port map( A => A_s(34), ZN => n854);
   U54 : INV_X1 port map( A => A_ns(34), ZN => n853);
   U55 : OAI221_X1 port map( B1 => n815, B2 => n856, C1 => n817, C2 => n857, A 
                           => n858, ZN => O_34_port);
   U56 : AOI22_X1 port map( A1 => A_ns(32), A2 => n814, B1 => A_s(32), B2 => 
                           n820, ZN => n858);
   U57 : INV_X1 port map( A => A_s(33), ZN => n857);
   U58 : INV_X1 port map( A => A_ns(33), ZN => n856);
   U59 : OAI221_X1 port map( B1 => n815, B2 => n859, C1 => n817, C2 => n860, A 
                           => n861, ZN => O_33_port);
   U60 : AOI22_X1 port map( A1 => A_ns(31), A2 => n814, B1 => A_s(31), B2 => 
                           n820, ZN => n861);
   U61 : INV_X1 port map( A => A_s(32), ZN => n860);
   U62 : INV_X1 port map( A => A_ns(32), ZN => n859);
   U63 : OAI221_X1 port map( B1 => n815, B2 => n862, C1 => n817, C2 => n863, A 
                           => n864, ZN => O_32_port);
   U64 : AOI22_X1 port map( A1 => A_ns(30), A2 => n814, B1 => A_s(30), B2 => 
                           n820, ZN => n864);
   U65 : INV_X1 port map( A => A_s(31), ZN => n863);
   U66 : INV_X1 port map( A => A_ns(31), ZN => n862);
   U67 : OAI221_X1 port map( B1 => n815, B2 => n865, C1 => n817, C2 => n866, A 
                           => n867, ZN => O_31_port);
   U68 : AOI22_X1 port map( A1 => A_ns(29), A2 => n814, B1 => A_s(29), B2 => 
                           n820, ZN => n867);
   U69 : INV_X1 port map( A => A_s(30), ZN => n866);
   U70 : INV_X1 port map( A => A_ns(30), ZN => n865);
   U71 : OAI221_X1 port map( B1 => n815, B2 => n868, C1 => n817, C2 => n869, A 
                           => n870, ZN => O_30_port);
   U72 : AOI22_X1 port map( A1 => A_ns(28), A2 => n814, B1 => A_s(28), B2 => 
                           n820, ZN => n870);
   U73 : INV_X1 port map( A => A_s(29), ZN => n869);
   U74 : INV_X1 port map( A => A_ns(29), ZN => n868);
   U75 : OAI221_X1 port map( B1 => n815, B2 => n871, C1 => n817, C2 => n872, A 
                           => n873, ZN => O_29_port);
   U76 : AOI22_X1 port map( A1 => A_ns(27), A2 => n814, B1 => A_s(27), B2 => 
                           n820, ZN => n873);
   U77 : INV_X1 port map( A => A_s(28), ZN => n872);
   U78 : INV_X1 port map( A => A_ns(28), ZN => n871);
   U79 : OAI221_X1 port map( B1 => n815, B2 => n874, C1 => n817, C2 => n875, A 
                           => n876, ZN => O_28_port);
   U80 : AOI22_X1 port map( A1 => A_ns(26), A2 => n814, B1 => A_s(26), B2 => 
                           n820, ZN => n876);
   U81 : INV_X1 port map( A => A_s(27), ZN => n875);
   U82 : INV_X1 port map( A => A_ns(27), ZN => n874);
   U83 : OAI221_X1 port map( B1 => n815, B2 => n877, C1 => n817, C2 => n878, A 
                           => n879, ZN => O_27_port);
   U84 : AOI22_X1 port map( A1 => A_ns(25), A2 => n814, B1 => A_s(25), B2 => 
                           n820, ZN => n879);
   U85 : INV_X1 port map( A => A_s(26), ZN => n878);
   U86 : INV_X1 port map( A => A_ns(26), ZN => n877);
   U87 : OAI221_X1 port map( B1 => n815, B2 => n880, C1 => n817, C2 => n881, A 
                           => n882, ZN => O_26_port);
   U88 : AOI22_X1 port map( A1 => A_ns(24), A2 => n814, B1 => A_s(24), B2 => 
                           n820, ZN => n882);
   U89 : INV_X1 port map( A => A_s(25), ZN => n881);
   U90 : INV_X1 port map( A => A_ns(25), ZN => n880);
   U91 : OAI221_X1 port map( B1 => n815, B2 => n883, C1 => n817, C2 => n884, A 
                           => n885, ZN => O_25_port);
   U92 : AOI22_X1 port map( A1 => A_ns(23), A2 => n814, B1 => A_s(23), B2 => 
                           n820, ZN => n885);
   U93 : INV_X1 port map( A => A_s(24), ZN => n884);
   U94 : INV_X1 port map( A => A_ns(24), ZN => n883);
   U95 : OAI221_X1 port map( B1 => n815, B2 => n886, C1 => n817, C2 => n887, A 
                           => n888, ZN => O_24_port);
   U96 : AOI22_X1 port map( A1 => A_ns(22), A2 => n814, B1 => A_s(22), B2 => 
                           n820, ZN => n888);
   U97 : INV_X1 port map( A => A_s(23), ZN => n887);
   U98 : INV_X1 port map( A => A_ns(23), ZN => n886);
   U99 : OAI221_X1 port map( B1 => n815, B2 => n889, C1 => n817, C2 => n890, A 
                           => n891, ZN => O_23_port);
   U100 : AOI22_X1 port map( A1 => A_ns(21), A2 => n814, B1 => A_s(21), B2 => 
                           n820, ZN => n891);
   U101 : INV_X1 port map( A => A_s(22), ZN => n890);
   U102 : INV_X1 port map( A => A_ns(22), ZN => n889);
   U103 : OAI221_X1 port map( B1 => n815, B2 => n892, C1 => n817, C2 => n893, A
                           => n894, ZN => O_22_port);
   U104 : AOI22_X1 port map( A1 => A_ns(20), A2 => n814, B1 => A_s(20), B2 => 
                           n820, ZN => n894);
   U105 : INV_X1 port map( A => A_s(21), ZN => n893);
   U106 : INV_X1 port map( A => A_ns(21), ZN => n892);
   U107 : OAI221_X1 port map( B1 => n815, B2 => n895, C1 => n817, C2 => n896, A
                           => n897, ZN => O_21_port);
   U108 : AOI22_X1 port map( A1 => A_ns(19), A2 => n814, B1 => A_s(19), B2 => 
                           n820, ZN => n897);
   U109 : INV_X1 port map( A => A_s(20), ZN => n896);
   U110 : INV_X1 port map( A => A_ns(20), ZN => n895);
   U111 : OAI221_X1 port map( B1 => n815, B2 => n898, C1 => n817, C2 => n899, A
                           => n900, ZN => O_20_port);
   U112 : AOI22_X1 port map( A1 => A_ns(18), A2 => n814, B1 => A_s(18), B2 => 
                           n820, ZN => n900);
   U113 : INV_X1 port map( A => A_s(19), ZN => n899);
   U114 : INV_X1 port map( A => A_ns(19), ZN => n898);
   U115 : OAI221_X1 port map( B1 => n815, B2 => n901, C1 => n817, C2 => n902, A
                           => n903, ZN => O_19_port);
   U116 : AOI22_X1 port map( A1 => A_ns(17), A2 => n814, B1 => A_s(17), B2 => 
                           n820, ZN => n903);
   U117 : INV_X1 port map( A => A_s(18), ZN => n902);
   U118 : INV_X1 port map( A => A_ns(18), ZN => n901);
   U119 : OAI221_X1 port map( B1 => n815, B2 => n904, C1 => n817, C2 => n905, A
                           => n906, ZN => O_18_port);
   U120 : AOI22_X1 port map( A1 => A_ns(16), A2 => n814, B1 => A_s(16), B2 => 
                           n820, ZN => n906);
   U121 : INV_X1 port map( A => A_s(17), ZN => n905);
   U122 : INV_X1 port map( A => A_ns(17), ZN => n904);
   U123 : OAI221_X1 port map( B1 => n815, B2 => n907, C1 => n817, C2 => n908, A
                           => n909, ZN => O_17_port);
   U124 : AOI22_X1 port map( A1 => A_ns(15), A2 => n814, B1 => A_s(15), B2 => 
                           n820, ZN => n909);
   U125 : INV_X1 port map( A => A_s(16), ZN => n908);
   U126 : INV_X1 port map( A => A_ns(16), ZN => n907);
   U127 : OAI221_X1 port map( B1 => n815, B2 => n910, C1 => n817, C2 => n911, A
                           => n912, ZN => O_16_port);
   U128 : AOI22_X1 port map( A1 => A_ns(14), A2 => n814, B1 => A_s(14), B2 => 
                           n820, ZN => n912);
   U129 : INV_X1 port map( A => A_s(15), ZN => n911);
   U130 : INV_X1 port map( A => A_ns(15), ZN => n910);
   U131 : OAI221_X1 port map( B1 => n815, B2 => n913, C1 => n817, C2 => n914, A
                           => n915, ZN => O_15_port);
   U132 : AOI22_X1 port map( A1 => A_ns(13), A2 => n814, B1 => A_s(13), B2 => 
                           n820, ZN => n915);
   U133 : INV_X1 port map( A => A_s(14), ZN => n914);
   U134 : INV_X1 port map( A => A_ns(14), ZN => n913);
   U135 : INV_X1 port map( A => n916, ZN => O_1_port);
   U136 : AOI22_X1 port map( A1 => n827, A2 => A_s(0), B1 => n826, B2 => 
                           A_ns(0), ZN => n916);
   U137 : OAI221_X1 port map( B1 => n815, B2 => n917, C1 => n817, C2 => n918, A
                           => n919, ZN => O_2_port);
   U138 : AOI22_X1 port map( A1 => A_ns(0), A2 => n814, B1 => A_s(0), B2 => 
                           n820, ZN => n919);
   U139 : INV_X1 port map( A => n920, ZN => O_3_port);
   U140 : AOI221_X1 port map( B1 => n826, B2 => A_ns(2), C1 => n827, C2 => 
                           A_s(2), A => n921, ZN => n920);
   U141 : OAI22_X1 port map( A1 => n917, A2 => n813, B1 => n918, B2 => n824, ZN
                           => n921);
   U142 : INV_X1 port map( A => A_s(1), ZN => n918);
   U143 : INV_X1 port map( A => A_ns(1), ZN => n917);
   U144 : OAI221_X1 port map( B1 => n815, B2 => n922, C1 => n817, C2 => n923, A
                           => n924, ZN => O_4_port);
   U145 : AOI22_X1 port map( A1 => A_ns(2), A2 => n814, B1 => A_s(2), B2 => 
                           n820, ZN => n924);
   U146 : INV_X1 port map( A => n925, ZN => O_5_port);
   U147 : AOI221_X1 port map( B1 => n826, B2 => A_ns(4), C1 => n827, C2 => 
                           A_s(4), A => n926, ZN => n925);
   U148 : OAI22_X1 port map( A1 => n922, A2 => n813, B1 => n923, B2 => n824, ZN
                           => n926);
   U149 : INV_X1 port map( A => A_s(3), ZN => n923);
   U150 : INV_X1 port map( A => A_ns(3), ZN => n922);
   U151 : OAI221_X1 port map( B1 => n815, B2 => n927, C1 => n817, C2 => n928, A
                           => n929, ZN => O_6_port);
   U152 : AOI22_X1 port map( A1 => A_ns(4), A2 => n814, B1 => A_s(4), B2 => 
                           n820, ZN => n929);
   U153 : INV_X1 port map( A => n930, ZN => O_7_port);
   U154 : AOI221_X1 port map( B1 => n826, B2 => A_ns(6), C1 => n827, C2 => 
                           A_s(6), A => n931, ZN => n930);
   U155 : OAI22_X1 port map( A1 => n927, A2 => n813, B1 => n928, B2 => n824, ZN
                           => n931);
   U156 : INV_X1 port map( A => A_s(5), ZN => n928);
   U157 : INV_X1 port map( A => A_ns(5), ZN => n927);
   U158 : OAI221_X1 port map( B1 => n815, B2 => n932, C1 => n817, C2 => n933, A
                           => n934, ZN => O_8_port);
   U159 : AOI22_X1 port map( A1 => A_ns(6), A2 => n814, B1 => A_s(6), B2 => 
                           n820, ZN => n934);
   U160 : INV_X1 port map( A => n935, ZN => O_9_port);
   U161 : AOI221_X1 port map( B1 => n826, B2 => A_ns(8), C1 => n827, C2 => 
                           A_s(8), A => n936, ZN => n935);
   U162 : OAI22_X1 port map( A1 => n932, A2 => n813, B1 => n933, B2 => n824, ZN
                           => n936);
   U163 : INV_X1 port map( A => A_s(7), ZN => n933);
   U164 : INV_X1 port map( A => A_ns(7), ZN => n932);
   U165 : OAI221_X1 port map( B1 => n815, B2 => n937, C1 => n817, C2 => n938, A
                           => n939, ZN => O_10_port);
   U166 : AOI22_X1 port map( A1 => A_ns(8), A2 => n814, B1 => A_s(8), B2 => 
                           n820, ZN => n939);
   U167 : INV_X1 port map( A => n940, ZN => O_11_port);
   U168 : AOI221_X1 port map( B1 => n826, B2 => A_ns(10), C1 => n827, C2 => 
                           A_s(10), A => n941, ZN => n940);
   U169 : OAI22_X1 port map( A1 => n937, A2 => n813, B1 => n938, B2 => n824, ZN
                           => n941);
   U170 : INV_X1 port map( A => A_s(9), ZN => n938);
   U171 : INV_X1 port map( A => A_ns(9), ZN => n937);
   U172 : OAI221_X1 port map( B1 => n815, B2 => n942, C1 => n817, C2 => n943, A
                           => n944, ZN => O_12_port);
   U173 : AOI22_X1 port map( A1 => A_ns(10), A2 => n814, B1 => A_s(10), B2 => 
                           n820, ZN => n944);
   U174 : INV_X1 port map( A => n945, ZN => O_13_port);
   U175 : AOI221_X1 port map( B1 => n826, B2 => A_ns(12), C1 => n827, C2 => 
                           A_s(12), A => n946, ZN => n945);
   U176 : OAI22_X1 port map( A1 => n942, A2 => n813, B1 => n943, B2 => n824, ZN
                           => n946);
   U177 : INV_X1 port map( A => A_s(11), ZN => n943);
   U178 : INV_X1 port map( A => A_ns(11), ZN => n942);
   U179 : INV_X1 port map( A => n817, ZN => n827);
   U180 : INV_X1 port map( A => n815, ZN => n826);
   U181 : OAI221_X1 port map( B1 => n815, B2 => n947, C1 => n817, C2 => n948, A
                           => n949, ZN => O_14_port);
   U182 : AOI22_X1 port map( A1 => A_ns(12), A2 => n814, B1 => A_s(12), B2 => 
                           n820, ZN => n949);
   U183 : NAND3_X1 port map( A1 => B(13), A2 => n950, A3 => B(14), ZN => n824);
   U184 : INV_X1 port map( A => A_s(13), ZN => n948);
   U185 : INV_X1 port map( A => A_ns(13), ZN => n947);
   U186 : INV_X1 port map( A => B(15), ZN => n950);
   U187 : XOR2_X1 port map( A => B(14), B => B(13), Z => n951);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT46_i12 is

   port( A_s, A_ns, B : in std_logic_vector (45 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (45 downto 0));

end BOOTHENC_NBIT46_i12;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT46_i12 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, n781, n782, n783, n784, n785, n786, n787, n788, n789, 
      n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, 
      n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, 
      n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, 
      n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, 
      n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, 
      n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, 
      n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, 
      n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, 
      n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, 
      n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, 
      n910, n911, n912, n913, n914, O_43_port, O_44_port, O_45_port, O_42_port,
      O_41_port, O_40_port, O_39_port, O_38_port, O_37_port, O_36_port, 
      O_35_port, O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, 
      O_29_port, O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, 
      O_23_port, O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, 
      O_17_port, O_16_port, O_15_port, O_14_port, O_13_port, O_1_port, O_2_port
      , O_3_port, O_4_port, O_5_port, O_6_port, O_7_port, O_8_port, O_9_port, 
      O_10_port, O_11_port, O_12_port : std_logic;

begin
   O <= ( O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, O_40_port, 
      O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, 
      O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, 
      O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, 
      O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, O_16_port, 
      O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, O_10_port, 
      O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, O_3_port, 
      O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), A_s(38), A_s(37), 
      A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), A_s(30), A_s(29), 
      A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), A_s(22), A_s(21), 
      A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), A_s(14), A_s(13), 
      A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), A_s(6), A_s(5), A_s(4)
      , A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, X_Logic0_port );
   A_nso <= ( A_ns(43), A_ns(42), A_ns(41), A_ns(40), A_ns(39), A_ns(38), 
      A_ns(37), A_ns(36), A_ns(35), A_ns(34), A_ns(33), A_ns(32), A_ns(31), 
      A_ns(30), A_ns(29), A_ns(28), A_ns(27), A_ns(26), A_ns(25), A_ns(24), 
      A_ns(23), A_ns(22), A_ns(21), A_ns(20), A_ns(19), A_ns(18), A_ns(17), 
      A_ns(16), A_ns(15), A_ns(14), A_ns(13), A_ns(12), A_ns(11), A_ns(10), 
      A_ns(9), A_ns(8), A_ns(7), A_ns(6), A_ns(5), A_ns(4), A_ns(3), A_ns(2), 
      A_ns(1), A_ns(0), X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : OR3_X1 port map( A1 => B(11), A2 => B(12), A3 => n913, ZN => n781);
   U3 : INV_X2 port map( A => n781, ZN => n782);
   U4 : NAND2_X2 port map( A1 => n914, A2 => n785, ZN => n783);
   U5 : INV_X2 port map( A => n792, ZN => n788);
   U6 : NAND2_X2 port map( A1 => n914, A2 => n913, ZN => n785);
   U7 : OAI221_X1 port map( B1 => n783, B2 => n784, C1 => n785, C2 => n786, A 
                           => n787, ZN => O_43_port);
   U8 : AOI22_X1 port map( A1 => A_ns(41), A2 => n782, B1 => A_s(41), B2 => 
                           n788, ZN => n787);
   U9 : INV_X1 port map( A => A_s(42), ZN => n786);
   U10 : INV_X1 port map( A => A_ns(42), ZN => n784);
   U11 : OAI221_X1 port map( B1 => n783, B2 => n789, C1 => n785, C2 => n790, A 
                           => n791, ZN => O_44_port);
   U12 : AOI22_X1 port map( A1 => A_ns(42), A2 => n782, B1 => A_s(42), B2 => 
                           n788, ZN => n791);
   U13 : OAI221_X1 port map( B1 => n781, B2 => n789, C1 => n792, C2 => n790, A 
                           => n793, ZN => O_45_port);
   U14 : AOI22_X1 port map( A1 => A_ns(44), A2 => n794, B1 => A_s(44), B2 => 
                           n795, ZN => n793);
   U15 : INV_X1 port map( A => A_s(43), ZN => n790);
   U16 : INV_X1 port map( A => A_ns(43), ZN => n789);
   U17 : OAI221_X1 port map( B1 => n781, B2 => n796, C1 => n792, C2 => n797, A 
                           => n798, ZN => O_42_port);
   U18 : AOI22_X1 port map( A1 => n794, A2 => A_ns(41), B1 => n795, B2 => 
                           A_s(41), ZN => n798);
   U19 : OAI221_X1 port map( B1 => n783, B2 => n796, C1 => n785, C2 => n797, A 
                           => n799, ZN => O_41_port);
   U20 : AOI22_X1 port map( A1 => A_ns(39), A2 => n782, B1 => A_s(39), B2 => 
                           n788, ZN => n799);
   U21 : INV_X1 port map( A => A_s(40), ZN => n797);
   U22 : INV_X1 port map( A => A_ns(40), ZN => n796);
   U23 : OAI221_X1 port map( B1 => n783, B2 => n800, C1 => n785, C2 => n801, A 
                           => n802, ZN => O_40_port);
   U24 : AOI22_X1 port map( A1 => A_ns(38), A2 => n782, B1 => A_s(38), B2 => 
                           n788, ZN => n802);
   U25 : INV_X1 port map( A => A_s(39), ZN => n801);
   U26 : INV_X1 port map( A => A_ns(39), ZN => n800);
   U27 : OAI221_X1 port map( B1 => n783, B2 => n803, C1 => n785, C2 => n804, A 
                           => n805, ZN => O_39_port);
   U28 : AOI22_X1 port map( A1 => A_ns(37), A2 => n782, B1 => A_s(37), B2 => 
                           n788, ZN => n805);
   U29 : INV_X1 port map( A => A_s(38), ZN => n804);
   U30 : INV_X1 port map( A => A_ns(38), ZN => n803);
   U31 : OAI221_X1 port map( B1 => n783, B2 => n806, C1 => n785, C2 => n807, A 
                           => n808, ZN => O_38_port);
   U32 : AOI22_X1 port map( A1 => A_ns(36), A2 => n782, B1 => A_s(36), B2 => 
                           n788, ZN => n808);
   U33 : INV_X1 port map( A => A_s(37), ZN => n807);
   U34 : INV_X1 port map( A => A_ns(37), ZN => n806);
   U35 : OAI221_X1 port map( B1 => n783, B2 => n809, C1 => n785, C2 => n810, A 
                           => n811, ZN => O_37_port);
   U36 : AOI22_X1 port map( A1 => A_ns(35), A2 => n782, B1 => A_s(35), B2 => 
                           n788, ZN => n811);
   U37 : INV_X1 port map( A => A_s(36), ZN => n810);
   U38 : INV_X1 port map( A => A_ns(36), ZN => n809);
   U39 : OAI221_X1 port map( B1 => n783, B2 => n812, C1 => n785, C2 => n813, A 
                           => n814, ZN => O_36_port);
   U40 : AOI22_X1 port map( A1 => A_ns(34), A2 => n782, B1 => A_s(34), B2 => 
                           n788, ZN => n814);
   U41 : INV_X1 port map( A => A_s(35), ZN => n813);
   U42 : INV_X1 port map( A => A_ns(35), ZN => n812);
   U43 : OAI221_X1 port map( B1 => n783, B2 => n815, C1 => n785, C2 => n816, A 
                           => n817, ZN => O_35_port);
   U44 : AOI22_X1 port map( A1 => A_ns(33), A2 => n782, B1 => A_s(33), B2 => 
                           n788, ZN => n817);
   U45 : INV_X1 port map( A => A_s(34), ZN => n816);
   U46 : INV_X1 port map( A => A_ns(34), ZN => n815);
   U47 : OAI221_X1 port map( B1 => n783, B2 => n818, C1 => n785, C2 => n819, A 
                           => n820, ZN => O_34_port);
   U48 : AOI22_X1 port map( A1 => A_ns(32), A2 => n782, B1 => A_s(32), B2 => 
                           n788, ZN => n820);
   U49 : INV_X1 port map( A => A_s(33), ZN => n819);
   U50 : INV_X1 port map( A => A_ns(33), ZN => n818);
   U51 : OAI221_X1 port map( B1 => n783, B2 => n821, C1 => n785, C2 => n822, A 
                           => n823, ZN => O_33_port);
   U52 : AOI22_X1 port map( A1 => A_ns(31), A2 => n782, B1 => A_s(31), B2 => 
                           n788, ZN => n823);
   U53 : INV_X1 port map( A => A_s(32), ZN => n822);
   U54 : INV_X1 port map( A => A_ns(32), ZN => n821);
   U55 : OAI221_X1 port map( B1 => n783, B2 => n824, C1 => n785, C2 => n825, A 
                           => n826, ZN => O_32_port);
   U56 : AOI22_X1 port map( A1 => A_ns(30), A2 => n782, B1 => A_s(30), B2 => 
                           n788, ZN => n826);
   U57 : INV_X1 port map( A => A_s(31), ZN => n825);
   U58 : INV_X1 port map( A => A_ns(31), ZN => n824);
   U59 : OAI221_X1 port map( B1 => n783, B2 => n827, C1 => n785, C2 => n828, A 
                           => n829, ZN => O_31_port);
   U60 : AOI22_X1 port map( A1 => A_ns(29), A2 => n782, B1 => A_s(29), B2 => 
                           n788, ZN => n829);
   U61 : INV_X1 port map( A => A_s(30), ZN => n828);
   U62 : INV_X1 port map( A => A_ns(30), ZN => n827);
   U63 : OAI221_X1 port map( B1 => n783, B2 => n830, C1 => n785, C2 => n831, A 
                           => n832, ZN => O_30_port);
   U64 : AOI22_X1 port map( A1 => A_ns(28), A2 => n782, B1 => A_s(28), B2 => 
                           n788, ZN => n832);
   U65 : INV_X1 port map( A => A_s(29), ZN => n831);
   U66 : INV_X1 port map( A => A_ns(29), ZN => n830);
   U67 : OAI221_X1 port map( B1 => n783, B2 => n833, C1 => n785, C2 => n834, A 
                           => n835, ZN => O_29_port);
   U68 : AOI22_X1 port map( A1 => A_ns(27), A2 => n782, B1 => A_s(27), B2 => 
                           n788, ZN => n835);
   U69 : INV_X1 port map( A => A_s(28), ZN => n834);
   U70 : INV_X1 port map( A => A_ns(28), ZN => n833);
   U71 : OAI221_X1 port map( B1 => n783, B2 => n836, C1 => n785, C2 => n837, A 
                           => n838, ZN => O_28_port);
   U72 : AOI22_X1 port map( A1 => A_ns(26), A2 => n782, B1 => A_s(26), B2 => 
                           n788, ZN => n838);
   U73 : INV_X1 port map( A => A_s(27), ZN => n837);
   U74 : INV_X1 port map( A => A_ns(27), ZN => n836);
   U75 : OAI221_X1 port map( B1 => n783, B2 => n839, C1 => n785, C2 => n840, A 
                           => n841, ZN => O_27_port);
   U76 : AOI22_X1 port map( A1 => A_ns(25), A2 => n782, B1 => A_s(25), B2 => 
                           n788, ZN => n841);
   U77 : INV_X1 port map( A => A_s(26), ZN => n840);
   U78 : INV_X1 port map( A => A_ns(26), ZN => n839);
   U79 : OAI221_X1 port map( B1 => n783, B2 => n842, C1 => n785, C2 => n843, A 
                           => n844, ZN => O_26_port);
   U80 : AOI22_X1 port map( A1 => A_ns(24), A2 => n782, B1 => A_s(24), B2 => 
                           n788, ZN => n844);
   U81 : INV_X1 port map( A => A_s(25), ZN => n843);
   U82 : INV_X1 port map( A => A_ns(25), ZN => n842);
   U83 : OAI221_X1 port map( B1 => n783, B2 => n845, C1 => n785, C2 => n846, A 
                           => n847, ZN => O_25_port);
   U84 : AOI22_X1 port map( A1 => A_ns(23), A2 => n782, B1 => A_s(23), B2 => 
                           n788, ZN => n847);
   U85 : INV_X1 port map( A => A_s(24), ZN => n846);
   U86 : INV_X1 port map( A => A_ns(24), ZN => n845);
   U87 : OAI221_X1 port map( B1 => n783, B2 => n848, C1 => n785, C2 => n849, A 
                           => n850, ZN => O_24_port);
   U88 : AOI22_X1 port map( A1 => A_ns(22), A2 => n782, B1 => A_s(22), B2 => 
                           n788, ZN => n850);
   U89 : INV_X1 port map( A => A_s(23), ZN => n849);
   U90 : INV_X1 port map( A => A_ns(23), ZN => n848);
   U91 : OAI221_X1 port map( B1 => n783, B2 => n851, C1 => n785, C2 => n852, A 
                           => n853, ZN => O_23_port);
   U92 : AOI22_X1 port map( A1 => A_ns(21), A2 => n782, B1 => A_s(21), B2 => 
                           n788, ZN => n853);
   U93 : INV_X1 port map( A => A_s(22), ZN => n852);
   U94 : INV_X1 port map( A => A_ns(22), ZN => n851);
   U95 : OAI221_X1 port map( B1 => n783, B2 => n854, C1 => n785, C2 => n855, A 
                           => n856, ZN => O_22_port);
   U96 : AOI22_X1 port map( A1 => A_ns(20), A2 => n782, B1 => A_s(20), B2 => 
                           n788, ZN => n856);
   U97 : INV_X1 port map( A => A_s(21), ZN => n855);
   U98 : INV_X1 port map( A => A_ns(21), ZN => n854);
   U99 : OAI221_X1 port map( B1 => n783, B2 => n857, C1 => n785, C2 => n858, A 
                           => n859, ZN => O_21_port);
   U100 : AOI22_X1 port map( A1 => A_ns(19), A2 => n782, B1 => A_s(19), B2 => 
                           n788, ZN => n859);
   U101 : INV_X1 port map( A => A_s(20), ZN => n858);
   U102 : INV_X1 port map( A => A_ns(20), ZN => n857);
   U103 : OAI221_X1 port map( B1 => n783, B2 => n860, C1 => n785, C2 => n861, A
                           => n862, ZN => O_20_port);
   U104 : AOI22_X1 port map( A1 => A_ns(18), A2 => n782, B1 => A_s(18), B2 => 
                           n788, ZN => n862);
   U105 : INV_X1 port map( A => A_s(19), ZN => n861);
   U106 : INV_X1 port map( A => A_ns(19), ZN => n860);
   U107 : OAI221_X1 port map( B1 => n783, B2 => n863, C1 => n785, C2 => n864, A
                           => n865, ZN => O_19_port);
   U108 : AOI22_X1 port map( A1 => A_ns(17), A2 => n782, B1 => A_s(17), B2 => 
                           n788, ZN => n865);
   U109 : INV_X1 port map( A => A_s(18), ZN => n864);
   U110 : INV_X1 port map( A => A_ns(18), ZN => n863);
   U111 : OAI221_X1 port map( B1 => n783, B2 => n866, C1 => n785, C2 => n867, A
                           => n868, ZN => O_18_port);
   U112 : AOI22_X1 port map( A1 => A_ns(16), A2 => n782, B1 => A_s(16), B2 => 
                           n788, ZN => n868);
   U113 : INV_X1 port map( A => A_s(17), ZN => n867);
   U114 : INV_X1 port map( A => A_ns(17), ZN => n866);
   U115 : OAI221_X1 port map( B1 => n783, B2 => n869, C1 => n785, C2 => n870, A
                           => n871, ZN => O_17_port);
   U116 : AOI22_X1 port map( A1 => A_ns(15), A2 => n782, B1 => A_s(15), B2 => 
                           n788, ZN => n871);
   U117 : INV_X1 port map( A => A_s(16), ZN => n870);
   U118 : INV_X1 port map( A => A_ns(16), ZN => n869);
   U119 : OAI221_X1 port map( B1 => n783, B2 => n872, C1 => n785, C2 => n873, A
                           => n874, ZN => O_16_port);
   U120 : AOI22_X1 port map( A1 => A_ns(14), A2 => n782, B1 => A_s(14), B2 => 
                           n788, ZN => n874);
   U121 : INV_X1 port map( A => A_s(15), ZN => n873);
   U122 : INV_X1 port map( A => A_ns(15), ZN => n872);
   U123 : OAI221_X1 port map( B1 => n783, B2 => n875, C1 => n785, C2 => n876, A
                           => n877, ZN => O_15_port);
   U124 : AOI22_X1 port map( A1 => A_ns(13), A2 => n782, B1 => A_s(13), B2 => 
                           n788, ZN => n877);
   U125 : INV_X1 port map( A => A_s(14), ZN => n876);
   U126 : INV_X1 port map( A => A_ns(14), ZN => n875);
   U127 : OAI221_X1 port map( B1 => n783, B2 => n878, C1 => n785, C2 => n879, A
                           => n880, ZN => O_14_port);
   U128 : AOI22_X1 port map( A1 => A_ns(12), A2 => n782, B1 => A_s(12), B2 => 
                           n788, ZN => n880);
   U129 : INV_X1 port map( A => A_s(13), ZN => n879);
   U130 : INV_X1 port map( A => A_ns(13), ZN => n878);
   U131 : OAI221_X1 port map( B1 => n783, B2 => n881, C1 => n785, C2 => n882, A
                           => n883, ZN => O_13_port);
   U132 : AOI22_X1 port map( A1 => A_ns(11), A2 => n782, B1 => A_s(11), B2 => 
                           n788, ZN => n883);
   U133 : INV_X1 port map( A => A_s(12), ZN => n882);
   U134 : INV_X1 port map( A => A_ns(12), ZN => n881);
   U135 : INV_X1 port map( A => n884, ZN => O_1_port);
   U136 : AOI22_X1 port map( A1 => n795, A2 => A_s(0), B1 => n794, B2 => 
                           A_ns(0), ZN => n884);
   U137 : OAI221_X1 port map( B1 => n783, B2 => n885, C1 => n785, C2 => n886, A
                           => n887, ZN => O_2_port);
   U138 : AOI22_X1 port map( A1 => A_ns(0), A2 => n782, B1 => A_s(0), B2 => 
                           n788, ZN => n887);
   U139 : INV_X1 port map( A => n888, ZN => O_3_port);
   U140 : AOI221_X1 port map( B1 => n794, B2 => A_ns(2), C1 => n795, C2 => 
                           A_s(2), A => n889, ZN => n888);
   U141 : OAI22_X1 port map( A1 => n885, A2 => n781, B1 => n886, B2 => n792, ZN
                           => n889);
   U142 : INV_X1 port map( A => A_s(1), ZN => n886);
   U143 : INV_X1 port map( A => A_ns(1), ZN => n885);
   U144 : OAI221_X1 port map( B1 => n783, B2 => n890, C1 => n785, C2 => n891, A
                           => n892, ZN => O_4_port);
   U145 : AOI22_X1 port map( A1 => A_ns(2), A2 => n782, B1 => A_s(2), B2 => 
                           n788, ZN => n892);
   U146 : INV_X1 port map( A => n893, ZN => O_5_port);
   U147 : AOI221_X1 port map( B1 => n794, B2 => A_ns(4), C1 => n795, C2 => 
                           A_s(4), A => n894, ZN => n893);
   U148 : OAI22_X1 port map( A1 => n890, A2 => n781, B1 => n891, B2 => n792, ZN
                           => n894);
   U149 : INV_X1 port map( A => A_s(3), ZN => n891);
   U150 : INV_X1 port map( A => A_ns(3), ZN => n890);
   U151 : OAI221_X1 port map( B1 => n783, B2 => n895, C1 => n785, C2 => n896, A
                           => n897, ZN => O_6_port);
   U152 : AOI22_X1 port map( A1 => A_ns(4), A2 => n782, B1 => A_s(4), B2 => 
                           n788, ZN => n897);
   U153 : INV_X1 port map( A => n898, ZN => O_7_port);
   U154 : AOI221_X1 port map( B1 => n794, B2 => A_ns(6), C1 => n795, C2 => 
                           A_s(6), A => n899, ZN => n898);
   U155 : OAI22_X1 port map( A1 => n895, A2 => n781, B1 => n896, B2 => n792, ZN
                           => n899);
   U156 : INV_X1 port map( A => A_s(5), ZN => n896);
   U157 : INV_X1 port map( A => A_ns(5), ZN => n895);
   U158 : OAI221_X1 port map( B1 => n783, B2 => n900, C1 => n785, C2 => n901, A
                           => n902, ZN => O_8_port);
   U159 : AOI22_X1 port map( A1 => A_ns(6), A2 => n782, B1 => A_s(6), B2 => 
                           n788, ZN => n902);
   U160 : INV_X1 port map( A => n903, ZN => O_9_port);
   U161 : AOI221_X1 port map( B1 => n794, B2 => A_ns(8), C1 => n795, C2 => 
                           A_s(8), A => n904, ZN => n903);
   U162 : OAI22_X1 port map( A1 => n900, A2 => n781, B1 => n901, B2 => n792, ZN
                           => n904);
   U163 : INV_X1 port map( A => A_s(7), ZN => n901);
   U164 : INV_X1 port map( A => A_ns(7), ZN => n900);
   U165 : OAI221_X1 port map( B1 => n783, B2 => n905, C1 => n785, C2 => n906, A
                           => n907, ZN => O_10_port);
   U166 : AOI22_X1 port map( A1 => A_ns(8), A2 => n782, B1 => A_s(8), B2 => 
                           n788, ZN => n907);
   U167 : INV_X1 port map( A => n908, ZN => O_11_port);
   U168 : AOI221_X1 port map( B1 => n794, B2 => A_ns(10), C1 => n795, C2 => 
                           A_s(10), A => n909, ZN => n908);
   U169 : OAI22_X1 port map( A1 => n905, A2 => n781, B1 => n906, B2 => n792, ZN
                           => n909);
   U170 : INV_X1 port map( A => A_s(9), ZN => n906);
   U171 : INV_X1 port map( A => A_ns(9), ZN => n905);
   U172 : INV_X1 port map( A => n785, ZN => n795);
   U173 : INV_X1 port map( A => n783, ZN => n794);
   U174 : OAI221_X1 port map( B1 => n783, B2 => n910, C1 => n785, C2 => n911, A
                           => n912, ZN => O_12_port);
   U175 : AOI22_X1 port map( A1 => A_ns(10), A2 => n782, B1 => A_s(10), B2 => 
                           n788, ZN => n912);
   U176 : NAND3_X1 port map( A1 => B(11), A2 => n913, A3 => B(12), ZN => n792);
   U177 : INV_X1 port map( A => A_s(11), ZN => n911);
   U178 : INV_X1 port map( A => A_ns(11), ZN => n910);
   U179 : INV_X1 port map( A => B(13), ZN => n913);
   U180 : XOR2_X1 port map( A => B(12), B => B(11), Z => n914);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT44_i10 is

   port( A_s, A_ns, B : in std_logic_vector (43 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (43 downto 0));

end BOOTHENC_NBIT44_i10;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT44_i10 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, n750, n751, n752, n753, n754, n755, n756, n757, n758, 
      n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, 
      n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, 
      n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, 
      n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, 
      n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, 
      n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, 
      n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, 
      n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, 
      n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, 
      n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, 
      n879, n880, O_42_port, O_41_port, O_43_port, O_40_port, O_39_port, 
      O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, O_33_port, 
      O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, O_27_port, 
      O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, O_21_port, 
      O_20_port, O_19_port, O_18_port, O_17_port, O_16_port, O_15_port, 
      O_14_port, O_13_port, O_12_port, O_11_port, O_1_port, O_2_port, O_3_port,
      O_4_port, O_5_port, O_6_port, O_7_port, O_8_port, O_9_port, O_10_port : 
      std_logic;

begin
   O <= ( O_43_port, O_42_port, O_41_port, O_40_port, O_39_port, O_38_port, 
      O_37_port, O_36_port, O_35_port, O_34_port, O_33_port, O_32_port, 
      O_31_port, O_30_port, O_29_port, O_28_port, O_27_port, O_26_port, 
      O_25_port, O_24_port, O_23_port, O_22_port, O_21_port, O_20_port, 
      O_19_port, O_18_port, O_17_port, O_16_port, O_15_port, O_14_port, 
      O_13_port, O_12_port, O_11_port, O_10_port, O_9_port, O_8_port, O_7_port,
      O_6_port, O_5_port, O_4_port, O_3_port, O_2_port, O_1_port, X_Logic0_port
      );
   A_so <= ( A_s(41), A_s(40), A_s(39), A_s(38), A_s(37), A_s(36), A_s(35), 
      A_s(34), A_s(33), A_s(32), A_s(31), A_s(30), A_s(29), A_s(28), A_s(27), 
      A_s(26), A_s(25), A_s(24), A_s(23), A_s(22), A_s(21), A_s(20), A_s(19), 
      A_s(18), A_s(17), A_s(16), A_s(15), A_s(14), A_s(13), A_s(12), A_s(11), 
      A_s(10), A_s(9), A_s(8), A_s(7), A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), 
      A_s(1), A_s(0), X_Logic0_port, X_Logic0_port );
   A_nso <= ( A_ns(41), A_ns(40), A_ns(39), A_ns(38), A_ns(37), A_ns(36), 
      A_ns(35), A_ns(34), A_ns(33), A_ns(32), A_ns(31), A_ns(30), A_ns(29), 
      A_ns(28), A_ns(27), A_ns(26), A_ns(25), A_ns(24), A_ns(23), A_ns(22), 
      A_ns(21), A_ns(20), A_ns(19), A_ns(18), A_ns(17), A_ns(16), A_ns(15), 
      A_ns(14), A_ns(13), A_ns(12), A_ns(11), A_ns(10), A_ns(9), A_ns(8), 
      A_ns(7), A_ns(6), A_ns(5), A_ns(4), A_ns(3), A_ns(2), A_ns(1), A_ns(0), 
      X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : OR3_X1 port map( A1 => B(10), A2 => B(9), A3 => n879, ZN => n750);
   U3 : INV_X2 port map( A => n750, ZN => n751);
   U4 : NAND2_X2 port map( A1 => n880, A2 => n754, ZN => n752);
   U5 : INV_X2 port map( A => n761, ZN => n757);
   U6 : NAND2_X2 port map( A1 => n880, A2 => n879, ZN => n754);
   U7 : OAI221_X1 port map( B1 => n752, B2 => n753, C1 => n754, C2 => n755, A 
                           => n756, ZN => O_42_port);
   U8 : AOI22_X1 port map( A1 => A_ns(40), A2 => n751, B1 => A_s(40), B2 => 
                           n757, ZN => n756);
   U9 : OAI221_X1 port map( B1 => n758, B2 => n752, C1 => n759, C2 => n754, A 
                           => n760, ZN => O_41_port);
   U10 : AOI22_X1 port map( A1 => A_ns(39), A2 => n751, B1 => A_s(39), B2 => 
                           n757, ZN => n760);
   U11 : INV_X1 port map( A => A_s(40), ZN => n759);
   U12 : INV_X1 port map( A => A_ns(40), ZN => n758);
   U13 : OAI221_X1 port map( B1 => n750, B2 => n753, C1 => n761, C2 => n755, A 
                           => n762, ZN => O_43_port);
   U14 : AOI22_X1 port map( A1 => A_ns(42), A2 => n763, B1 => A_s(42), B2 => 
                           n764, ZN => n762);
   U15 : INV_X1 port map( A => A_s(41), ZN => n755);
   U16 : INV_X1 port map( A => A_ns(41), ZN => n753);
   U17 : OAI221_X1 port map( B1 => n752, B2 => n765, C1 => n754, C2 => n766, A 
                           => n767, ZN => O_40_port);
   U18 : AOI22_X1 port map( A1 => A_ns(38), A2 => n751, B1 => A_s(38), B2 => 
                           n757, ZN => n767);
   U19 : INV_X1 port map( A => A_s(39), ZN => n766);
   U20 : INV_X1 port map( A => A_ns(39), ZN => n765);
   U21 : OAI221_X1 port map( B1 => n752, B2 => n768, C1 => n754, C2 => n769, A 
                           => n770, ZN => O_39_port);
   U22 : AOI22_X1 port map( A1 => A_ns(37), A2 => n751, B1 => A_s(37), B2 => 
                           n757, ZN => n770);
   U23 : INV_X1 port map( A => A_s(38), ZN => n769);
   U24 : INV_X1 port map( A => A_ns(38), ZN => n768);
   U25 : OAI221_X1 port map( B1 => n752, B2 => n771, C1 => n754, C2 => n772, A 
                           => n773, ZN => O_38_port);
   U26 : AOI22_X1 port map( A1 => A_ns(36), A2 => n751, B1 => A_s(36), B2 => 
                           n757, ZN => n773);
   U27 : INV_X1 port map( A => A_s(37), ZN => n772);
   U28 : INV_X1 port map( A => A_ns(37), ZN => n771);
   U29 : OAI221_X1 port map( B1 => n752, B2 => n774, C1 => n754, C2 => n775, A 
                           => n776, ZN => O_37_port);
   U30 : AOI22_X1 port map( A1 => A_ns(35), A2 => n751, B1 => A_s(35), B2 => 
                           n757, ZN => n776);
   U31 : INV_X1 port map( A => A_s(36), ZN => n775);
   U32 : INV_X1 port map( A => A_ns(36), ZN => n774);
   U33 : OAI221_X1 port map( B1 => n752, B2 => n777, C1 => n754, C2 => n778, A 
                           => n779, ZN => O_36_port);
   U34 : AOI22_X1 port map( A1 => A_ns(34), A2 => n751, B1 => A_s(34), B2 => 
                           n757, ZN => n779);
   U35 : INV_X1 port map( A => A_s(35), ZN => n778);
   U36 : INV_X1 port map( A => A_ns(35), ZN => n777);
   U37 : OAI221_X1 port map( B1 => n752, B2 => n780, C1 => n754, C2 => n781, A 
                           => n782, ZN => O_35_port);
   U38 : AOI22_X1 port map( A1 => A_ns(33), A2 => n751, B1 => A_s(33), B2 => 
                           n757, ZN => n782);
   U39 : INV_X1 port map( A => A_s(34), ZN => n781);
   U40 : INV_X1 port map( A => A_ns(34), ZN => n780);
   U41 : OAI221_X1 port map( B1 => n752, B2 => n783, C1 => n754, C2 => n784, A 
                           => n785, ZN => O_34_port);
   U42 : AOI22_X1 port map( A1 => A_ns(32), A2 => n751, B1 => A_s(32), B2 => 
                           n757, ZN => n785);
   U43 : INV_X1 port map( A => A_s(33), ZN => n784);
   U44 : INV_X1 port map( A => A_ns(33), ZN => n783);
   U45 : OAI221_X1 port map( B1 => n752, B2 => n786, C1 => n754, C2 => n787, A 
                           => n788, ZN => O_33_port);
   U46 : AOI22_X1 port map( A1 => A_ns(31), A2 => n751, B1 => A_s(31), B2 => 
                           n757, ZN => n788);
   U47 : INV_X1 port map( A => A_s(32), ZN => n787);
   U48 : INV_X1 port map( A => A_ns(32), ZN => n786);
   U49 : OAI221_X1 port map( B1 => n752, B2 => n789, C1 => n754, C2 => n790, A 
                           => n791, ZN => O_32_port);
   U50 : AOI22_X1 port map( A1 => A_ns(30), A2 => n751, B1 => A_s(30), B2 => 
                           n757, ZN => n791);
   U51 : INV_X1 port map( A => A_s(31), ZN => n790);
   U52 : INV_X1 port map( A => A_ns(31), ZN => n789);
   U53 : OAI221_X1 port map( B1 => n752, B2 => n792, C1 => n754, C2 => n793, A 
                           => n794, ZN => O_31_port);
   U54 : AOI22_X1 port map( A1 => A_ns(29), A2 => n751, B1 => A_s(29), B2 => 
                           n757, ZN => n794);
   U55 : INV_X1 port map( A => A_s(30), ZN => n793);
   U56 : INV_X1 port map( A => A_ns(30), ZN => n792);
   U57 : OAI221_X1 port map( B1 => n752, B2 => n795, C1 => n754, C2 => n796, A 
                           => n797, ZN => O_30_port);
   U58 : AOI22_X1 port map( A1 => A_ns(28), A2 => n751, B1 => A_s(28), B2 => 
                           n757, ZN => n797);
   U59 : INV_X1 port map( A => A_s(29), ZN => n796);
   U60 : INV_X1 port map( A => A_ns(29), ZN => n795);
   U61 : OAI221_X1 port map( B1 => n752, B2 => n798, C1 => n754, C2 => n799, A 
                           => n800, ZN => O_29_port);
   U62 : AOI22_X1 port map( A1 => A_ns(27), A2 => n751, B1 => A_s(27), B2 => 
                           n757, ZN => n800);
   U63 : INV_X1 port map( A => A_s(28), ZN => n799);
   U64 : INV_X1 port map( A => A_ns(28), ZN => n798);
   U65 : OAI221_X1 port map( B1 => n752, B2 => n801, C1 => n754, C2 => n802, A 
                           => n803, ZN => O_28_port);
   U66 : AOI22_X1 port map( A1 => A_ns(26), A2 => n751, B1 => A_s(26), B2 => 
                           n757, ZN => n803);
   U67 : INV_X1 port map( A => A_s(27), ZN => n802);
   U68 : INV_X1 port map( A => A_ns(27), ZN => n801);
   U69 : OAI221_X1 port map( B1 => n752, B2 => n804, C1 => n754, C2 => n805, A 
                           => n806, ZN => O_27_port);
   U70 : AOI22_X1 port map( A1 => A_ns(25), A2 => n751, B1 => A_s(25), B2 => 
                           n757, ZN => n806);
   U71 : INV_X1 port map( A => A_s(26), ZN => n805);
   U72 : INV_X1 port map( A => A_ns(26), ZN => n804);
   U73 : OAI221_X1 port map( B1 => n752, B2 => n807, C1 => n754, C2 => n808, A 
                           => n809, ZN => O_26_port);
   U74 : AOI22_X1 port map( A1 => A_ns(24), A2 => n751, B1 => A_s(24), B2 => 
                           n757, ZN => n809);
   U75 : INV_X1 port map( A => A_s(25), ZN => n808);
   U76 : INV_X1 port map( A => A_ns(25), ZN => n807);
   U77 : OAI221_X1 port map( B1 => n752, B2 => n810, C1 => n754, C2 => n811, A 
                           => n812, ZN => O_25_port);
   U78 : AOI22_X1 port map( A1 => A_ns(23), A2 => n751, B1 => A_s(23), B2 => 
                           n757, ZN => n812);
   U79 : INV_X1 port map( A => A_s(24), ZN => n811);
   U80 : INV_X1 port map( A => A_ns(24), ZN => n810);
   U81 : OAI221_X1 port map( B1 => n752, B2 => n813, C1 => n754, C2 => n814, A 
                           => n815, ZN => O_24_port);
   U82 : AOI22_X1 port map( A1 => A_ns(22), A2 => n751, B1 => A_s(22), B2 => 
                           n757, ZN => n815);
   U83 : INV_X1 port map( A => A_s(23), ZN => n814);
   U84 : INV_X1 port map( A => A_ns(23), ZN => n813);
   U85 : OAI221_X1 port map( B1 => n752, B2 => n816, C1 => n754, C2 => n817, A 
                           => n818, ZN => O_23_port);
   U86 : AOI22_X1 port map( A1 => A_ns(21), A2 => n751, B1 => A_s(21), B2 => 
                           n757, ZN => n818);
   U87 : INV_X1 port map( A => A_s(22), ZN => n817);
   U88 : INV_X1 port map( A => A_ns(22), ZN => n816);
   U89 : OAI221_X1 port map( B1 => n752, B2 => n819, C1 => n754, C2 => n820, A 
                           => n821, ZN => O_22_port);
   U90 : AOI22_X1 port map( A1 => A_ns(20), A2 => n751, B1 => A_s(20), B2 => 
                           n757, ZN => n821);
   U91 : INV_X1 port map( A => A_s(21), ZN => n820);
   U92 : INV_X1 port map( A => A_ns(21), ZN => n819);
   U93 : OAI221_X1 port map( B1 => n752, B2 => n822, C1 => n754, C2 => n823, A 
                           => n824, ZN => O_21_port);
   U94 : AOI22_X1 port map( A1 => A_ns(19), A2 => n751, B1 => A_s(19), B2 => 
                           n757, ZN => n824);
   U95 : INV_X1 port map( A => A_s(20), ZN => n823);
   U96 : INV_X1 port map( A => A_ns(20), ZN => n822);
   U97 : OAI221_X1 port map( B1 => n752, B2 => n825, C1 => n754, C2 => n826, A 
                           => n827, ZN => O_20_port);
   U98 : AOI22_X1 port map( A1 => A_ns(18), A2 => n751, B1 => A_s(18), B2 => 
                           n757, ZN => n827);
   U99 : INV_X1 port map( A => A_s(19), ZN => n826);
   U100 : INV_X1 port map( A => A_ns(19), ZN => n825);
   U101 : OAI221_X1 port map( B1 => n752, B2 => n828, C1 => n754, C2 => n829, A
                           => n830, ZN => O_19_port);
   U102 : AOI22_X1 port map( A1 => A_ns(17), A2 => n751, B1 => A_s(17), B2 => 
                           n757, ZN => n830);
   U103 : INV_X1 port map( A => A_s(18), ZN => n829);
   U104 : INV_X1 port map( A => A_ns(18), ZN => n828);
   U105 : OAI221_X1 port map( B1 => n752, B2 => n831, C1 => n754, C2 => n832, A
                           => n833, ZN => O_18_port);
   U106 : AOI22_X1 port map( A1 => A_ns(16), A2 => n751, B1 => A_s(16), B2 => 
                           n757, ZN => n833);
   U107 : INV_X1 port map( A => A_s(17), ZN => n832);
   U108 : INV_X1 port map( A => A_ns(17), ZN => n831);
   U109 : OAI221_X1 port map( B1 => n752, B2 => n834, C1 => n754, C2 => n835, A
                           => n836, ZN => O_17_port);
   U110 : AOI22_X1 port map( A1 => A_ns(15), A2 => n751, B1 => A_s(15), B2 => 
                           n757, ZN => n836);
   U111 : INV_X1 port map( A => A_s(16), ZN => n835);
   U112 : INV_X1 port map( A => A_ns(16), ZN => n834);
   U113 : OAI221_X1 port map( B1 => n752, B2 => n837, C1 => n754, C2 => n838, A
                           => n839, ZN => O_16_port);
   U114 : AOI22_X1 port map( A1 => A_ns(14), A2 => n751, B1 => A_s(14), B2 => 
                           n757, ZN => n839);
   U115 : INV_X1 port map( A => A_s(15), ZN => n838);
   U116 : INV_X1 port map( A => A_ns(15), ZN => n837);
   U117 : OAI221_X1 port map( B1 => n752, B2 => n840, C1 => n754, C2 => n841, A
                           => n842, ZN => O_15_port);
   U118 : AOI22_X1 port map( A1 => A_ns(13), A2 => n751, B1 => A_s(13), B2 => 
                           n757, ZN => n842);
   U119 : INV_X1 port map( A => A_s(14), ZN => n841);
   U120 : INV_X1 port map( A => A_ns(14), ZN => n840);
   U121 : OAI221_X1 port map( B1 => n752, B2 => n843, C1 => n754, C2 => n844, A
                           => n845, ZN => O_14_port);
   U122 : AOI22_X1 port map( A1 => A_ns(12), A2 => n751, B1 => A_s(12), B2 => 
                           n757, ZN => n845);
   U123 : INV_X1 port map( A => A_s(13), ZN => n844);
   U124 : INV_X1 port map( A => A_ns(13), ZN => n843);
   U125 : OAI221_X1 port map( B1 => n752, B2 => n846, C1 => n754, C2 => n847, A
                           => n848, ZN => O_13_port);
   U126 : AOI22_X1 port map( A1 => A_ns(11), A2 => n751, B1 => A_s(11), B2 => 
                           n757, ZN => n848);
   U127 : INV_X1 port map( A => A_s(12), ZN => n847);
   U128 : INV_X1 port map( A => A_ns(12), ZN => n846);
   U129 : OAI221_X1 port map( B1 => n752, B2 => n849, C1 => n754, C2 => n850, A
                           => n851, ZN => O_12_port);
   U130 : AOI22_X1 port map( A1 => A_ns(10), A2 => n751, B1 => A_s(10), B2 => 
                           n757, ZN => n851);
   U131 : INV_X1 port map( A => A_s(11), ZN => n850);
   U132 : INV_X1 port map( A => A_ns(11), ZN => n849);
   U133 : OAI221_X1 port map( B1 => n752, B2 => n852, C1 => n754, C2 => n853, A
                           => n854, ZN => O_11_port);
   U134 : AOI22_X1 port map( A1 => A_ns(9), A2 => n751, B1 => A_s(9), B2 => 
                           n757, ZN => n854);
   U135 : INV_X1 port map( A => A_s(10), ZN => n853);
   U136 : INV_X1 port map( A => A_ns(10), ZN => n852);
   U137 : INV_X1 port map( A => n855, ZN => O_1_port);
   U138 : AOI22_X1 port map( A1 => n764, A2 => A_s(0), B1 => n763, B2 => 
                           A_ns(0), ZN => n855);
   U139 : OAI221_X1 port map( B1 => n752, B2 => n856, C1 => n754, C2 => n857, A
                           => n858, ZN => O_2_port);
   U140 : AOI22_X1 port map( A1 => A_ns(0), A2 => n751, B1 => A_s(0), B2 => 
                           n757, ZN => n858);
   U141 : INV_X1 port map( A => n859, ZN => O_3_port);
   U142 : AOI221_X1 port map( B1 => n763, B2 => A_ns(2), C1 => n764, C2 => 
                           A_s(2), A => n860, ZN => n859);
   U143 : OAI22_X1 port map( A1 => n856, A2 => n750, B1 => n857, B2 => n761, ZN
                           => n860);
   U144 : INV_X1 port map( A => A_s(1), ZN => n857);
   U145 : INV_X1 port map( A => A_ns(1), ZN => n856);
   U146 : OAI221_X1 port map( B1 => n752, B2 => n861, C1 => n754, C2 => n862, A
                           => n863, ZN => O_4_port);
   U147 : AOI22_X1 port map( A1 => A_ns(2), A2 => n751, B1 => A_s(2), B2 => 
                           n757, ZN => n863);
   U148 : INV_X1 port map( A => n864, ZN => O_5_port);
   U149 : AOI221_X1 port map( B1 => n763, B2 => A_ns(4), C1 => n764, C2 => 
                           A_s(4), A => n865, ZN => n864);
   U150 : OAI22_X1 port map( A1 => n861, A2 => n750, B1 => n862, B2 => n761, ZN
                           => n865);
   U151 : INV_X1 port map( A => A_s(3), ZN => n862);
   U152 : INV_X1 port map( A => A_ns(3), ZN => n861);
   U153 : OAI221_X1 port map( B1 => n752, B2 => n866, C1 => n754, C2 => n867, A
                           => n868, ZN => O_6_port);
   U154 : AOI22_X1 port map( A1 => A_ns(4), A2 => n751, B1 => A_s(4), B2 => 
                           n757, ZN => n868);
   U155 : INV_X1 port map( A => n869, ZN => O_7_port);
   U156 : AOI221_X1 port map( B1 => n763, B2 => A_ns(6), C1 => n764, C2 => 
                           A_s(6), A => n870, ZN => n869);
   U157 : OAI22_X1 port map( A1 => n866, A2 => n750, B1 => n867, B2 => n761, ZN
                           => n870);
   U158 : INV_X1 port map( A => A_s(5), ZN => n867);
   U159 : INV_X1 port map( A => A_ns(5), ZN => n866);
   U160 : OAI221_X1 port map( B1 => n752, B2 => n871, C1 => n754, C2 => n872, A
                           => n873, ZN => O_8_port);
   U161 : AOI22_X1 port map( A1 => A_ns(6), A2 => n751, B1 => A_s(6), B2 => 
                           n757, ZN => n873);
   U162 : INV_X1 port map( A => n874, ZN => O_9_port);
   U163 : AOI221_X1 port map( B1 => n763, B2 => A_ns(8), C1 => n764, C2 => 
                           A_s(8), A => n875, ZN => n874);
   U164 : OAI22_X1 port map( A1 => n871, A2 => n750, B1 => n872, B2 => n761, ZN
                           => n875);
   U165 : INV_X1 port map( A => A_s(7), ZN => n872);
   U166 : INV_X1 port map( A => A_ns(7), ZN => n871);
   U167 : INV_X1 port map( A => n754, ZN => n764);
   U168 : INV_X1 port map( A => n752, ZN => n763);
   U169 : OAI221_X1 port map( B1 => n752, B2 => n876, C1 => n754, C2 => n877, A
                           => n878, ZN => O_10_port);
   U170 : AOI22_X1 port map( A1 => A_ns(8), A2 => n751, B1 => A_s(8), B2 => 
                           n757, ZN => n878);
   U171 : NAND3_X1 port map( A1 => B(10), A2 => n879, A3 => B(9), ZN => n761);
   U172 : INV_X1 port map( A => A_s(9), ZN => n877);
   U173 : INV_X1 port map( A => A_ns(9), ZN => n876);
   U174 : INV_X1 port map( A => B(11), ZN => n879);
   U175 : XOR2_X1 port map( A => B(9), B => B(10), Z => n880);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT42_i8 is

   port( A_s, A_ns, B : in std_logic_vector (41 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (41 downto 0));

end BOOTHENC_NBIT42_i8;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT42_i8 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, n712, n713, n714, n715, n716, n717, n718, n719, n720, 
      n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, 
      n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, 
      n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, 
      n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, 
      n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, 
      n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, 
      n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, 
      n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, 
      n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, 
      n829, n830, n831, n832, n833, n834, n835, n836, n837, O_40_port, 
      O_39_port, O_41_port, O_38_port, O_37_port, O_36_port, O_35_port, 
      O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, 
      O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, 
      O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, 
      O_16_port, O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, 
      O_10_port, O_9_port, O_1_port, O_2_port, O_3_port, O_4_port, O_5_port, 
      O_6_port, O_7_port, O_8_port : std_logic;

begin
   O <= ( O_41_port, O_40_port, O_39_port, O_38_port, O_37_port, O_36_port, 
      O_35_port, O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, 
      O_29_port, O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, 
      O_23_port, O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, 
      O_17_port, O_16_port, O_15_port, O_14_port, O_13_port, O_12_port, 
      O_11_port, O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, 
      O_4_port, O_3_port, O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(39), A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), 
      A_s(32), A_s(31), A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), 
      A_s(24), A_s(23), A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), 
      A_s(16), A_s(15), A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), 
      A_s(8), A_s(7), A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), 
      X_Logic0_port, X_Logic0_port );
   A_nso <= ( A_ns(39), A_ns(38), A_ns(37), A_ns(36), A_ns(35), A_ns(34), 
      A_ns(33), A_ns(32), A_ns(31), A_ns(30), A_ns(29), A_ns(28), A_ns(27), 
      A_ns(26), A_ns(25), A_ns(24), A_ns(23), A_ns(22), A_ns(21), A_ns(20), 
      A_ns(19), A_ns(18), A_ns(17), A_ns(16), A_ns(15), A_ns(14), A_ns(13), 
      A_ns(12), A_ns(11), A_ns(10), A_ns(9), A_ns(8), A_ns(7), A_ns(6), A_ns(5)
      , A_ns(4), A_ns(3), A_ns(2), A_ns(1), A_ns(0), X_Logic0_port, 
      X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : OR3_X1 port map( A1 => B(7), A2 => B(8), A3 => n836, ZN => n712);
   U3 : INV_X2 port map( A => n712, ZN => n713);
   U4 : NAND2_X2 port map( A1 => n837, A2 => n716, ZN => n714);
   U5 : INV_X2 port map( A => n723, ZN => n719);
   U6 : NAND2_X2 port map( A1 => n837, A2 => n836, ZN => n716);
   U7 : OAI221_X1 port map( B1 => n714, B2 => n715, C1 => n716, C2 => n717, A 
                           => n718, ZN => O_40_port);
   U8 : AOI22_X1 port map( A1 => A_ns(38), A2 => n713, B1 => A_s(38), B2 => 
                           n719, ZN => n718);
   U9 : OAI221_X1 port map( B1 => n720, B2 => n714, C1 => n721, C2 => n716, A 
                           => n722, ZN => O_39_port);
   U10 : AOI22_X1 port map( A1 => A_ns(37), A2 => n713, B1 => A_s(37), B2 => 
                           n719, ZN => n722);
   U11 : INV_X1 port map( A => A_s(38), ZN => n721);
   U12 : INV_X1 port map( A => A_ns(38), ZN => n720);
   U13 : OAI221_X1 port map( B1 => n712, B2 => n715, C1 => n723, C2 => n717, A 
                           => n724, ZN => O_41_port);
   U14 : AOI22_X1 port map( A1 => A_ns(40), A2 => n725, B1 => A_s(40), B2 => 
                           n726, ZN => n724);
   U15 : INV_X1 port map( A => A_s(39), ZN => n717);
   U16 : INV_X1 port map( A => A_ns(39), ZN => n715);
   U17 : OAI221_X1 port map( B1 => n714, B2 => n727, C1 => n716, C2 => n728, A 
                           => n729, ZN => O_38_port);
   U18 : AOI22_X1 port map( A1 => A_ns(36), A2 => n713, B1 => A_s(36), B2 => 
                           n719, ZN => n729);
   U19 : INV_X1 port map( A => A_s(37), ZN => n728);
   U20 : INV_X1 port map( A => A_ns(37), ZN => n727);
   U21 : OAI221_X1 port map( B1 => n714, B2 => n730, C1 => n716, C2 => n731, A 
                           => n732, ZN => O_37_port);
   U22 : AOI22_X1 port map( A1 => A_ns(35), A2 => n713, B1 => A_s(35), B2 => 
                           n719, ZN => n732);
   U23 : INV_X1 port map( A => A_s(36), ZN => n731);
   U24 : INV_X1 port map( A => A_ns(36), ZN => n730);
   U25 : OAI221_X1 port map( B1 => n714, B2 => n733, C1 => n716, C2 => n734, A 
                           => n735, ZN => O_36_port);
   U26 : AOI22_X1 port map( A1 => A_ns(34), A2 => n713, B1 => A_s(34), B2 => 
                           n719, ZN => n735);
   U27 : INV_X1 port map( A => A_s(35), ZN => n734);
   U28 : INV_X1 port map( A => A_ns(35), ZN => n733);
   U29 : OAI221_X1 port map( B1 => n714, B2 => n736, C1 => n716, C2 => n737, A 
                           => n738, ZN => O_35_port);
   U30 : AOI22_X1 port map( A1 => A_ns(33), A2 => n713, B1 => A_s(33), B2 => 
                           n719, ZN => n738);
   U31 : INV_X1 port map( A => A_s(34), ZN => n737);
   U32 : INV_X1 port map( A => A_ns(34), ZN => n736);
   U33 : OAI221_X1 port map( B1 => n714, B2 => n739, C1 => n716, C2 => n740, A 
                           => n741, ZN => O_34_port);
   U34 : AOI22_X1 port map( A1 => A_ns(32), A2 => n713, B1 => A_s(32), B2 => 
                           n719, ZN => n741);
   U35 : INV_X1 port map( A => A_s(33), ZN => n740);
   U36 : INV_X1 port map( A => A_ns(33), ZN => n739);
   U37 : OAI221_X1 port map( B1 => n714, B2 => n742, C1 => n716, C2 => n743, A 
                           => n744, ZN => O_33_port);
   U38 : AOI22_X1 port map( A1 => A_ns(31), A2 => n713, B1 => A_s(31), B2 => 
                           n719, ZN => n744);
   U39 : INV_X1 port map( A => A_s(32), ZN => n743);
   U40 : INV_X1 port map( A => A_ns(32), ZN => n742);
   U41 : OAI221_X1 port map( B1 => n714, B2 => n745, C1 => n716, C2 => n746, A 
                           => n747, ZN => O_32_port);
   U42 : AOI22_X1 port map( A1 => A_ns(30), A2 => n713, B1 => A_s(30), B2 => 
                           n719, ZN => n747);
   U43 : INV_X1 port map( A => A_s(31), ZN => n746);
   U44 : INV_X1 port map( A => A_ns(31), ZN => n745);
   U45 : OAI221_X1 port map( B1 => n714, B2 => n748, C1 => n716, C2 => n749, A 
                           => n750, ZN => O_31_port);
   U46 : AOI22_X1 port map( A1 => A_ns(29), A2 => n713, B1 => A_s(29), B2 => 
                           n719, ZN => n750);
   U47 : INV_X1 port map( A => A_s(30), ZN => n749);
   U48 : INV_X1 port map( A => A_ns(30), ZN => n748);
   U49 : OAI221_X1 port map( B1 => n714, B2 => n751, C1 => n716, C2 => n752, A 
                           => n753, ZN => O_30_port);
   U50 : AOI22_X1 port map( A1 => A_ns(28), A2 => n713, B1 => A_s(28), B2 => 
                           n719, ZN => n753);
   U51 : INV_X1 port map( A => A_s(29), ZN => n752);
   U52 : INV_X1 port map( A => A_ns(29), ZN => n751);
   U53 : OAI221_X1 port map( B1 => n714, B2 => n754, C1 => n716, C2 => n755, A 
                           => n756, ZN => O_29_port);
   U54 : AOI22_X1 port map( A1 => A_ns(27), A2 => n713, B1 => A_s(27), B2 => 
                           n719, ZN => n756);
   U55 : INV_X1 port map( A => A_s(28), ZN => n755);
   U56 : INV_X1 port map( A => A_ns(28), ZN => n754);
   U57 : OAI221_X1 port map( B1 => n714, B2 => n757, C1 => n716, C2 => n758, A 
                           => n759, ZN => O_28_port);
   U58 : AOI22_X1 port map( A1 => A_ns(26), A2 => n713, B1 => A_s(26), B2 => 
                           n719, ZN => n759);
   U59 : INV_X1 port map( A => A_s(27), ZN => n758);
   U60 : INV_X1 port map( A => A_ns(27), ZN => n757);
   U61 : OAI221_X1 port map( B1 => n714, B2 => n760, C1 => n716, C2 => n761, A 
                           => n762, ZN => O_27_port);
   U62 : AOI22_X1 port map( A1 => A_ns(25), A2 => n713, B1 => A_s(25), B2 => 
                           n719, ZN => n762);
   U63 : INV_X1 port map( A => A_s(26), ZN => n761);
   U64 : INV_X1 port map( A => A_ns(26), ZN => n760);
   U65 : OAI221_X1 port map( B1 => n714, B2 => n763, C1 => n716, C2 => n764, A 
                           => n765, ZN => O_26_port);
   U66 : AOI22_X1 port map( A1 => A_ns(24), A2 => n713, B1 => A_s(24), B2 => 
                           n719, ZN => n765);
   U67 : INV_X1 port map( A => A_s(25), ZN => n764);
   U68 : INV_X1 port map( A => A_ns(25), ZN => n763);
   U69 : OAI221_X1 port map( B1 => n714, B2 => n766, C1 => n716, C2 => n767, A 
                           => n768, ZN => O_25_port);
   U70 : AOI22_X1 port map( A1 => A_ns(23), A2 => n713, B1 => A_s(23), B2 => 
                           n719, ZN => n768);
   U71 : INV_X1 port map( A => A_s(24), ZN => n767);
   U72 : INV_X1 port map( A => A_ns(24), ZN => n766);
   U73 : OAI221_X1 port map( B1 => n714, B2 => n769, C1 => n716, C2 => n770, A 
                           => n771, ZN => O_24_port);
   U74 : AOI22_X1 port map( A1 => A_ns(22), A2 => n713, B1 => A_s(22), B2 => 
                           n719, ZN => n771);
   U75 : INV_X1 port map( A => A_s(23), ZN => n770);
   U76 : INV_X1 port map( A => A_ns(23), ZN => n769);
   U77 : OAI221_X1 port map( B1 => n714, B2 => n772, C1 => n716, C2 => n773, A 
                           => n774, ZN => O_23_port);
   U78 : AOI22_X1 port map( A1 => A_ns(21), A2 => n713, B1 => A_s(21), B2 => 
                           n719, ZN => n774);
   U79 : INV_X1 port map( A => A_s(22), ZN => n773);
   U80 : INV_X1 port map( A => A_ns(22), ZN => n772);
   U81 : OAI221_X1 port map( B1 => n714, B2 => n775, C1 => n716, C2 => n776, A 
                           => n777, ZN => O_22_port);
   U82 : AOI22_X1 port map( A1 => A_ns(20), A2 => n713, B1 => A_s(20), B2 => 
                           n719, ZN => n777);
   U83 : INV_X1 port map( A => A_s(21), ZN => n776);
   U84 : INV_X1 port map( A => A_ns(21), ZN => n775);
   U85 : OAI221_X1 port map( B1 => n714, B2 => n778, C1 => n716, C2 => n779, A 
                           => n780, ZN => O_21_port);
   U86 : AOI22_X1 port map( A1 => A_ns(19), A2 => n713, B1 => A_s(19), B2 => 
                           n719, ZN => n780);
   U87 : INV_X1 port map( A => A_s(20), ZN => n779);
   U88 : INV_X1 port map( A => A_ns(20), ZN => n778);
   U89 : OAI221_X1 port map( B1 => n714, B2 => n781, C1 => n716, C2 => n782, A 
                           => n783, ZN => O_20_port);
   U90 : AOI22_X1 port map( A1 => A_ns(18), A2 => n713, B1 => A_s(18), B2 => 
                           n719, ZN => n783);
   U91 : INV_X1 port map( A => A_s(19), ZN => n782);
   U92 : INV_X1 port map( A => A_ns(19), ZN => n781);
   U93 : OAI221_X1 port map( B1 => n714, B2 => n784, C1 => n716, C2 => n785, A 
                           => n786, ZN => O_19_port);
   U94 : AOI22_X1 port map( A1 => A_ns(17), A2 => n713, B1 => A_s(17), B2 => 
                           n719, ZN => n786);
   U95 : INV_X1 port map( A => A_s(18), ZN => n785);
   U96 : INV_X1 port map( A => A_ns(18), ZN => n784);
   U97 : OAI221_X1 port map( B1 => n714, B2 => n787, C1 => n716, C2 => n788, A 
                           => n789, ZN => O_18_port);
   U98 : AOI22_X1 port map( A1 => A_ns(16), A2 => n713, B1 => A_s(16), B2 => 
                           n719, ZN => n789);
   U99 : INV_X1 port map( A => A_s(17), ZN => n788);
   U100 : INV_X1 port map( A => A_ns(17), ZN => n787);
   U101 : OAI221_X1 port map( B1 => n714, B2 => n790, C1 => n716, C2 => n791, A
                           => n792, ZN => O_17_port);
   U102 : AOI22_X1 port map( A1 => A_ns(15), A2 => n713, B1 => A_s(15), B2 => 
                           n719, ZN => n792);
   U103 : INV_X1 port map( A => A_s(16), ZN => n791);
   U104 : INV_X1 port map( A => A_ns(16), ZN => n790);
   U105 : OAI221_X1 port map( B1 => n714, B2 => n793, C1 => n716, C2 => n794, A
                           => n795, ZN => O_16_port);
   U106 : AOI22_X1 port map( A1 => A_ns(14), A2 => n713, B1 => A_s(14), B2 => 
                           n719, ZN => n795);
   U107 : INV_X1 port map( A => A_s(15), ZN => n794);
   U108 : INV_X1 port map( A => A_ns(15), ZN => n793);
   U109 : OAI221_X1 port map( B1 => n714, B2 => n796, C1 => n716, C2 => n797, A
                           => n798, ZN => O_15_port);
   U110 : AOI22_X1 port map( A1 => A_ns(13), A2 => n713, B1 => A_s(13), B2 => 
                           n719, ZN => n798);
   U111 : INV_X1 port map( A => A_s(14), ZN => n797);
   U112 : INV_X1 port map( A => A_ns(14), ZN => n796);
   U113 : OAI221_X1 port map( B1 => n714, B2 => n799, C1 => n716, C2 => n800, A
                           => n801, ZN => O_14_port);
   U114 : AOI22_X1 port map( A1 => A_ns(12), A2 => n713, B1 => A_s(12), B2 => 
                           n719, ZN => n801);
   U115 : INV_X1 port map( A => A_s(13), ZN => n800);
   U116 : INV_X1 port map( A => A_ns(13), ZN => n799);
   U117 : OAI221_X1 port map( B1 => n714, B2 => n802, C1 => n716, C2 => n803, A
                           => n804, ZN => O_13_port);
   U118 : AOI22_X1 port map( A1 => A_ns(11), A2 => n713, B1 => A_s(11), B2 => 
                           n719, ZN => n804);
   U119 : INV_X1 port map( A => A_s(12), ZN => n803);
   U120 : INV_X1 port map( A => A_ns(12), ZN => n802);
   U121 : OAI221_X1 port map( B1 => n714, B2 => n805, C1 => n716, C2 => n806, A
                           => n807, ZN => O_12_port);
   U122 : AOI22_X1 port map( A1 => A_ns(10), A2 => n713, B1 => A_s(10), B2 => 
                           n719, ZN => n807);
   U123 : INV_X1 port map( A => A_s(11), ZN => n806);
   U124 : INV_X1 port map( A => A_ns(11), ZN => n805);
   U125 : OAI221_X1 port map( B1 => n714, B2 => n808, C1 => n716, C2 => n809, A
                           => n810, ZN => O_11_port);
   U126 : AOI22_X1 port map( A1 => A_ns(9), A2 => n713, B1 => A_s(9), B2 => 
                           n719, ZN => n810);
   U127 : INV_X1 port map( A => A_s(10), ZN => n809);
   U128 : INV_X1 port map( A => A_ns(10), ZN => n808);
   U129 : OAI221_X1 port map( B1 => n714, B2 => n811, C1 => n716, C2 => n812, A
                           => n813, ZN => O_10_port);
   U130 : AOI22_X1 port map( A1 => A_ns(8), A2 => n713, B1 => A_s(8), B2 => 
                           n719, ZN => n813);
   U131 : INV_X1 port map( A => A_s(9), ZN => n812);
   U132 : INV_X1 port map( A => A_ns(9), ZN => n811);
   U133 : OAI221_X1 port map( B1 => n714, B2 => n814, C1 => n716, C2 => n815, A
                           => n816, ZN => O_9_port);
   U134 : AOI22_X1 port map( A1 => A_ns(7), A2 => n713, B1 => A_s(7), B2 => 
                           n719, ZN => n816);
   U135 : INV_X1 port map( A => A_s(8), ZN => n815);
   U136 : INV_X1 port map( A => A_ns(8), ZN => n814);
   U137 : INV_X1 port map( A => n817, ZN => O_1_port);
   U138 : AOI22_X1 port map( A1 => n726, A2 => A_s(0), B1 => n725, B2 => 
                           A_ns(0), ZN => n817);
   U139 : OAI221_X1 port map( B1 => n714, B2 => n818, C1 => n716, C2 => n819, A
                           => n820, ZN => O_2_port);
   U140 : AOI22_X1 port map( A1 => A_ns(0), A2 => n713, B1 => A_s(0), B2 => 
                           n719, ZN => n820);
   U141 : INV_X1 port map( A => n821, ZN => O_3_port);
   U142 : AOI221_X1 port map( B1 => n725, B2 => A_ns(2), C1 => n726, C2 => 
                           A_s(2), A => n822, ZN => n821);
   U143 : OAI22_X1 port map( A1 => n818, A2 => n712, B1 => n819, B2 => n723, ZN
                           => n822);
   U144 : INV_X1 port map( A => A_s(1), ZN => n819);
   U145 : INV_X1 port map( A => A_ns(1), ZN => n818);
   U146 : OAI221_X1 port map( B1 => n714, B2 => n823, C1 => n716, C2 => n824, A
                           => n825, ZN => O_4_port);
   U147 : AOI22_X1 port map( A1 => A_ns(2), A2 => n713, B1 => A_s(2), B2 => 
                           n719, ZN => n825);
   U148 : INV_X1 port map( A => n826, ZN => O_5_port);
   U149 : AOI221_X1 port map( B1 => n725, B2 => A_ns(4), C1 => n726, C2 => 
                           A_s(4), A => n827, ZN => n826);
   U150 : OAI22_X1 port map( A1 => n823, A2 => n712, B1 => n824, B2 => n723, ZN
                           => n827);
   U151 : INV_X1 port map( A => A_s(3), ZN => n824);
   U152 : INV_X1 port map( A => A_ns(3), ZN => n823);
   U153 : OAI221_X1 port map( B1 => n714, B2 => n828, C1 => n716, C2 => n829, A
                           => n830, ZN => O_6_port);
   U154 : AOI22_X1 port map( A1 => A_ns(4), A2 => n713, B1 => A_s(4), B2 => 
                           n719, ZN => n830);
   U155 : INV_X1 port map( A => n831, ZN => O_7_port);
   U156 : AOI221_X1 port map( B1 => n725, B2 => A_ns(6), C1 => n726, C2 => 
                           A_s(6), A => n832, ZN => n831);
   U157 : OAI22_X1 port map( A1 => n828, A2 => n712, B1 => n829, B2 => n723, ZN
                           => n832);
   U158 : INV_X1 port map( A => A_s(5), ZN => n829);
   U159 : INV_X1 port map( A => A_ns(5), ZN => n828);
   U160 : INV_X1 port map( A => n716, ZN => n726);
   U161 : INV_X1 port map( A => n714, ZN => n725);
   U162 : OAI221_X1 port map( B1 => n714, B2 => n833, C1 => n716, C2 => n834, A
                           => n835, ZN => O_8_port);
   U163 : AOI22_X1 port map( A1 => A_ns(6), A2 => n713, B1 => A_s(6), B2 => 
                           n719, ZN => n835);
   U164 : NAND3_X1 port map( A1 => B(7), A2 => n836, A3 => B(8), ZN => n723);
   U165 : INV_X1 port map( A => A_s(7), ZN => n834);
   U166 : INV_X1 port map( A => A_ns(7), ZN => n833);
   U167 : INV_X1 port map( A => B(9), ZN => n836);
   U168 : XOR2_X1 port map( A => B(8), B => B(7), Z => n837);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT40_i6 is

   port( A_s, A_ns, B : in std_logic_vector (39 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (39 downto 0));

end BOOTHENC_NBIT40_i6;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT40_i6 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, n671, n672, n673, n674, n675, n676, n677, n678, n679, 
      n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, 
      n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, 
      n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, 
      n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, 
      n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, 
      n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, 
      n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, 
      n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, 
      n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, 
      n788, n789, n790, n791, n792, O_38_port, O_37_port, O_39_port, O_36_port,
      O_35_port, O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, 
      O_29_port, O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, 
      O_23_port, O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, 
      O_17_port, O_16_port, O_15_port, O_14_port, O_13_port, O_12_port, 
      O_11_port, O_10_port, O_9_port, O_8_port, O_7_port, O_1_port, O_2_port, 
      O_3_port, O_4_port, O_5_port, O_6_port : std_logic;

begin
   O <= ( O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, 
      O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, 
      O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, 
      O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, O_16_port, 
      O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, O_10_port, 
      O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, O_3_port, 
      O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   A_nso <= ( A_ns(37), A_ns(36), A_ns(35), A_ns(34), A_ns(33), A_ns(32), 
      A_ns(31), A_ns(30), A_ns(29), A_ns(28), A_ns(27), A_ns(26), A_ns(25), 
      A_ns(24), A_ns(23), A_ns(22), A_ns(21), A_ns(20), A_ns(19), A_ns(18), 
      A_ns(17), A_ns(16), A_ns(15), A_ns(14), A_ns(13), A_ns(12), A_ns(11), 
      A_ns(10), A_ns(9), A_ns(8), A_ns(7), A_ns(6), A_ns(5), A_ns(4), A_ns(3), 
      A_ns(2), A_ns(1), A_ns(0), X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : NAND2_X2 port map( A1 => n792, A2 => n791, ZN => n674);
   U3 : INV_X2 port map( A => n683, ZN => n678);
   U4 : NAND2_X2 port map( A1 => n792, A2 => n674, ZN => n672);
   U5 : INV_X2 port map( A => n682, ZN => n671);
   U6 : OAI221_X1 port map( B1 => n672, B2 => n673, C1 => n674, C2 => n675, A 
                           => n676, ZN => O_38_port);
   U7 : AOI22_X1 port map( A1 => A_ns(36), A2 => n671, B1 => A_s(36), B2 => 
                           n678, ZN => n676);
   U8 : OAI221_X1 port map( B1 => n679, B2 => n672, C1 => n680, C2 => n674, A 
                           => n681, ZN => O_37_port);
   U9 : AOI22_X1 port map( A1 => A_ns(35), A2 => n671, B1 => A_s(35), B2 => 
                           n678, ZN => n681);
   U10 : INV_X1 port map( A => A_s(36), ZN => n680);
   U11 : INV_X1 port map( A => A_ns(36), ZN => n679);
   U12 : OAI221_X1 port map( B1 => n682, B2 => n673, C1 => n683, C2 => n675, A 
                           => n684, ZN => O_39_port);
   U13 : AOI22_X1 port map( A1 => A_ns(38), A2 => n685, B1 => A_s(38), B2 => 
                           n686, ZN => n684);
   U14 : INV_X1 port map( A => A_s(37), ZN => n675);
   U15 : INV_X1 port map( A => A_ns(37), ZN => n673);
   U16 : OAI221_X1 port map( B1 => n672, B2 => n687, C1 => n674, C2 => n688, A 
                           => n689, ZN => O_36_port);
   U17 : AOI22_X1 port map( A1 => A_ns(34), A2 => n671, B1 => A_s(34), B2 => 
                           n678, ZN => n689);
   U18 : INV_X1 port map( A => A_s(35), ZN => n688);
   U19 : INV_X1 port map( A => A_ns(35), ZN => n687);
   U20 : OAI221_X1 port map( B1 => n672, B2 => n690, C1 => n674, C2 => n691, A 
                           => n692, ZN => O_35_port);
   U21 : AOI22_X1 port map( A1 => A_ns(33), A2 => n671, B1 => A_s(33), B2 => 
                           n678, ZN => n692);
   U22 : INV_X1 port map( A => A_s(34), ZN => n691);
   U23 : INV_X1 port map( A => A_ns(34), ZN => n690);
   U24 : OAI221_X1 port map( B1 => n672, B2 => n693, C1 => n674, C2 => n694, A 
                           => n695, ZN => O_34_port);
   U25 : AOI22_X1 port map( A1 => A_ns(32), A2 => n671, B1 => A_s(32), B2 => 
                           n678, ZN => n695);
   U26 : INV_X1 port map( A => A_s(33), ZN => n694);
   U27 : INV_X1 port map( A => A_ns(33), ZN => n693);
   U28 : OAI221_X1 port map( B1 => n672, B2 => n696, C1 => n674, C2 => n697, A 
                           => n698, ZN => O_33_port);
   U29 : AOI22_X1 port map( A1 => A_ns(31), A2 => n671, B1 => A_s(31), B2 => 
                           n678, ZN => n698);
   U30 : INV_X1 port map( A => A_s(32), ZN => n697);
   U31 : INV_X1 port map( A => A_ns(32), ZN => n696);
   U32 : OAI221_X1 port map( B1 => n672, B2 => n699, C1 => n674, C2 => n700, A 
                           => n701, ZN => O_32_port);
   U33 : AOI22_X1 port map( A1 => A_ns(30), A2 => n671, B1 => A_s(30), B2 => 
                           n678, ZN => n701);
   U34 : INV_X1 port map( A => A_s(31), ZN => n700);
   U35 : INV_X1 port map( A => A_ns(31), ZN => n699);
   U36 : OAI221_X1 port map( B1 => n672, B2 => n702, C1 => n674, C2 => n703, A 
                           => n704, ZN => O_31_port);
   U37 : AOI22_X1 port map( A1 => A_ns(29), A2 => n671, B1 => A_s(29), B2 => 
                           n678, ZN => n704);
   U38 : INV_X1 port map( A => A_s(30), ZN => n703);
   U39 : INV_X1 port map( A => A_ns(30), ZN => n702);
   U40 : OAI221_X1 port map( B1 => n672, B2 => n705, C1 => n674, C2 => n706, A 
                           => n707, ZN => O_30_port);
   U41 : AOI22_X1 port map( A1 => A_ns(28), A2 => n671, B1 => A_s(28), B2 => 
                           n678, ZN => n707);
   U42 : INV_X1 port map( A => A_s(29), ZN => n706);
   U43 : INV_X1 port map( A => A_ns(29), ZN => n705);
   U44 : OAI221_X1 port map( B1 => n672, B2 => n708, C1 => n674, C2 => n709, A 
                           => n710, ZN => O_29_port);
   U45 : AOI22_X1 port map( A1 => A_ns(27), A2 => n671, B1 => A_s(27), B2 => 
                           n678, ZN => n710);
   U46 : INV_X1 port map( A => A_s(28), ZN => n709);
   U47 : INV_X1 port map( A => A_ns(28), ZN => n708);
   U48 : OAI221_X1 port map( B1 => n672, B2 => n711, C1 => n674, C2 => n712, A 
                           => n713, ZN => O_28_port);
   U49 : AOI22_X1 port map( A1 => A_ns(26), A2 => n671, B1 => A_s(26), B2 => 
                           n678, ZN => n713);
   U50 : INV_X1 port map( A => A_s(27), ZN => n712);
   U51 : INV_X1 port map( A => A_ns(27), ZN => n711);
   U52 : OAI221_X1 port map( B1 => n672, B2 => n714, C1 => n674, C2 => n715, A 
                           => n716, ZN => O_27_port);
   U53 : AOI22_X1 port map( A1 => A_ns(25), A2 => n671, B1 => A_s(25), B2 => 
                           n678, ZN => n716);
   U54 : INV_X1 port map( A => A_s(26), ZN => n715);
   U55 : INV_X1 port map( A => A_ns(26), ZN => n714);
   U56 : OAI221_X1 port map( B1 => n672, B2 => n717, C1 => n674, C2 => n718, A 
                           => n719, ZN => O_26_port);
   U57 : AOI22_X1 port map( A1 => A_ns(24), A2 => n671, B1 => A_s(24), B2 => 
                           n678, ZN => n719);
   U58 : INV_X1 port map( A => A_s(25), ZN => n718);
   U59 : INV_X1 port map( A => A_ns(25), ZN => n717);
   U60 : OAI221_X1 port map( B1 => n672, B2 => n720, C1 => n674, C2 => n721, A 
                           => n722, ZN => O_25_port);
   U61 : AOI22_X1 port map( A1 => A_ns(23), A2 => n671, B1 => A_s(23), B2 => 
                           n678, ZN => n722);
   U62 : INV_X1 port map( A => A_s(24), ZN => n721);
   U63 : INV_X1 port map( A => A_ns(24), ZN => n720);
   U64 : OAI221_X1 port map( B1 => n672, B2 => n723, C1 => n674, C2 => n724, A 
                           => n725, ZN => O_24_port);
   U65 : AOI22_X1 port map( A1 => A_ns(22), A2 => n671, B1 => A_s(22), B2 => 
                           n678, ZN => n725);
   U66 : INV_X1 port map( A => A_s(23), ZN => n724);
   U67 : INV_X1 port map( A => A_ns(23), ZN => n723);
   U68 : OAI221_X1 port map( B1 => n672, B2 => n726, C1 => n674, C2 => n727, A 
                           => n728, ZN => O_23_port);
   U69 : AOI22_X1 port map( A1 => A_ns(21), A2 => n671, B1 => A_s(21), B2 => 
                           n678, ZN => n728);
   U70 : INV_X1 port map( A => A_s(22), ZN => n727);
   U71 : INV_X1 port map( A => A_ns(22), ZN => n726);
   U72 : OAI221_X1 port map( B1 => n672, B2 => n729, C1 => n674, C2 => n730, A 
                           => n731, ZN => O_22_port);
   U73 : AOI22_X1 port map( A1 => A_ns(20), A2 => n671, B1 => A_s(20), B2 => 
                           n678, ZN => n731);
   U74 : INV_X1 port map( A => A_s(21), ZN => n730);
   U75 : INV_X1 port map( A => A_ns(21), ZN => n729);
   U76 : OAI221_X1 port map( B1 => n672, B2 => n732, C1 => n674, C2 => n733, A 
                           => n734, ZN => O_21_port);
   U77 : AOI22_X1 port map( A1 => A_ns(19), A2 => n671, B1 => A_s(19), B2 => 
                           n678, ZN => n734);
   U78 : INV_X1 port map( A => A_s(20), ZN => n733);
   U79 : INV_X1 port map( A => A_ns(20), ZN => n732);
   U80 : OAI221_X1 port map( B1 => n672, B2 => n735, C1 => n674, C2 => n736, A 
                           => n737, ZN => O_20_port);
   U81 : AOI22_X1 port map( A1 => A_ns(18), A2 => n671, B1 => A_s(18), B2 => 
                           n678, ZN => n737);
   U82 : INV_X1 port map( A => A_s(19), ZN => n736);
   U83 : INV_X1 port map( A => A_ns(19), ZN => n735);
   U84 : OAI221_X1 port map( B1 => n672, B2 => n738, C1 => n674, C2 => n739, A 
                           => n740, ZN => O_19_port);
   U85 : AOI22_X1 port map( A1 => A_ns(17), A2 => n671, B1 => A_s(17), B2 => 
                           n678, ZN => n740);
   U86 : INV_X1 port map( A => A_s(18), ZN => n739);
   U87 : INV_X1 port map( A => A_ns(18), ZN => n738);
   U88 : OAI221_X1 port map( B1 => n672, B2 => n741, C1 => n674, C2 => n742, A 
                           => n743, ZN => O_18_port);
   U89 : AOI22_X1 port map( A1 => A_ns(16), A2 => n671, B1 => A_s(16), B2 => 
                           n678, ZN => n743);
   U90 : INV_X1 port map( A => A_s(17), ZN => n742);
   U91 : INV_X1 port map( A => A_ns(17), ZN => n741);
   U92 : OAI221_X1 port map( B1 => n672, B2 => n744, C1 => n674, C2 => n745, A 
                           => n746, ZN => O_17_port);
   U93 : AOI22_X1 port map( A1 => A_ns(15), A2 => n671, B1 => A_s(15), B2 => 
                           n678, ZN => n746);
   U94 : INV_X1 port map( A => A_s(16), ZN => n745);
   U95 : INV_X1 port map( A => A_ns(16), ZN => n744);
   U96 : OAI221_X1 port map( B1 => n672, B2 => n747, C1 => n674, C2 => n748, A 
                           => n749, ZN => O_16_port);
   U97 : AOI22_X1 port map( A1 => A_ns(14), A2 => n671, B1 => A_s(14), B2 => 
                           n678, ZN => n749);
   U98 : INV_X1 port map( A => A_s(15), ZN => n748);
   U99 : INV_X1 port map( A => A_ns(15), ZN => n747);
   U100 : OAI221_X1 port map( B1 => n672, B2 => n750, C1 => n674, C2 => n751, A
                           => n752, ZN => O_15_port);
   U101 : AOI22_X1 port map( A1 => A_ns(13), A2 => n671, B1 => A_s(13), B2 => 
                           n678, ZN => n752);
   U102 : INV_X1 port map( A => A_s(14), ZN => n751);
   U103 : INV_X1 port map( A => A_ns(14), ZN => n750);
   U104 : OAI221_X1 port map( B1 => n672, B2 => n753, C1 => n674, C2 => n754, A
                           => n755, ZN => O_14_port);
   U105 : AOI22_X1 port map( A1 => A_ns(12), A2 => n671, B1 => A_s(12), B2 => 
                           n678, ZN => n755);
   U106 : INV_X1 port map( A => A_s(13), ZN => n754);
   U107 : INV_X1 port map( A => A_ns(13), ZN => n753);
   U108 : OAI221_X1 port map( B1 => n672, B2 => n756, C1 => n674, C2 => n757, A
                           => n758, ZN => O_13_port);
   U109 : AOI22_X1 port map( A1 => A_ns(11), A2 => n671, B1 => A_s(11), B2 => 
                           n678, ZN => n758);
   U110 : INV_X1 port map( A => A_s(12), ZN => n757);
   U111 : INV_X1 port map( A => A_ns(12), ZN => n756);
   U112 : OAI221_X1 port map( B1 => n672, B2 => n759, C1 => n674, C2 => n760, A
                           => n761, ZN => O_12_port);
   U113 : AOI22_X1 port map( A1 => A_ns(10), A2 => n671, B1 => A_s(10), B2 => 
                           n678, ZN => n761);
   U114 : INV_X1 port map( A => A_s(11), ZN => n760);
   U115 : INV_X1 port map( A => A_ns(11), ZN => n759);
   U116 : OAI221_X1 port map( B1 => n672, B2 => n762, C1 => n674, C2 => n763, A
                           => n764, ZN => O_11_port);
   U117 : AOI22_X1 port map( A1 => A_ns(9), A2 => n671, B1 => A_s(9), B2 => 
                           n678, ZN => n764);
   U118 : INV_X1 port map( A => A_s(10), ZN => n763);
   U119 : INV_X1 port map( A => A_ns(10), ZN => n762);
   U120 : OAI221_X1 port map( B1 => n672, B2 => n765, C1 => n674, C2 => n766, A
                           => n767, ZN => O_10_port);
   U121 : AOI22_X1 port map( A1 => A_ns(8), A2 => n671, B1 => A_s(8), B2 => 
                           n678, ZN => n767);
   U122 : INV_X1 port map( A => A_s(9), ZN => n766);
   U123 : INV_X1 port map( A => A_ns(9), ZN => n765);
   U124 : OAI221_X1 port map( B1 => n672, B2 => n768, C1 => n674, C2 => n769, A
                           => n770, ZN => O_9_port);
   U125 : AOI22_X1 port map( A1 => A_ns(7), A2 => n677, B1 => A_s(7), B2 => 
                           n678, ZN => n770);
   U126 : INV_X1 port map( A => A_s(8), ZN => n769);
   U127 : INV_X1 port map( A => A_ns(8), ZN => n768);
   U128 : OAI221_X1 port map( B1 => n672, B2 => n771, C1 => n674, C2 => n772, A
                           => n773, ZN => O_8_port);
   U129 : AOI22_X1 port map( A1 => A_ns(6), A2 => n677, B1 => A_s(6), B2 => 
                           n678, ZN => n773);
   U130 : INV_X1 port map( A => A_s(7), ZN => n772);
   U131 : INV_X1 port map( A => A_ns(7), ZN => n771);
   U132 : OAI221_X1 port map( B1 => n672, B2 => n774, C1 => n674, C2 => n775, A
                           => n776, ZN => O_7_port);
   U133 : AOI22_X1 port map( A1 => A_ns(5), A2 => n677, B1 => A_s(5), B2 => 
                           n678, ZN => n776);
   U134 : INV_X1 port map( A => A_s(6), ZN => n775);
   U135 : INV_X1 port map( A => A_ns(6), ZN => n774);
   U136 : INV_X1 port map( A => n777, ZN => O_1_port);
   U137 : AOI22_X1 port map( A1 => n686, A2 => A_s(0), B1 => n685, B2 => 
                           A_ns(0), ZN => n777);
   U138 : OAI221_X1 port map( B1 => n672, B2 => n778, C1 => n674, C2 => n779, A
                           => n780, ZN => O_2_port);
   U139 : AOI22_X1 port map( A1 => A_ns(0), A2 => n677, B1 => A_s(0), B2 => 
                           n678, ZN => n780);
   U140 : INV_X1 port map( A => n781, ZN => O_3_port);
   U141 : AOI221_X1 port map( B1 => n685, B2 => A_ns(2), C1 => n686, C2 => 
                           A_s(2), A => n782, ZN => n781);
   U142 : OAI22_X1 port map( A1 => n778, A2 => n682, B1 => n779, B2 => n683, ZN
                           => n782);
   U143 : INV_X1 port map( A => A_s(1), ZN => n779);
   U144 : INV_X1 port map( A => A_ns(1), ZN => n778);
   U145 : OAI221_X1 port map( B1 => n672, B2 => n783, C1 => n674, C2 => n784, A
                           => n785, ZN => O_4_port);
   U146 : AOI22_X1 port map( A1 => A_ns(2), A2 => n677, B1 => A_s(2), B2 => 
                           n678, ZN => n785);
   U147 : INV_X1 port map( A => n786, ZN => O_5_port);
   U148 : AOI221_X1 port map( B1 => n685, B2 => A_ns(4), C1 => n686, C2 => 
                           A_s(4), A => n787, ZN => n786);
   U149 : OAI22_X1 port map( A1 => n783, A2 => n682, B1 => n784, B2 => n683, ZN
                           => n787);
   U150 : INV_X1 port map( A => A_s(3), ZN => n784);
   U151 : INV_X1 port map( A => n677, ZN => n682);
   U152 : INV_X1 port map( A => A_ns(3), ZN => n783);
   U153 : INV_X1 port map( A => n674, ZN => n686);
   U154 : INV_X1 port map( A => n672, ZN => n685);
   U155 : OAI221_X1 port map( B1 => n672, B2 => n788, C1 => n674, C2 => n789, A
                           => n790, ZN => O_6_port);
   U156 : AOI22_X1 port map( A1 => A_ns(4), A2 => n677, B1 => A_s(4), B2 => 
                           n678, ZN => n790);
   U157 : NAND3_X1 port map( A1 => B(5), A2 => n791, A3 => B(6), ZN => n683);
   U158 : NOR3_X1 port map( A1 => B(5), A2 => B(6), A3 => n791, ZN => n677);
   U159 : INV_X1 port map( A => A_s(5), ZN => n789);
   U160 : INV_X1 port map( A => A_ns(5), ZN => n788);
   U161 : INV_X1 port map( A => B(7), ZN => n791);
   U162 : XOR2_X1 port map( A => B(6), B => B(5), Z => n792);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT38_i4 is

   port( A_s, A_ns, B : in std_logic_vector (37 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (37 downto 0));

end BOOTHENC_NBIT38_i4;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT38_i4 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, n633, n634, n635, n636, n637, n638, n639, n640, n641, 
      n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, 
      n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, 
      n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, 
      n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, 
      n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, 
      n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, 
      n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, 
      n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, 
      n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, 
      O_36_port, O_35_port, O_37_port, O_34_port, O_33_port, O_32_port, 
      O_31_port, O_30_port, O_29_port, O_28_port, O_27_port, O_26_port, 
      O_25_port, O_24_port, O_23_port, O_22_port, O_21_port, O_20_port, 
      O_19_port, O_18_port, O_17_port, O_16_port, O_15_port, O_14_port, 
      O_13_port, O_12_port, O_11_port, O_10_port, O_9_port, O_8_port, O_7_port,
      O_6_port, O_5_port, O_1_port, O_2_port, O_3_port, O_4_port : std_logic;

begin
   O <= ( O_37_port, O_36_port, O_35_port, O_34_port, O_33_port, O_32_port, 
      O_31_port, O_30_port, O_29_port, O_28_port, O_27_port, O_26_port, 
      O_25_port, O_24_port, O_23_port, O_22_port, O_21_port, O_20_port, 
      O_19_port, O_18_port, O_17_port, O_16_port, O_15_port, O_14_port, 
      O_13_port, O_12_port, O_11_port, O_10_port, O_9_port, O_8_port, O_7_port,
      O_6_port, O_5_port, O_4_port, O_3_port, O_2_port, O_1_port, X_Logic0_port
      );
   A_so <= ( A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), A_s(30), A_s(29), 
      A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), A_s(22), A_s(21), 
      A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), A_s(14), A_s(13), 
      A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), A_s(6), A_s(5), A_s(4)
      , A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, X_Logic0_port );
   A_nso <= ( A_ns(35), A_ns(34), A_ns(33), A_ns(32), A_ns(31), A_ns(30), 
      A_ns(29), A_ns(28), A_ns(27), A_ns(26), A_ns(25), A_ns(24), A_ns(23), 
      A_ns(22), A_ns(21), A_ns(20), A_ns(19), A_ns(18), A_ns(17), A_ns(16), 
      A_ns(15), A_ns(14), A_ns(13), A_ns(12), A_ns(11), A_ns(10), A_ns(9), 
      A_ns(8), A_ns(7), A_ns(6), A_ns(5), A_ns(4), A_ns(3), A_ns(2), A_ns(1), 
      A_ns(0), X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : NAND2_X2 port map( A1 => n749, A2 => n636, ZN => n634);
   U3 : NAND2_X2 port map( A1 => n749, A2 => n748, ZN => n636);
   U4 : INV_X2 port map( A => n645, ZN => n640);
   U5 : INV_X2 port map( A => n644, ZN => n633);
   U6 : OAI221_X1 port map( B1 => n634, B2 => n635, C1 => n636, C2 => n637, A 
                           => n638, ZN => O_36_port);
   U7 : AOI22_X1 port map( A1 => A_ns(34), A2 => n633, B1 => A_s(34), B2 => 
                           n640, ZN => n638);
   U8 : OAI221_X1 port map( B1 => n641, B2 => n634, C1 => n642, C2 => n636, A 
                           => n643, ZN => O_35_port);
   U9 : AOI22_X1 port map( A1 => A_ns(33), A2 => n633, B1 => A_s(33), B2 => 
                           n640, ZN => n643);
   U10 : INV_X1 port map( A => A_s(34), ZN => n642);
   U11 : INV_X1 port map( A => A_ns(34), ZN => n641);
   U12 : OAI221_X1 port map( B1 => n644, B2 => n635, C1 => n645, C2 => n637, A 
                           => n646, ZN => O_37_port);
   U13 : AOI22_X1 port map( A1 => A_ns(36), A2 => n647, B1 => A_s(36), B2 => 
                           n648, ZN => n646);
   U14 : INV_X1 port map( A => A_s(35), ZN => n637);
   U15 : INV_X1 port map( A => A_ns(35), ZN => n635);
   U16 : OAI221_X1 port map( B1 => n634, B2 => n649, C1 => n636, C2 => n650, A 
                           => n651, ZN => O_34_port);
   U17 : AOI22_X1 port map( A1 => A_ns(32), A2 => n633, B1 => A_s(32), B2 => 
                           n640, ZN => n651);
   U18 : INV_X1 port map( A => A_s(33), ZN => n650);
   U19 : INV_X1 port map( A => A_ns(33), ZN => n649);
   U20 : OAI221_X1 port map( B1 => n634, B2 => n652, C1 => n636, C2 => n653, A 
                           => n654, ZN => O_33_port);
   U21 : AOI22_X1 port map( A1 => A_ns(31), A2 => n633, B1 => A_s(31), B2 => 
                           n640, ZN => n654);
   U22 : INV_X1 port map( A => A_s(32), ZN => n653);
   U23 : INV_X1 port map( A => A_ns(32), ZN => n652);
   U24 : OAI221_X1 port map( B1 => n634, B2 => n655, C1 => n636, C2 => n656, A 
                           => n657, ZN => O_32_port);
   U25 : AOI22_X1 port map( A1 => A_ns(30), A2 => n633, B1 => A_s(30), B2 => 
                           n640, ZN => n657);
   U26 : INV_X1 port map( A => A_s(31), ZN => n656);
   U27 : INV_X1 port map( A => A_ns(31), ZN => n655);
   U28 : OAI221_X1 port map( B1 => n634, B2 => n658, C1 => n636, C2 => n659, A 
                           => n660, ZN => O_31_port);
   U29 : AOI22_X1 port map( A1 => A_ns(29), A2 => n633, B1 => A_s(29), B2 => 
                           n640, ZN => n660);
   U30 : INV_X1 port map( A => A_s(30), ZN => n659);
   U31 : INV_X1 port map( A => A_ns(30), ZN => n658);
   U32 : OAI221_X1 port map( B1 => n634, B2 => n661, C1 => n636, C2 => n662, A 
                           => n663, ZN => O_30_port);
   U33 : AOI22_X1 port map( A1 => A_ns(28), A2 => n633, B1 => A_s(28), B2 => 
                           n640, ZN => n663);
   U34 : INV_X1 port map( A => A_s(29), ZN => n662);
   U35 : INV_X1 port map( A => A_ns(29), ZN => n661);
   U36 : OAI221_X1 port map( B1 => n634, B2 => n664, C1 => n636, C2 => n665, A 
                           => n666, ZN => O_29_port);
   U37 : AOI22_X1 port map( A1 => A_ns(27), A2 => n633, B1 => A_s(27), B2 => 
                           n640, ZN => n666);
   U38 : INV_X1 port map( A => A_s(28), ZN => n665);
   U39 : INV_X1 port map( A => A_ns(28), ZN => n664);
   U40 : OAI221_X1 port map( B1 => n634, B2 => n667, C1 => n636, C2 => n668, A 
                           => n669, ZN => O_28_port);
   U41 : AOI22_X1 port map( A1 => A_ns(26), A2 => n633, B1 => A_s(26), B2 => 
                           n640, ZN => n669);
   U42 : INV_X1 port map( A => A_s(27), ZN => n668);
   U43 : INV_X1 port map( A => A_ns(27), ZN => n667);
   U44 : OAI221_X1 port map( B1 => n634, B2 => n670, C1 => n636, C2 => n671, A 
                           => n672, ZN => O_27_port);
   U45 : AOI22_X1 port map( A1 => A_ns(25), A2 => n633, B1 => A_s(25), B2 => 
                           n640, ZN => n672);
   U46 : INV_X1 port map( A => A_s(26), ZN => n671);
   U47 : INV_X1 port map( A => A_ns(26), ZN => n670);
   U48 : OAI221_X1 port map( B1 => n634, B2 => n673, C1 => n636, C2 => n674, A 
                           => n675, ZN => O_26_port);
   U49 : AOI22_X1 port map( A1 => A_ns(24), A2 => n633, B1 => A_s(24), B2 => 
                           n640, ZN => n675);
   U50 : INV_X1 port map( A => A_s(25), ZN => n674);
   U51 : INV_X1 port map( A => A_ns(25), ZN => n673);
   U52 : OAI221_X1 port map( B1 => n634, B2 => n676, C1 => n636, C2 => n677, A 
                           => n678, ZN => O_25_port);
   U53 : AOI22_X1 port map( A1 => A_ns(23), A2 => n633, B1 => A_s(23), B2 => 
                           n640, ZN => n678);
   U54 : INV_X1 port map( A => A_s(24), ZN => n677);
   U55 : INV_X1 port map( A => A_ns(24), ZN => n676);
   U56 : OAI221_X1 port map( B1 => n634, B2 => n679, C1 => n636, C2 => n680, A 
                           => n681, ZN => O_24_port);
   U57 : AOI22_X1 port map( A1 => A_ns(22), A2 => n633, B1 => A_s(22), B2 => 
                           n640, ZN => n681);
   U58 : INV_X1 port map( A => A_s(23), ZN => n680);
   U59 : INV_X1 port map( A => A_ns(23), ZN => n679);
   U60 : OAI221_X1 port map( B1 => n634, B2 => n682, C1 => n636, C2 => n683, A 
                           => n684, ZN => O_23_port);
   U61 : AOI22_X1 port map( A1 => A_ns(21), A2 => n633, B1 => A_s(21), B2 => 
                           n640, ZN => n684);
   U62 : INV_X1 port map( A => A_s(22), ZN => n683);
   U63 : INV_X1 port map( A => A_ns(22), ZN => n682);
   U64 : OAI221_X1 port map( B1 => n634, B2 => n685, C1 => n636, C2 => n686, A 
                           => n687, ZN => O_22_port);
   U65 : AOI22_X1 port map( A1 => A_ns(20), A2 => n633, B1 => A_s(20), B2 => 
                           n640, ZN => n687);
   U66 : INV_X1 port map( A => A_s(21), ZN => n686);
   U67 : INV_X1 port map( A => A_ns(21), ZN => n685);
   U68 : OAI221_X1 port map( B1 => n634, B2 => n688, C1 => n636, C2 => n689, A 
                           => n690, ZN => O_21_port);
   U69 : AOI22_X1 port map( A1 => A_ns(19), A2 => n633, B1 => A_s(19), B2 => 
                           n640, ZN => n690);
   U70 : INV_X1 port map( A => A_s(20), ZN => n689);
   U71 : INV_X1 port map( A => A_ns(20), ZN => n688);
   U72 : OAI221_X1 port map( B1 => n634, B2 => n691, C1 => n636, C2 => n692, A 
                           => n693, ZN => O_20_port);
   U73 : AOI22_X1 port map( A1 => A_ns(18), A2 => n633, B1 => A_s(18), B2 => 
                           n640, ZN => n693);
   U74 : INV_X1 port map( A => A_s(19), ZN => n692);
   U75 : INV_X1 port map( A => A_ns(19), ZN => n691);
   U76 : OAI221_X1 port map( B1 => n634, B2 => n694, C1 => n636, C2 => n695, A 
                           => n696, ZN => O_19_port);
   U77 : AOI22_X1 port map( A1 => A_ns(17), A2 => n633, B1 => A_s(17), B2 => 
                           n640, ZN => n696);
   U78 : INV_X1 port map( A => A_s(18), ZN => n695);
   U79 : INV_X1 port map( A => A_ns(18), ZN => n694);
   U80 : OAI221_X1 port map( B1 => n634, B2 => n697, C1 => n636, C2 => n698, A 
                           => n699, ZN => O_18_port);
   U81 : AOI22_X1 port map( A1 => A_ns(16), A2 => n633, B1 => A_s(16), B2 => 
                           n640, ZN => n699);
   U82 : INV_X1 port map( A => A_s(17), ZN => n698);
   U83 : INV_X1 port map( A => A_ns(17), ZN => n697);
   U84 : OAI221_X1 port map( B1 => n634, B2 => n700, C1 => n636, C2 => n701, A 
                           => n702, ZN => O_17_port);
   U85 : AOI22_X1 port map( A1 => A_ns(15), A2 => n633, B1 => A_s(15), B2 => 
                           n640, ZN => n702);
   U86 : INV_X1 port map( A => A_s(16), ZN => n701);
   U87 : INV_X1 port map( A => A_ns(16), ZN => n700);
   U88 : OAI221_X1 port map( B1 => n634, B2 => n703, C1 => n636, C2 => n704, A 
                           => n705, ZN => O_16_port);
   U89 : AOI22_X1 port map( A1 => A_ns(14), A2 => n633, B1 => A_s(14), B2 => 
                           n640, ZN => n705);
   U90 : INV_X1 port map( A => A_s(15), ZN => n704);
   U91 : INV_X1 port map( A => A_ns(15), ZN => n703);
   U92 : OAI221_X1 port map( B1 => n634, B2 => n706, C1 => n636, C2 => n707, A 
                           => n708, ZN => O_15_port);
   U93 : AOI22_X1 port map( A1 => A_ns(13), A2 => n633, B1 => A_s(13), B2 => 
                           n640, ZN => n708);
   U94 : INV_X1 port map( A => A_s(14), ZN => n707);
   U95 : INV_X1 port map( A => A_ns(14), ZN => n706);
   U96 : OAI221_X1 port map( B1 => n634, B2 => n709, C1 => n636, C2 => n710, A 
                           => n711, ZN => O_14_port);
   U97 : AOI22_X1 port map( A1 => A_ns(12), A2 => n633, B1 => A_s(12), B2 => 
                           n640, ZN => n711);
   U98 : INV_X1 port map( A => A_s(13), ZN => n710);
   U99 : INV_X1 port map( A => A_ns(13), ZN => n709);
   U100 : OAI221_X1 port map( B1 => n634, B2 => n712, C1 => n636, C2 => n713, A
                           => n714, ZN => O_13_port);
   U101 : AOI22_X1 port map( A1 => A_ns(11), A2 => n633, B1 => A_s(11), B2 => 
                           n640, ZN => n714);
   U102 : INV_X1 port map( A => A_s(12), ZN => n713);
   U103 : INV_X1 port map( A => A_ns(12), ZN => n712);
   U104 : OAI221_X1 port map( B1 => n634, B2 => n715, C1 => n636, C2 => n716, A
                           => n717, ZN => O_12_port);
   U105 : AOI22_X1 port map( A1 => A_ns(10), A2 => n633, B1 => A_s(10), B2 => 
                           n640, ZN => n717);
   U106 : INV_X1 port map( A => A_s(11), ZN => n716);
   U107 : INV_X1 port map( A => A_ns(11), ZN => n715);
   U108 : OAI221_X1 port map( B1 => n634, B2 => n718, C1 => n636, C2 => n719, A
                           => n720, ZN => O_11_port);
   U109 : AOI22_X1 port map( A1 => A_ns(9), A2 => n633, B1 => A_s(9), B2 => 
                           n640, ZN => n720);
   U110 : INV_X1 port map( A => A_s(10), ZN => n719);
   U111 : INV_X1 port map( A => A_ns(10), ZN => n718);
   U112 : OAI221_X1 port map( B1 => n634, B2 => n721, C1 => n636, C2 => n722, A
                           => n723, ZN => O_10_port);
   U113 : AOI22_X1 port map( A1 => A_ns(8), A2 => n633, B1 => A_s(8), B2 => 
                           n640, ZN => n723);
   U114 : INV_X1 port map( A => A_s(9), ZN => n722);
   U115 : INV_X1 port map( A => A_ns(9), ZN => n721);
   U116 : OAI221_X1 port map( B1 => n634, B2 => n724, C1 => n636, C2 => n725, A
                           => n726, ZN => O_9_port);
   U117 : AOI22_X1 port map( A1 => A_ns(7), A2 => n633, B1 => A_s(7), B2 => 
                           n640, ZN => n726);
   U118 : INV_X1 port map( A => A_s(8), ZN => n725);
   U119 : INV_X1 port map( A => A_ns(8), ZN => n724);
   U120 : OAI221_X1 port map( B1 => n634, B2 => n727, C1 => n636, C2 => n728, A
                           => n729, ZN => O_8_port);
   U121 : AOI22_X1 port map( A1 => A_ns(6), A2 => n633, B1 => A_s(6), B2 => 
                           n640, ZN => n729);
   U122 : INV_X1 port map( A => A_s(7), ZN => n728);
   U123 : INV_X1 port map( A => A_ns(7), ZN => n727);
   U124 : OAI221_X1 port map( B1 => n634, B2 => n730, C1 => n636, C2 => n731, A
                           => n732, ZN => O_7_port);
   U125 : AOI22_X1 port map( A1 => A_ns(5), A2 => n639, B1 => A_s(5), B2 => 
                           n640, ZN => n732);
   U126 : INV_X1 port map( A => A_s(6), ZN => n731);
   U127 : INV_X1 port map( A => A_ns(6), ZN => n730);
   U128 : OAI221_X1 port map( B1 => n634, B2 => n733, C1 => n636, C2 => n734, A
                           => n735, ZN => O_6_port);
   U129 : AOI22_X1 port map( A1 => A_ns(4), A2 => n639, B1 => A_s(4), B2 => 
                           n640, ZN => n735);
   U130 : INV_X1 port map( A => A_s(5), ZN => n734);
   U131 : INV_X1 port map( A => A_ns(5), ZN => n733);
   U132 : OAI221_X1 port map( B1 => n634, B2 => n736, C1 => n636, C2 => n737, A
                           => n738, ZN => O_5_port);
   U133 : AOI22_X1 port map( A1 => A_ns(3), A2 => n639, B1 => A_s(3), B2 => 
                           n640, ZN => n738);
   U134 : INV_X1 port map( A => A_s(4), ZN => n737);
   U135 : INV_X1 port map( A => A_ns(4), ZN => n736);
   U136 : INV_X1 port map( A => n739, ZN => O_1_port);
   U137 : AOI22_X1 port map( A1 => n648, A2 => A_s(0), B1 => n647, B2 => 
                           A_ns(0), ZN => n739);
   U138 : OAI221_X1 port map( B1 => n634, B2 => n740, C1 => n636, C2 => n741, A
                           => n742, ZN => O_2_port);
   U139 : AOI22_X1 port map( A1 => A_ns(0), A2 => n639, B1 => A_s(0), B2 => 
                           n640, ZN => n742);
   U140 : INV_X1 port map( A => n743, ZN => O_3_port);
   U141 : AOI221_X1 port map( B1 => n647, B2 => A_ns(2), C1 => n648, C2 => 
                           A_s(2), A => n744, ZN => n743);
   U142 : OAI22_X1 port map( A1 => n740, A2 => n644, B1 => n741, B2 => n645, ZN
                           => n744);
   U143 : INV_X1 port map( A => A_s(1), ZN => n741);
   U144 : INV_X1 port map( A => n639, ZN => n644);
   U145 : INV_X1 port map( A => A_ns(1), ZN => n740);
   U146 : INV_X1 port map( A => n636, ZN => n648);
   U147 : INV_X1 port map( A => n634, ZN => n647);
   U148 : OAI221_X1 port map( B1 => n634, B2 => n745, C1 => n636, C2 => n746, A
                           => n747, ZN => O_4_port);
   U149 : AOI22_X1 port map( A1 => A_ns(2), A2 => n639, B1 => A_s(2), B2 => 
                           n640, ZN => n747);
   U150 : NAND3_X1 port map( A1 => B(3), A2 => n748, A3 => B(4), ZN => n645);
   U151 : NOR3_X1 port map( A1 => B(3), A2 => B(4), A3 => n748, ZN => n639);
   U152 : INV_X1 port map( A => A_s(3), ZN => n746);
   U153 : INV_X1 port map( A => A_ns(3), ZN => n745);
   U154 : INV_X1 port map( A => B(5), ZN => n748);
   U155 : XOR2_X1 port map( A => B(4), B => B(3), Z => n749);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT36_i2 is

   port( A_s, A_ns, B : in std_logic_vector (35 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (35 downto 0));

end BOOTHENC_NBIT36_i2;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT36_i2 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, O_7_port, O_4_port, O_2_port, O_35_port, O_33_port, 
      O_31_port, O_29_port, O_27_port, O_25_port, O_23_port, O_21_port, 
      O_19_port, O_17_port, O_15_port, O_13_port, O_11_port, O_10_port, 
      O_9_port, O_5_port, n571, n572, n573, n574, n575, n576, n577, n578, n579,
      n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, 
      n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, 
      n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, 
      n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, 
      n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, 
      n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, 
      n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, 
      n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, 
      n676, n677, n678, n679, n680, n681, O_34_port, O_32_port, O_30_port, 
      O_28_port, O_26_port, O_24_port, O_22_port, O_20_port, O_18_port, 
      O_16_port, O_14_port, O_12_port, O_8_port, O_6_port, O_3_port, O_1_port :
      std_logic;

begin
   O <= ( O_35_port, O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, 
      O_29_port, O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, 
      O_23_port, O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, 
      O_17_port, O_16_port, O_15_port, O_14_port, O_13_port, O_12_port, 
      O_11_port, O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, 
      O_4_port, O_3_port, O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(33), A_s(32), A_s(31), A_s(30), A_s(29), A_s(28), A_s(27), 
      A_s(26), A_s(25), A_s(24), A_s(23), A_s(22), A_s(21), A_s(20), A_s(19), 
      A_s(18), A_s(17), A_s(16), A_s(15), A_s(14), A_s(13), A_s(12), A_s(11), 
      A_s(10), A_s(9), A_s(8), A_s(7), A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), 
      A_s(1), A_s(0), X_Logic0_port, X_Logic0_port );
   A_nso <= ( A_ns(33), A_ns(32), A_ns(31), A_ns(30), A_ns(29), A_ns(28), 
      A_ns(27), A_ns(26), A_ns(25), A_ns(24), A_ns(23), A_ns(22), A_ns(21), 
      A_ns(20), A_ns(19), A_ns(18), A_ns(17), A_ns(16), A_ns(15), A_ns(14), 
      A_ns(13), A_ns(12), A_ns(11), A_ns(10), A_ns(9), A_ns(8), A_ns(7), 
      A_ns(6), A_ns(5), A_ns(4), A_ns(3), A_ns(2), A_ns(1), A_ns(0), 
      X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : OR3_X1 port map( A1 => B(1), A2 => B(2), A3 => n681, ZN => n571);
   U3 : NAND3_X2 port map( A1 => B(2), A2 => n681, A3 => B(1), ZN => n575);
   U4 : INV_X2 port map( A => n571, ZN => n572);
   U5 : INV_X2 port map( A => n622, ZN => n578);
   U6 : NAND2_X2 port map( A1 => B(3), A2 => n680, ZN => n573);
   U7 : OAI221_X1 port map( B1 => n573, B2 => n574, C1 => n575, C2 => n576, A 
                           => n577, ZN => O_34_port);
   U8 : AOI22_X1 port map( A1 => A_ns(32), A2 => n572, B1 => A_s(33), B2 => 
                           n578, ZN => n577);
   U9 : INV_X1 port map( A => A_s(32), ZN => n576);
   U10 : INV_X1 port map( A => A_ns(33), ZN => n574);
   U11 : OAI221_X1 port map( B1 => n573, B2 => n579, C1 => n575, C2 => n580, A 
                           => n581, ZN => O_32_port);
   U12 : AOI22_X1 port map( A1 => A_ns(30), A2 => n572, B1 => A_s(31), B2 => 
                           n578, ZN => n581);
   U13 : INV_X1 port map( A => A_s(30), ZN => n580);
   U14 : INV_X1 port map( A => A_ns(31), ZN => n579);
   U15 : OAI221_X1 port map( B1 => n573, B2 => n582, C1 => n575, C2 => n583, A 
                           => n584, ZN => O_30_port);
   U16 : AOI22_X1 port map( A1 => A_ns(28), A2 => n572, B1 => A_s(29), B2 => 
                           n578, ZN => n584);
   U17 : INV_X1 port map( A => A_s(28), ZN => n583);
   U18 : INV_X1 port map( A => A_ns(29), ZN => n582);
   U19 : OAI221_X1 port map( B1 => n573, B2 => n585, C1 => n575, C2 => n586, A 
                           => n587, ZN => O_28_port);
   U20 : AOI22_X1 port map( A1 => A_ns(26), A2 => n572, B1 => A_s(27), B2 => 
                           n578, ZN => n587);
   U21 : INV_X1 port map( A => A_s(26), ZN => n586);
   U22 : INV_X1 port map( A => A_ns(27), ZN => n585);
   U23 : OAI221_X1 port map( B1 => n573, B2 => n588, C1 => n575, C2 => n589, A 
                           => n590, ZN => O_26_port);
   U24 : AOI22_X1 port map( A1 => A_ns(24), A2 => n572, B1 => A_s(25), B2 => 
                           n578, ZN => n590);
   U25 : INV_X1 port map( A => A_s(24), ZN => n589);
   U26 : INV_X1 port map( A => A_ns(25), ZN => n588);
   U27 : OAI221_X1 port map( B1 => n573, B2 => n591, C1 => n575, C2 => n592, A 
                           => n593, ZN => O_24_port);
   U28 : AOI22_X1 port map( A1 => A_ns(22), A2 => n572, B1 => A_s(23), B2 => 
                           n578, ZN => n593);
   U29 : INV_X1 port map( A => A_s(22), ZN => n592);
   U30 : INV_X1 port map( A => A_ns(23), ZN => n591);
   U31 : OAI221_X1 port map( B1 => n573, B2 => n594, C1 => n575, C2 => n595, A 
                           => n596, ZN => O_22_port);
   U32 : AOI22_X1 port map( A1 => A_ns(20), A2 => n572, B1 => A_s(21), B2 => 
                           n578, ZN => n596);
   U33 : INV_X1 port map( A => A_s(20), ZN => n595);
   U34 : INV_X1 port map( A => A_ns(21), ZN => n594);
   U35 : OAI221_X1 port map( B1 => n573, B2 => n597, C1 => n575, C2 => n598, A 
                           => n599, ZN => O_20_port);
   U36 : AOI22_X1 port map( A1 => A_ns(18), A2 => n572, B1 => A_s(19), B2 => 
                           n578, ZN => n599);
   U37 : INV_X1 port map( A => A_s(18), ZN => n598);
   U38 : INV_X1 port map( A => A_ns(19), ZN => n597);
   U39 : OAI221_X1 port map( B1 => n573, B2 => n600, C1 => n575, C2 => n601, A 
                           => n602, ZN => O_18_port);
   U40 : AOI22_X1 port map( A1 => A_ns(16), A2 => n572, B1 => A_s(17), B2 => 
                           n578, ZN => n602);
   U41 : INV_X1 port map( A => A_s(16), ZN => n601);
   U42 : INV_X1 port map( A => A_ns(17), ZN => n600);
   U43 : OAI221_X1 port map( B1 => n573, B2 => n603, C1 => n575, C2 => n604, A 
                           => n605, ZN => O_16_port);
   U44 : AOI22_X1 port map( A1 => A_ns(14), A2 => n572, B1 => A_s(15), B2 => 
                           n578, ZN => n605);
   U45 : INV_X1 port map( A => A_s(14), ZN => n604);
   U46 : INV_X1 port map( A => A_ns(15), ZN => n603);
   U47 : OAI221_X1 port map( B1 => n573, B2 => n606, C1 => n575, C2 => n607, A 
                           => n608, ZN => O_14_port);
   U48 : AOI22_X1 port map( A1 => A_ns(12), A2 => n572, B1 => A_s(13), B2 => 
                           n578, ZN => n608);
   U49 : INV_X1 port map( A => A_s(12), ZN => n607);
   U50 : INV_X1 port map( A => A_ns(13), ZN => n606);
   U51 : OAI221_X1 port map( B1 => n573, B2 => n609, C1 => n575, C2 => n610, A 
                           => n611, ZN => O_12_port);
   U52 : AOI22_X1 port map( A1 => A_ns(10), A2 => n572, B1 => A_s(11), B2 => 
                           n578, ZN => n611);
   U53 : INV_X1 port map( A => A_s(10), ZN => n610);
   U54 : INV_X1 port map( A => A_ns(11), ZN => n609);
   U55 : OAI221_X1 port map( B1 => n573, B2 => n612, C1 => n575, C2 => n613, A 
                           => n614, ZN => O_8_port);
   U56 : AOI22_X1 port map( A1 => A_ns(6), A2 => n572, B1 => A_s(7), B2 => n578
                           , ZN => n614);
   U57 : INV_X1 port map( A => A_s(6), ZN => n613);
   U58 : INV_X1 port map( A => A_ns(7), ZN => n612);
   U59 : OAI221_X1 port map( B1 => n573, B2 => n615, C1 => n575, C2 => n616, A 
                           => n617, ZN => O_6_port);
   U60 : AOI22_X1 port map( A1 => A_ns(4), A2 => n572, B1 => A_s(5), B2 => n578
                           , ZN => n617);
   U61 : INV_X1 port map( A => A_s(4), ZN => n616);
   U62 : INV_X1 port map( A => A_ns(5), ZN => n615);
   U63 : OAI221_X1 port map( B1 => n573, B2 => n618, C1 => n575, C2 => n619, A 
                           => n620, ZN => O_3_port);
   U64 : AOI22_X1 port map( A1 => A_ns(1), A2 => n572, B1 => A_s(2), B2 => n578
                           , ZN => n620);
   U65 : INV_X1 port map( A => A_s(1), ZN => n619);
   U66 : INV_X1 port map( A => A_ns(2), ZN => n618);
   U67 : OAI22_X1 port map( A1 => n573, A2 => n621, B1 => n622, B2 => n623, ZN 
                           => O_1_port);
   U68 : INV_X1 port map( A => A_ns(0), ZN => n621);
   U69 : OAI221_X1 port map( B1 => n573, B2 => n624, C1 => n575, C2 => n625, A 
                           => n626, ZN => O_9_port);
   U70 : AOI22_X1 port map( A1 => A_ns(7), A2 => n572, B1 => A_s(8), B2 => n578
                           , ZN => n626);
   U71 : INV_X1 port map( A => A_s(7), ZN => n625);
   U72 : INV_X1 port map( A => A_ns(8), ZN => n624);
   U73 : OAI221_X1 port map( B1 => n573, B2 => n627, C1 => n575, C2 => n628, A 
                           => n629, ZN => O_7_port);
   U74 : AOI22_X1 port map( A1 => A_ns(5), A2 => n572, B1 => A_s(6), B2 => n578
                           , ZN => n629);
   U75 : INV_X1 port map( A => A_s(5), ZN => n628);
   U76 : INV_X1 port map( A => A_ns(6), ZN => n627);
   U77 : OAI221_X1 port map( B1 => n573, B2 => n630, C1 => n575, C2 => n631, A 
                           => n632, ZN => O_5_port);
   U78 : AOI22_X1 port map( A1 => A_ns(3), A2 => n572, B1 => A_s(4), B2 => n578
                           , ZN => n632);
   U79 : INV_X1 port map( A => A_s(3), ZN => n631);
   U80 : INV_X1 port map( A => A_ns(4), ZN => n630);
   U81 : OAI221_X1 port map( B1 => n573, B2 => n633, C1 => n575, C2 => n634, A 
                           => n635, ZN => O_4_port);
   U82 : AOI22_X1 port map( A1 => A_ns(2), A2 => n572, B1 => A_s(3), B2 => n578
                           , ZN => n635);
   U83 : INV_X1 port map( A => A_s(2), ZN => n634);
   U84 : INV_X1 port map( A => A_ns(3), ZN => n633);
   U85 : OAI221_X1 port map( B1 => n573, B2 => n636, C1 => n637, C2 => n575, A 
                           => n638, ZN => O_35_port);
   U86 : AOI22_X1 port map( A1 => A_ns(33), A2 => n572, B1 => A_s(34), B2 => 
                           n578, ZN => n638);
   U87 : INV_X1 port map( A => A_s(33), ZN => n637);
   U88 : INV_X1 port map( A => A_ns(34), ZN => n636);
   U89 : OAI221_X1 port map( B1 => n639, B2 => n573, C1 => n575, C2 => n640, A 
                           => n641, ZN => O_33_port);
   U90 : AOI22_X1 port map( A1 => A_ns(31), A2 => n572, B1 => A_s(32), B2 => 
                           n578, ZN => n641);
   U91 : INV_X1 port map( A => A_s(31), ZN => n640);
   U92 : INV_X1 port map( A => A_ns(32), ZN => n639);
   U93 : OAI221_X1 port map( B1 => n573, B2 => n642, C1 => n575, C2 => n643, A 
                           => n644, ZN => O_31_port);
   U94 : AOI22_X1 port map( A1 => A_ns(29), A2 => n572, B1 => A_s(30), B2 => 
                           n578, ZN => n644);
   U95 : INV_X1 port map( A => A_s(29), ZN => n643);
   U96 : INV_X1 port map( A => A_ns(30), ZN => n642);
   U97 : OAI221_X1 port map( B1 => n573, B2 => n645, C1 => n575, C2 => n623, A 
                           => n646, ZN => O_2_port);
   U98 : AOI22_X1 port map( A1 => A_ns(0), A2 => n572, B1 => A_s(1), B2 => n578
                           , ZN => n646);
   U99 : INV_X1 port map( A => A_s(0), ZN => n623);
   U100 : INV_X1 port map( A => A_ns(1), ZN => n645);
   U101 : OAI221_X1 port map( B1 => n573, B2 => n647, C1 => n575, C2 => n648, A
                           => n649, ZN => O_29_port);
   U102 : AOI22_X1 port map( A1 => A_ns(27), A2 => n572, B1 => A_s(28), B2 => 
                           n578, ZN => n649);
   U103 : INV_X1 port map( A => A_s(27), ZN => n648);
   U104 : INV_X1 port map( A => A_ns(28), ZN => n647);
   U105 : OAI221_X1 port map( B1 => n573, B2 => n650, C1 => n575, C2 => n651, A
                           => n652, ZN => O_27_port);
   U106 : AOI22_X1 port map( A1 => A_ns(25), A2 => n572, B1 => A_s(26), B2 => 
                           n578, ZN => n652);
   U107 : INV_X1 port map( A => A_s(25), ZN => n651);
   U108 : INV_X1 port map( A => A_ns(26), ZN => n650);
   U109 : OAI221_X1 port map( B1 => n573, B2 => n653, C1 => n575, C2 => n654, A
                           => n655, ZN => O_25_port);
   U110 : AOI22_X1 port map( A1 => A_ns(23), A2 => n572, B1 => A_s(24), B2 => 
                           n578, ZN => n655);
   U111 : INV_X1 port map( A => A_s(23), ZN => n654);
   U112 : INV_X1 port map( A => A_ns(24), ZN => n653);
   U113 : OAI221_X1 port map( B1 => n573, B2 => n656, C1 => n575, C2 => n657, A
                           => n658, ZN => O_23_port);
   U114 : AOI22_X1 port map( A1 => A_ns(21), A2 => n572, B1 => A_s(22), B2 => 
                           n578, ZN => n658);
   U115 : INV_X1 port map( A => A_s(21), ZN => n657);
   U116 : INV_X1 port map( A => A_ns(22), ZN => n656);
   U117 : OAI221_X1 port map( B1 => n573, B2 => n659, C1 => n575, C2 => n660, A
                           => n661, ZN => O_21_port);
   U118 : AOI22_X1 port map( A1 => A_ns(19), A2 => n572, B1 => A_s(20), B2 => 
                           n578, ZN => n661);
   U119 : INV_X1 port map( A => A_s(19), ZN => n660);
   U120 : INV_X1 port map( A => A_ns(20), ZN => n659);
   U121 : OAI221_X1 port map( B1 => n573, B2 => n662, C1 => n575, C2 => n663, A
                           => n664, ZN => O_19_port);
   U122 : AOI22_X1 port map( A1 => A_ns(17), A2 => n572, B1 => A_s(18), B2 => 
                           n578, ZN => n664);
   U123 : INV_X1 port map( A => A_s(17), ZN => n663);
   U124 : INV_X1 port map( A => A_ns(18), ZN => n662);
   U125 : OAI221_X1 port map( B1 => n573, B2 => n665, C1 => n575, C2 => n666, A
                           => n667, ZN => O_17_port);
   U126 : AOI22_X1 port map( A1 => A_ns(15), A2 => n572, B1 => A_s(16), B2 => 
                           n578, ZN => n667);
   U127 : INV_X1 port map( A => A_s(15), ZN => n666);
   U128 : INV_X1 port map( A => A_ns(16), ZN => n665);
   U129 : OAI221_X1 port map( B1 => n573, B2 => n668, C1 => n575, C2 => n669, A
                           => n670, ZN => O_15_port);
   U130 : AOI22_X1 port map( A1 => A_ns(13), A2 => n572, B1 => A_s(14), B2 => 
                           n578, ZN => n670);
   U131 : INV_X1 port map( A => A_s(13), ZN => n669);
   U132 : INV_X1 port map( A => A_ns(14), ZN => n668);
   U133 : OAI221_X1 port map( B1 => n573, B2 => n671, C1 => n575, C2 => n672, A
                           => n673, ZN => O_13_port);
   U134 : AOI22_X1 port map( A1 => A_ns(11), A2 => n572, B1 => A_s(12), B2 => 
                           n578, ZN => n673);
   U135 : INV_X1 port map( A => A_s(11), ZN => n672);
   U136 : INV_X1 port map( A => A_ns(12), ZN => n671);
   U137 : OAI221_X1 port map( B1 => n573, B2 => n674, C1 => n575, C2 => n675, A
                           => n676, ZN => O_11_port);
   U138 : AOI22_X1 port map( A1 => A_ns(9), A2 => n572, B1 => A_s(10), B2 => 
                           n578, ZN => n676);
   U139 : INV_X1 port map( A => A_s(9), ZN => n675);
   U140 : INV_X1 port map( A => A_ns(10), ZN => n674);
   U141 : OAI221_X1 port map( B1 => n573, B2 => n677, C1 => n575, C2 => n678, A
                           => n679, ZN => O_10_port);
   U142 : AOI22_X1 port map( A1 => A_ns(8), A2 => n572, B1 => A_s(9), B2 => 
                           n578, ZN => n679);
   U143 : NAND2_X1 port map( A1 => n680, A2 => n681, ZN => n622);
   U144 : INV_X1 port map( A => A_s(8), ZN => n678);
   U145 : INV_X1 port map( A => B(3), ZN => n681);
   U146 : INV_X1 port map( A => A_ns(9), ZN => n677);
   U147 : XOR2_X1 port map( A => B(1), B => B(2), Z => n680);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHENC_NBIT34_i0 is

   port( A_s, A_ns, B : in std_logic_vector (33 downto 0);  O, A_so, A_nso : 
         out std_logic_vector (33 downto 0));

end BOOTHENC_NBIT34_i0;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT34_i0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, n356, n357, n358, n359, n360, n361, n362, n363, n364, 
      n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, 
      n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, 
      n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, 
      n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, 
      n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, 
      n425, n426, n427, n428 : std_logic;

begin
   A_so <= ( A_s(32), A_s(31), A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), 
      A_s(25), A_s(24), A_s(23), A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), 
      A_s(17), A_s(16), A_s(15), A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), 
      A_s(9), A_s(8), A_s(7), A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), 
      A_s(0), X_Logic0_port );
   A_nso <= ( A_ns(32), A_ns(31), A_ns(30), A_ns(29), A_ns(28), A_ns(27), 
      A_ns(26), A_ns(25), A_ns(24), A_ns(23), A_ns(22), A_ns(21), A_ns(20), 
      A_ns(19), A_ns(18), A_ns(17), A_ns(16), A_ns(15), A_ns(14), A_ns(13), 
      A_ns(12), A_ns(11), A_ns(10), A_ns(9), A_ns(8), A_ns(7), A_ns(6), A_ns(5)
      , A_ns(4), A_ns(3), A_ns(2), A_ns(1), A_ns(0), X_Logic0_port );
   
   X_Logic0_port <= '0';
   U3 : NAND2_X2 port map( A1 => B(0), A2 => B(1), ZN => n358);
   U4 : INV_X2 port map( A => n375, ZN => n361);
   U5 : OR2_X2 port map( A1 => n427, A2 => B(0), ZN => n356);
   U6 : OAI221_X1 port map( B1 => n356, B2 => n357, C1 => n358, C2 => n359, A 
                           => n360, ZN => O(9));
   U7 : NAND2_X1 port map( A1 => A_s(9), A2 => n361, ZN => n360);
   U8 : OAI221_X1 port map( B1 => n356, B2 => n362, C1 => n357, C2 => n358, A 
                           => n363, ZN => O(8));
   U9 : NAND2_X1 port map( A1 => A_s(8), A2 => n361, ZN => n363);
   U10 : INV_X1 port map( A => A_ns(8), ZN => n357);
   U11 : OAI221_X1 port map( B1 => n356, B2 => n364, C1 => n358, C2 => n362, A 
                           => n365, ZN => O(7));
   U12 : NAND2_X1 port map( A1 => A_s(7), A2 => n361, ZN => n365);
   U13 : INV_X1 port map( A => A_ns(7), ZN => n362);
   U14 : OAI221_X1 port map( B1 => n356, B2 => n366, C1 => n358, C2 => n364, A 
                           => n367, ZN => O(6));
   U15 : NAND2_X1 port map( A1 => A_s(6), A2 => n361, ZN => n367);
   U16 : INV_X1 port map( A => A_ns(6), ZN => n364);
   U17 : OAI221_X1 port map( B1 => n356, B2 => n368, C1 => n358, C2 => n366, A 
                           => n369, ZN => O(5));
   U18 : NAND2_X1 port map( A1 => A_s(5), A2 => n361, ZN => n369);
   U19 : INV_X1 port map( A => A_ns(5), ZN => n366);
   U20 : OAI221_X1 port map( B1 => n356, B2 => n370, C1 => n358, C2 => n368, A 
                           => n371, ZN => O(4));
   U21 : NAND2_X1 port map( A1 => A_s(4), A2 => n361, ZN => n371);
   U22 : INV_X1 port map( A => A_ns(4), ZN => n368);
   U23 : OAI221_X1 port map( B1 => n356, B2 => n372, C1 => n358, C2 => n370, A 
                           => n373, ZN => O(3));
   U24 : NAND2_X1 port map( A1 => A_s(3), A2 => n361, ZN => n373);
   U25 : INV_X1 port map( A => A_ns(3), ZN => n370);
   U26 : OAI222_X1 port map( A1 => n374, A2 => n375, B1 => n376, B2 => n356, C1
                           => n377, C2 => n358, ZN => O(33));
   U27 : INV_X1 port map( A => A_ns(33), ZN => n377);
   U28 : INV_X1 port map( A => A_s(33), ZN => n374);
   U29 : OAI221_X1 port map( B1 => n356, B2 => n378, C1 => n358, C2 => n376, A 
                           => n379, ZN => O(32));
   U30 : NAND2_X1 port map( A1 => A_s(32), A2 => n361, ZN => n379);
   U31 : INV_X1 port map( A => A_ns(32), ZN => n376);
   U32 : OAI221_X1 port map( B1 => n356, B2 => n380, C1 => n358, C2 => n378, A 
                           => n381, ZN => O(31));
   U33 : NAND2_X1 port map( A1 => A_s(31), A2 => n361, ZN => n381);
   U34 : INV_X1 port map( A => A_ns(31), ZN => n378);
   U35 : OAI221_X1 port map( B1 => n356, B2 => n382, C1 => n358, C2 => n380, A 
                           => n383, ZN => O(30));
   U36 : NAND2_X1 port map( A1 => A_s(30), A2 => n361, ZN => n383);
   U37 : INV_X1 port map( A => A_ns(30), ZN => n380);
   U38 : OAI221_X1 port map( B1 => n356, B2 => n384, C1 => n358, C2 => n372, A 
                           => n385, ZN => O(2));
   U39 : NAND2_X1 port map( A1 => A_s(2), A2 => n361, ZN => n385);
   U40 : INV_X1 port map( A => A_ns(2), ZN => n372);
   U41 : OAI221_X1 port map( B1 => n356, B2 => n386, C1 => n358, C2 => n382, A 
                           => n387, ZN => O(29));
   U42 : NAND2_X1 port map( A1 => A_s(29), A2 => n361, ZN => n387);
   U43 : INV_X1 port map( A => A_ns(29), ZN => n382);
   U44 : OAI221_X1 port map( B1 => n356, B2 => n388, C1 => n358, C2 => n386, A 
                           => n389, ZN => O(28));
   U45 : NAND2_X1 port map( A1 => A_s(28), A2 => n361, ZN => n389);
   U46 : INV_X1 port map( A => A_ns(28), ZN => n386);
   U47 : OAI221_X1 port map( B1 => n356, B2 => n390, C1 => n358, C2 => n388, A 
                           => n391, ZN => O(27));
   U48 : NAND2_X1 port map( A1 => A_s(27), A2 => n361, ZN => n391);
   U49 : INV_X1 port map( A => A_ns(27), ZN => n388);
   U50 : OAI221_X1 port map( B1 => n356, B2 => n392, C1 => n358, C2 => n390, A 
                           => n393, ZN => O(26));
   U51 : NAND2_X1 port map( A1 => A_s(26), A2 => n361, ZN => n393);
   U52 : INV_X1 port map( A => A_ns(26), ZN => n390);
   U53 : OAI221_X1 port map( B1 => n356, B2 => n394, C1 => n358, C2 => n392, A 
                           => n395, ZN => O(25));
   U54 : NAND2_X1 port map( A1 => A_s(25), A2 => n361, ZN => n395);
   U55 : INV_X1 port map( A => A_ns(25), ZN => n392);
   U56 : OAI221_X1 port map( B1 => n356, B2 => n396, C1 => n358, C2 => n394, A 
                           => n397, ZN => O(24));
   U57 : NAND2_X1 port map( A1 => A_s(24), A2 => n361, ZN => n397);
   U58 : INV_X1 port map( A => A_ns(24), ZN => n394);
   U59 : OAI221_X1 port map( B1 => n356, B2 => n398, C1 => n358, C2 => n396, A 
                           => n399, ZN => O(23));
   U60 : NAND2_X1 port map( A1 => A_s(23), A2 => n361, ZN => n399);
   U61 : INV_X1 port map( A => A_ns(23), ZN => n396);
   U62 : OAI221_X1 port map( B1 => n356, B2 => n400, C1 => n358, C2 => n398, A 
                           => n401, ZN => O(22));
   U63 : NAND2_X1 port map( A1 => A_s(22), A2 => n361, ZN => n401);
   U64 : INV_X1 port map( A => A_ns(22), ZN => n398);
   U65 : OAI221_X1 port map( B1 => n356, B2 => n402, C1 => n358, C2 => n400, A 
                           => n403, ZN => O(21));
   U66 : NAND2_X1 port map( A1 => A_s(21), A2 => n361, ZN => n403);
   U67 : INV_X1 port map( A => A_ns(21), ZN => n400);
   U68 : OAI221_X1 port map( B1 => n356, B2 => n404, C1 => n358, C2 => n402, A 
                           => n405, ZN => O(20));
   U69 : NAND2_X1 port map( A1 => A_s(20), A2 => n361, ZN => n405);
   U70 : INV_X1 port map( A => A_ns(20), ZN => n402);
   U71 : OAI221_X1 port map( B1 => n356, B2 => n406, C1 => n358, C2 => n384, A 
                           => n407, ZN => O(1));
   U72 : NAND2_X1 port map( A1 => A_s(1), A2 => n361, ZN => n407);
   U73 : INV_X1 port map( A => A_ns(1), ZN => n384);
   U74 : OAI221_X1 port map( B1 => n356, B2 => n408, C1 => n358, C2 => n404, A 
                           => n409, ZN => O(19));
   U75 : NAND2_X1 port map( A1 => A_s(19), A2 => n361, ZN => n409);
   U76 : INV_X1 port map( A => A_ns(19), ZN => n404);
   U77 : OAI221_X1 port map( B1 => n356, B2 => n410, C1 => n358, C2 => n408, A 
                           => n411, ZN => O(18));
   U78 : NAND2_X1 port map( A1 => A_s(18), A2 => n361, ZN => n411);
   U79 : INV_X1 port map( A => A_ns(18), ZN => n408);
   U80 : OAI221_X1 port map( B1 => n356, B2 => n412, C1 => n358, C2 => n410, A 
                           => n413, ZN => O(17));
   U81 : NAND2_X1 port map( A1 => A_s(17), A2 => n361, ZN => n413);
   U82 : INV_X1 port map( A => A_ns(17), ZN => n410);
   U83 : OAI221_X1 port map( B1 => n356, B2 => n414, C1 => n358, C2 => n412, A 
                           => n415, ZN => O(16));
   U84 : NAND2_X1 port map( A1 => A_s(16), A2 => n361, ZN => n415);
   U85 : INV_X1 port map( A => A_ns(16), ZN => n412);
   U86 : OAI221_X1 port map( B1 => n356, B2 => n416, C1 => n358, C2 => n414, A 
                           => n417, ZN => O(15));
   U87 : NAND2_X1 port map( A1 => A_s(15), A2 => n361, ZN => n417);
   U88 : INV_X1 port map( A => A_ns(15), ZN => n414);
   U89 : OAI221_X1 port map( B1 => n356, B2 => n418, C1 => n358, C2 => n416, A 
                           => n419, ZN => O(14));
   U90 : NAND2_X1 port map( A1 => A_s(14), A2 => n361, ZN => n419);
   U91 : INV_X1 port map( A => A_ns(14), ZN => n416);
   U92 : OAI221_X1 port map( B1 => n356, B2 => n420, C1 => n358, C2 => n418, A 
                           => n421, ZN => O(13));
   U93 : NAND2_X1 port map( A1 => A_s(13), A2 => n361, ZN => n421);
   U94 : INV_X1 port map( A => A_ns(13), ZN => n418);
   U95 : OAI221_X1 port map( B1 => n356, B2 => n422, C1 => n358, C2 => n420, A 
                           => n423, ZN => O(12));
   U96 : NAND2_X1 port map( A1 => A_s(12), A2 => n361, ZN => n423);
   U97 : INV_X1 port map( A => A_ns(12), ZN => n420);
   U98 : OAI221_X1 port map( B1 => n356, B2 => n424, C1 => n358, C2 => n422, A 
                           => n425, ZN => O(11));
   U99 : NAND2_X1 port map( A1 => A_s(11), A2 => n361, ZN => n425);
   U100 : INV_X1 port map( A => A_ns(11), ZN => n422);
   U101 : OAI221_X1 port map( B1 => n356, B2 => n359, C1 => n358, C2 => n424, A
                           => n426, ZN => O(10));
   U102 : NAND2_X1 port map( A1 => A_s(10), A2 => n361, ZN => n426);
   U103 : INV_X1 port map( A => A_ns(10), ZN => n424);
   U104 : INV_X1 port map( A => A_ns(9), ZN => n359);
   U105 : OAI22_X1 port map( A1 => n375, A2 => n428, B1 => n358, B2 => n406, ZN
                           => O(0));
   U106 : INV_X1 port map( A => A_ns(0), ZN => n406);
   U107 : INV_X1 port map( A => A_s(0), ZN => n428);
   U108 : NAND2_X1 port map( A1 => B(0), A2 => n427, ZN => n375);
   U109 : INV_X1 port map( A => B(1), ZN => n427);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32.all;

entity BOOTHMUL_NBIT32 is

   port( A, B : in std_logic_vector (31 downto 0);  S : out std_logic_vector 
         (63 downto 0));

end BOOTHMUL_NBIT32;

architecture SYN_BEHAVIOURAL of BOOTHMUL_NBIT32 is

   component BOOTHMUL_NBIT32_DW01_sub_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component RCA_NBIT64
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT62
      port( A, B : in std_logic_vector (61 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (61 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT60
      port( A, B : in std_logic_vector (59 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (59 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT58
      port( A, B : in std_logic_vector (57 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (57 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT56
      port( A, B : in std_logic_vector (55 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (55 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT54
      port( A, B : in std_logic_vector (53 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (53 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT52
      port( A, B : in std_logic_vector (51 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (51 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT50
      port( A, B : in std_logic_vector (49 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (49 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT48
      port( A, B : in std_logic_vector (47 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (47 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT46
      port( A, B : in std_logic_vector (45 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (45 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT44
      port( A, B : in std_logic_vector (43 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (43 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT42
      port( A, B : in std_logic_vector (41 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (41 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT40
      port( A, B : in std_logic_vector (39 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (39 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT38
      port( A, B : in std_logic_vector (37 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (37 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT36
      port( A, B : in std_logic_vector (35 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (35 downto 0);  Co : out std_logic);
   end component;
   
   component BOOTHENC_NBIT64_i30
      port( A_s, A_ns, B : in std_logic_vector (63 downto 0);  O, A_so, A_nso :
            out std_logic_vector (63 downto 0));
   end component;
   
   component BOOTHENC_NBIT62_i28
      port( A_s, A_ns, B : in std_logic_vector (61 downto 0);  O, A_so, A_nso :
            out std_logic_vector (61 downto 0));
   end component;
   
   component BOOTHENC_NBIT60_i26
      port( A_s, A_ns, B : in std_logic_vector (59 downto 0);  O, A_so, A_nso :
            out std_logic_vector (59 downto 0));
   end component;
   
   component BOOTHENC_NBIT58_i24
      port( A_s, A_ns, B : in std_logic_vector (57 downto 0);  O, A_so, A_nso :
            out std_logic_vector (57 downto 0));
   end component;
   
   component BOOTHENC_NBIT56_i22
      port( A_s, A_ns, B : in std_logic_vector (55 downto 0);  O, A_so, A_nso :
            out std_logic_vector (55 downto 0));
   end component;
   
   component BOOTHENC_NBIT54_i20
      port( A_s, A_ns, B : in std_logic_vector (53 downto 0);  O, A_so, A_nso :
            out std_logic_vector (53 downto 0));
   end component;
   
   component BOOTHENC_NBIT52_i18
      port( A_s, A_ns, B : in std_logic_vector (51 downto 0);  O, A_so, A_nso :
            out std_logic_vector (51 downto 0));
   end component;
   
   component BOOTHENC_NBIT50_i16
      port( A_s, A_ns, B : in std_logic_vector (49 downto 0);  O, A_so, A_nso :
            out std_logic_vector (49 downto 0));
   end component;
   
   component BOOTHENC_NBIT48_i14
      port( A_s, A_ns, B : in std_logic_vector (47 downto 0);  O, A_so, A_nso :
            out std_logic_vector (47 downto 0));
   end component;
   
   component BOOTHENC_NBIT46_i12
      port( A_s, A_ns, B : in std_logic_vector (45 downto 0);  O, A_so, A_nso :
            out std_logic_vector (45 downto 0));
   end component;
   
   component BOOTHENC_NBIT44_i10
      port( A_s, A_ns, B : in std_logic_vector (43 downto 0);  O, A_so, A_nso :
            out std_logic_vector (43 downto 0));
   end component;
   
   component BOOTHENC_NBIT42_i8
      port( A_s, A_ns, B : in std_logic_vector (41 downto 0);  O, A_so, A_nso :
            out std_logic_vector (41 downto 0));
   end component;
   
   component BOOTHENC_NBIT40_i6
      port( A_s, A_ns, B : in std_logic_vector (39 downto 0);  O, A_so, A_nso :
            out std_logic_vector (39 downto 0));
   end component;
   
   component BOOTHENC_NBIT38_i4
      port( A_s, A_ns, B : in std_logic_vector (37 downto 0);  O, A_so, A_nso :
            out std_logic_vector (37 downto 0));
   end component;
   
   component BOOTHENC_NBIT36_i2
      port( A_s, A_ns, B : in std_logic_vector (35 downto 0);  O, A_so, A_nso :
            out std_logic_vector (35 downto 0));
   end component;
   
   component BOOTHENC_NBIT34_i0
      port( A_s, A_ns, B : in std_logic_vector (33 downto 0);  O, A_so, A_nso :
            out std_logic_vector (33 downto 0));
   end component;
   
   signal X_Logic0_port, A_n_65, A_n_30_port, A_n_29_port, A_n_28_port, 
      A_n_27_port, A_n_26_port, A_n_25_port, A_n_24_port, A_n_23_port, 
      A_n_22_port, A_n_21_port, A_n_20_port, A_n_19_port, A_n_18_port, 
      A_n_17_port, A_n_16_port, A_n_15_port, A_n_14_port, A_n_13_port, 
      A_n_12_port, A_n_11_port, A_n_10_port, A_n_9_port, A_n_8_port, A_n_7_port
      , A_n_6_port, A_n_5_port, A_n_4_port, A_n_3_port, A_n_2_port, A_n_1_port,
      A_n_0_port, SHIFT_1_31_port, SHIFT_1_30_port, SHIFT_1_29_port, 
      SHIFT_1_28_port, SHIFT_1_27_port, SHIFT_1_26_port, SHIFT_1_25_port, 
      SHIFT_1_24_port, SHIFT_1_23_port, SHIFT_1_22_port, SHIFT_1_21_port, 
      SHIFT_1_20_port, SHIFT_1_19_port, SHIFT_1_18_port, SHIFT_1_17_port, 
      SHIFT_1_16_port, SHIFT_1_15_port, SHIFT_1_14_port, SHIFT_1_13_port, 
      SHIFT_1_12_port, SHIFT_1_11_port, SHIFT_1_10_port, SHIFT_1_9_port, 
      SHIFT_1_8_port, SHIFT_1_7_port, SHIFT_1_6_port, SHIFT_1_5_port, 
      SHIFT_1_4_port, SHIFT_1_3_port, SHIFT_1_2_port, SHIFT_1_1_port, 
      SHIFT_1_0_port, SHIFT_15_61_port, SHIFT_15_60_port, SHIFT_15_59_port, 
      SHIFT_15_58_port, SHIFT_15_57_port, SHIFT_15_56_port, SHIFT_15_55_port, 
      SHIFT_15_54_port, SHIFT_15_53_port, SHIFT_15_52_port, SHIFT_15_51_port, 
      SHIFT_15_50_port, SHIFT_15_49_port, SHIFT_15_48_port, SHIFT_15_47_port, 
      SHIFT_15_46_port, SHIFT_15_45_port, SHIFT_15_44_port, SHIFT_15_43_port, 
      SHIFT_15_42_port, SHIFT_15_41_port, SHIFT_15_40_port, SHIFT_15_39_port, 
      SHIFT_15_38_port, SHIFT_15_37_port, SHIFT_15_36_port, SHIFT_15_35_port, 
      SHIFT_15_34_port, SHIFT_15_33_port, SHIFT_15_32_port, SHIFT_15_31_port, 
      SHIFT_15_30_port, SHIFT_15_29_port, SHIFT_15_28_port, SHIFT_15_27_port, 
      SHIFT_15_26_port, SHIFT_15_25_port, SHIFT_15_24_port, SHIFT_15_23_port, 
      SHIFT_15_22_port, SHIFT_15_21_port, SHIFT_15_20_port, SHIFT_15_19_port, 
      SHIFT_15_18_port, SHIFT_15_17_port, SHIFT_15_16_port, SHIFT_15_15_port, 
      SHIFT_15_14_port, SHIFT_15_13_port, SHIFT_15_12_port, SHIFT_15_11_port, 
      SHIFT_15_10_port, SHIFT_15_9_port, SHIFT_15_8_port, SHIFT_15_7_port, 
      SHIFT_15_6_port, SHIFT_15_5_port, SHIFT_15_4_port, SHIFT_15_3_port, 
      SHIFT_15_2_port, SHIFT_15_1_port, SHIFT_15_0_port, SHIFT_14_59_port, 
      SHIFT_14_58_port, SHIFT_14_57_port, SHIFT_14_56_port, SHIFT_14_55_port, 
      SHIFT_14_54_port, SHIFT_14_53_port, SHIFT_14_52_port, SHIFT_14_51_port, 
      SHIFT_14_50_port, SHIFT_14_49_port, SHIFT_14_48_port, SHIFT_14_47_port, 
      SHIFT_14_46_port, SHIFT_14_45_port, SHIFT_14_44_port, SHIFT_14_43_port, 
      SHIFT_14_42_port, SHIFT_14_41_port, SHIFT_14_40_port, SHIFT_14_39_port, 
      SHIFT_14_38_port, SHIFT_14_37_port, SHIFT_14_36_port, SHIFT_14_35_port, 
      SHIFT_14_34_port, SHIFT_14_33_port, SHIFT_14_32_port, SHIFT_14_31_port, 
      SHIFT_14_30_port, SHIFT_14_29_port, SHIFT_14_28_port, SHIFT_14_27_port, 
      SHIFT_14_26_port, SHIFT_14_25_port, SHIFT_14_24_port, SHIFT_14_23_port, 
      SHIFT_14_22_port, SHIFT_14_21_port, SHIFT_14_20_port, SHIFT_14_19_port, 
      SHIFT_14_18_port, SHIFT_14_17_port, SHIFT_14_16_port, SHIFT_14_15_port, 
      SHIFT_14_14_port, SHIFT_14_13_port, SHIFT_14_12_port, SHIFT_14_11_port, 
      SHIFT_14_10_port, SHIFT_14_9_port, SHIFT_14_8_port, SHIFT_14_7_port, 
      SHIFT_14_6_port, SHIFT_14_5_port, SHIFT_14_4_port, SHIFT_14_3_port, 
      SHIFT_14_2_port, SHIFT_14_1_port, SHIFT_14_0_port, SHIFT_13_57_port, 
      SHIFT_13_56_port, SHIFT_13_55_port, SHIFT_13_54_port, SHIFT_13_53_port, 
      SHIFT_13_52_port, SHIFT_13_51_port, SHIFT_13_50_port, SHIFT_13_49_port, 
      SHIFT_13_48_port, SHIFT_13_47_port, SHIFT_13_46_port, SHIFT_13_45_port, 
      SHIFT_13_44_port, SHIFT_13_43_port, SHIFT_13_42_port, SHIFT_13_41_port, 
      SHIFT_13_40_port, SHIFT_13_39_port, SHIFT_13_38_port, SHIFT_13_37_port, 
      SHIFT_13_36_port, SHIFT_13_35_port, SHIFT_13_34_port, SHIFT_13_33_port, 
      SHIFT_13_32_port, SHIFT_13_31_port, SHIFT_13_30_port, SHIFT_13_29_port, 
      SHIFT_13_28_port, SHIFT_13_27_port, SHIFT_13_26_port, SHIFT_13_25_port, 
      SHIFT_13_24_port, SHIFT_13_23_port, SHIFT_13_22_port, SHIFT_13_21_port, 
      SHIFT_13_20_port, SHIFT_13_19_port, SHIFT_13_18_port, SHIFT_13_17_port, 
      SHIFT_13_16_port, SHIFT_13_15_port, SHIFT_13_14_port, SHIFT_13_13_port, 
      SHIFT_13_12_port, SHIFT_13_11_port, SHIFT_13_10_port, SHIFT_13_9_port, 
      SHIFT_13_8_port, SHIFT_13_7_port, SHIFT_13_6_port, SHIFT_13_5_port, 
      SHIFT_13_4_port, SHIFT_13_3_port, SHIFT_13_2_port, SHIFT_13_1_port, 
      SHIFT_13_0_port, SHIFT_12_55_port, SHIFT_12_54_port, SHIFT_12_53_port, 
      SHIFT_12_52_port, SHIFT_12_51_port, SHIFT_12_50_port, SHIFT_12_49_port, 
      SHIFT_12_48_port, SHIFT_12_47_port, SHIFT_12_46_port, SHIFT_12_45_port, 
      SHIFT_12_44_port, SHIFT_12_43_port, SHIFT_12_42_port, SHIFT_12_41_port, 
      SHIFT_12_40_port, SHIFT_12_39_port, SHIFT_12_38_port, SHIFT_12_37_port, 
      SHIFT_12_36_port, SHIFT_12_35_port, SHIFT_12_34_port, SHIFT_12_33_port, 
      SHIFT_12_32_port, SHIFT_12_31_port, SHIFT_12_30_port, SHIFT_12_29_port, 
      SHIFT_12_28_port, SHIFT_12_27_port, SHIFT_12_26_port, SHIFT_12_25_port, 
      SHIFT_12_24_port, SHIFT_12_23_port, SHIFT_12_22_port, SHIFT_12_21_port, 
      SHIFT_12_20_port, SHIFT_12_19_port, SHIFT_12_18_port, SHIFT_12_17_port, 
      SHIFT_12_16_port, SHIFT_12_15_port, SHIFT_12_14_port, SHIFT_12_13_port, 
      SHIFT_12_12_port, SHIFT_12_11_port, SHIFT_12_10_port, SHIFT_12_9_port, 
      SHIFT_12_8_port, SHIFT_12_7_port, SHIFT_12_6_port, SHIFT_12_5_port, 
      SHIFT_12_4_port, SHIFT_12_3_port, SHIFT_12_2_port, SHIFT_12_1_port, 
      SHIFT_12_0_port, SHIFT_11_53_port, SHIFT_11_52_port, SHIFT_11_51_port, 
      SHIFT_11_50_port, SHIFT_11_49_port, SHIFT_11_48_port, SHIFT_11_47_port, 
      SHIFT_11_46_port, SHIFT_11_45_port, SHIFT_11_44_port, SHIFT_11_43_port, 
      SHIFT_11_42_port, SHIFT_11_41_port, SHIFT_11_40_port, SHIFT_11_39_port, 
      SHIFT_11_38_port, SHIFT_11_37_port, SHIFT_11_36_port, SHIFT_11_35_port, 
      SHIFT_11_34_port, SHIFT_11_33_port, SHIFT_11_32_port, SHIFT_11_31_port, 
      SHIFT_11_30_port, SHIFT_11_29_port, SHIFT_11_28_port, SHIFT_11_27_port, 
      SHIFT_11_26_port, SHIFT_11_25_port, SHIFT_11_24_port, SHIFT_11_23_port, 
      SHIFT_11_22_port, SHIFT_11_21_port, SHIFT_11_20_port, SHIFT_11_19_port, 
      SHIFT_11_18_port, SHIFT_11_17_port, SHIFT_11_16_port, SHIFT_11_15_port, 
      SHIFT_11_14_port, SHIFT_11_13_port, SHIFT_11_12_port, SHIFT_11_11_port, 
      SHIFT_11_10_port, SHIFT_11_9_port, SHIFT_11_8_port, SHIFT_11_7_port, 
      SHIFT_11_6_port, SHIFT_11_5_port, SHIFT_11_4_port, SHIFT_11_3_port, 
      SHIFT_11_2_port, SHIFT_11_1_port, SHIFT_11_0_port, SHIFT_10_51_port, 
      SHIFT_10_50_port, SHIFT_10_49_port, SHIFT_10_48_port, SHIFT_10_47_port, 
      SHIFT_10_46_port, SHIFT_10_45_port, SHIFT_10_44_port, SHIFT_10_43_port, 
      SHIFT_10_42_port, SHIFT_10_41_port, SHIFT_10_40_port, SHIFT_10_39_port, 
      SHIFT_10_38_port, SHIFT_10_37_port, SHIFT_10_36_port, SHIFT_10_35_port, 
      SHIFT_10_34_port, SHIFT_10_33_port, SHIFT_10_32_port, SHIFT_10_31_port, 
      SHIFT_10_30_port, SHIFT_10_29_port, SHIFT_10_28_port, SHIFT_10_27_port, 
      SHIFT_10_26_port, SHIFT_10_25_port, SHIFT_10_24_port, SHIFT_10_23_port, 
      SHIFT_10_22_port, SHIFT_10_21_port, SHIFT_10_20_port, SHIFT_10_19_port, 
      SHIFT_10_18_port, SHIFT_10_17_port, SHIFT_10_16_port, SHIFT_10_15_port, 
      SHIFT_10_14_port, SHIFT_10_13_port, SHIFT_10_12_port, SHIFT_10_11_port, 
      SHIFT_10_10_port, SHIFT_10_9_port, SHIFT_10_8_port, SHIFT_10_7_port, 
      SHIFT_10_6_port, SHIFT_10_5_port, SHIFT_10_4_port, SHIFT_10_3_port, 
      SHIFT_10_2_port, SHIFT_10_1_port, SHIFT_10_0_port, SHIFT_9_49_port, 
      SHIFT_9_48_port, SHIFT_9_47_port, SHIFT_9_46_port, SHIFT_9_45_port, 
      SHIFT_9_44_port, SHIFT_9_43_port, SHIFT_9_42_port, SHIFT_9_41_port, 
      SHIFT_9_40_port, SHIFT_9_39_port, SHIFT_9_38_port, SHIFT_9_37_port, 
      SHIFT_9_36_port, SHIFT_9_35_port, SHIFT_9_34_port, SHIFT_9_33_port, 
      SHIFT_9_32_port, SHIFT_9_31_port, SHIFT_9_30_port, SHIFT_9_29_port, 
      SHIFT_9_28_port, SHIFT_9_27_port, SHIFT_9_26_port, SHIFT_9_25_port, 
      SHIFT_9_24_port, SHIFT_9_23_port, SHIFT_9_22_port, SHIFT_9_21_port, 
      SHIFT_9_20_port, SHIFT_9_19_port, SHIFT_9_18_port, SHIFT_9_17_port, 
      SHIFT_9_16_port, SHIFT_9_15_port, SHIFT_9_14_port, SHIFT_9_13_port, 
      SHIFT_9_12_port, SHIFT_9_11_port, SHIFT_9_10_port, SHIFT_9_9_port, 
      SHIFT_9_8_port, SHIFT_9_7_port, SHIFT_9_6_port, SHIFT_9_5_port, 
      SHIFT_9_4_port, SHIFT_9_3_port, SHIFT_9_2_port, SHIFT_9_1_port, 
      SHIFT_9_0_port, SHIFT_8_47_port, SHIFT_8_46_port, SHIFT_8_45_port, 
      SHIFT_8_44_port, SHIFT_8_43_port, SHIFT_8_42_port, SHIFT_8_41_port, 
      SHIFT_8_40_port, SHIFT_8_39_port, SHIFT_8_38_port, SHIFT_8_37_port, 
      SHIFT_8_36_port, SHIFT_8_35_port, SHIFT_8_34_port, SHIFT_8_33_port, 
      SHIFT_8_32_port, SHIFT_8_31_port, SHIFT_8_30_port, SHIFT_8_29_port, 
      SHIFT_8_28_port, SHIFT_8_27_port, SHIFT_8_26_port, SHIFT_8_25_port, 
      SHIFT_8_24_port, SHIFT_8_23_port, SHIFT_8_22_port, SHIFT_8_21_port, 
      SHIFT_8_20_port, SHIFT_8_19_port, SHIFT_8_18_port, SHIFT_8_17_port, 
      SHIFT_8_16_port, SHIFT_8_15_port, SHIFT_8_14_port, SHIFT_8_13_port, 
      SHIFT_8_12_port, SHIFT_8_11_port, SHIFT_8_10_port, SHIFT_8_9_port, 
      SHIFT_8_8_port, SHIFT_8_7_port, SHIFT_8_6_port, SHIFT_8_5_port, 
      SHIFT_8_4_port, SHIFT_8_3_port, SHIFT_8_2_port, SHIFT_8_1_port, 
      SHIFT_8_0_port, SHIFT_7_45_port, SHIFT_7_44_port, SHIFT_7_43_port, 
      SHIFT_7_42_port, SHIFT_7_41_port, SHIFT_7_40_port, SHIFT_7_39_port, 
      SHIFT_7_38_port, SHIFT_7_37_port, SHIFT_7_36_port, SHIFT_7_35_port, 
      SHIFT_7_34_port, SHIFT_7_33_port, SHIFT_7_32_port, SHIFT_7_31_port, 
      SHIFT_7_30_port, SHIFT_7_29_port, SHIFT_7_28_port, SHIFT_7_27_port, 
      SHIFT_7_26_port, SHIFT_7_25_port, SHIFT_7_24_port, SHIFT_7_23_port, 
      SHIFT_7_22_port, SHIFT_7_21_port, SHIFT_7_20_port, SHIFT_7_19_port, 
      SHIFT_7_18_port, SHIFT_7_17_port, SHIFT_7_16_port, SHIFT_7_15_port, 
      SHIFT_7_14_port, SHIFT_7_13_port, SHIFT_7_12_port, SHIFT_7_11_port, 
      SHIFT_7_10_port, SHIFT_7_9_port, SHIFT_7_8_port, SHIFT_7_7_port, 
      SHIFT_7_6_port, SHIFT_7_5_port, SHIFT_7_4_port, SHIFT_7_3_port, 
      SHIFT_7_2_port, SHIFT_7_1_port, SHIFT_7_0_port, SHIFT_6_43_port, 
      SHIFT_6_42_port, SHIFT_6_41_port, SHIFT_6_40_port, SHIFT_6_39_port, 
      SHIFT_6_38_port, SHIFT_6_37_port, SHIFT_6_36_port, SHIFT_6_35_port, 
      SHIFT_6_34_port, SHIFT_6_33_port, SHIFT_6_32_port, SHIFT_6_31_port, 
      SHIFT_6_30_port, SHIFT_6_29_port, SHIFT_6_28_port, SHIFT_6_27_port, 
      SHIFT_6_26_port, SHIFT_6_25_port, SHIFT_6_24_port, SHIFT_6_23_port, 
      SHIFT_6_22_port, SHIFT_6_21_port, SHIFT_6_20_port, SHIFT_6_19_port, 
      SHIFT_6_18_port, SHIFT_6_17_port, SHIFT_6_16_port, SHIFT_6_15_port, 
      SHIFT_6_14_port, SHIFT_6_13_port, SHIFT_6_12_port, SHIFT_6_11_port, 
      SHIFT_6_10_port, SHIFT_6_9_port, SHIFT_6_8_port, SHIFT_6_7_port, 
      SHIFT_6_6_port, SHIFT_6_5_port, SHIFT_6_4_port, SHIFT_6_3_port, 
      SHIFT_6_2_port, SHIFT_6_1_port, SHIFT_6_0_port, SHIFT_5_41_port, 
      SHIFT_5_40_port, SHIFT_5_39_port, SHIFT_5_38_port, SHIFT_5_37_port, 
      SHIFT_5_36_port, SHIFT_5_35_port, SHIFT_5_34_port, SHIFT_5_33_port, 
      SHIFT_5_32_port, SHIFT_5_31_port, SHIFT_5_30_port, SHIFT_5_29_port, 
      SHIFT_5_28_port, SHIFT_5_27_port, SHIFT_5_26_port, SHIFT_5_25_port, 
      SHIFT_5_24_port, SHIFT_5_23_port, SHIFT_5_22_port, SHIFT_5_21_port, 
      SHIFT_5_20_port, SHIFT_5_19_port, SHIFT_5_18_port, SHIFT_5_17_port, 
      SHIFT_5_16_port, SHIFT_5_15_port, SHIFT_5_14_port, SHIFT_5_13_port, 
      SHIFT_5_12_port, SHIFT_5_11_port, SHIFT_5_10_port, SHIFT_5_9_port, 
      SHIFT_5_8_port, SHIFT_5_7_port, SHIFT_5_6_port, SHIFT_5_5_port, 
      SHIFT_5_4_port, SHIFT_5_3_port, SHIFT_5_2_port, SHIFT_5_1_port, 
      SHIFT_5_0_port, SHIFT_4_39_port, SHIFT_4_38_port, SHIFT_4_37_port, 
      SHIFT_4_36_port, SHIFT_4_35_port, SHIFT_4_34_port, SHIFT_4_33_port, 
      SHIFT_4_32_port, SHIFT_4_31_port, SHIFT_4_30_port, SHIFT_4_29_port, 
      SHIFT_4_28_port, SHIFT_4_27_port, SHIFT_4_26_port, SHIFT_4_25_port, 
      SHIFT_4_24_port, SHIFT_4_23_port, SHIFT_4_22_port, SHIFT_4_21_port, 
      SHIFT_4_20_port, SHIFT_4_19_port, SHIFT_4_18_port, SHIFT_4_17_port, 
      SHIFT_4_16_port, SHIFT_4_15_port, SHIFT_4_14_port, SHIFT_4_13_port, 
      SHIFT_4_12_port, SHIFT_4_11_port, SHIFT_4_10_port, SHIFT_4_9_port, 
      SHIFT_4_8_port, SHIFT_4_7_port, SHIFT_4_6_port, SHIFT_4_5_port, 
      SHIFT_4_4_port, SHIFT_4_3_port, SHIFT_4_2_port, SHIFT_4_1_port, 
      SHIFT_4_0_port, SHIFT_3_37_port, SHIFT_3_36_port, SHIFT_3_35_port, 
      SHIFT_3_34_port, SHIFT_3_33_port, SHIFT_3_32_port, SHIFT_3_31_port, 
      SHIFT_3_30_port, SHIFT_3_29_port, SHIFT_3_28_port, SHIFT_3_27_port, 
      SHIFT_3_26_port, SHIFT_3_25_port, SHIFT_3_24_port, SHIFT_3_23_port, 
      SHIFT_3_22_port, SHIFT_3_21_port, SHIFT_3_20_port, SHIFT_3_19_port, 
      SHIFT_3_18_port, SHIFT_3_17_port, SHIFT_3_16_port, SHIFT_3_15_port, 
      SHIFT_3_14_port, SHIFT_3_13_port, SHIFT_3_12_port, SHIFT_3_11_port, 
      SHIFT_3_10_port, SHIFT_3_9_port, SHIFT_3_8_port, SHIFT_3_7_port, 
      SHIFT_3_6_port, SHIFT_3_5_port, SHIFT_3_4_port, SHIFT_3_3_port, 
      SHIFT_3_2_port, SHIFT_3_1_port, SHIFT_3_0_port, SHIFT_2_35_port, 
      SHIFT_2_34_port, SHIFT_2_33_port, SHIFT_2_32_port, SHIFT_2_31_port, 
      SHIFT_2_30_port, SHIFT_2_29_port, SHIFT_2_28_port, SHIFT_2_27_port, 
      SHIFT_2_26_port, SHIFT_2_25_port, SHIFT_2_24_port, SHIFT_2_23_port, 
      SHIFT_2_22_port, SHIFT_2_21_port, SHIFT_2_20_port, SHIFT_2_19_port, 
      SHIFT_2_18_port, SHIFT_2_17_port, SHIFT_2_16_port, SHIFT_2_15_port, 
      SHIFT_2_14_port, SHIFT_2_13_port, SHIFT_2_12_port, SHIFT_2_11_port, 
      SHIFT_2_10_port, SHIFT_2_9_port, SHIFT_2_8_port, SHIFT_2_7_port, 
      SHIFT_2_6_port, SHIFT_2_5_port, SHIFT_2_4_port, SHIFT_2_3_port, 
      SHIFT_2_2_port, SHIFT_2_1_port, SHIFT_2_0_port, SHIFT_1_33_port, 
      SHIFT_1_32_port, SHIFT_n_1_31_port, SHIFT_n_1_30_port, SHIFT_n_1_29_port,
      SHIFT_n_1_28_port, SHIFT_n_1_27_port, SHIFT_n_1_26_port, 
      SHIFT_n_1_25_port, SHIFT_n_1_24_port, SHIFT_n_1_23_port, 
      SHIFT_n_1_22_port, SHIFT_n_1_21_port, SHIFT_n_1_20_port, 
      SHIFT_n_1_19_port, SHIFT_n_1_18_port, SHIFT_n_1_17_port, 
      SHIFT_n_1_16_port, SHIFT_n_1_15_port, SHIFT_n_1_14_port, 
      SHIFT_n_1_13_port, SHIFT_n_1_12_port, SHIFT_n_1_11_port, 
      SHIFT_n_1_10_port, SHIFT_n_1_9_port, SHIFT_n_1_8_port, SHIFT_n_1_7_port, 
      SHIFT_n_1_6_port, SHIFT_n_1_5_port, SHIFT_n_1_4_port, SHIFT_n_1_3_port, 
      SHIFT_n_1_2_port, SHIFT_n_1_1_port, SHIFT_n_1_0_port, SHIFT_n_15_61_port,
      SHIFT_n_15_60_port, SHIFT_n_15_59_port, SHIFT_n_15_58_port, 
      SHIFT_n_15_57_port, SHIFT_n_15_56_port, SHIFT_n_15_55_port, 
      SHIFT_n_15_54_port, SHIFT_n_15_53_port, SHIFT_n_15_52_port, 
      SHIFT_n_15_51_port, SHIFT_n_15_50_port, SHIFT_n_15_49_port, 
      SHIFT_n_15_48_port, SHIFT_n_15_47_port, SHIFT_n_15_46_port, 
      SHIFT_n_15_45_port, SHIFT_n_15_44_port, SHIFT_n_15_43_port, 
      SHIFT_n_15_42_port, SHIFT_n_15_41_port, SHIFT_n_15_40_port, 
      SHIFT_n_15_39_port, SHIFT_n_15_38_port, SHIFT_n_15_37_port, 
      SHIFT_n_15_36_port, SHIFT_n_15_35_port, SHIFT_n_15_34_port, 
      SHIFT_n_15_33_port, SHIFT_n_15_32_port, SHIFT_n_15_31_port, 
      SHIFT_n_15_30_port, SHIFT_n_15_29_port, SHIFT_n_15_28_port, 
      SHIFT_n_15_27_port, SHIFT_n_15_26_port, SHIFT_n_15_25_port, 
      SHIFT_n_15_24_port, SHIFT_n_15_23_port, SHIFT_n_15_22_port, 
      SHIFT_n_15_21_port, SHIFT_n_15_20_port, SHIFT_n_15_19_port, 
      SHIFT_n_15_18_port, SHIFT_n_15_17_port, SHIFT_n_15_16_port, 
      SHIFT_n_15_15_port, SHIFT_n_15_14_port, SHIFT_n_15_13_port, 
      SHIFT_n_15_12_port, SHIFT_n_15_11_port, SHIFT_n_15_10_port, 
      SHIFT_n_15_9_port, SHIFT_n_15_8_port, SHIFT_n_15_7_port, 
      SHIFT_n_15_6_port, SHIFT_n_15_5_port, SHIFT_n_15_4_port, 
      SHIFT_n_15_3_port, SHIFT_n_15_2_port, SHIFT_n_15_1_port, 
      SHIFT_n_15_0_port, SHIFT_n_14_59_port, SHIFT_n_14_58_port, 
      SHIFT_n_14_57_port, SHIFT_n_14_56_port, SHIFT_n_14_55_port, 
      SHIFT_n_14_54_port, SHIFT_n_14_53_port, SHIFT_n_14_52_port, 
      SHIFT_n_14_51_port, SHIFT_n_14_50_port, SHIFT_n_14_49_port, 
      SHIFT_n_14_48_port, SHIFT_n_14_47_port, SHIFT_n_14_46_port, 
      SHIFT_n_14_45_port, SHIFT_n_14_44_port, SHIFT_n_14_43_port, 
      SHIFT_n_14_42_port, SHIFT_n_14_41_port, SHIFT_n_14_40_port, 
      SHIFT_n_14_39_port, SHIFT_n_14_38_port, SHIFT_n_14_37_port, 
      SHIFT_n_14_36_port, SHIFT_n_14_35_port, SHIFT_n_14_34_port, 
      SHIFT_n_14_33_port, SHIFT_n_14_32_port, SHIFT_n_14_31_port, 
      SHIFT_n_14_30_port, SHIFT_n_14_29_port, SHIFT_n_14_28_port, 
      SHIFT_n_14_27_port, SHIFT_n_14_26_port, SHIFT_n_14_25_port, 
      SHIFT_n_14_24_port, SHIFT_n_14_23_port, SHIFT_n_14_22_port, 
      SHIFT_n_14_21_port, SHIFT_n_14_20_port, SHIFT_n_14_19_port, 
      SHIFT_n_14_18_port, SHIFT_n_14_17_port, SHIFT_n_14_16_port, 
      SHIFT_n_14_15_port, SHIFT_n_14_14_port, SHIFT_n_14_13_port, 
      SHIFT_n_14_12_port, SHIFT_n_14_11_port, SHIFT_n_14_10_port, 
      SHIFT_n_14_9_port, SHIFT_n_14_8_port, SHIFT_n_14_7_port, 
      SHIFT_n_14_6_port, SHIFT_n_14_5_port, SHIFT_n_14_4_port, 
      SHIFT_n_14_3_port, SHIFT_n_14_2_port, SHIFT_n_14_1_port, 
      SHIFT_n_14_0_port, SHIFT_n_13_57_port, SHIFT_n_13_56_port, 
      SHIFT_n_13_55_port, SHIFT_n_13_54_port, SHIFT_n_13_53_port, 
      SHIFT_n_13_52_port, SHIFT_n_13_51_port, SHIFT_n_13_50_port, 
      SHIFT_n_13_49_port, SHIFT_n_13_48_port, SHIFT_n_13_47_port, 
      SHIFT_n_13_46_port, SHIFT_n_13_45_port, SHIFT_n_13_44_port, 
      SHIFT_n_13_43_port, SHIFT_n_13_42_port, SHIFT_n_13_41_port, 
      SHIFT_n_13_40_port, SHIFT_n_13_39_port, SHIFT_n_13_38_port, 
      SHIFT_n_13_37_port, SHIFT_n_13_36_port, SHIFT_n_13_35_port, 
      SHIFT_n_13_34_port, SHIFT_n_13_33_port, SHIFT_n_13_32_port, 
      SHIFT_n_13_31_port, SHIFT_n_13_30_port, SHIFT_n_13_29_port, 
      SHIFT_n_13_28_port, SHIFT_n_13_27_port, SHIFT_n_13_26_port, 
      SHIFT_n_13_25_port, SHIFT_n_13_24_port, SHIFT_n_13_23_port, 
      SHIFT_n_13_22_port, SHIFT_n_13_21_port, SHIFT_n_13_20_port, 
      SHIFT_n_13_19_port, SHIFT_n_13_18_port, SHIFT_n_13_17_port, 
      SHIFT_n_13_16_port, SHIFT_n_13_15_port, SHIFT_n_13_14_port, 
      SHIFT_n_13_13_port, SHIFT_n_13_12_port, SHIFT_n_13_11_port, 
      SHIFT_n_13_10_port, SHIFT_n_13_9_port, SHIFT_n_13_8_port, 
      SHIFT_n_13_7_port, SHIFT_n_13_6_port, SHIFT_n_13_5_port, 
      SHIFT_n_13_4_port, SHIFT_n_13_3_port, SHIFT_n_13_2_port, 
      SHIFT_n_13_1_port, SHIFT_n_13_0_port, SHIFT_n_12_55_port, 
      SHIFT_n_12_54_port, SHIFT_n_12_53_port, SHIFT_n_12_52_port, 
      SHIFT_n_12_51_port, SHIFT_n_12_50_port, SHIFT_n_12_49_port, 
      SHIFT_n_12_48_port, SHIFT_n_12_47_port, SHIFT_n_12_46_port, 
      SHIFT_n_12_45_port, SHIFT_n_12_44_port, SHIFT_n_12_43_port, 
      SHIFT_n_12_42_port, SHIFT_n_12_41_port, SHIFT_n_12_40_port, 
      SHIFT_n_12_39_port, SHIFT_n_12_38_port, SHIFT_n_12_37_port, 
      SHIFT_n_12_36_port, SHIFT_n_12_35_port, SHIFT_n_12_34_port, 
      SHIFT_n_12_33_port, SHIFT_n_12_32_port, SHIFT_n_12_31_port, 
      SHIFT_n_12_30_port, SHIFT_n_12_29_port, SHIFT_n_12_28_port, 
      SHIFT_n_12_27_port, SHIFT_n_12_26_port, SHIFT_n_12_25_port, 
      SHIFT_n_12_24_port, SHIFT_n_12_23_port, SHIFT_n_12_22_port, 
      SHIFT_n_12_21_port, SHIFT_n_12_20_port, SHIFT_n_12_19_port, 
      SHIFT_n_12_18_port, SHIFT_n_12_17_port, SHIFT_n_12_16_port, 
      SHIFT_n_12_15_port, SHIFT_n_12_14_port, SHIFT_n_12_13_port, 
      SHIFT_n_12_12_port, SHIFT_n_12_11_port, SHIFT_n_12_10_port, 
      SHIFT_n_12_9_port, SHIFT_n_12_8_port, SHIFT_n_12_7_port, 
      SHIFT_n_12_6_port, SHIFT_n_12_5_port, SHIFT_n_12_4_port, 
      SHIFT_n_12_3_port, SHIFT_n_12_2_port, SHIFT_n_12_1_port, 
      SHIFT_n_12_0_port, SHIFT_n_11_53_port, SHIFT_n_11_52_port, 
      SHIFT_n_11_51_port, SHIFT_n_11_50_port, SHIFT_n_11_49_port, 
      SHIFT_n_11_48_port, SHIFT_n_11_47_port, SHIFT_n_11_46_port, 
      SHIFT_n_11_45_port, SHIFT_n_11_44_port, SHIFT_n_11_43_port, 
      SHIFT_n_11_42_port, SHIFT_n_11_41_port, SHIFT_n_11_40_port, 
      SHIFT_n_11_39_port, SHIFT_n_11_38_port, SHIFT_n_11_37_port, 
      SHIFT_n_11_36_port, SHIFT_n_11_35_port, SHIFT_n_11_34_port, 
      SHIFT_n_11_33_port, SHIFT_n_11_32_port, SHIFT_n_11_31_port, 
      SHIFT_n_11_30_port, SHIFT_n_11_29_port, SHIFT_n_11_28_port, 
      SHIFT_n_11_27_port, SHIFT_n_11_26_port, SHIFT_n_11_25_port, 
      SHIFT_n_11_24_port, SHIFT_n_11_23_port, SHIFT_n_11_22_port, 
      SHIFT_n_11_21_port, SHIFT_n_11_20_port, SHIFT_n_11_19_port, 
      SHIFT_n_11_18_port, SHIFT_n_11_17_port, SHIFT_n_11_16_port, 
      SHIFT_n_11_15_port, SHIFT_n_11_14_port, SHIFT_n_11_13_port, 
      SHIFT_n_11_12_port, SHIFT_n_11_11_port, SHIFT_n_11_10_port, 
      SHIFT_n_11_9_port, SHIFT_n_11_8_port, SHIFT_n_11_7_port, 
      SHIFT_n_11_6_port, SHIFT_n_11_5_port, SHIFT_n_11_4_port, 
      SHIFT_n_11_3_port, SHIFT_n_11_2_port, SHIFT_n_11_1_port, 
      SHIFT_n_11_0_port, SHIFT_n_10_51_port, SHIFT_n_10_50_port, 
      SHIFT_n_10_49_port, SHIFT_n_10_48_port, SHIFT_n_10_47_port, 
      SHIFT_n_10_46_port, SHIFT_n_10_45_port, SHIFT_n_10_44_port, 
      SHIFT_n_10_43_port, SHIFT_n_10_42_port, SHIFT_n_10_41_port, 
      SHIFT_n_10_40_port, SHIFT_n_10_39_port, SHIFT_n_10_38_port, 
      SHIFT_n_10_37_port, SHIFT_n_10_36_port, SHIFT_n_10_35_port, 
      SHIFT_n_10_34_port, SHIFT_n_10_33_port, SHIFT_n_10_32_port, 
      SHIFT_n_10_31_port, SHIFT_n_10_30_port, SHIFT_n_10_29_port, 
      SHIFT_n_10_28_port, SHIFT_n_10_27_port, SHIFT_n_10_26_port, 
      SHIFT_n_10_25_port, SHIFT_n_10_24_port, SHIFT_n_10_23_port, 
      SHIFT_n_10_22_port, SHIFT_n_10_21_port, SHIFT_n_10_20_port, 
      SHIFT_n_10_19_port, SHIFT_n_10_18_port, SHIFT_n_10_17_port, 
      SHIFT_n_10_16_port, SHIFT_n_10_15_port, SHIFT_n_10_14_port, 
      SHIFT_n_10_13_port, SHIFT_n_10_12_port, SHIFT_n_10_11_port, 
      SHIFT_n_10_10_port, SHIFT_n_10_9_port, SHIFT_n_10_8_port, 
      SHIFT_n_10_7_port, SHIFT_n_10_6_port, SHIFT_n_10_5_port, 
      SHIFT_n_10_4_port, SHIFT_n_10_3_port, SHIFT_n_10_2_port, 
      SHIFT_n_10_1_port, SHIFT_n_10_0_port, SHIFT_n_9_49_port, 
      SHIFT_n_9_48_port, SHIFT_n_9_47_port, SHIFT_n_9_46_port, 
      SHIFT_n_9_45_port, SHIFT_n_9_44_port, SHIFT_n_9_43_port, 
      SHIFT_n_9_42_port, SHIFT_n_9_41_port, SHIFT_n_9_40_port, 
      SHIFT_n_9_39_port, SHIFT_n_9_38_port, SHIFT_n_9_37_port, 
      SHIFT_n_9_36_port, SHIFT_n_9_35_port, SHIFT_n_9_34_port, 
      SHIFT_n_9_33_port, SHIFT_n_9_32_port, SHIFT_n_9_31_port, 
      SHIFT_n_9_30_port, SHIFT_n_9_29_port, SHIFT_n_9_28_port, 
      SHIFT_n_9_27_port, SHIFT_n_9_26_port, SHIFT_n_9_25_port, 
      SHIFT_n_9_24_port, SHIFT_n_9_23_port, SHIFT_n_9_22_port, 
      SHIFT_n_9_21_port, SHIFT_n_9_20_port, SHIFT_n_9_19_port, 
      SHIFT_n_9_18_port, SHIFT_n_9_17_port, SHIFT_n_9_16_port, 
      SHIFT_n_9_15_port, SHIFT_n_9_14_port, SHIFT_n_9_13_port, 
      SHIFT_n_9_12_port, SHIFT_n_9_11_port, SHIFT_n_9_10_port, SHIFT_n_9_9_port
      , SHIFT_n_9_8_port, SHIFT_n_9_7_port, SHIFT_n_9_6_port, SHIFT_n_9_5_port,
      SHIFT_n_9_4_port, SHIFT_n_9_3_port, SHIFT_n_9_2_port, SHIFT_n_9_1_port, 
      SHIFT_n_9_0_port, SHIFT_n_8_47_port, SHIFT_n_8_46_port, SHIFT_n_8_45_port
      , SHIFT_n_8_44_port, SHIFT_n_8_43_port, SHIFT_n_8_42_port, 
      SHIFT_n_8_41_port, SHIFT_n_8_40_port, SHIFT_n_8_39_port, 
      SHIFT_n_8_38_port, SHIFT_n_8_37_port, SHIFT_n_8_36_port, 
      SHIFT_n_8_35_port, SHIFT_n_8_34_port, SHIFT_n_8_33_port, 
      SHIFT_n_8_32_port, SHIFT_n_8_31_port, SHIFT_n_8_30_port, 
      SHIFT_n_8_29_port, SHIFT_n_8_28_port, SHIFT_n_8_27_port, 
      SHIFT_n_8_26_port, SHIFT_n_8_25_port, SHIFT_n_8_24_port, 
      SHIFT_n_8_23_port, SHIFT_n_8_22_port, SHIFT_n_8_21_port, 
      SHIFT_n_8_20_port, SHIFT_n_8_19_port, SHIFT_n_8_18_port, 
      SHIFT_n_8_17_port, SHIFT_n_8_16_port, SHIFT_n_8_15_port, 
      SHIFT_n_8_14_port, SHIFT_n_8_13_port, SHIFT_n_8_12_port, 
      SHIFT_n_8_11_port, SHIFT_n_8_10_port, SHIFT_n_8_9_port, SHIFT_n_8_8_port,
      SHIFT_n_8_7_port, SHIFT_n_8_6_port, SHIFT_n_8_5_port, SHIFT_n_8_4_port, 
      SHIFT_n_8_3_port, SHIFT_n_8_2_port, SHIFT_n_8_1_port, SHIFT_n_8_0_port, 
      SHIFT_n_7_45_port, SHIFT_n_7_44_port, SHIFT_n_7_43_port, 
      SHIFT_n_7_42_port, SHIFT_n_7_41_port, SHIFT_n_7_40_port, 
      SHIFT_n_7_39_port, SHIFT_n_7_38_port, SHIFT_n_7_37_port, 
      SHIFT_n_7_36_port, SHIFT_n_7_35_port, SHIFT_n_7_34_port, 
      SHIFT_n_7_33_port, SHIFT_n_7_32_port, SHIFT_n_7_31_port, 
      SHIFT_n_7_30_port, SHIFT_n_7_29_port, SHIFT_n_7_28_port, 
      SHIFT_n_7_27_port, SHIFT_n_7_26_port, SHIFT_n_7_25_port, 
      SHIFT_n_7_24_port, SHIFT_n_7_23_port, SHIFT_n_7_22_port, 
      SHIFT_n_7_21_port, SHIFT_n_7_20_port, SHIFT_n_7_19_port, 
      SHIFT_n_7_18_port, SHIFT_n_7_17_port, SHIFT_n_7_16_port, 
      SHIFT_n_7_15_port, SHIFT_n_7_14_port, SHIFT_n_7_13_port, 
      SHIFT_n_7_12_port, SHIFT_n_7_11_port, SHIFT_n_7_10_port, SHIFT_n_7_9_port
      , SHIFT_n_7_8_port, SHIFT_n_7_7_port, SHIFT_n_7_6_port, SHIFT_n_7_5_port,
      SHIFT_n_7_4_port, SHIFT_n_7_3_port, SHIFT_n_7_2_port, SHIFT_n_7_1_port, 
      SHIFT_n_7_0_port, SHIFT_n_6_43_port, SHIFT_n_6_42_port, SHIFT_n_6_41_port
      , SHIFT_n_6_40_port, SHIFT_n_6_39_port, SHIFT_n_6_38_port, 
      SHIFT_n_6_37_port, SHIFT_n_6_36_port, SHIFT_n_6_35_port, 
      SHIFT_n_6_34_port, SHIFT_n_6_33_port, SHIFT_n_6_32_port, 
      SHIFT_n_6_31_port, SHIFT_n_6_30_port, SHIFT_n_6_29_port, 
      SHIFT_n_6_28_port, SHIFT_n_6_27_port, SHIFT_n_6_26_port, 
      SHIFT_n_6_25_port, SHIFT_n_6_24_port, SHIFT_n_6_23_port, 
      SHIFT_n_6_22_port, SHIFT_n_6_21_port, SHIFT_n_6_20_port, 
      SHIFT_n_6_19_port, SHIFT_n_6_18_port, SHIFT_n_6_17_port, 
      SHIFT_n_6_16_port, SHIFT_n_6_15_port, SHIFT_n_6_14_port, 
      SHIFT_n_6_13_port, SHIFT_n_6_12_port, SHIFT_n_6_11_port, 
      SHIFT_n_6_10_port, SHIFT_n_6_9_port, SHIFT_n_6_8_port, SHIFT_n_6_7_port, 
      SHIFT_n_6_6_port, SHIFT_n_6_5_port, SHIFT_n_6_4_port, SHIFT_n_6_3_port, 
      SHIFT_n_6_2_port, SHIFT_n_6_1_port, SHIFT_n_6_0_port, SHIFT_n_5_41_port, 
      SHIFT_n_5_40_port, SHIFT_n_5_39_port, SHIFT_n_5_38_port, 
      SHIFT_n_5_37_port, SHIFT_n_5_36_port, SHIFT_n_5_35_port, 
      SHIFT_n_5_34_port, SHIFT_n_5_33_port, SHIFT_n_5_32_port, 
      SHIFT_n_5_31_port, SHIFT_n_5_30_port, SHIFT_n_5_29_port, 
      SHIFT_n_5_28_port, SHIFT_n_5_27_port, SHIFT_n_5_26_port, 
      SHIFT_n_5_25_port, SHIFT_n_5_24_port, SHIFT_n_5_23_port, 
      SHIFT_n_5_22_port, SHIFT_n_5_21_port, SHIFT_n_5_20_port, 
      SHIFT_n_5_19_port, SHIFT_n_5_18_port, SHIFT_n_5_17_port, 
      SHIFT_n_5_16_port, SHIFT_n_5_15_port, SHIFT_n_5_14_port, 
      SHIFT_n_5_13_port, SHIFT_n_5_12_port, SHIFT_n_5_11_port, 
      SHIFT_n_5_10_port, SHIFT_n_5_9_port, SHIFT_n_5_8_port, SHIFT_n_5_7_port, 
      SHIFT_n_5_6_port, SHIFT_n_5_5_port, SHIFT_n_5_4_port, SHIFT_n_5_3_port, 
      SHIFT_n_5_2_port, SHIFT_n_5_1_port, SHIFT_n_5_0_port, SHIFT_n_4_39_port, 
      SHIFT_n_4_38_port, SHIFT_n_4_37_port, SHIFT_n_4_36_port, 
      SHIFT_n_4_35_port, SHIFT_n_4_34_port, SHIFT_n_4_33_port, 
      SHIFT_n_4_32_port, SHIFT_n_4_31_port, SHIFT_n_4_30_port, 
      SHIFT_n_4_29_port, SHIFT_n_4_28_port, SHIFT_n_4_27_port, 
      SHIFT_n_4_26_port, SHIFT_n_4_25_port, SHIFT_n_4_24_port, 
      SHIFT_n_4_23_port, SHIFT_n_4_22_port, SHIFT_n_4_21_port, 
      SHIFT_n_4_20_port, SHIFT_n_4_19_port, SHIFT_n_4_18_port, 
      SHIFT_n_4_17_port, SHIFT_n_4_16_port, SHIFT_n_4_15_port, 
      SHIFT_n_4_14_port, SHIFT_n_4_13_port, SHIFT_n_4_12_port, 
      SHIFT_n_4_11_port, SHIFT_n_4_10_port, SHIFT_n_4_9_port, SHIFT_n_4_8_port,
      SHIFT_n_4_7_port, SHIFT_n_4_6_port, SHIFT_n_4_5_port, SHIFT_n_4_4_port, 
      SHIFT_n_4_3_port, SHIFT_n_4_2_port, SHIFT_n_4_1_port, SHIFT_n_4_0_port, 
      SHIFT_n_3_37_port, SHIFT_n_3_36_port, SHIFT_n_3_35_port, 
      SHIFT_n_3_34_port, SHIFT_n_3_33_port, SHIFT_n_3_32_port, 
      SHIFT_n_3_31_port, SHIFT_n_3_30_port, SHIFT_n_3_29_port, 
      SHIFT_n_3_28_port, SHIFT_n_3_27_port, SHIFT_n_3_26_port, 
      SHIFT_n_3_25_port, SHIFT_n_3_24_port, SHIFT_n_3_23_port, 
      SHIFT_n_3_22_port, SHIFT_n_3_21_port, SHIFT_n_3_20_port, 
      SHIFT_n_3_19_port, SHIFT_n_3_18_port, SHIFT_n_3_17_port, 
      SHIFT_n_3_16_port, SHIFT_n_3_15_port, SHIFT_n_3_14_port, 
      SHIFT_n_3_13_port, SHIFT_n_3_12_port, SHIFT_n_3_11_port, 
      SHIFT_n_3_10_port, SHIFT_n_3_9_port, SHIFT_n_3_8_port, SHIFT_n_3_7_port, 
      SHIFT_n_3_6_port, SHIFT_n_3_5_port, SHIFT_n_3_4_port, SHIFT_n_3_3_port, 
      SHIFT_n_3_2_port, SHIFT_n_3_1_port, SHIFT_n_3_0_port, SHIFT_n_2_35_port, 
      SHIFT_n_2_34_port, SHIFT_n_2_33_port, SHIFT_n_2_32_port, 
      SHIFT_n_2_31_port, SHIFT_n_2_30_port, SHIFT_n_2_29_port, 
      SHIFT_n_2_28_port, SHIFT_n_2_27_port, SHIFT_n_2_26_port, 
      SHIFT_n_2_25_port, SHIFT_n_2_24_port, SHIFT_n_2_23_port, 
      SHIFT_n_2_22_port, SHIFT_n_2_21_port, SHIFT_n_2_20_port, 
      SHIFT_n_2_19_port, SHIFT_n_2_18_port, SHIFT_n_2_17_port, 
      SHIFT_n_2_16_port, SHIFT_n_2_15_port, SHIFT_n_2_14_port, 
      SHIFT_n_2_13_port, SHIFT_n_2_12_port, SHIFT_n_2_11_port, 
      SHIFT_n_2_10_port, SHIFT_n_2_9_port, SHIFT_n_2_8_port, SHIFT_n_2_7_port, 
      SHIFT_n_2_6_port, SHIFT_n_2_5_port, SHIFT_n_2_4_port, SHIFT_n_2_3_port, 
      SHIFT_n_2_2_port, SHIFT_n_2_1_port, SHIFT_n_2_0_port, SHIFT_n_1_33_port, 
      SHIFT_n_1_32_port, OTMP_8_15_port, OTMP_8_14_port, OTMP_8_13_port, 
      OTMP_8_12_port, OTMP_8_11_port, OTMP_8_10_port, OTMP_8_9_port, 
      OTMP_8_8_port, OTMP_8_7_port, OTMP_8_6_port, OTMP_8_5_port, OTMP_8_4_port
      , OTMP_8_3_port, OTMP_8_2_port, OTMP_8_1_port, OTMP_8_0_port, 
      OTMP_7_47_port, OTMP_7_46_port, OTMP_7_45_port, OTMP_7_44_port, 
      OTMP_7_43_port, OTMP_7_42_port, OTMP_7_41_port, OTMP_7_40_port, 
      OTMP_7_39_port, OTMP_7_38_port, OTMP_7_37_port, OTMP_7_36_port, 
      OTMP_7_35_port, OTMP_7_34_port, OTMP_7_33_port, OTMP_7_32_port, 
      OTMP_7_31_port, OTMP_7_30_port, OTMP_7_29_port, OTMP_7_28_port, 
      OTMP_7_27_port, OTMP_7_26_port, OTMP_7_25_port, OTMP_7_24_port, 
      OTMP_7_23_port, OTMP_7_22_port, OTMP_7_21_port, OTMP_7_20_port, 
      OTMP_7_19_port, OTMP_7_18_port, OTMP_7_17_port, OTMP_7_16_port, 
      OTMP_7_15_port, OTMP_7_14_port, OTMP_7_13_port, OTMP_7_12_port, 
      OTMP_7_11_port, OTMP_7_10_port, OTMP_7_9_port, OTMP_7_8_port, 
      OTMP_7_7_port, OTMP_7_6_port, OTMP_7_5_port, OTMP_7_4_port, OTMP_7_3_port
      , OTMP_7_2_port, OTMP_7_1_port, OTMP_7_0_port, OTMP_6_45_port, 
      OTMP_6_44_port, OTMP_6_43_port, OTMP_6_42_port, OTMP_6_41_port, 
      OTMP_6_40_port, OTMP_6_39_port, OTMP_6_38_port, OTMP_6_37_port, 
      OTMP_6_36_port, OTMP_6_35_port, OTMP_6_34_port, OTMP_6_33_port, 
      OTMP_6_32_port, OTMP_6_31_port, OTMP_6_30_port, OTMP_6_29_port, 
      OTMP_6_28_port, OTMP_6_27_port, OTMP_6_26_port, OTMP_6_25_port, 
      OTMP_6_24_port, OTMP_6_23_port, OTMP_6_22_port, OTMP_6_21_port, 
      OTMP_6_20_port, OTMP_6_19_port, OTMP_6_18_port, OTMP_6_17_port, 
      OTMP_6_16_port, OTMP_6_15_port, OTMP_6_14_port, OTMP_6_13_port, 
      OTMP_6_12_port, OTMP_6_11_port, OTMP_6_10_port, OTMP_6_9_port, 
      OTMP_6_8_port, OTMP_6_7_port, OTMP_6_6_port, OTMP_6_5_port, OTMP_6_4_port
      , OTMP_6_3_port, OTMP_6_2_port, OTMP_6_1_port, OTMP_6_0_port, 
      OTMP_5_43_port, OTMP_5_42_port, OTMP_5_41_port, OTMP_5_40_port, 
      OTMP_5_39_port, OTMP_5_38_port, OTMP_5_37_port, OTMP_5_36_port, 
      OTMP_5_35_port, OTMP_5_34_port, OTMP_5_33_port, OTMP_5_32_port, 
      OTMP_5_31_port, OTMP_5_30_port, OTMP_5_29_port, OTMP_5_28_port, 
      OTMP_5_27_port, OTMP_5_26_port, OTMP_5_25_port, OTMP_5_24_port, 
      OTMP_5_23_port, OTMP_5_22_port, OTMP_5_21_port, OTMP_5_20_port, 
      OTMP_5_19_port, OTMP_5_18_port, OTMP_5_17_port, OTMP_5_16_port, 
      OTMP_5_15_port, OTMP_5_14_port, OTMP_5_13_port, OTMP_5_12_port, 
      OTMP_5_11_port, OTMP_5_10_port, OTMP_5_9_port, OTMP_5_8_port, 
      OTMP_5_7_port, OTMP_5_6_port, OTMP_5_5_port, OTMP_5_4_port, OTMP_5_3_port
      , OTMP_5_2_port, OTMP_5_1_port, OTMP_5_0_port, OTMP_4_41_port, 
      OTMP_4_40_port, OTMP_4_39_port, OTMP_4_38_port, OTMP_4_37_port, 
      OTMP_4_36_port, OTMP_4_35_port, OTMP_4_34_port, OTMP_4_33_port, 
      OTMP_4_32_port, OTMP_4_31_port, OTMP_4_30_port, OTMP_4_29_port, 
      OTMP_4_28_port, OTMP_4_27_port, OTMP_4_26_port, OTMP_4_25_port, 
      OTMP_4_24_port, OTMP_4_23_port, OTMP_4_22_port, OTMP_4_21_port, 
      OTMP_4_20_port, OTMP_4_19_port, OTMP_4_18_port, OTMP_4_17_port, 
      OTMP_4_16_port, OTMP_4_15_port, OTMP_4_14_port, OTMP_4_13_port, 
      OTMP_4_12_port, OTMP_4_11_port, OTMP_4_10_port, OTMP_4_9_port, 
      OTMP_4_8_port, OTMP_4_7_port, OTMP_4_6_port, OTMP_4_5_port, OTMP_4_4_port
      , OTMP_4_3_port, OTMP_4_2_port, OTMP_4_1_port, OTMP_4_0_port, 
      OTMP_3_39_port, OTMP_3_38_port, OTMP_3_37_port, OTMP_3_36_port, 
      OTMP_3_35_port, OTMP_3_34_port, OTMP_3_33_port, OTMP_3_32_port, 
      OTMP_3_31_port, OTMP_3_30_port, OTMP_3_29_port, OTMP_3_28_port, 
      OTMP_3_27_port, OTMP_3_26_port, OTMP_3_25_port, OTMP_3_24_port, 
      OTMP_3_23_port, OTMP_3_22_port, OTMP_3_21_port, OTMP_3_20_port, 
      OTMP_3_19_port, OTMP_3_18_port, OTMP_3_17_port, OTMP_3_16_port, 
      OTMP_3_15_port, OTMP_3_14_port, OTMP_3_13_port, OTMP_3_12_port, 
      OTMP_3_11_port, OTMP_3_10_port, OTMP_3_9_port, OTMP_3_8_port, 
      OTMP_3_7_port, OTMP_3_6_port, OTMP_3_5_port, OTMP_3_4_port, OTMP_3_3_port
      , OTMP_3_2_port, OTMP_3_1_port, OTMP_3_0_port, OTMP_2_37_port, 
      OTMP_2_36_port, OTMP_2_35_port, OTMP_2_34_port, OTMP_2_33_port, 
      OTMP_2_32_port, OTMP_2_31_port, OTMP_2_30_port, OTMP_2_29_port, 
      OTMP_2_28_port, OTMP_2_27_port, OTMP_2_26_port, OTMP_2_25_port, 
      OTMP_2_24_port, OTMP_2_23_port, OTMP_2_22_port, OTMP_2_21_port, 
      OTMP_2_20_port, OTMP_2_19_port, OTMP_2_18_port, OTMP_2_17_port, 
      OTMP_2_16_port, OTMP_2_15_port, OTMP_2_14_port, OTMP_2_13_port, 
      OTMP_2_12_port, OTMP_2_11_port, OTMP_2_10_port, OTMP_2_9_port, 
      OTMP_2_8_port, OTMP_2_7_port, OTMP_2_6_port, OTMP_2_5_port, OTMP_2_4_port
      , OTMP_2_3_port, OTMP_2_2_port, OTMP_2_1_port, OTMP_2_0_port, 
      OTMP_1_35_port, OTMP_1_34_port, OTMP_1_33_port, OTMP_1_32_port, 
      OTMP_1_31_port, OTMP_1_30_port, OTMP_1_29_port, OTMP_1_28_port, 
      OTMP_1_27_port, OTMP_1_26_port, OTMP_1_25_port, OTMP_1_24_port, 
      OTMP_1_23_port, OTMP_1_22_port, OTMP_1_21_port, OTMP_1_20_port, 
      OTMP_1_19_port, OTMP_1_18_port, OTMP_1_17_port, OTMP_1_16_port, 
      OTMP_1_15_port, OTMP_1_14_port, OTMP_1_13_port, OTMP_1_12_port, 
      OTMP_1_11_port, OTMP_1_10_port, OTMP_1_9_port, OTMP_1_8_port, 
      OTMP_1_7_port, OTMP_1_6_port, OTMP_1_5_port, OTMP_1_4_port, OTMP_1_3_port
      , OTMP_1_2_port, OTMP_1_1_port, OTMP_1_0_port, OTMP_0_34_port, 
      OTMP_0_32_port, OTMP_0_31_port, OTMP_0_30_port, OTMP_0_29_port, 
      OTMP_0_28_port, OTMP_0_27_port, OTMP_0_26_port, OTMP_0_25_port, 
      OTMP_0_24_port, OTMP_0_23_port, OTMP_0_22_port, OTMP_0_21_port, 
      OTMP_0_20_port, OTMP_0_19_port, OTMP_0_18_port, OTMP_0_17_port, 
      OTMP_0_16_port, OTMP_0_15_port, OTMP_0_14_port, OTMP_0_13_port, 
      OTMP_0_12_port, OTMP_0_11_port, OTMP_0_10_port, OTMP_0_9_port, 
      OTMP_0_8_port, OTMP_0_7_port, OTMP_0_6_port, OTMP_0_5_port, OTMP_0_4_port
      , OTMP_0_3_port, OTMP_0_2_port, OTMP_0_1_port, OTMP_0_0_port, 
      OTMP_15_63_port, OTMP_15_62_port, OTMP_15_61_port, OTMP_15_60_port, 
      OTMP_15_59_port, OTMP_15_58_port, OTMP_15_57_port, OTMP_15_56_port, 
      OTMP_15_55_port, OTMP_15_54_port, OTMP_15_53_port, OTMP_15_52_port, 
      OTMP_15_51_port, OTMP_15_50_port, OTMP_15_49_port, OTMP_15_48_port, 
      OTMP_15_47_port, OTMP_15_46_port, OTMP_15_45_port, OTMP_15_44_port, 
      OTMP_15_43_port, OTMP_15_42_port, OTMP_15_41_port, OTMP_15_40_port, 
      OTMP_15_39_port, OTMP_15_38_port, OTMP_15_37_port, OTMP_15_36_port, 
      OTMP_15_35_port, OTMP_15_34_port, OTMP_15_33_port, OTMP_15_32_port, 
      OTMP_15_31_port, OTMP_15_30_port, OTMP_15_29_port, OTMP_15_28_port, 
      OTMP_15_27_port, OTMP_15_26_port, OTMP_15_25_port, OTMP_15_24_port, 
      OTMP_15_23_port, OTMP_15_22_port, OTMP_15_21_port, OTMP_15_20_port, 
      OTMP_15_19_port, OTMP_15_18_port, OTMP_15_17_port, OTMP_15_16_port, 
      OTMP_15_15_port, OTMP_15_14_port, OTMP_15_13_port, OTMP_15_12_port, 
      OTMP_15_11_port, OTMP_15_10_port, OTMP_15_9_port, OTMP_15_8_port, 
      OTMP_15_7_port, OTMP_15_6_port, OTMP_15_5_port, OTMP_15_4_port, 
      OTMP_15_3_port, OTMP_15_2_port, OTMP_15_1_port, OTMP_15_0_port, 
      OTMP_14_61_port, OTMP_14_60_port, OTMP_14_59_port, OTMP_14_58_port, 
      OTMP_14_57_port, OTMP_14_56_port, OTMP_14_55_port, OTMP_14_54_port, 
      OTMP_14_53_port, OTMP_14_52_port, OTMP_14_51_port, OTMP_14_50_port, 
      OTMP_14_49_port, OTMP_14_48_port, OTMP_14_47_port, OTMP_14_46_port, 
      OTMP_14_45_port, OTMP_14_44_port, OTMP_14_43_port, OTMP_14_42_port, 
      OTMP_14_41_port, OTMP_14_40_port, OTMP_14_39_port, OTMP_14_38_port, 
      OTMP_14_37_port, OTMP_14_36_port, OTMP_14_35_port, OTMP_14_34_port, 
      OTMP_14_33_port, OTMP_14_32_port, OTMP_14_31_port, OTMP_14_30_port, 
      OTMP_14_29_port, OTMP_14_28_port, OTMP_14_27_port, OTMP_14_26_port, 
      OTMP_14_25_port, OTMP_14_24_port, OTMP_14_23_port, OTMP_14_22_port, 
      OTMP_14_21_port, OTMP_14_20_port, OTMP_14_19_port, OTMP_14_18_port, 
      OTMP_14_17_port, OTMP_14_16_port, OTMP_14_15_port, OTMP_14_14_port, 
      OTMP_14_13_port, OTMP_14_12_port, OTMP_14_11_port, OTMP_14_10_port, 
      OTMP_14_9_port, OTMP_14_8_port, OTMP_14_7_port, OTMP_14_6_port, 
      OTMP_14_5_port, OTMP_14_4_port, OTMP_14_3_port, OTMP_14_2_port, 
      OTMP_14_1_port, OTMP_14_0_port, OTMP_13_59_port, OTMP_13_58_port, 
      OTMP_13_57_port, OTMP_13_56_port, OTMP_13_55_port, OTMP_13_54_port, 
      OTMP_13_53_port, OTMP_13_52_port, OTMP_13_51_port, OTMP_13_50_port, 
      OTMP_13_49_port, OTMP_13_48_port, OTMP_13_47_port, OTMP_13_46_port, 
      OTMP_13_45_port, OTMP_13_44_port, OTMP_13_43_port, OTMP_13_42_port, 
      OTMP_13_41_port, OTMP_13_40_port, OTMP_13_39_port, OTMP_13_38_port, 
      OTMP_13_37_port, OTMP_13_36_port, OTMP_13_35_port, OTMP_13_34_port, 
      OTMP_13_33_port, OTMP_13_32_port, OTMP_13_31_port, OTMP_13_30_port, 
      OTMP_13_29_port, OTMP_13_28_port, OTMP_13_27_port, OTMP_13_26_port, 
      OTMP_13_25_port, OTMP_13_24_port, OTMP_13_23_port, OTMP_13_22_port, 
      OTMP_13_21_port, OTMP_13_20_port, OTMP_13_19_port, OTMP_13_18_port, 
      OTMP_13_17_port, OTMP_13_16_port, OTMP_13_15_port, OTMP_13_14_port, 
      OTMP_13_13_port, OTMP_13_12_port, OTMP_13_11_port, OTMP_13_10_port, 
      OTMP_13_9_port, OTMP_13_8_port, OTMP_13_7_port, OTMP_13_6_port, 
      OTMP_13_5_port, OTMP_13_4_port, OTMP_13_3_port, OTMP_13_2_port, 
      OTMP_13_1_port, OTMP_13_0_port, OTMP_12_57_port, OTMP_12_56_port, 
      OTMP_12_55_port, OTMP_12_54_port, OTMP_12_53_port, OTMP_12_52_port, 
      OTMP_12_51_port, OTMP_12_50_port, OTMP_12_49_port, OTMP_12_48_port, 
      OTMP_12_47_port, OTMP_12_46_port, OTMP_12_45_port, OTMP_12_44_port, 
      OTMP_12_43_port, OTMP_12_42_port, OTMP_12_41_port, OTMP_12_40_port, 
      OTMP_12_39_port, OTMP_12_38_port, OTMP_12_37_port, OTMP_12_36_port, 
      OTMP_12_35_port, OTMP_12_34_port, OTMP_12_33_port, OTMP_12_32_port, 
      OTMP_12_31_port, OTMP_12_30_port, OTMP_12_29_port, OTMP_12_28_port, 
      OTMP_12_27_port, OTMP_12_26_port, OTMP_12_25_port, OTMP_12_24_port, 
      OTMP_12_23_port, OTMP_12_22_port, OTMP_12_21_port, OTMP_12_20_port, 
      OTMP_12_19_port, OTMP_12_18_port, OTMP_12_17_port, OTMP_12_16_port, 
      OTMP_12_15_port, OTMP_12_14_port, OTMP_12_13_port, OTMP_12_12_port, 
      OTMP_12_11_port, OTMP_12_10_port, OTMP_12_9_port, OTMP_12_8_port, 
      OTMP_12_7_port, OTMP_12_6_port, OTMP_12_5_port, OTMP_12_4_port, 
      OTMP_12_3_port, OTMP_12_2_port, OTMP_12_1_port, OTMP_12_0_port, 
      OTMP_11_55_port, OTMP_11_54_port, OTMP_11_53_port, OTMP_11_52_port, 
      OTMP_11_51_port, OTMP_11_50_port, OTMP_11_49_port, OTMP_11_48_port, 
      OTMP_11_47_port, OTMP_11_46_port, OTMP_11_45_port, OTMP_11_44_port, 
      OTMP_11_43_port, OTMP_11_42_port, OTMP_11_41_port, OTMP_11_40_port, 
      OTMP_11_39_port, OTMP_11_38_port, OTMP_11_37_port, OTMP_11_36_port, 
      OTMP_11_35_port, OTMP_11_34_port, OTMP_11_33_port, OTMP_11_32_port, 
      OTMP_11_31_port, OTMP_11_30_port, OTMP_11_29_port, OTMP_11_28_port, 
      OTMP_11_27_port, OTMP_11_26_port, OTMP_11_25_port, OTMP_11_24_port, 
      OTMP_11_23_port, OTMP_11_22_port, OTMP_11_21_port, OTMP_11_20_port, 
      OTMP_11_19_port, OTMP_11_18_port, OTMP_11_17_port, OTMP_11_16_port, 
      OTMP_11_15_port, OTMP_11_14_port, OTMP_11_13_port, OTMP_11_12_port, 
      OTMP_11_11_port, OTMP_11_10_port, OTMP_11_9_port, OTMP_11_8_port, 
      OTMP_11_7_port, OTMP_11_6_port, OTMP_11_5_port, OTMP_11_4_port, 
      OTMP_11_3_port, OTMP_11_2_port, OTMP_11_1_port, OTMP_11_0_port, 
      OTMP_10_53_port, OTMP_10_52_port, OTMP_10_51_port, OTMP_10_50_port, 
      OTMP_10_49_port, OTMP_10_48_port, OTMP_10_47_port, OTMP_10_46_port, 
      OTMP_10_45_port, OTMP_10_44_port, OTMP_10_43_port, OTMP_10_42_port, 
      OTMP_10_41_port, OTMP_10_40_port, OTMP_10_39_port, OTMP_10_38_port, 
      OTMP_10_37_port, OTMP_10_36_port, OTMP_10_35_port, OTMP_10_34_port, 
      OTMP_10_33_port, OTMP_10_32_port, OTMP_10_31_port, OTMP_10_30_port, 
      OTMP_10_29_port, OTMP_10_28_port, OTMP_10_27_port, OTMP_10_26_port, 
      OTMP_10_25_port, OTMP_10_24_port, OTMP_10_23_port, OTMP_10_22_port, 
      OTMP_10_21_port, OTMP_10_20_port, OTMP_10_19_port, OTMP_10_18_port, 
      OTMP_10_17_port, OTMP_10_16_port, OTMP_10_15_port, OTMP_10_14_port, 
      OTMP_10_13_port, OTMP_10_12_port, OTMP_10_11_port, OTMP_10_10_port, 
      OTMP_10_9_port, OTMP_10_8_port, OTMP_10_7_port, OTMP_10_6_port, 
      OTMP_10_5_port, OTMP_10_4_port, OTMP_10_3_port, OTMP_10_2_port, 
      OTMP_10_1_port, OTMP_10_0_port, OTMP_9_51_port, OTMP_9_50_port, 
      OTMP_9_49_port, OTMP_9_48_port, OTMP_9_47_port, OTMP_9_46_port, 
      OTMP_9_45_port, OTMP_9_44_port, OTMP_9_43_port, OTMP_9_42_port, 
      OTMP_9_41_port, OTMP_9_40_port, OTMP_9_39_port, OTMP_9_38_port, 
      OTMP_9_37_port, OTMP_9_36_port, OTMP_9_35_port, OTMP_9_34_port, 
      OTMP_9_33_port, OTMP_9_32_port, OTMP_9_31_port, OTMP_9_30_port, 
      OTMP_9_29_port, OTMP_9_28_port, OTMP_9_27_port, OTMP_9_26_port, 
      OTMP_9_25_port, OTMP_9_24_port, OTMP_9_23_port, OTMP_9_22_port, 
      OTMP_9_21_port, OTMP_9_20_port, OTMP_9_19_port, OTMP_9_18_port, 
      OTMP_9_17_port, OTMP_9_16_port, OTMP_9_15_port, OTMP_9_14_port, 
      OTMP_9_13_port, OTMP_9_12_port, OTMP_9_11_port, OTMP_9_10_port, 
      OTMP_9_9_port, OTMP_9_8_port, OTMP_9_7_port, OTMP_9_6_port, OTMP_9_5_port
      , OTMP_9_4_port, OTMP_9_3_port, OTMP_9_2_port, OTMP_9_1_port, 
      OTMP_9_0_port, OTMP_8_49_port, OTMP_8_48_port, OTMP_8_47_port, 
      OTMP_8_46_port, OTMP_8_45_port, OTMP_8_44_port, OTMP_8_43_port, 
      OTMP_8_42_port, OTMP_8_41_port, OTMP_8_40_port, OTMP_8_39_port, 
      OTMP_8_38_port, OTMP_8_37_port, OTMP_8_36_port, OTMP_8_35_port, 
      OTMP_8_34_port, OTMP_8_33_port, OTMP_8_32_port, OTMP_8_31_port, 
      OTMP_8_30_port, OTMP_8_29_port, OTMP_8_28_port, OTMP_8_27_port, 
      OTMP_8_26_port, OTMP_8_25_port, OTMP_8_24_port, OTMP_8_23_port, 
      OTMP_8_22_port, OTMP_8_21_port, OTMP_8_20_port, OTMP_8_19_port, 
      OTMP_8_18_port, OTMP_8_17_port, OTMP_8_16_port, PTMP_8_15_port, 
      PTMP_8_14_port, PTMP_8_13_port, PTMP_8_12_port, PTMP_8_11_port, 
      PTMP_8_10_port, PTMP_8_9_port, PTMP_8_8_port, PTMP_8_7_port, 
      PTMP_8_6_port, PTMP_8_5_port, PTMP_8_4_port, PTMP_8_3_port, PTMP_8_2_port
      , PTMP_8_1_port, PTMP_8_0_port, PTMP_7_49_port, PTMP_7_48_port, 
      PTMP_7_47_port, PTMP_7_46_port, PTMP_7_45_port, PTMP_7_44_port, 
      PTMP_7_43_port, PTMP_7_42_port, PTMP_7_41_port, PTMP_7_40_port, 
      PTMP_7_39_port, PTMP_7_38_port, PTMP_7_37_port, PTMP_7_36_port, 
      PTMP_7_35_port, PTMP_7_34_port, PTMP_7_33_port, PTMP_7_32_port, 
      PTMP_7_31_port, PTMP_7_30_port, PTMP_7_29_port, PTMP_7_28_port, 
      PTMP_7_27_port, PTMP_7_26_port, PTMP_7_25_port, PTMP_7_24_port, 
      PTMP_7_23_port, PTMP_7_22_port, PTMP_7_21_port, PTMP_7_20_port, 
      PTMP_7_19_port, PTMP_7_18_port, PTMP_7_17_port, PTMP_7_16_port, 
      PTMP_7_15_port, PTMP_7_14_port, PTMP_7_13_port, PTMP_7_12_port, 
      PTMP_7_11_port, PTMP_7_10_port, PTMP_7_9_port, PTMP_7_8_port, 
      PTMP_7_7_port, PTMP_7_6_port, PTMP_7_5_port, PTMP_7_4_port, PTMP_7_3_port
      , PTMP_7_2_port, PTMP_7_1_port, PTMP_7_0_port, PTMP_6_47_port, 
      PTMP_6_46_port, PTMP_6_45_port, PTMP_6_44_port, PTMP_6_43_port, 
      PTMP_6_42_port, PTMP_6_41_port, PTMP_6_40_port, PTMP_6_39_port, 
      PTMP_6_38_port, PTMP_6_37_port, PTMP_6_36_port, PTMP_6_35_port, 
      PTMP_6_34_port, PTMP_6_33_port, PTMP_6_32_port, PTMP_6_31_port, 
      PTMP_6_30_port, PTMP_6_29_port, PTMP_6_28_port, PTMP_6_27_port, 
      PTMP_6_26_port, PTMP_6_25_port, PTMP_6_24_port, PTMP_6_23_port, 
      PTMP_6_22_port, PTMP_6_21_port, PTMP_6_20_port, PTMP_6_19_port, 
      PTMP_6_18_port, PTMP_6_17_port, PTMP_6_16_port, PTMP_6_15_port, 
      PTMP_6_14_port, PTMP_6_13_port, PTMP_6_12_port, PTMP_6_11_port, 
      PTMP_6_10_port, PTMP_6_9_port, PTMP_6_8_port, PTMP_6_7_port, 
      PTMP_6_6_port, PTMP_6_5_port, PTMP_6_4_port, PTMP_6_3_port, PTMP_6_2_port
      , PTMP_6_1_port, PTMP_6_0_port, PTMP_5_45_port, PTMP_5_44_port, 
      PTMP_5_43_port, PTMP_5_42_port, PTMP_5_41_port, PTMP_5_40_port, 
      PTMP_5_39_port, PTMP_5_38_port, PTMP_5_37_port, PTMP_5_36_port, 
      PTMP_5_35_port, PTMP_5_34_port, PTMP_5_33_port, PTMP_5_32_port, 
      PTMP_5_31_port, PTMP_5_30_port, PTMP_5_29_port, PTMP_5_28_port, 
      PTMP_5_27_port, PTMP_5_26_port, PTMP_5_25_port, PTMP_5_24_port, 
      PTMP_5_23_port, PTMP_5_22_port, PTMP_5_21_port, PTMP_5_20_port, 
      PTMP_5_19_port, PTMP_5_18_port, PTMP_5_17_port, PTMP_5_16_port, 
      PTMP_5_15_port, PTMP_5_14_port, PTMP_5_13_port, PTMP_5_12_port, 
      PTMP_5_11_port, PTMP_5_10_port, PTMP_5_9_port, PTMP_5_8_port, 
      PTMP_5_7_port, PTMP_5_6_port, PTMP_5_5_port, PTMP_5_4_port, PTMP_5_3_port
      , PTMP_5_2_port, PTMP_5_1_port, PTMP_5_0_port, PTMP_4_43_port, 
      PTMP_4_42_port, PTMP_4_41_port, PTMP_4_40_port, PTMP_4_39_port, 
      PTMP_4_38_port, PTMP_4_37_port, PTMP_4_36_port, PTMP_4_35_port, 
      PTMP_4_34_port, PTMP_4_33_port, PTMP_4_32_port, PTMP_4_31_port, 
      PTMP_4_30_port, PTMP_4_29_port, PTMP_4_28_port, PTMP_4_27_port, 
      PTMP_4_26_port, PTMP_4_25_port, PTMP_4_24_port, PTMP_4_23_port, 
      PTMP_4_22_port, PTMP_4_21_port, PTMP_4_20_port, PTMP_4_19_port, 
      PTMP_4_18_port, PTMP_4_17_port, PTMP_4_16_port, PTMP_4_15_port, 
      PTMP_4_14_port, PTMP_4_13_port, PTMP_4_12_port, PTMP_4_11_port, 
      PTMP_4_10_port, PTMP_4_9_port, PTMP_4_8_port, PTMP_4_7_port, 
      PTMP_4_6_port, PTMP_4_5_port, PTMP_4_4_port, PTMP_4_3_port, PTMP_4_2_port
      , PTMP_4_1_port, PTMP_4_0_port, PTMP_3_41_port, PTMP_3_40_port, 
      PTMP_3_39_port, PTMP_3_38_port, PTMP_3_37_port, PTMP_3_36_port, 
      PTMP_3_35_port, PTMP_3_34_port, PTMP_3_33_port, PTMP_3_32_port, 
      PTMP_3_31_port, PTMP_3_30_port, PTMP_3_29_port, PTMP_3_28_port, 
      PTMP_3_27_port, PTMP_3_26_port, PTMP_3_25_port, PTMP_3_24_port, 
      PTMP_3_23_port, PTMP_3_22_port, PTMP_3_21_port, PTMP_3_20_port, 
      PTMP_3_19_port, PTMP_3_18_port, PTMP_3_17_port, PTMP_3_16_port, 
      PTMP_3_15_port, PTMP_3_14_port, PTMP_3_13_port, PTMP_3_12_port, 
      PTMP_3_11_port, PTMP_3_10_port, PTMP_3_9_port, PTMP_3_8_port, 
      PTMP_3_7_port, PTMP_3_6_port, PTMP_3_5_port, PTMP_3_4_port, PTMP_3_3_port
      , PTMP_3_2_port, PTMP_3_1_port, PTMP_3_0_port, PTMP_2_39_port, 
      PTMP_2_38_port, PTMP_2_37_port, PTMP_2_36_port, PTMP_2_35_port, 
      PTMP_2_34_port, PTMP_2_33_port, PTMP_2_32_port, PTMP_2_31_port, 
      PTMP_2_30_port, PTMP_2_29_port, PTMP_2_28_port, PTMP_2_27_port, 
      PTMP_2_26_port, PTMP_2_25_port, PTMP_2_24_port, PTMP_2_23_port, 
      PTMP_2_22_port, PTMP_2_21_port, PTMP_2_20_port, PTMP_2_19_port, 
      PTMP_2_18_port, PTMP_2_17_port, PTMP_2_16_port, PTMP_2_15_port, 
      PTMP_2_14_port, PTMP_2_13_port, PTMP_2_12_port, PTMP_2_11_port, 
      PTMP_2_10_port, PTMP_2_9_port, PTMP_2_8_port, PTMP_2_7_port, 
      PTMP_2_6_port, PTMP_2_5_port, PTMP_2_4_port, PTMP_2_3_port, PTMP_2_2_port
      , PTMP_2_1_port, PTMP_2_0_port, PTMP_1_37_port, PTMP_1_36_port, 
      PTMP_1_35_port, PTMP_1_34_port, PTMP_1_33_port, PTMP_1_32_port, 
      PTMP_1_31_port, PTMP_1_30_port, PTMP_1_29_port, PTMP_1_28_port, 
      PTMP_1_27_port, PTMP_1_26_port, PTMP_1_25_port, PTMP_1_24_port, 
      PTMP_1_23_port, PTMP_1_22_port, PTMP_1_21_port, PTMP_1_20_port, 
      PTMP_1_19_port, PTMP_1_18_port, PTMP_1_17_port, PTMP_1_16_port, 
      PTMP_1_15_port, PTMP_1_14_port, PTMP_1_13_port, PTMP_1_12_port, 
      PTMP_1_11_port, PTMP_1_10_port, PTMP_1_9_port, PTMP_1_8_port, 
      PTMP_1_7_port, PTMP_1_6_port, PTMP_1_5_port, PTMP_1_4_port, PTMP_1_3_port
      , PTMP_1_2_port, PTMP_1_1_port, PTMP_1_0_port, PTMP_0_36_port, 
      PTMP_0_34_port, PTMP_0_33_port, PTMP_0_32_port, PTMP_0_31_port, 
      PTMP_0_30_port, PTMP_0_29_port, PTMP_0_28_port, PTMP_0_27_port, 
      PTMP_0_26_port, PTMP_0_25_port, PTMP_0_24_port, PTMP_0_23_port, 
      PTMP_0_22_port, PTMP_0_21_port, PTMP_0_20_port, PTMP_0_19_port, 
      PTMP_0_18_port, PTMP_0_17_port, PTMP_0_16_port, PTMP_0_15_port, 
      PTMP_0_14_port, PTMP_0_13_port, PTMP_0_12_port, PTMP_0_11_port, 
      PTMP_0_10_port, PTMP_0_9_port, PTMP_0_8_port, PTMP_0_7_port, 
      PTMP_0_6_port, PTMP_0_5_port, PTMP_0_4_port, PTMP_0_3_port, PTMP_0_2_port
      , PTMP_0_1_port, PTMP_0_0_port, PTMP_13_61_port, PTMP_13_60_port, 
      PTMP_13_59_port, PTMP_13_58_port, PTMP_13_57_port, PTMP_13_56_port, 
      PTMP_13_55_port, PTMP_13_54_port, PTMP_13_53_port, PTMP_13_52_port, 
      PTMP_13_51_port, PTMP_13_50_port, PTMP_13_49_port, PTMP_13_48_port, 
      PTMP_13_47_port, PTMP_13_46_port, PTMP_13_45_port, PTMP_13_44_port, 
      PTMP_13_43_port, PTMP_13_42_port, PTMP_13_41_port, PTMP_13_40_port, 
      PTMP_13_39_port, PTMP_13_38_port, PTMP_13_37_port, PTMP_13_36_port, 
      PTMP_13_35_port, PTMP_13_34_port, PTMP_13_33_port, PTMP_13_32_port, 
      PTMP_13_31_port, PTMP_13_30_port, PTMP_13_29_port, PTMP_13_28_port, 
      PTMP_13_27_port, PTMP_13_26_port, PTMP_13_25_port, PTMP_13_24_port, 
      PTMP_13_23_port, PTMP_13_22_port, PTMP_13_21_port, PTMP_13_20_port, 
      PTMP_13_19_port, PTMP_13_18_port, PTMP_13_17_port, PTMP_13_16_port, 
      PTMP_13_15_port, PTMP_13_14_port, PTMP_13_13_port, PTMP_13_12_port, 
      PTMP_13_11_port, PTMP_13_10_port, PTMP_13_9_port, PTMP_13_8_port, 
      PTMP_13_7_port, PTMP_13_6_port, PTMP_13_5_port, PTMP_13_4_port, 
      PTMP_13_3_port, PTMP_13_2_port, PTMP_13_1_port, PTMP_13_0_port, 
      PTMP_12_59_port, PTMP_12_58_port, PTMP_12_57_port, PTMP_12_56_port, 
      PTMP_12_55_port, PTMP_12_54_port, PTMP_12_53_port, PTMP_12_52_port, 
      PTMP_12_51_port, PTMP_12_50_port, PTMP_12_49_port, PTMP_12_48_port, 
      PTMP_12_47_port, PTMP_12_46_port, PTMP_12_45_port, PTMP_12_44_port, 
      PTMP_12_43_port, PTMP_12_42_port, PTMP_12_41_port, PTMP_12_40_port, 
      PTMP_12_39_port, PTMP_12_38_port, PTMP_12_37_port, PTMP_12_36_port, 
      PTMP_12_35_port, PTMP_12_34_port, PTMP_12_33_port, PTMP_12_32_port, 
      PTMP_12_31_port, PTMP_12_30_port, PTMP_12_29_port, PTMP_12_28_port, 
      PTMP_12_27_port, PTMP_12_26_port, PTMP_12_25_port, PTMP_12_24_port, 
      PTMP_12_23_port, PTMP_12_22_port, PTMP_12_21_port, PTMP_12_20_port, 
      PTMP_12_19_port, PTMP_12_18_port, PTMP_12_17_port, PTMP_12_16_port, 
      PTMP_12_15_port, PTMP_12_14_port, PTMP_12_13_port, PTMP_12_12_port, 
      PTMP_12_11_port, PTMP_12_10_port, PTMP_12_9_port, PTMP_12_8_port, 
      PTMP_12_7_port, PTMP_12_6_port, PTMP_12_5_port, PTMP_12_4_port, 
      PTMP_12_3_port, PTMP_12_2_port, PTMP_12_1_port, PTMP_12_0_port, 
      PTMP_11_57_port, PTMP_11_56_port, PTMP_11_55_port, PTMP_11_54_port, 
      PTMP_11_53_port, PTMP_11_52_port, PTMP_11_51_port, PTMP_11_50_port, 
      PTMP_11_49_port, PTMP_11_48_port, PTMP_11_47_port, PTMP_11_46_port, 
      PTMP_11_45_port, PTMP_11_44_port, PTMP_11_43_port, PTMP_11_42_port, 
      PTMP_11_41_port, PTMP_11_40_port, PTMP_11_39_port, PTMP_11_38_port, 
      PTMP_11_37_port, PTMP_11_36_port, PTMP_11_35_port, PTMP_11_34_port, 
      PTMP_11_33_port, PTMP_11_32_port, PTMP_11_31_port, PTMP_11_30_port, 
      PTMP_11_29_port, PTMP_11_28_port, PTMP_11_27_port, PTMP_11_26_port, 
      PTMP_11_25_port, PTMP_11_24_port, PTMP_11_23_port, PTMP_11_22_port, 
      PTMP_11_21_port, PTMP_11_20_port, PTMP_11_19_port, PTMP_11_18_port, 
      PTMP_11_17_port, PTMP_11_16_port, PTMP_11_15_port, PTMP_11_14_port, 
      PTMP_11_13_port, PTMP_11_12_port, PTMP_11_11_port, PTMP_11_10_port, 
      PTMP_11_9_port, PTMP_11_8_port, PTMP_11_7_port, PTMP_11_6_port, 
      PTMP_11_5_port, PTMP_11_4_port, PTMP_11_3_port, PTMP_11_2_port, 
      PTMP_11_1_port, PTMP_11_0_port, PTMP_10_55_port, PTMP_10_54_port, 
      PTMP_10_53_port, PTMP_10_52_port, PTMP_10_51_port, PTMP_10_50_port, 
      PTMP_10_49_port, PTMP_10_48_port, PTMP_10_47_port, PTMP_10_46_port, 
      PTMP_10_45_port, PTMP_10_44_port, PTMP_10_43_port, PTMP_10_42_port, 
      PTMP_10_41_port, PTMP_10_40_port, PTMP_10_39_port, PTMP_10_38_port, 
      PTMP_10_37_port, PTMP_10_36_port, PTMP_10_35_port, PTMP_10_34_port, 
      PTMP_10_33_port, PTMP_10_32_port, PTMP_10_31_port, PTMP_10_30_port, 
      PTMP_10_29_port, PTMP_10_28_port, PTMP_10_27_port, PTMP_10_26_port, 
      PTMP_10_25_port, PTMP_10_24_port, PTMP_10_23_port, PTMP_10_22_port, 
      PTMP_10_21_port, PTMP_10_20_port, PTMP_10_19_port, PTMP_10_18_port, 
      PTMP_10_17_port, PTMP_10_16_port, PTMP_10_15_port, PTMP_10_14_port, 
      PTMP_10_13_port, PTMP_10_12_port, PTMP_10_11_port, PTMP_10_10_port, 
      PTMP_10_9_port, PTMP_10_8_port, PTMP_10_7_port, PTMP_10_6_port, 
      PTMP_10_5_port, PTMP_10_4_port, PTMP_10_3_port, PTMP_10_2_port, 
      PTMP_10_1_port, PTMP_10_0_port, PTMP_9_53_port, PTMP_9_52_port, 
      PTMP_9_51_port, PTMP_9_50_port, PTMP_9_49_port, PTMP_9_48_port, 
      PTMP_9_47_port, PTMP_9_46_port, PTMP_9_45_port, PTMP_9_44_port, 
      PTMP_9_43_port, PTMP_9_42_port, PTMP_9_41_port, PTMP_9_40_port, 
      PTMP_9_39_port, PTMP_9_38_port, PTMP_9_37_port, PTMP_9_36_port, 
      PTMP_9_35_port, PTMP_9_34_port, PTMP_9_33_port, PTMP_9_32_port, 
      PTMP_9_31_port, PTMP_9_30_port, PTMP_9_29_port, PTMP_9_28_port, 
      PTMP_9_27_port, PTMP_9_26_port, PTMP_9_25_port, PTMP_9_24_port, 
      PTMP_9_23_port, PTMP_9_22_port, PTMP_9_21_port, PTMP_9_20_port, 
      PTMP_9_19_port, PTMP_9_18_port, PTMP_9_17_port, PTMP_9_16_port, 
      PTMP_9_15_port, PTMP_9_14_port, PTMP_9_13_port, PTMP_9_12_port, 
      PTMP_9_11_port, PTMP_9_10_port, PTMP_9_9_port, PTMP_9_8_port, 
      PTMP_9_7_port, PTMP_9_6_port, PTMP_9_5_port, PTMP_9_4_port, PTMP_9_3_port
      , PTMP_9_2_port, PTMP_9_1_port, PTMP_9_0_port, PTMP_8_51_port, 
      PTMP_8_50_port, PTMP_8_49_port, PTMP_8_48_port, PTMP_8_47_port, 
      PTMP_8_46_port, PTMP_8_45_port, PTMP_8_44_port, PTMP_8_43_port, 
      PTMP_8_42_port, PTMP_8_41_port, PTMP_8_40_port, PTMP_8_39_port, 
      PTMP_8_38_port, PTMP_8_37_port, PTMP_8_36_port, PTMP_8_35_port, 
      PTMP_8_34_port, PTMP_8_33_port, PTMP_8_32_port, PTMP_8_31_port, 
      PTMP_8_30_port, PTMP_8_29_port, PTMP_8_28_port, PTMP_8_27_port, 
      PTMP_8_26_port, PTMP_8_25_port, PTMP_8_24_port, PTMP_8_23_port, 
      PTMP_8_22_port, PTMP_8_21_port, PTMP_8_20_port, PTMP_8_19_port, 
      PTMP_8_18_port, PTMP_8_17_port, PTMP_8_16_port, n1, n2, n_1080, n_1081, 
      n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, 
      n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, 
      n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, 
      n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, 
      n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, 
      n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, 
      n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, 
      n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, 
      n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, 
      n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, 
      n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, 
      n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, 
      n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, 
      n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, 
      n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, 
      n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, 
      n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, 
      n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, 
      n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, 
      n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, 
      n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, 
      n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, 
      n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, 
      n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296 : 
      std_logic;

begin
   
   X_Logic0_port <= '0';
   n1 <= '0';
   n2 <= '0';
   ENC1 : BOOTHENC_NBIT34_i0 port map( A_s(33) => A(31), A_s(32) => A(31), 
                           A_s(31) => A(31), A_s(30) => A(30), A_s(29) => A(29)
                           , A_s(28) => A(28), A_s(27) => A(27), A_s(26) => 
                           A(26), A_s(25) => A(25), A_s(24) => A(24), A_s(23) 
                           => A(23), A_s(22) => A(22), A_s(21) => A(21), 
                           A_s(20) => A(20), A_s(19) => A(19), A_s(18) => A(18)
                           , A_s(17) => A(17), A_s(16) => A(16), A_s(15) => 
                           A(15), A_s(14) => A(14), A_s(13) => A(13), A_s(12) 
                           => A(12), A_s(11) => A(11), A_s(10) => A(10), A_s(9)
                           => A(9), A_s(8) => A(8), A_s(7) => A(7), A_s(6) => 
                           A(6), A_s(5) => A(5), A_s(4) => A(4), A_s(3) => A(3)
                           , A_s(2) => A(2), A_s(1) => A(1), A_s(0) => A(0), 
                           A_ns(33) => A_n_65, A_ns(32) => A_n_65, A_ns(31) => 
                           A_n_65, A_ns(30) => A_n_30_port, A_ns(29) => 
                           A_n_29_port, A_ns(28) => A_n_28_port, A_ns(27) => 
                           A_n_27_port, A_ns(26) => A_n_26_port, A_ns(25) => 
                           A_n_25_port, A_ns(24) => A_n_24_port, A_ns(23) => 
                           A_n_23_port, A_ns(22) => A_n_22_port, A_ns(21) => 
                           A_n_21_port, A_ns(20) => A_n_20_port, A_ns(19) => 
                           A_n_19_port, A_ns(18) => A_n_18_port, A_ns(17) => 
                           A_n_17_port, A_ns(16) => A_n_16_port, A_ns(15) => 
                           A_n_15_port, A_ns(14) => A_n_14_port, A_ns(13) => 
                           A_n_13_port, A_ns(12) => A_n_12_port, A_ns(11) => 
                           A_n_11_port, A_ns(10) => A_n_10_port, A_ns(9) => 
                           A_n_9_port, A_ns(8) => A_n_8_port, A_ns(7) => 
                           A_n_7_port, A_ns(6) => A_n_6_port, A_ns(5) => 
                           A_n_5_port, A_ns(4) => A_n_4_port, A_ns(3) => 
                           A_n_3_port, A_ns(2) => A_n_2_port, A_ns(1) => 
                           A_n_1_port, A_ns(0) => A_n_0_port, B(33) => B(31), 
                           B(32) => B(31), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), O(33) => OTMP_0_34_port, O(32) 
                           => OTMP_0_32_port, O(31) => OTMP_0_31_port, O(30) =>
                           OTMP_0_30_port, O(29) => OTMP_0_29_port, O(28) => 
                           OTMP_0_28_port, O(27) => OTMP_0_27_port, O(26) => 
                           OTMP_0_26_port, O(25) => OTMP_0_25_port, O(24) => 
                           OTMP_0_24_port, O(23) => OTMP_0_23_port, O(22) => 
                           OTMP_0_22_port, O(21) => OTMP_0_21_port, O(20) => 
                           OTMP_0_20_port, O(19) => OTMP_0_19_port, O(18) => 
                           OTMP_0_18_port, O(17) => OTMP_0_17_port, O(16) => 
                           OTMP_0_16_port, O(15) => OTMP_0_15_port, O(14) => 
                           OTMP_0_14_port, O(13) => OTMP_0_13_port, O(12) => 
                           OTMP_0_12_port, O(11) => OTMP_0_11_port, O(10) => 
                           OTMP_0_10_port, O(9) => OTMP_0_9_port, O(8) => 
                           OTMP_0_8_port, O(7) => OTMP_0_7_port, O(6) => 
                           OTMP_0_6_port, O(5) => OTMP_0_5_port, O(4) => 
                           OTMP_0_4_port, O(3) => OTMP_0_3_port, O(2) => 
                           OTMP_0_2_port, O(1) => OTMP_0_1_port, O(0) => 
                           OTMP_0_0_port, A_so(33) => SHIFT_1_33_port, A_so(32)
                           => SHIFT_1_32_port, A_so(31) => SHIFT_1_31_port, 
                           A_so(30) => SHIFT_1_30_port, A_so(29) => 
                           SHIFT_1_29_port, A_so(28) => SHIFT_1_28_port, 
                           A_so(27) => SHIFT_1_27_port, A_so(26) => 
                           SHIFT_1_26_port, A_so(25) => SHIFT_1_25_port, 
                           A_so(24) => SHIFT_1_24_port, A_so(23) => 
                           SHIFT_1_23_port, A_so(22) => SHIFT_1_22_port, 
                           A_so(21) => SHIFT_1_21_port, A_so(20) => 
                           SHIFT_1_20_port, A_so(19) => SHIFT_1_19_port, 
                           A_so(18) => SHIFT_1_18_port, A_so(17) => 
                           SHIFT_1_17_port, A_so(16) => SHIFT_1_16_port, 
                           A_so(15) => SHIFT_1_15_port, A_so(14) => 
                           SHIFT_1_14_port, A_so(13) => SHIFT_1_13_port, 
                           A_so(12) => SHIFT_1_12_port, A_so(11) => 
                           SHIFT_1_11_port, A_so(10) => SHIFT_1_10_port, 
                           A_so(9) => SHIFT_1_9_port, A_so(8) => SHIFT_1_8_port
                           , A_so(7) => SHIFT_1_7_port, A_so(6) => 
                           SHIFT_1_6_port, A_so(5) => SHIFT_1_5_port, A_so(4) 
                           => SHIFT_1_4_port, A_so(3) => SHIFT_1_3_port, 
                           A_so(2) => SHIFT_1_2_port, A_so(1) => SHIFT_1_1_port
                           , A_so(0) => n_1080, A_nso(33) => SHIFT_n_1_33_port,
                           A_nso(32) => SHIFT_n_1_32_port, A_nso(31) => 
                           SHIFT_n_1_31_port, A_nso(30) => SHIFT_n_1_30_port, 
                           A_nso(29) => SHIFT_n_1_29_port, A_nso(28) => 
                           SHIFT_n_1_28_port, A_nso(27) => SHIFT_n_1_27_port, 
                           A_nso(26) => SHIFT_n_1_26_port, A_nso(25) => 
                           SHIFT_n_1_25_port, A_nso(24) => SHIFT_n_1_24_port, 
                           A_nso(23) => SHIFT_n_1_23_port, A_nso(22) => 
                           SHIFT_n_1_22_port, A_nso(21) => SHIFT_n_1_21_port, 
                           A_nso(20) => SHIFT_n_1_20_port, A_nso(19) => 
                           SHIFT_n_1_19_port, A_nso(18) => SHIFT_n_1_18_port, 
                           A_nso(17) => SHIFT_n_1_17_port, A_nso(16) => 
                           SHIFT_n_1_16_port, A_nso(15) => SHIFT_n_1_15_port, 
                           A_nso(14) => SHIFT_n_1_14_port, A_nso(13) => 
                           SHIFT_n_1_13_port, A_nso(12) => SHIFT_n_1_12_port, 
                           A_nso(11) => SHIFT_n_1_11_port, A_nso(10) => 
                           SHIFT_n_1_10_port, A_nso(9) => SHIFT_n_1_9_port, 
                           A_nso(8) => SHIFT_n_1_8_port, A_nso(7) => 
                           SHIFT_n_1_7_port, A_nso(6) => SHIFT_n_1_6_port, 
                           A_nso(5) => SHIFT_n_1_5_port, A_nso(4) => 
                           SHIFT_n_1_4_port, A_nso(3) => SHIFT_n_1_3_port, 
                           A_nso(2) => SHIFT_n_1_2_port, A_nso(1) => 
                           SHIFT_n_1_1_port, A_nso(0) => n_1081);
   ENC_1 : BOOTHENC_NBIT36_i2 port map( A_s(35) => SHIFT_1_33_port, A_s(34) => 
                           SHIFT_1_33_port, A_s(33) => SHIFT_1_33_port, A_s(32)
                           => SHIFT_1_32_port, A_s(31) => SHIFT_1_31_port, 
                           A_s(30) => SHIFT_1_30_port, A_s(29) => 
                           SHIFT_1_29_port, A_s(28) => SHIFT_1_28_port, A_s(27)
                           => SHIFT_1_27_port, A_s(26) => SHIFT_1_26_port, 
                           A_s(25) => SHIFT_1_25_port, A_s(24) => 
                           SHIFT_1_24_port, A_s(23) => SHIFT_1_23_port, A_s(22)
                           => SHIFT_1_22_port, A_s(21) => SHIFT_1_21_port, 
                           A_s(20) => SHIFT_1_20_port, A_s(19) => 
                           SHIFT_1_19_port, A_s(18) => SHIFT_1_18_port, A_s(17)
                           => SHIFT_1_17_port, A_s(16) => SHIFT_1_16_port, 
                           A_s(15) => SHIFT_1_15_port, A_s(14) => 
                           SHIFT_1_14_port, A_s(13) => SHIFT_1_13_port, A_s(12)
                           => SHIFT_1_12_port, A_s(11) => SHIFT_1_11_port, 
                           A_s(10) => SHIFT_1_10_port, A_s(9) => SHIFT_1_9_port
                           , A_s(8) => SHIFT_1_8_port, A_s(7) => SHIFT_1_7_port
                           , A_s(6) => SHIFT_1_6_port, A_s(5) => SHIFT_1_5_port
                           , A_s(4) => SHIFT_1_4_port, A_s(3) => SHIFT_1_3_port
                           , A_s(2) => SHIFT_1_2_port, A_s(1) => SHIFT_1_1_port
                           , A_s(0) => SHIFT_1_0_port, A_ns(35) => 
                           SHIFT_n_1_33_port, A_ns(34) => SHIFT_n_1_33_port, 
                           A_ns(33) => SHIFT_n_1_33_port, A_ns(32) => 
                           SHIFT_n_1_32_port, A_ns(31) => SHIFT_n_1_31_port, 
                           A_ns(30) => SHIFT_n_1_30_port, A_ns(29) => 
                           SHIFT_n_1_29_port, A_ns(28) => SHIFT_n_1_28_port, 
                           A_ns(27) => SHIFT_n_1_27_port, A_ns(26) => 
                           SHIFT_n_1_26_port, A_ns(25) => SHIFT_n_1_25_port, 
                           A_ns(24) => SHIFT_n_1_24_port, A_ns(23) => 
                           SHIFT_n_1_23_port, A_ns(22) => SHIFT_n_1_22_port, 
                           A_ns(21) => SHIFT_n_1_21_port, A_ns(20) => 
                           SHIFT_n_1_20_port, A_ns(19) => SHIFT_n_1_19_port, 
                           A_ns(18) => SHIFT_n_1_18_port, A_ns(17) => 
                           SHIFT_n_1_17_port, A_ns(16) => SHIFT_n_1_16_port, 
                           A_ns(15) => SHIFT_n_1_15_port, A_ns(14) => 
                           SHIFT_n_1_14_port, A_ns(13) => SHIFT_n_1_13_port, 
                           A_ns(12) => SHIFT_n_1_12_port, A_ns(11) => 
                           SHIFT_n_1_11_port, A_ns(10) => SHIFT_n_1_10_port, 
                           A_ns(9) => SHIFT_n_1_9_port, A_ns(8) => 
                           SHIFT_n_1_8_port, A_ns(7) => SHIFT_n_1_7_port, 
                           A_ns(6) => SHIFT_n_1_6_port, A_ns(5) => 
                           SHIFT_n_1_5_port, A_ns(4) => SHIFT_n_1_4_port, 
                           A_ns(3) => SHIFT_n_1_3_port, A_ns(2) => 
                           SHIFT_n_1_2_port, A_ns(1) => SHIFT_n_1_1_port, 
                           A_ns(0) => SHIFT_n_1_0_port, B(35) => B(31), B(34) 
                           => B(31), B(33) => B(31), B(32) => B(31), B(31) => 
                           B(31), B(30) => B(30), B(29) => B(29), B(28) => 
                           B(28), B(27) => B(27), B(26) => B(26), B(25) => 
                           B(25), B(24) => B(24), B(23) => B(23), B(22) => 
                           B(22), B(21) => B(21), B(20) => B(20), B(19) => 
                           B(19), B(18) => B(18), B(17) => B(17), B(16) => 
                           B(16), B(15) => B(15), B(14) => B(14), B(13) => 
                           B(13), B(12) => B(12), B(11) => B(11), B(10) => 
                           B(10), B(9) => B(9), B(8) => B(8), B(7) => B(7), 
                           B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3) => 
                           B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), 
                           O(35) => OTMP_1_35_port, O(34) => OTMP_1_34_port, 
                           O(33) => OTMP_1_33_port, O(32) => OTMP_1_32_port, 
                           O(31) => OTMP_1_31_port, O(30) => OTMP_1_30_port, 
                           O(29) => OTMP_1_29_port, O(28) => OTMP_1_28_port, 
                           O(27) => OTMP_1_27_port, O(26) => OTMP_1_26_port, 
                           O(25) => OTMP_1_25_port, O(24) => OTMP_1_24_port, 
                           O(23) => OTMP_1_23_port, O(22) => OTMP_1_22_port, 
                           O(21) => OTMP_1_21_port, O(20) => OTMP_1_20_port, 
                           O(19) => OTMP_1_19_port, O(18) => OTMP_1_18_port, 
                           O(17) => OTMP_1_17_port, O(16) => OTMP_1_16_port, 
                           O(15) => OTMP_1_15_port, O(14) => OTMP_1_14_port, 
                           O(13) => OTMP_1_13_port, O(12) => OTMP_1_12_port, 
                           O(11) => OTMP_1_11_port, O(10) => OTMP_1_10_port, 
                           O(9) => OTMP_1_9_port, O(8) => OTMP_1_8_port, O(7) 
                           => OTMP_1_7_port, O(6) => OTMP_1_6_port, O(5) => 
                           OTMP_1_5_port, O(4) => OTMP_1_4_port, O(3) => 
                           OTMP_1_3_port, O(2) => OTMP_1_2_port, O(1) => 
                           OTMP_1_1_port, O(0) => n_1082, A_so(35) => 
                           SHIFT_2_35_port, A_so(34) => SHIFT_2_34_port, 
                           A_so(33) => SHIFT_2_33_port, A_so(32) => 
                           SHIFT_2_32_port, A_so(31) => SHIFT_2_31_port, 
                           A_so(30) => SHIFT_2_30_port, A_so(29) => 
                           SHIFT_2_29_port, A_so(28) => SHIFT_2_28_port, 
                           A_so(27) => SHIFT_2_27_port, A_so(26) => 
                           SHIFT_2_26_port, A_so(25) => SHIFT_2_25_port, 
                           A_so(24) => SHIFT_2_24_port, A_so(23) => 
                           SHIFT_2_23_port, A_so(22) => SHIFT_2_22_port, 
                           A_so(21) => SHIFT_2_21_port, A_so(20) => 
                           SHIFT_2_20_port, A_so(19) => SHIFT_2_19_port, 
                           A_so(18) => SHIFT_2_18_port, A_so(17) => 
                           SHIFT_2_17_port, A_so(16) => SHIFT_2_16_port, 
                           A_so(15) => SHIFT_2_15_port, A_so(14) => 
                           SHIFT_2_14_port, A_so(13) => SHIFT_2_13_port, 
                           A_so(12) => SHIFT_2_12_port, A_so(11) => 
                           SHIFT_2_11_port, A_so(10) => SHIFT_2_10_port, 
                           A_so(9) => SHIFT_2_9_port, A_so(8) => SHIFT_2_8_port
                           , A_so(7) => SHIFT_2_7_port, A_so(6) => 
                           SHIFT_2_6_port, A_so(5) => SHIFT_2_5_port, A_so(4) 
                           => SHIFT_2_4_port, A_so(3) => SHIFT_2_3_port, 
                           A_so(2) => SHIFT_2_2_port, A_so(1) => n_1083, 
                           A_so(0) => n_1084, A_nso(35) => SHIFT_n_2_35_port, 
                           A_nso(34) => SHIFT_n_2_34_port, A_nso(33) => 
                           SHIFT_n_2_33_port, A_nso(32) => SHIFT_n_2_32_port, 
                           A_nso(31) => SHIFT_n_2_31_port, A_nso(30) => 
                           SHIFT_n_2_30_port, A_nso(29) => SHIFT_n_2_29_port, 
                           A_nso(28) => SHIFT_n_2_28_port, A_nso(27) => 
                           SHIFT_n_2_27_port, A_nso(26) => SHIFT_n_2_26_port, 
                           A_nso(25) => SHIFT_n_2_25_port, A_nso(24) => 
                           SHIFT_n_2_24_port, A_nso(23) => SHIFT_n_2_23_port, 
                           A_nso(22) => SHIFT_n_2_22_port, A_nso(21) => 
                           SHIFT_n_2_21_port, A_nso(20) => SHIFT_n_2_20_port, 
                           A_nso(19) => SHIFT_n_2_19_port, A_nso(18) => 
                           SHIFT_n_2_18_port, A_nso(17) => SHIFT_n_2_17_port, 
                           A_nso(16) => SHIFT_n_2_16_port, A_nso(15) => 
                           SHIFT_n_2_15_port, A_nso(14) => SHIFT_n_2_14_port, 
                           A_nso(13) => SHIFT_n_2_13_port, A_nso(12) => 
                           SHIFT_n_2_12_port, A_nso(11) => SHIFT_n_2_11_port, 
                           A_nso(10) => SHIFT_n_2_10_port, A_nso(9) => 
                           SHIFT_n_2_9_port, A_nso(8) => SHIFT_n_2_8_port, 
                           A_nso(7) => SHIFT_n_2_7_port, A_nso(6) => 
                           SHIFT_n_2_6_port, A_nso(5) => SHIFT_n_2_5_port, 
                           A_nso(4) => SHIFT_n_2_4_port, A_nso(3) => 
                           SHIFT_n_2_3_port, A_nso(2) => SHIFT_n_2_2_port, 
                           A_nso(1) => n_1085, A_nso(0) => n_1086);
   ENC_2 : BOOTHENC_NBIT38_i4 port map( A_s(37) => SHIFT_2_35_port, A_s(36) => 
                           SHIFT_2_35_port, A_s(35) => SHIFT_2_35_port, A_s(34)
                           => SHIFT_2_34_port, A_s(33) => SHIFT_2_33_port, 
                           A_s(32) => SHIFT_2_32_port, A_s(31) => 
                           SHIFT_2_31_port, A_s(30) => SHIFT_2_30_port, A_s(29)
                           => SHIFT_2_29_port, A_s(28) => SHIFT_2_28_port, 
                           A_s(27) => SHIFT_2_27_port, A_s(26) => 
                           SHIFT_2_26_port, A_s(25) => SHIFT_2_25_port, A_s(24)
                           => SHIFT_2_24_port, A_s(23) => SHIFT_2_23_port, 
                           A_s(22) => SHIFT_2_22_port, A_s(21) => 
                           SHIFT_2_21_port, A_s(20) => SHIFT_2_20_port, A_s(19)
                           => SHIFT_2_19_port, A_s(18) => SHIFT_2_18_port, 
                           A_s(17) => SHIFT_2_17_port, A_s(16) => 
                           SHIFT_2_16_port, A_s(15) => SHIFT_2_15_port, A_s(14)
                           => SHIFT_2_14_port, A_s(13) => SHIFT_2_13_port, 
                           A_s(12) => SHIFT_2_12_port, A_s(11) => 
                           SHIFT_2_11_port, A_s(10) => SHIFT_2_10_port, A_s(9) 
                           => SHIFT_2_9_port, A_s(8) => SHIFT_2_8_port, A_s(7) 
                           => SHIFT_2_7_port, A_s(6) => SHIFT_2_6_port, A_s(5) 
                           => SHIFT_2_5_port, A_s(4) => SHIFT_2_4_port, A_s(3) 
                           => SHIFT_2_3_port, A_s(2) => SHIFT_2_2_port, A_s(1) 
                           => SHIFT_2_1_port, A_s(0) => SHIFT_2_0_port, 
                           A_ns(37) => SHIFT_n_2_35_port, A_ns(36) => 
                           SHIFT_n_2_35_port, A_ns(35) => SHIFT_n_2_35_port, 
                           A_ns(34) => SHIFT_n_2_34_port, A_ns(33) => 
                           SHIFT_n_2_33_port, A_ns(32) => SHIFT_n_2_32_port, 
                           A_ns(31) => SHIFT_n_2_31_port, A_ns(30) => 
                           SHIFT_n_2_30_port, A_ns(29) => SHIFT_n_2_29_port, 
                           A_ns(28) => SHIFT_n_2_28_port, A_ns(27) => 
                           SHIFT_n_2_27_port, A_ns(26) => SHIFT_n_2_26_port, 
                           A_ns(25) => SHIFT_n_2_25_port, A_ns(24) => 
                           SHIFT_n_2_24_port, A_ns(23) => SHIFT_n_2_23_port, 
                           A_ns(22) => SHIFT_n_2_22_port, A_ns(21) => 
                           SHIFT_n_2_21_port, A_ns(20) => SHIFT_n_2_20_port, 
                           A_ns(19) => SHIFT_n_2_19_port, A_ns(18) => 
                           SHIFT_n_2_18_port, A_ns(17) => SHIFT_n_2_17_port, 
                           A_ns(16) => SHIFT_n_2_16_port, A_ns(15) => 
                           SHIFT_n_2_15_port, A_ns(14) => SHIFT_n_2_14_port, 
                           A_ns(13) => SHIFT_n_2_13_port, A_ns(12) => 
                           SHIFT_n_2_12_port, A_ns(11) => SHIFT_n_2_11_port, 
                           A_ns(10) => SHIFT_n_2_10_port, A_ns(9) => 
                           SHIFT_n_2_9_port, A_ns(8) => SHIFT_n_2_8_port, 
                           A_ns(7) => SHIFT_n_2_7_port, A_ns(6) => 
                           SHIFT_n_2_6_port, A_ns(5) => SHIFT_n_2_5_port, 
                           A_ns(4) => SHIFT_n_2_4_port, A_ns(3) => 
                           SHIFT_n_2_3_port, A_ns(2) => SHIFT_n_2_2_port, 
                           A_ns(1) => SHIFT_n_2_1_port, A_ns(0) => 
                           SHIFT_n_2_0_port, B(37) => B(31), B(36) => B(31), 
                           B(35) => B(31), B(34) => B(31), B(33) => B(31), 
                           B(32) => B(31), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), O(37) => OTMP_2_37_port, O(36) 
                           => OTMP_2_36_port, O(35) => OTMP_2_35_port, O(34) =>
                           OTMP_2_34_port, O(33) => OTMP_2_33_port, O(32) => 
                           OTMP_2_32_port, O(31) => OTMP_2_31_port, O(30) => 
                           OTMP_2_30_port, O(29) => OTMP_2_29_port, O(28) => 
                           OTMP_2_28_port, O(27) => OTMP_2_27_port, O(26) => 
                           OTMP_2_26_port, O(25) => OTMP_2_25_port, O(24) => 
                           OTMP_2_24_port, O(23) => OTMP_2_23_port, O(22) => 
                           OTMP_2_22_port, O(21) => OTMP_2_21_port, O(20) => 
                           OTMP_2_20_port, O(19) => OTMP_2_19_port, O(18) => 
                           OTMP_2_18_port, O(17) => OTMP_2_17_port, O(16) => 
                           OTMP_2_16_port, O(15) => OTMP_2_15_port, O(14) => 
                           OTMP_2_14_port, O(13) => OTMP_2_13_port, O(12) => 
                           OTMP_2_12_port, O(11) => OTMP_2_11_port, O(10) => 
                           OTMP_2_10_port, O(9) => OTMP_2_9_port, O(8) => 
                           OTMP_2_8_port, O(7) => OTMP_2_7_port, O(6) => 
                           OTMP_2_6_port, O(5) => OTMP_2_5_port, O(4) => 
                           OTMP_2_4_port, O(3) => OTMP_2_3_port, O(2) => 
                           OTMP_2_2_port, O(1) => OTMP_2_1_port, O(0) => n_1087
                           , A_so(37) => SHIFT_3_37_port, A_so(36) => 
                           SHIFT_3_36_port, A_so(35) => SHIFT_3_35_port, 
                           A_so(34) => SHIFT_3_34_port, A_so(33) => 
                           SHIFT_3_33_port, A_so(32) => SHIFT_3_32_port, 
                           A_so(31) => SHIFT_3_31_port, A_so(30) => 
                           SHIFT_3_30_port, A_so(29) => SHIFT_3_29_port, 
                           A_so(28) => SHIFT_3_28_port, A_so(27) => 
                           SHIFT_3_27_port, A_so(26) => SHIFT_3_26_port, 
                           A_so(25) => SHIFT_3_25_port, A_so(24) => 
                           SHIFT_3_24_port, A_so(23) => SHIFT_3_23_port, 
                           A_so(22) => SHIFT_3_22_port, A_so(21) => 
                           SHIFT_3_21_port, A_so(20) => SHIFT_3_20_port, 
                           A_so(19) => SHIFT_3_19_port, A_so(18) => 
                           SHIFT_3_18_port, A_so(17) => SHIFT_3_17_port, 
                           A_so(16) => SHIFT_3_16_port, A_so(15) => 
                           SHIFT_3_15_port, A_so(14) => SHIFT_3_14_port, 
                           A_so(13) => SHIFT_3_13_port, A_so(12) => 
                           SHIFT_3_12_port, A_so(11) => SHIFT_3_11_port, 
                           A_so(10) => SHIFT_3_10_port, A_so(9) => 
                           SHIFT_3_9_port, A_so(8) => SHIFT_3_8_port, A_so(7) 
                           => SHIFT_3_7_port, A_so(6) => SHIFT_3_6_port, 
                           A_so(5) => SHIFT_3_5_port, A_so(4) => SHIFT_3_4_port
                           , A_so(3) => SHIFT_3_3_port, A_so(2) => 
                           SHIFT_3_2_port, A_so(1) => n_1088, A_so(0) => n_1089
                           , A_nso(37) => SHIFT_n_3_37_port, A_nso(36) => 
                           SHIFT_n_3_36_port, A_nso(35) => SHIFT_n_3_35_port, 
                           A_nso(34) => SHIFT_n_3_34_port, A_nso(33) => 
                           SHIFT_n_3_33_port, A_nso(32) => SHIFT_n_3_32_port, 
                           A_nso(31) => SHIFT_n_3_31_port, A_nso(30) => 
                           SHIFT_n_3_30_port, A_nso(29) => SHIFT_n_3_29_port, 
                           A_nso(28) => SHIFT_n_3_28_port, A_nso(27) => 
                           SHIFT_n_3_27_port, A_nso(26) => SHIFT_n_3_26_port, 
                           A_nso(25) => SHIFT_n_3_25_port, A_nso(24) => 
                           SHIFT_n_3_24_port, A_nso(23) => SHIFT_n_3_23_port, 
                           A_nso(22) => SHIFT_n_3_22_port, A_nso(21) => 
                           SHIFT_n_3_21_port, A_nso(20) => SHIFT_n_3_20_port, 
                           A_nso(19) => SHIFT_n_3_19_port, A_nso(18) => 
                           SHIFT_n_3_18_port, A_nso(17) => SHIFT_n_3_17_port, 
                           A_nso(16) => SHIFT_n_3_16_port, A_nso(15) => 
                           SHIFT_n_3_15_port, A_nso(14) => SHIFT_n_3_14_port, 
                           A_nso(13) => SHIFT_n_3_13_port, A_nso(12) => 
                           SHIFT_n_3_12_port, A_nso(11) => SHIFT_n_3_11_port, 
                           A_nso(10) => SHIFT_n_3_10_port, A_nso(9) => 
                           SHIFT_n_3_9_port, A_nso(8) => SHIFT_n_3_8_port, 
                           A_nso(7) => SHIFT_n_3_7_port, A_nso(6) => 
                           SHIFT_n_3_6_port, A_nso(5) => SHIFT_n_3_5_port, 
                           A_nso(4) => SHIFT_n_3_4_port, A_nso(3) => 
                           SHIFT_n_3_3_port, A_nso(2) => SHIFT_n_3_2_port, 
                           A_nso(1) => n_1090, A_nso(0) => n_1091);
   ENC_3 : BOOTHENC_NBIT40_i6 port map( A_s(39) => SHIFT_3_37_port, A_s(38) => 
                           SHIFT_3_37_port, A_s(37) => SHIFT_3_37_port, A_s(36)
                           => SHIFT_3_36_port, A_s(35) => SHIFT_3_35_port, 
                           A_s(34) => SHIFT_3_34_port, A_s(33) => 
                           SHIFT_3_33_port, A_s(32) => SHIFT_3_32_port, A_s(31)
                           => SHIFT_3_31_port, A_s(30) => SHIFT_3_30_port, 
                           A_s(29) => SHIFT_3_29_port, A_s(28) => 
                           SHIFT_3_28_port, A_s(27) => SHIFT_3_27_port, A_s(26)
                           => SHIFT_3_26_port, A_s(25) => SHIFT_3_25_port, 
                           A_s(24) => SHIFT_3_24_port, A_s(23) => 
                           SHIFT_3_23_port, A_s(22) => SHIFT_3_22_port, A_s(21)
                           => SHIFT_3_21_port, A_s(20) => SHIFT_3_20_port, 
                           A_s(19) => SHIFT_3_19_port, A_s(18) => 
                           SHIFT_3_18_port, A_s(17) => SHIFT_3_17_port, A_s(16)
                           => SHIFT_3_16_port, A_s(15) => SHIFT_3_15_port, 
                           A_s(14) => SHIFT_3_14_port, A_s(13) => 
                           SHIFT_3_13_port, A_s(12) => SHIFT_3_12_port, A_s(11)
                           => SHIFT_3_11_port, A_s(10) => SHIFT_3_10_port, 
                           A_s(9) => SHIFT_3_9_port, A_s(8) => SHIFT_3_8_port, 
                           A_s(7) => SHIFT_3_7_port, A_s(6) => SHIFT_3_6_port, 
                           A_s(5) => SHIFT_3_5_port, A_s(4) => SHIFT_3_4_port, 
                           A_s(3) => SHIFT_3_3_port, A_s(2) => SHIFT_3_2_port, 
                           A_s(1) => SHIFT_3_1_port, A_s(0) => SHIFT_3_0_port, 
                           A_ns(39) => SHIFT_n_3_37_port, A_ns(38) => 
                           SHIFT_n_3_37_port, A_ns(37) => SHIFT_n_3_37_port, 
                           A_ns(36) => SHIFT_n_3_36_port, A_ns(35) => 
                           SHIFT_n_3_35_port, A_ns(34) => SHIFT_n_3_34_port, 
                           A_ns(33) => SHIFT_n_3_33_port, A_ns(32) => 
                           SHIFT_n_3_32_port, A_ns(31) => SHIFT_n_3_31_port, 
                           A_ns(30) => SHIFT_n_3_30_port, A_ns(29) => 
                           SHIFT_n_3_29_port, A_ns(28) => SHIFT_n_3_28_port, 
                           A_ns(27) => SHIFT_n_3_27_port, A_ns(26) => 
                           SHIFT_n_3_26_port, A_ns(25) => SHIFT_n_3_25_port, 
                           A_ns(24) => SHIFT_n_3_24_port, A_ns(23) => 
                           SHIFT_n_3_23_port, A_ns(22) => SHIFT_n_3_22_port, 
                           A_ns(21) => SHIFT_n_3_21_port, A_ns(20) => 
                           SHIFT_n_3_20_port, A_ns(19) => SHIFT_n_3_19_port, 
                           A_ns(18) => SHIFT_n_3_18_port, A_ns(17) => 
                           SHIFT_n_3_17_port, A_ns(16) => SHIFT_n_3_16_port, 
                           A_ns(15) => SHIFT_n_3_15_port, A_ns(14) => 
                           SHIFT_n_3_14_port, A_ns(13) => SHIFT_n_3_13_port, 
                           A_ns(12) => SHIFT_n_3_12_port, A_ns(11) => 
                           SHIFT_n_3_11_port, A_ns(10) => SHIFT_n_3_10_port, 
                           A_ns(9) => SHIFT_n_3_9_port, A_ns(8) => 
                           SHIFT_n_3_8_port, A_ns(7) => SHIFT_n_3_7_port, 
                           A_ns(6) => SHIFT_n_3_6_port, A_ns(5) => 
                           SHIFT_n_3_5_port, A_ns(4) => SHIFT_n_3_4_port, 
                           A_ns(3) => SHIFT_n_3_3_port, A_ns(2) => 
                           SHIFT_n_3_2_port, A_ns(1) => SHIFT_n_3_1_port, 
                           A_ns(0) => SHIFT_n_3_0_port, B(39) => B(31), B(38) 
                           => B(31), B(37) => B(31), B(36) => B(31), B(35) => 
                           B(31), B(34) => B(31), B(33) => B(31), B(32) => 
                           B(31), B(31) => B(31), B(30) => B(30), B(29) => 
                           B(29), B(28) => B(28), B(27) => B(27), B(26) => 
                           B(26), B(25) => B(25), B(24) => B(24), B(23) => 
                           B(23), B(22) => B(22), B(21) => B(21), B(20) => 
                           B(20), B(19) => B(19), B(18) => B(18), B(17) => 
                           B(17), B(16) => B(16), B(15) => B(15), B(14) => 
                           B(14), B(13) => B(13), B(12) => B(12), B(11) => 
                           B(11), B(10) => B(10), B(9) => B(9), B(8) => B(8), 
                           B(7) => B(7), B(6) => B(6), B(5) => B(5), B(4) => 
                           B(4), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), O(39) => OTMP_3_39_port, O(38) => 
                           OTMP_3_38_port, O(37) => OTMP_3_37_port, O(36) => 
                           OTMP_3_36_port, O(35) => OTMP_3_35_port, O(34) => 
                           OTMP_3_34_port, O(33) => OTMP_3_33_port, O(32) => 
                           OTMP_3_32_port, O(31) => OTMP_3_31_port, O(30) => 
                           OTMP_3_30_port, O(29) => OTMP_3_29_port, O(28) => 
                           OTMP_3_28_port, O(27) => OTMP_3_27_port, O(26) => 
                           OTMP_3_26_port, O(25) => OTMP_3_25_port, O(24) => 
                           OTMP_3_24_port, O(23) => OTMP_3_23_port, O(22) => 
                           OTMP_3_22_port, O(21) => OTMP_3_21_port, O(20) => 
                           OTMP_3_20_port, O(19) => OTMP_3_19_port, O(18) => 
                           OTMP_3_18_port, O(17) => OTMP_3_17_port, O(16) => 
                           OTMP_3_16_port, O(15) => OTMP_3_15_port, O(14) => 
                           OTMP_3_14_port, O(13) => OTMP_3_13_port, O(12) => 
                           OTMP_3_12_port, O(11) => OTMP_3_11_port, O(10) => 
                           OTMP_3_10_port, O(9) => OTMP_3_9_port, O(8) => 
                           OTMP_3_8_port, O(7) => OTMP_3_7_port, O(6) => 
                           OTMP_3_6_port, O(5) => OTMP_3_5_port, O(4) => 
                           OTMP_3_4_port, O(3) => OTMP_3_3_port, O(2) => 
                           OTMP_3_2_port, O(1) => OTMP_3_1_port, O(0) => n_1092
                           , A_so(39) => SHIFT_4_39_port, A_so(38) => 
                           SHIFT_4_38_port, A_so(37) => SHIFT_4_37_port, 
                           A_so(36) => SHIFT_4_36_port, A_so(35) => 
                           SHIFT_4_35_port, A_so(34) => SHIFT_4_34_port, 
                           A_so(33) => SHIFT_4_33_port, A_so(32) => 
                           SHIFT_4_32_port, A_so(31) => SHIFT_4_31_port, 
                           A_so(30) => SHIFT_4_30_port, A_so(29) => 
                           SHIFT_4_29_port, A_so(28) => SHIFT_4_28_port, 
                           A_so(27) => SHIFT_4_27_port, A_so(26) => 
                           SHIFT_4_26_port, A_so(25) => SHIFT_4_25_port, 
                           A_so(24) => SHIFT_4_24_port, A_so(23) => 
                           SHIFT_4_23_port, A_so(22) => SHIFT_4_22_port, 
                           A_so(21) => SHIFT_4_21_port, A_so(20) => 
                           SHIFT_4_20_port, A_so(19) => SHIFT_4_19_port, 
                           A_so(18) => SHIFT_4_18_port, A_so(17) => 
                           SHIFT_4_17_port, A_so(16) => SHIFT_4_16_port, 
                           A_so(15) => SHIFT_4_15_port, A_so(14) => 
                           SHIFT_4_14_port, A_so(13) => SHIFT_4_13_port, 
                           A_so(12) => SHIFT_4_12_port, A_so(11) => 
                           SHIFT_4_11_port, A_so(10) => SHIFT_4_10_port, 
                           A_so(9) => SHIFT_4_9_port, A_so(8) => SHIFT_4_8_port
                           , A_so(7) => SHIFT_4_7_port, A_so(6) => 
                           SHIFT_4_6_port, A_so(5) => SHIFT_4_5_port, A_so(4) 
                           => SHIFT_4_4_port, A_so(3) => SHIFT_4_3_port, 
                           A_so(2) => SHIFT_4_2_port, A_so(1) => n_1093, 
                           A_so(0) => n_1094, A_nso(39) => SHIFT_n_4_39_port, 
                           A_nso(38) => SHIFT_n_4_38_port, A_nso(37) => 
                           SHIFT_n_4_37_port, A_nso(36) => SHIFT_n_4_36_port, 
                           A_nso(35) => SHIFT_n_4_35_port, A_nso(34) => 
                           SHIFT_n_4_34_port, A_nso(33) => SHIFT_n_4_33_port, 
                           A_nso(32) => SHIFT_n_4_32_port, A_nso(31) => 
                           SHIFT_n_4_31_port, A_nso(30) => SHIFT_n_4_30_port, 
                           A_nso(29) => SHIFT_n_4_29_port, A_nso(28) => 
                           SHIFT_n_4_28_port, A_nso(27) => SHIFT_n_4_27_port, 
                           A_nso(26) => SHIFT_n_4_26_port, A_nso(25) => 
                           SHIFT_n_4_25_port, A_nso(24) => SHIFT_n_4_24_port, 
                           A_nso(23) => SHIFT_n_4_23_port, A_nso(22) => 
                           SHIFT_n_4_22_port, A_nso(21) => SHIFT_n_4_21_port, 
                           A_nso(20) => SHIFT_n_4_20_port, A_nso(19) => 
                           SHIFT_n_4_19_port, A_nso(18) => SHIFT_n_4_18_port, 
                           A_nso(17) => SHIFT_n_4_17_port, A_nso(16) => 
                           SHIFT_n_4_16_port, A_nso(15) => SHIFT_n_4_15_port, 
                           A_nso(14) => SHIFT_n_4_14_port, A_nso(13) => 
                           SHIFT_n_4_13_port, A_nso(12) => SHIFT_n_4_12_port, 
                           A_nso(11) => SHIFT_n_4_11_port, A_nso(10) => 
                           SHIFT_n_4_10_port, A_nso(9) => SHIFT_n_4_9_port, 
                           A_nso(8) => SHIFT_n_4_8_port, A_nso(7) => 
                           SHIFT_n_4_7_port, A_nso(6) => SHIFT_n_4_6_port, 
                           A_nso(5) => SHIFT_n_4_5_port, A_nso(4) => 
                           SHIFT_n_4_4_port, A_nso(3) => SHIFT_n_4_3_port, 
                           A_nso(2) => SHIFT_n_4_2_port, A_nso(1) => n_1095, 
                           A_nso(0) => n_1096);
   ENC_4 : BOOTHENC_NBIT42_i8 port map( A_s(41) => SHIFT_4_39_port, A_s(40) => 
                           SHIFT_4_39_port, A_s(39) => SHIFT_4_39_port, A_s(38)
                           => SHIFT_4_38_port, A_s(37) => SHIFT_4_37_port, 
                           A_s(36) => SHIFT_4_36_port, A_s(35) => 
                           SHIFT_4_35_port, A_s(34) => SHIFT_4_34_port, A_s(33)
                           => SHIFT_4_33_port, A_s(32) => SHIFT_4_32_port, 
                           A_s(31) => SHIFT_4_31_port, A_s(30) => 
                           SHIFT_4_30_port, A_s(29) => SHIFT_4_29_port, A_s(28)
                           => SHIFT_4_28_port, A_s(27) => SHIFT_4_27_port, 
                           A_s(26) => SHIFT_4_26_port, A_s(25) => 
                           SHIFT_4_25_port, A_s(24) => SHIFT_4_24_port, A_s(23)
                           => SHIFT_4_23_port, A_s(22) => SHIFT_4_22_port, 
                           A_s(21) => SHIFT_4_21_port, A_s(20) => 
                           SHIFT_4_20_port, A_s(19) => SHIFT_4_19_port, A_s(18)
                           => SHIFT_4_18_port, A_s(17) => SHIFT_4_17_port, 
                           A_s(16) => SHIFT_4_16_port, A_s(15) => 
                           SHIFT_4_15_port, A_s(14) => SHIFT_4_14_port, A_s(13)
                           => SHIFT_4_13_port, A_s(12) => SHIFT_4_12_port, 
                           A_s(11) => SHIFT_4_11_port, A_s(10) => 
                           SHIFT_4_10_port, A_s(9) => SHIFT_4_9_port, A_s(8) =>
                           SHIFT_4_8_port, A_s(7) => SHIFT_4_7_port, A_s(6) => 
                           SHIFT_4_6_port, A_s(5) => SHIFT_4_5_port, A_s(4) => 
                           SHIFT_4_4_port, A_s(3) => SHIFT_4_3_port, A_s(2) => 
                           SHIFT_4_2_port, A_s(1) => SHIFT_4_1_port, A_s(0) => 
                           SHIFT_4_0_port, A_ns(41) => SHIFT_n_4_39_port, 
                           A_ns(40) => SHIFT_n_4_39_port, A_ns(39) => 
                           SHIFT_n_4_39_port, A_ns(38) => SHIFT_n_4_38_port, 
                           A_ns(37) => SHIFT_n_4_37_port, A_ns(36) => 
                           SHIFT_n_4_36_port, A_ns(35) => SHIFT_n_4_35_port, 
                           A_ns(34) => SHIFT_n_4_34_port, A_ns(33) => 
                           SHIFT_n_4_33_port, A_ns(32) => SHIFT_n_4_32_port, 
                           A_ns(31) => SHIFT_n_4_31_port, A_ns(30) => 
                           SHIFT_n_4_30_port, A_ns(29) => SHIFT_n_4_29_port, 
                           A_ns(28) => SHIFT_n_4_28_port, A_ns(27) => 
                           SHIFT_n_4_27_port, A_ns(26) => SHIFT_n_4_26_port, 
                           A_ns(25) => SHIFT_n_4_25_port, A_ns(24) => 
                           SHIFT_n_4_24_port, A_ns(23) => SHIFT_n_4_23_port, 
                           A_ns(22) => SHIFT_n_4_22_port, A_ns(21) => 
                           SHIFT_n_4_21_port, A_ns(20) => SHIFT_n_4_20_port, 
                           A_ns(19) => SHIFT_n_4_19_port, A_ns(18) => 
                           SHIFT_n_4_18_port, A_ns(17) => SHIFT_n_4_17_port, 
                           A_ns(16) => SHIFT_n_4_16_port, A_ns(15) => 
                           SHIFT_n_4_15_port, A_ns(14) => SHIFT_n_4_14_port, 
                           A_ns(13) => SHIFT_n_4_13_port, A_ns(12) => 
                           SHIFT_n_4_12_port, A_ns(11) => SHIFT_n_4_11_port, 
                           A_ns(10) => SHIFT_n_4_10_port, A_ns(9) => 
                           SHIFT_n_4_9_port, A_ns(8) => SHIFT_n_4_8_port, 
                           A_ns(7) => SHIFT_n_4_7_port, A_ns(6) => 
                           SHIFT_n_4_6_port, A_ns(5) => SHIFT_n_4_5_port, 
                           A_ns(4) => SHIFT_n_4_4_port, A_ns(3) => 
                           SHIFT_n_4_3_port, A_ns(2) => SHIFT_n_4_2_port, 
                           A_ns(1) => SHIFT_n_4_1_port, A_ns(0) => 
                           SHIFT_n_4_0_port, B(41) => B(31), B(40) => B(31), 
                           B(39) => B(31), B(38) => B(31), B(37) => B(31), 
                           B(36) => B(31), B(35) => B(31), B(34) => B(31), 
                           B(33) => B(31), B(32) => B(31), B(31) => B(31), 
                           B(30) => B(30), B(29) => B(29), B(28) => B(28), 
                           B(27) => B(27), B(26) => B(26), B(25) => B(25), 
                           B(24) => B(24), B(23) => B(23), B(22) => B(22), 
                           B(21) => B(21), B(20) => B(20), B(19) => B(19), 
                           B(18) => B(18), B(17) => B(17), B(16) => B(16), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => B(0), O(41) => 
                           OTMP_4_41_port, O(40) => OTMP_4_40_port, O(39) => 
                           OTMP_4_39_port, O(38) => OTMP_4_38_port, O(37) => 
                           OTMP_4_37_port, O(36) => OTMP_4_36_port, O(35) => 
                           OTMP_4_35_port, O(34) => OTMP_4_34_port, O(33) => 
                           OTMP_4_33_port, O(32) => OTMP_4_32_port, O(31) => 
                           OTMP_4_31_port, O(30) => OTMP_4_30_port, O(29) => 
                           OTMP_4_29_port, O(28) => OTMP_4_28_port, O(27) => 
                           OTMP_4_27_port, O(26) => OTMP_4_26_port, O(25) => 
                           OTMP_4_25_port, O(24) => OTMP_4_24_port, O(23) => 
                           OTMP_4_23_port, O(22) => OTMP_4_22_port, O(21) => 
                           OTMP_4_21_port, O(20) => OTMP_4_20_port, O(19) => 
                           OTMP_4_19_port, O(18) => OTMP_4_18_port, O(17) => 
                           OTMP_4_17_port, O(16) => OTMP_4_16_port, O(15) => 
                           OTMP_4_15_port, O(14) => OTMP_4_14_port, O(13) => 
                           OTMP_4_13_port, O(12) => OTMP_4_12_port, O(11) => 
                           OTMP_4_11_port, O(10) => OTMP_4_10_port, O(9) => 
                           OTMP_4_9_port, O(8) => OTMP_4_8_port, O(7) => 
                           OTMP_4_7_port, O(6) => OTMP_4_6_port, O(5) => 
                           OTMP_4_5_port, O(4) => OTMP_4_4_port, O(3) => 
                           OTMP_4_3_port, O(2) => OTMP_4_2_port, O(1) => 
                           OTMP_4_1_port, O(0) => n_1097, A_so(41) => 
                           SHIFT_5_41_port, A_so(40) => SHIFT_5_40_port, 
                           A_so(39) => SHIFT_5_39_port, A_so(38) => 
                           SHIFT_5_38_port, A_so(37) => SHIFT_5_37_port, 
                           A_so(36) => SHIFT_5_36_port, A_so(35) => 
                           SHIFT_5_35_port, A_so(34) => SHIFT_5_34_port, 
                           A_so(33) => SHIFT_5_33_port, A_so(32) => 
                           SHIFT_5_32_port, A_so(31) => SHIFT_5_31_port, 
                           A_so(30) => SHIFT_5_30_port, A_so(29) => 
                           SHIFT_5_29_port, A_so(28) => SHIFT_5_28_port, 
                           A_so(27) => SHIFT_5_27_port, A_so(26) => 
                           SHIFT_5_26_port, A_so(25) => SHIFT_5_25_port, 
                           A_so(24) => SHIFT_5_24_port, A_so(23) => 
                           SHIFT_5_23_port, A_so(22) => SHIFT_5_22_port, 
                           A_so(21) => SHIFT_5_21_port, A_so(20) => 
                           SHIFT_5_20_port, A_so(19) => SHIFT_5_19_port, 
                           A_so(18) => SHIFT_5_18_port, A_so(17) => 
                           SHIFT_5_17_port, A_so(16) => SHIFT_5_16_port, 
                           A_so(15) => SHIFT_5_15_port, A_so(14) => 
                           SHIFT_5_14_port, A_so(13) => SHIFT_5_13_port, 
                           A_so(12) => SHIFT_5_12_port, A_so(11) => 
                           SHIFT_5_11_port, A_so(10) => SHIFT_5_10_port, 
                           A_so(9) => SHIFT_5_9_port, A_so(8) => SHIFT_5_8_port
                           , A_so(7) => SHIFT_5_7_port, A_so(6) => 
                           SHIFT_5_6_port, A_so(5) => SHIFT_5_5_port, A_so(4) 
                           => SHIFT_5_4_port, A_so(3) => SHIFT_5_3_port, 
                           A_so(2) => SHIFT_5_2_port, A_so(1) => n_1098, 
                           A_so(0) => n_1099, A_nso(41) => SHIFT_n_5_41_port, 
                           A_nso(40) => SHIFT_n_5_40_port, A_nso(39) => 
                           SHIFT_n_5_39_port, A_nso(38) => SHIFT_n_5_38_port, 
                           A_nso(37) => SHIFT_n_5_37_port, A_nso(36) => 
                           SHIFT_n_5_36_port, A_nso(35) => SHIFT_n_5_35_port, 
                           A_nso(34) => SHIFT_n_5_34_port, A_nso(33) => 
                           SHIFT_n_5_33_port, A_nso(32) => SHIFT_n_5_32_port, 
                           A_nso(31) => SHIFT_n_5_31_port, A_nso(30) => 
                           SHIFT_n_5_30_port, A_nso(29) => SHIFT_n_5_29_port, 
                           A_nso(28) => SHIFT_n_5_28_port, A_nso(27) => 
                           SHIFT_n_5_27_port, A_nso(26) => SHIFT_n_5_26_port, 
                           A_nso(25) => SHIFT_n_5_25_port, A_nso(24) => 
                           SHIFT_n_5_24_port, A_nso(23) => SHIFT_n_5_23_port, 
                           A_nso(22) => SHIFT_n_5_22_port, A_nso(21) => 
                           SHIFT_n_5_21_port, A_nso(20) => SHIFT_n_5_20_port, 
                           A_nso(19) => SHIFT_n_5_19_port, A_nso(18) => 
                           SHIFT_n_5_18_port, A_nso(17) => SHIFT_n_5_17_port, 
                           A_nso(16) => SHIFT_n_5_16_port, A_nso(15) => 
                           SHIFT_n_5_15_port, A_nso(14) => SHIFT_n_5_14_port, 
                           A_nso(13) => SHIFT_n_5_13_port, A_nso(12) => 
                           SHIFT_n_5_12_port, A_nso(11) => SHIFT_n_5_11_port, 
                           A_nso(10) => SHIFT_n_5_10_port, A_nso(9) => 
                           SHIFT_n_5_9_port, A_nso(8) => SHIFT_n_5_8_port, 
                           A_nso(7) => SHIFT_n_5_7_port, A_nso(6) => 
                           SHIFT_n_5_6_port, A_nso(5) => SHIFT_n_5_5_port, 
                           A_nso(4) => SHIFT_n_5_4_port, A_nso(3) => 
                           SHIFT_n_5_3_port, A_nso(2) => SHIFT_n_5_2_port, 
                           A_nso(1) => n_1100, A_nso(0) => n_1101);
   ENC_5 : BOOTHENC_NBIT44_i10 port map( A_s(43) => SHIFT_5_41_port, A_s(42) =>
                           SHIFT_5_41_port, A_s(41) => SHIFT_5_41_port, A_s(40)
                           => SHIFT_5_40_port, A_s(39) => SHIFT_5_39_port, 
                           A_s(38) => SHIFT_5_38_port, A_s(37) => 
                           SHIFT_5_37_port, A_s(36) => SHIFT_5_36_port, A_s(35)
                           => SHIFT_5_35_port, A_s(34) => SHIFT_5_34_port, 
                           A_s(33) => SHIFT_5_33_port, A_s(32) => 
                           SHIFT_5_32_port, A_s(31) => SHIFT_5_31_port, A_s(30)
                           => SHIFT_5_30_port, A_s(29) => SHIFT_5_29_port, 
                           A_s(28) => SHIFT_5_28_port, A_s(27) => 
                           SHIFT_5_27_port, A_s(26) => SHIFT_5_26_port, A_s(25)
                           => SHIFT_5_25_port, A_s(24) => SHIFT_5_24_port, 
                           A_s(23) => SHIFT_5_23_port, A_s(22) => 
                           SHIFT_5_22_port, A_s(21) => SHIFT_5_21_port, A_s(20)
                           => SHIFT_5_20_port, A_s(19) => SHIFT_5_19_port, 
                           A_s(18) => SHIFT_5_18_port, A_s(17) => 
                           SHIFT_5_17_port, A_s(16) => SHIFT_5_16_port, A_s(15)
                           => SHIFT_5_15_port, A_s(14) => SHIFT_5_14_port, 
                           A_s(13) => SHIFT_5_13_port, A_s(12) => 
                           SHIFT_5_12_port, A_s(11) => SHIFT_5_11_port, A_s(10)
                           => SHIFT_5_10_port, A_s(9) => SHIFT_5_9_port, A_s(8)
                           => SHIFT_5_8_port, A_s(7) => SHIFT_5_7_port, A_s(6) 
                           => SHIFT_5_6_port, A_s(5) => SHIFT_5_5_port, A_s(4) 
                           => SHIFT_5_4_port, A_s(3) => SHIFT_5_3_port, A_s(2) 
                           => SHIFT_5_2_port, A_s(1) => SHIFT_5_1_port, A_s(0) 
                           => SHIFT_5_0_port, A_ns(43) => SHIFT_n_5_41_port, 
                           A_ns(42) => SHIFT_n_5_41_port, A_ns(41) => 
                           SHIFT_n_5_41_port, A_ns(40) => SHIFT_n_5_40_port, 
                           A_ns(39) => SHIFT_n_5_39_port, A_ns(38) => 
                           SHIFT_n_5_38_port, A_ns(37) => SHIFT_n_5_37_port, 
                           A_ns(36) => SHIFT_n_5_36_port, A_ns(35) => 
                           SHIFT_n_5_35_port, A_ns(34) => SHIFT_n_5_34_port, 
                           A_ns(33) => SHIFT_n_5_33_port, A_ns(32) => 
                           SHIFT_n_5_32_port, A_ns(31) => SHIFT_n_5_31_port, 
                           A_ns(30) => SHIFT_n_5_30_port, A_ns(29) => 
                           SHIFT_n_5_29_port, A_ns(28) => SHIFT_n_5_28_port, 
                           A_ns(27) => SHIFT_n_5_27_port, A_ns(26) => 
                           SHIFT_n_5_26_port, A_ns(25) => SHIFT_n_5_25_port, 
                           A_ns(24) => SHIFT_n_5_24_port, A_ns(23) => 
                           SHIFT_n_5_23_port, A_ns(22) => SHIFT_n_5_22_port, 
                           A_ns(21) => SHIFT_n_5_21_port, A_ns(20) => 
                           SHIFT_n_5_20_port, A_ns(19) => SHIFT_n_5_19_port, 
                           A_ns(18) => SHIFT_n_5_18_port, A_ns(17) => 
                           SHIFT_n_5_17_port, A_ns(16) => SHIFT_n_5_16_port, 
                           A_ns(15) => SHIFT_n_5_15_port, A_ns(14) => 
                           SHIFT_n_5_14_port, A_ns(13) => SHIFT_n_5_13_port, 
                           A_ns(12) => SHIFT_n_5_12_port, A_ns(11) => 
                           SHIFT_n_5_11_port, A_ns(10) => SHIFT_n_5_10_port, 
                           A_ns(9) => SHIFT_n_5_9_port, A_ns(8) => 
                           SHIFT_n_5_8_port, A_ns(7) => SHIFT_n_5_7_port, 
                           A_ns(6) => SHIFT_n_5_6_port, A_ns(5) => 
                           SHIFT_n_5_5_port, A_ns(4) => SHIFT_n_5_4_port, 
                           A_ns(3) => SHIFT_n_5_3_port, A_ns(2) => 
                           SHIFT_n_5_2_port, A_ns(1) => SHIFT_n_5_1_port, 
                           A_ns(0) => SHIFT_n_5_0_port, B(43) => B(31), B(42) 
                           => B(31), B(41) => B(31), B(40) => B(31), B(39) => 
                           B(31), B(38) => B(31), B(37) => B(31), B(36) => 
                           B(31), B(35) => B(31), B(34) => B(31), B(33) => 
                           B(31), B(32) => B(31), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), O(43) => OTMP_5_43_port, 
                           O(42) => OTMP_5_42_port, O(41) => OTMP_5_41_port, 
                           O(40) => OTMP_5_40_port, O(39) => OTMP_5_39_port, 
                           O(38) => OTMP_5_38_port, O(37) => OTMP_5_37_port, 
                           O(36) => OTMP_5_36_port, O(35) => OTMP_5_35_port, 
                           O(34) => OTMP_5_34_port, O(33) => OTMP_5_33_port, 
                           O(32) => OTMP_5_32_port, O(31) => OTMP_5_31_port, 
                           O(30) => OTMP_5_30_port, O(29) => OTMP_5_29_port, 
                           O(28) => OTMP_5_28_port, O(27) => OTMP_5_27_port, 
                           O(26) => OTMP_5_26_port, O(25) => OTMP_5_25_port, 
                           O(24) => OTMP_5_24_port, O(23) => OTMP_5_23_port, 
                           O(22) => OTMP_5_22_port, O(21) => OTMP_5_21_port, 
                           O(20) => OTMP_5_20_port, O(19) => OTMP_5_19_port, 
                           O(18) => OTMP_5_18_port, O(17) => OTMP_5_17_port, 
                           O(16) => OTMP_5_16_port, O(15) => OTMP_5_15_port, 
                           O(14) => OTMP_5_14_port, O(13) => OTMP_5_13_port, 
                           O(12) => OTMP_5_12_port, O(11) => OTMP_5_11_port, 
                           O(10) => OTMP_5_10_port, O(9) => OTMP_5_9_port, O(8)
                           => OTMP_5_8_port, O(7) => OTMP_5_7_port, O(6) => 
                           OTMP_5_6_port, O(5) => OTMP_5_5_port, O(4) => 
                           OTMP_5_4_port, O(3) => OTMP_5_3_port, O(2) => 
                           OTMP_5_2_port, O(1) => OTMP_5_1_port, O(0) => n_1102
                           , A_so(43) => SHIFT_6_43_port, A_so(42) => 
                           SHIFT_6_42_port, A_so(41) => SHIFT_6_41_port, 
                           A_so(40) => SHIFT_6_40_port, A_so(39) => 
                           SHIFT_6_39_port, A_so(38) => SHIFT_6_38_port, 
                           A_so(37) => SHIFT_6_37_port, A_so(36) => 
                           SHIFT_6_36_port, A_so(35) => SHIFT_6_35_port, 
                           A_so(34) => SHIFT_6_34_port, A_so(33) => 
                           SHIFT_6_33_port, A_so(32) => SHIFT_6_32_port, 
                           A_so(31) => SHIFT_6_31_port, A_so(30) => 
                           SHIFT_6_30_port, A_so(29) => SHIFT_6_29_port, 
                           A_so(28) => SHIFT_6_28_port, A_so(27) => 
                           SHIFT_6_27_port, A_so(26) => SHIFT_6_26_port, 
                           A_so(25) => SHIFT_6_25_port, A_so(24) => 
                           SHIFT_6_24_port, A_so(23) => SHIFT_6_23_port, 
                           A_so(22) => SHIFT_6_22_port, A_so(21) => 
                           SHIFT_6_21_port, A_so(20) => SHIFT_6_20_port, 
                           A_so(19) => SHIFT_6_19_port, A_so(18) => 
                           SHIFT_6_18_port, A_so(17) => SHIFT_6_17_port, 
                           A_so(16) => SHIFT_6_16_port, A_so(15) => 
                           SHIFT_6_15_port, A_so(14) => SHIFT_6_14_port, 
                           A_so(13) => SHIFT_6_13_port, A_so(12) => 
                           SHIFT_6_12_port, A_so(11) => SHIFT_6_11_port, 
                           A_so(10) => SHIFT_6_10_port, A_so(9) => 
                           SHIFT_6_9_port, A_so(8) => SHIFT_6_8_port, A_so(7) 
                           => SHIFT_6_7_port, A_so(6) => SHIFT_6_6_port, 
                           A_so(5) => SHIFT_6_5_port, A_so(4) => SHIFT_6_4_port
                           , A_so(3) => SHIFT_6_3_port, A_so(2) => 
                           SHIFT_6_2_port, A_so(1) => n_1103, A_so(0) => n_1104
                           , A_nso(43) => SHIFT_n_6_43_port, A_nso(42) => 
                           SHIFT_n_6_42_port, A_nso(41) => SHIFT_n_6_41_port, 
                           A_nso(40) => SHIFT_n_6_40_port, A_nso(39) => 
                           SHIFT_n_6_39_port, A_nso(38) => SHIFT_n_6_38_port, 
                           A_nso(37) => SHIFT_n_6_37_port, A_nso(36) => 
                           SHIFT_n_6_36_port, A_nso(35) => SHIFT_n_6_35_port, 
                           A_nso(34) => SHIFT_n_6_34_port, A_nso(33) => 
                           SHIFT_n_6_33_port, A_nso(32) => SHIFT_n_6_32_port, 
                           A_nso(31) => SHIFT_n_6_31_port, A_nso(30) => 
                           SHIFT_n_6_30_port, A_nso(29) => SHIFT_n_6_29_port, 
                           A_nso(28) => SHIFT_n_6_28_port, A_nso(27) => 
                           SHIFT_n_6_27_port, A_nso(26) => SHIFT_n_6_26_port, 
                           A_nso(25) => SHIFT_n_6_25_port, A_nso(24) => 
                           SHIFT_n_6_24_port, A_nso(23) => SHIFT_n_6_23_port, 
                           A_nso(22) => SHIFT_n_6_22_port, A_nso(21) => 
                           SHIFT_n_6_21_port, A_nso(20) => SHIFT_n_6_20_port, 
                           A_nso(19) => SHIFT_n_6_19_port, A_nso(18) => 
                           SHIFT_n_6_18_port, A_nso(17) => SHIFT_n_6_17_port, 
                           A_nso(16) => SHIFT_n_6_16_port, A_nso(15) => 
                           SHIFT_n_6_15_port, A_nso(14) => SHIFT_n_6_14_port, 
                           A_nso(13) => SHIFT_n_6_13_port, A_nso(12) => 
                           SHIFT_n_6_12_port, A_nso(11) => SHIFT_n_6_11_port, 
                           A_nso(10) => SHIFT_n_6_10_port, A_nso(9) => 
                           SHIFT_n_6_9_port, A_nso(8) => SHIFT_n_6_8_port, 
                           A_nso(7) => SHIFT_n_6_7_port, A_nso(6) => 
                           SHIFT_n_6_6_port, A_nso(5) => SHIFT_n_6_5_port, 
                           A_nso(4) => SHIFT_n_6_4_port, A_nso(3) => 
                           SHIFT_n_6_3_port, A_nso(2) => SHIFT_n_6_2_port, 
                           A_nso(1) => n_1105, A_nso(0) => n_1106);
   ENC_6 : BOOTHENC_NBIT46_i12 port map( A_s(45) => SHIFT_6_43_port, A_s(44) =>
                           SHIFT_6_43_port, A_s(43) => SHIFT_6_43_port, A_s(42)
                           => SHIFT_6_42_port, A_s(41) => SHIFT_6_41_port, 
                           A_s(40) => SHIFT_6_40_port, A_s(39) => 
                           SHIFT_6_39_port, A_s(38) => SHIFT_6_38_port, A_s(37)
                           => SHIFT_6_37_port, A_s(36) => SHIFT_6_36_port, 
                           A_s(35) => SHIFT_6_35_port, A_s(34) => 
                           SHIFT_6_34_port, A_s(33) => SHIFT_6_33_port, A_s(32)
                           => SHIFT_6_32_port, A_s(31) => SHIFT_6_31_port, 
                           A_s(30) => SHIFT_6_30_port, A_s(29) => 
                           SHIFT_6_29_port, A_s(28) => SHIFT_6_28_port, A_s(27)
                           => SHIFT_6_27_port, A_s(26) => SHIFT_6_26_port, 
                           A_s(25) => SHIFT_6_25_port, A_s(24) => 
                           SHIFT_6_24_port, A_s(23) => SHIFT_6_23_port, A_s(22)
                           => SHIFT_6_22_port, A_s(21) => SHIFT_6_21_port, 
                           A_s(20) => SHIFT_6_20_port, A_s(19) => 
                           SHIFT_6_19_port, A_s(18) => SHIFT_6_18_port, A_s(17)
                           => SHIFT_6_17_port, A_s(16) => SHIFT_6_16_port, 
                           A_s(15) => SHIFT_6_15_port, A_s(14) => 
                           SHIFT_6_14_port, A_s(13) => SHIFT_6_13_port, A_s(12)
                           => SHIFT_6_12_port, A_s(11) => SHIFT_6_11_port, 
                           A_s(10) => SHIFT_6_10_port, A_s(9) => SHIFT_6_9_port
                           , A_s(8) => SHIFT_6_8_port, A_s(7) => SHIFT_6_7_port
                           , A_s(6) => SHIFT_6_6_port, A_s(5) => SHIFT_6_5_port
                           , A_s(4) => SHIFT_6_4_port, A_s(3) => SHIFT_6_3_port
                           , A_s(2) => SHIFT_6_2_port, A_s(1) => SHIFT_6_1_port
                           , A_s(0) => SHIFT_6_0_port, A_ns(45) => 
                           SHIFT_n_6_43_port, A_ns(44) => SHIFT_n_6_43_port, 
                           A_ns(43) => SHIFT_n_6_43_port, A_ns(42) => 
                           SHIFT_n_6_42_port, A_ns(41) => SHIFT_n_6_41_port, 
                           A_ns(40) => SHIFT_n_6_40_port, A_ns(39) => 
                           SHIFT_n_6_39_port, A_ns(38) => SHIFT_n_6_38_port, 
                           A_ns(37) => SHIFT_n_6_37_port, A_ns(36) => 
                           SHIFT_n_6_36_port, A_ns(35) => SHIFT_n_6_35_port, 
                           A_ns(34) => SHIFT_n_6_34_port, A_ns(33) => 
                           SHIFT_n_6_33_port, A_ns(32) => SHIFT_n_6_32_port, 
                           A_ns(31) => SHIFT_n_6_31_port, A_ns(30) => 
                           SHIFT_n_6_30_port, A_ns(29) => SHIFT_n_6_29_port, 
                           A_ns(28) => SHIFT_n_6_28_port, A_ns(27) => 
                           SHIFT_n_6_27_port, A_ns(26) => SHIFT_n_6_26_port, 
                           A_ns(25) => SHIFT_n_6_25_port, A_ns(24) => 
                           SHIFT_n_6_24_port, A_ns(23) => SHIFT_n_6_23_port, 
                           A_ns(22) => SHIFT_n_6_22_port, A_ns(21) => 
                           SHIFT_n_6_21_port, A_ns(20) => SHIFT_n_6_20_port, 
                           A_ns(19) => SHIFT_n_6_19_port, A_ns(18) => 
                           SHIFT_n_6_18_port, A_ns(17) => SHIFT_n_6_17_port, 
                           A_ns(16) => SHIFT_n_6_16_port, A_ns(15) => 
                           SHIFT_n_6_15_port, A_ns(14) => SHIFT_n_6_14_port, 
                           A_ns(13) => SHIFT_n_6_13_port, A_ns(12) => 
                           SHIFT_n_6_12_port, A_ns(11) => SHIFT_n_6_11_port, 
                           A_ns(10) => SHIFT_n_6_10_port, A_ns(9) => 
                           SHIFT_n_6_9_port, A_ns(8) => SHIFT_n_6_8_port, 
                           A_ns(7) => SHIFT_n_6_7_port, A_ns(6) => 
                           SHIFT_n_6_6_port, A_ns(5) => SHIFT_n_6_5_port, 
                           A_ns(4) => SHIFT_n_6_4_port, A_ns(3) => 
                           SHIFT_n_6_3_port, A_ns(2) => SHIFT_n_6_2_port, 
                           A_ns(1) => SHIFT_n_6_1_port, A_ns(0) => 
                           SHIFT_n_6_0_port, B(45) => B(31), B(44) => B(31), 
                           B(43) => B(31), B(42) => B(31), B(41) => B(31), 
                           B(40) => B(31), B(39) => B(31), B(38) => B(31), 
                           B(37) => B(31), B(36) => B(31), B(35) => B(31), 
                           B(34) => B(31), B(33) => B(31), B(32) => B(31), 
                           B(31) => B(31), B(30) => B(30), B(29) => B(29), 
                           B(28) => B(28), B(27) => B(27), B(26) => B(26), 
                           B(25) => B(25), B(24) => B(24), B(23) => B(23), 
                           B(22) => B(22), B(21) => B(21), B(20) => B(20), 
                           B(19) => B(19), B(18) => B(18), B(17) => B(17), 
                           B(16) => B(16), B(15) => B(15), B(14) => B(14), 
                           B(13) => B(13), B(12) => B(12), B(11) => B(11), 
                           B(10) => B(10), B(9) => B(9), B(8) => B(8), B(7) => 
                           B(7), B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3)
                           => B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), 
                           O(45) => OTMP_6_45_port, O(44) => OTMP_6_44_port, 
                           O(43) => OTMP_6_43_port, O(42) => OTMP_6_42_port, 
                           O(41) => OTMP_6_41_port, O(40) => OTMP_6_40_port, 
                           O(39) => OTMP_6_39_port, O(38) => OTMP_6_38_port, 
                           O(37) => OTMP_6_37_port, O(36) => OTMP_6_36_port, 
                           O(35) => OTMP_6_35_port, O(34) => OTMP_6_34_port, 
                           O(33) => OTMP_6_33_port, O(32) => OTMP_6_32_port, 
                           O(31) => OTMP_6_31_port, O(30) => OTMP_6_30_port, 
                           O(29) => OTMP_6_29_port, O(28) => OTMP_6_28_port, 
                           O(27) => OTMP_6_27_port, O(26) => OTMP_6_26_port, 
                           O(25) => OTMP_6_25_port, O(24) => OTMP_6_24_port, 
                           O(23) => OTMP_6_23_port, O(22) => OTMP_6_22_port, 
                           O(21) => OTMP_6_21_port, O(20) => OTMP_6_20_port, 
                           O(19) => OTMP_6_19_port, O(18) => OTMP_6_18_port, 
                           O(17) => OTMP_6_17_port, O(16) => OTMP_6_16_port, 
                           O(15) => OTMP_6_15_port, O(14) => OTMP_6_14_port, 
                           O(13) => OTMP_6_13_port, O(12) => OTMP_6_12_port, 
                           O(11) => OTMP_6_11_port, O(10) => OTMP_6_10_port, 
                           O(9) => OTMP_6_9_port, O(8) => OTMP_6_8_port, O(7) 
                           => OTMP_6_7_port, O(6) => OTMP_6_6_port, O(5) => 
                           OTMP_6_5_port, O(4) => OTMP_6_4_port, O(3) => 
                           OTMP_6_3_port, O(2) => OTMP_6_2_port, O(1) => 
                           OTMP_6_1_port, O(0) => n_1107, A_so(45) => 
                           SHIFT_7_45_port, A_so(44) => SHIFT_7_44_port, 
                           A_so(43) => SHIFT_7_43_port, A_so(42) => 
                           SHIFT_7_42_port, A_so(41) => SHIFT_7_41_port, 
                           A_so(40) => SHIFT_7_40_port, A_so(39) => 
                           SHIFT_7_39_port, A_so(38) => SHIFT_7_38_port, 
                           A_so(37) => SHIFT_7_37_port, A_so(36) => 
                           SHIFT_7_36_port, A_so(35) => SHIFT_7_35_port, 
                           A_so(34) => SHIFT_7_34_port, A_so(33) => 
                           SHIFT_7_33_port, A_so(32) => SHIFT_7_32_port, 
                           A_so(31) => SHIFT_7_31_port, A_so(30) => 
                           SHIFT_7_30_port, A_so(29) => SHIFT_7_29_port, 
                           A_so(28) => SHIFT_7_28_port, A_so(27) => 
                           SHIFT_7_27_port, A_so(26) => SHIFT_7_26_port, 
                           A_so(25) => SHIFT_7_25_port, A_so(24) => 
                           SHIFT_7_24_port, A_so(23) => SHIFT_7_23_port, 
                           A_so(22) => SHIFT_7_22_port, A_so(21) => 
                           SHIFT_7_21_port, A_so(20) => SHIFT_7_20_port, 
                           A_so(19) => SHIFT_7_19_port, A_so(18) => 
                           SHIFT_7_18_port, A_so(17) => SHIFT_7_17_port, 
                           A_so(16) => SHIFT_7_16_port, A_so(15) => 
                           SHIFT_7_15_port, A_so(14) => SHIFT_7_14_port, 
                           A_so(13) => SHIFT_7_13_port, A_so(12) => 
                           SHIFT_7_12_port, A_so(11) => SHIFT_7_11_port, 
                           A_so(10) => SHIFT_7_10_port, A_so(9) => 
                           SHIFT_7_9_port, A_so(8) => SHIFT_7_8_port, A_so(7) 
                           => SHIFT_7_7_port, A_so(6) => SHIFT_7_6_port, 
                           A_so(5) => SHIFT_7_5_port, A_so(4) => SHIFT_7_4_port
                           , A_so(3) => SHIFT_7_3_port, A_so(2) => 
                           SHIFT_7_2_port, A_so(1) => n_1108, A_so(0) => n_1109
                           , A_nso(45) => SHIFT_n_7_45_port, A_nso(44) => 
                           SHIFT_n_7_44_port, A_nso(43) => SHIFT_n_7_43_port, 
                           A_nso(42) => SHIFT_n_7_42_port, A_nso(41) => 
                           SHIFT_n_7_41_port, A_nso(40) => SHIFT_n_7_40_port, 
                           A_nso(39) => SHIFT_n_7_39_port, A_nso(38) => 
                           SHIFT_n_7_38_port, A_nso(37) => SHIFT_n_7_37_port, 
                           A_nso(36) => SHIFT_n_7_36_port, A_nso(35) => 
                           SHIFT_n_7_35_port, A_nso(34) => SHIFT_n_7_34_port, 
                           A_nso(33) => SHIFT_n_7_33_port, A_nso(32) => 
                           SHIFT_n_7_32_port, A_nso(31) => SHIFT_n_7_31_port, 
                           A_nso(30) => SHIFT_n_7_30_port, A_nso(29) => 
                           SHIFT_n_7_29_port, A_nso(28) => SHIFT_n_7_28_port, 
                           A_nso(27) => SHIFT_n_7_27_port, A_nso(26) => 
                           SHIFT_n_7_26_port, A_nso(25) => SHIFT_n_7_25_port, 
                           A_nso(24) => SHIFT_n_7_24_port, A_nso(23) => 
                           SHIFT_n_7_23_port, A_nso(22) => SHIFT_n_7_22_port, 
                           A_nso(21) => SHIFT_n_7_21_port, A_nso(20) => 
                           SHIFT_n_7_20_port, A_nso(19) => SHIFT_n_7_19_port, 
                           A_nso(18) => SHIFT_n_7_18_port, A_nso(17) => 
                           SHIFT_n_7_17_port, A_nso(16) => SHIFT_n_7_16_port, 
                           A_nso(15) => SHIFT_n_7_15_port, A_nso(14) => 
                           SHIFT_n_7_14_port, A_nso(13) => SHIFT_n_7_13_port, 
                           A_nso(12) => SHIFT_n_7_12_port, A_nso(11) => 
                           SHIFT_n_7_11_port, A_nso(10) => SHIFT_n_7_10_port, 
                           A_nso(9) => SHIFT_n_7_9_port, A_nso(8) => 
                           SHIFT_n_7_8_port, A_nso(7) => SHIFT_n_7_7_port, 
                           A_nso(6) => SHIFT_n_7_6_port, A_nso(5) => 
                           SHIFT_n_7_5_port, A_nso(4) => SHIFT_n_7_4_port, 
                           A_nso(3) => SHIFT_n_7_3_port, A_nso(2) => 
                           SHIFT_n_7_2_port, A_nso(1) => n_1110, A_nso(0) => 
                           n_1111);
   ENC_7 : BOOTHENC_NBIT48_i14 port map( A_s(47) => SHIFT_7_45_port, A_s(46) =>
                           SHIFT_7_45_port, A_s(45) => SHIFT_7_45_port, A_s(44)
                           => SHIFT_7_44_port, A_s(43) => SHIFT_7_43_port, 
                           A_s(42) => SHIFT_7_42_port, A_s(41) => 
                           SHIFT_7_41_port, A_s(40) => SHIFT_7_40_port, A_s(39)
                           => SHIFT_7_39_port, A_s(38) => SHIFT_7_38_port, 
                           A_s(37) => SHIFT_7_37_port, A_s(36) => 
                           SHIFT_7_36_port, A_s(35) => SHIFT_7_35_port, A_s(34)
                           => SHIFT_7_34_port, A_s(33) => SHIFT_7_33_port, 
                           A_s(32) => SHIFT_7_32_port, A_s(31) => 
                           SHIFT_7_31_port, A_s(30) => SHIFT_7_30_port, A_s(29)
                           => SHIFT_7_29_port, A_s(28) => SHIFT_7_28_port, 
                           A_s(27) => SHIFT_7_27_port, A_s(26) => 
                           SHIFT_7_26_port, A_s(25) => SHIFT_7_25_port, A_s(24)
                           => SHIFT_7_24_port, A_s(23) => SHIFT_7_23_port, 
                           A_s(22) => SHIFT_7_22_port, A_s(21) => 
                           SHIFT_7_21_port, A_s(20) => SHIFT_7_20_port, A_s(19)
                           => SHIFT_7_19_port, A_s(18) => SHIFT_7_18_port, 
                           A_s(17) => SHIFT_7_17_port, A_s(16) => 
                           SHIFT_7_16_port, A_s(15) => SHIFT_7_15_port, A_s(14)
                           => SHIFT_7_14_port, A_s(13) => SHIFT_7_13_port, 
                           A_s(12) => SHIFT_7_12_port, A_s(11) => 
                           SHIFT_7_11_port, A_s(10) => SHIFT_7_10_port, A_s(9) 
                           => SHIFT_7_9_port, A_s(8) => SHIFT_7_8_port, A_s(7) 
                           => SHIFT_7_7_port, A_s(6) => SHIFT_7_6_port, A_s(5) 
                           => SHIFT_7_5_port, A_s(4) => SHIFT_7_4_port, A_s(3) 
                           => SHIFT_7_3_port, A_s(2) => SHIFT_7_2_port, A_s(1) 
                           => SHIFT_7_1_port, A_s(0) => SHIFT_7_0_port, 
                           A_ns(47) => SHIFT_n_7_45_port, A_ns(46) => 
                           SHIFT_n_7_45_port, A_ns(45) => SHIFT_n_7_45_port, 
                           A_ns(44) => SHIFT_n_7_44_port, A_ns(43) => 
                           SHIFT_n_7_43_port, A_ns(42) => SHIFT_n_7_42_port, 
                           A_ns(41) => SHIFT_n_7_41_port, A_ns(40) => 
                           SHIFT_n_7_40_port, A_ns(39) => SHIFT_n_7_39_port, 
                           A_ns(38) => SHIFT_n_7_38_port, A_ns(37) => 
                           SHIFT_n_7_37_port, A_ns(36) => SHIFT_n_7_36_port, 
                           A_ns(35) => SHIFT_n_7_35_port, A_ns(34) => 
                           SHIFT_n_7_34_port, A_ns(33) => SHIFT_n_7_33_port, 
                           A_ns(32) => SHIFT_n_7_32_port, A_ns(31) => 
                           SHIFT_n_7_31_port, A_ns(30) => SHIFT_n_7_30_port, 
                           A_ns(29) => SHIFT_n_7_29_port, A_ns(28) => 
                           SHIFT_n_7_28_port, A_ns(27) => SHIFT_n_7_27_port, 
                           A_ns(26) => SHIFT_n_7_26_port, A_ns(25) => 
                           SHIFT_n_7_25_port, A_ns(24) => SHIFT_n_7_24_port, 
                           A_ns(23) => SHIFT_n_7_23_port, A_ns(22) => 
                           SHIFT_n_7_22_port, A_ns(21) => SHIFT_n_7_21_port, 
                           A_ns(20) => SHIFT_n_7_20_port, A_ns(19) => 
                           SHIFT_n_7_19_port, A_ns(18) => SHIFT_n_7_18_port, 
                           A_ns(17) => SHIFT_n_7_17_port, A_ns(16) => 
                           SHIFT_n_7_16_port, A_ns(15) => SHIFT_n_7_15_port, 
                           A_ns(14) => SHIFT_n_7_14_port, A_ns(13) => 
                           SHIFT_n_7_13_port, A_ns(12) => SHIFT_n_7_12_port, 
                           A_ns(11) => SHIFT_n_7_11_port, A_ns(10) => 
                           SHIFT_n_7_10_port, A_ns(9) => SHIFT_n_7_9_port, 
                           A_ns(8) => SHIFT_n_7_8_port, A_ns(7) => 
                           SHIFT_n_7_7_port, A_ns(6) => SHIFT_n_7_6_port, 
                           A_ns(5) => SHIFT_n_7_5_port, A_ns(4) => 
                           SHIFT_n_7_4_port, A_ns(3) => SHIFT_n_7_3_port, 
                           A_ns(2) => SHIFT_n_7_2_port, A_ns(1) => 
                           SHIFT_n_7_1_port, A_ns(0) => SHIFT_n_7_0_port, B(47)
                           => B(31), B(46) => B(31), B(45) => B(31), B(44) => 
                           B(31), B(43) => B(31), B(42) => B(31), B(41) => 
                           B(31), B(40) => B(31), B(39) => B(31), B(38) => 
                           B(31), B(37) => B(31), B(36) => B(31), B(35) => 
                           B(31), B(34) => B(31), B(33) => B(31), B(32) => 
                           B(31), B(31) => B(31), B(30) => B(30), B(29) => 
                           B(29), B(28) => B(28), B(27) => B(27), B(26) => 
                           B(26), B(25) => B(25), B(24) => B(24), B(23) => 
                           B(23), B(22) => B(22), B(21) => B(21), B(20) => 
                           B(20), B(19) => B(19), B(18) => B(18), B(17) => 
                           B(17), B(16) => B(16), B(15) => B(15), B(14) => 
                           B(14), B(13) => B(13), B(12) => B(12), B(11) => 
                           B(11), B(10) => B(10), B(9) => B(9), B(8) => B(8), 
                           B(7) => B(7), B(6) => B(6), B(5) => B(5), B(4) => 
                           B(4), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), O(47) => OTMP_7_47_port, O(46) => 
                           OTMP_7_46_port, O(45) => OTMP_7_45_port, O(44) => 
                           OTMP_7_44_port, O(43) => OTMP_7_43_port, O(42) => 
                           OTMP_7_42_port, O(41) => OTMP_7_41_port, O(40) => 
                           OTMP_7_40_port, O(39) => OTMP_7_39_port, O(38) => 
                           OTMP_7_38_port, O(37) => OTMP_7_37_port, O(36) => 
                           OTMP_7_36_port, O(35) => OTMP_7_35_port, O(34) => 
                           OTMP_7_34_port, O(33) => OTMP_7_33_port, O(32) => 
                           OTMP_7_32_port, O(31) => OTMP_7_31_port, O(30) => 
                           OTMP_7_30_port, O(29) => OTMP_7_29_port, O(28) => 
                           OTMP_7_28_port, O(27) => OTMP_7_27_port, O(26) => 
                           OTMP_7_26_port, O(25) => OTMP_7_25_port, O(24) => 
                           OTMP_7_24_port, O(23) => OTMP_7_23_port, O(22) => 
                           OTMP_7_22_port, O(21) => OTMP_7_21_port, O(20) => 
                           OTMP_7_20_port, O(19) => OTMP_7_19_port, O(18) => 
                           OTMP_7_18_port, O(17) => OTMP_7_17_port, O(16) => 
                           OTMP_7_16_port, O(15) => OTMP_7_15_port, O(14) => 
                           OTMP_7_14_port, O(13) => OTMP_7_13_port, O(12) => 
                           OTMP_7_12_port, O(11) => OTMP_7_11_port, O(10) => 
                           OTMP_7_10_port, O(9) => OTMP_7_9_port, O(8) => 
                           OTMP_7_8_port, O(7) => OTMP_7_7_port, O(6) => 
                           OTMP_7_6_port, O(5) => OTMP_7_5_port, O(4) => 
                           OTMP_7_4_port, O(3) => OTMP_7_3_port, O(2) => 
                           OTMP_7_2_port, O(1) => OTMP_7_1_port, O(0) => n_1112
                           , A_so(47) => SHIFT_8_47_port, A_so(46) => 
                           SHIFT_8_46_port, A_so(45) => SHIFT_8_45_port, 
                           A_so(44) => SHIFT_8_44_port, A_so(43) => 
                           SHIFT_8_43_port, A_so(42) => SHIFT_8_42_port, 
                           A_so(41) => SHIFT_8_41_port, A_so(40) => 
                           SHIFT_8_40_port, A_so(39) => SHIFT_8_39_port, 
                           A_so(38) => SHIFT_8_38_port, A_so(37) => 
                           SHIFT_8_37_port, A_so(36) => SHIFT_8_36_port, 
                           A_so(35) => SHIFT_8_35_port, A_so(34) => 
                           SHIFT_8_34_port, A_so(33) => SHIFT_8_33_port, 
                           A_so(32) => SHIFT_8_32_port, A_so(31) => 
                           SHIFT_8_31_port, A_so(30) => SHIFT_8_30_port, 
                           A_so(29) => SHIFT_8_29_port, A_so(28) => 
                           SHIFT_8_28_port, A_so(27) => SHIFT_8_27_port, 
                           A_so(26) => SHIFT_8_26_port, A_so(25) => 
                           SHIFT_8_25_port, A_so(24) => SHIFT_8_24_port, 
                           A_so(23) => SHIFT_8_23_port, A_so(22) => 
                           SHIFT_8_22_port, A_so(21) => SHIFT_8_21_port, 
                           A_so(20) => SHIFT_8_20_port, A_so(19) => 
                           SHIFT_8_19_port, A_so(18) => SHIFT_8_18_port, 
                           A_so(17) => SHIFT_8_17_port, A_so(16) => 
                           SHIFT_8_16_port, A_so(15) => SHIFT_8_15_port, 
                           A_so(14) => SHIFT_8_14_port, A_so(13) => 
                           SHIFT_8_13_port, A_so(12) => SHIFT_8_12_port, 
                           A_so(11) => SHIFT_8_11_port, A_so(10) => 
                           SHIFT_8_10_port, A_so(9) => SHIFT_8_9_port, A_so(8) 
                           => SHIFT_8_8_port, A_so(7) => SHIFT_8_7_port, 
                           A_so(6) => SHIFT_8_6_port, A_so(5) => SHIFT_8_5_port
                           , A_so(4) => SHIFT_8_4_port, A_so(3) => 
                           SHIFT_8_3_port, A_so(2) => SHIFT_8_2_port, A_so(1) 
                           => n_1113, A_so(0) => n_1114, A_nso(47) => 
                           SHIFT_n_8_47_port, A_nso(46) => SHIFT_n_8_46_port, 
                           A_nso(45) => SHIFT_n_8_45_port, A_nso(44) => 
                           SHIFT_n_8_44_port, A_nso(43) => SHIFT_n_8_43_port, 
                           A_nso(42) => SHIFT_n_8_42_port, A_nso(41) => 
                           SHIFT_n_8_41_port, A_nso(40) => SHIFT_n_8_40_port, 
                           A_nso(39) => SHIFT_n_8_39_port, A_nso(38) => 
                           SHIFT_n_8_38_port, A_nso(37) => SHIFT_n_8_37_port, 
                           A_nso(36) => SHIFT_n_8_36_port, A_nso(35) => 
                           SHIFT_n_8_35_port, A_nso(34) => SHIFT_n_8_34_port, 
                           A_nso(33) => SHIFT_n_8_33_port, A_nso(32) => 
                           SHIFT_n_8_32_port, A_nso(31) => SHIFT_n_8_31_port, 
                           A_nso(30) => SHIFT_n_8_30_port, A_nso(29) => 
                           SHIFT_n_8_29_port, A_nso(28) => SHIFT_n_8_28_port, 
                           A_nso(27) => SHIFT_n_8_27_port, A_nso(26) => 
                           SHIFT_n_8_26_port, A_nso(25) => SHIFT_n_8_25_port, 
                           A_nso(24) => SHIFT_n_8_24_port, A_nso(23) => 
                           SHIFT_n_8_23_port, A_nso(22) => SHIFT_n_8_22_port, 
                           A_nso(21) => SHIFT_n_8_21_port, A_nso(20) => 
                           SHIFT_n_8_20_port, A_nso(19) => SHIFT_n_8_19_port, 
                           A_nso(18) => SHIFT_n_8_18_port, A_nso(17) => 
                           SHIFT_n_8_17_port, A_nso(16) => SHIFT_n_8_16_port, 
                           A_nso(15) => SHIFT_n_8_15_port, A_nso(14) => 
                           SHIFT_n_8_14_port, A_nso(13) => SHIFT_n_8_13_port, 
                           A_nso(12) => SHIFT_n_8_12_port, A_nso(11) => 
                           SHIFT_n_8_11_port, A_nso(10) => SHIFT_n_8_10_port, 
                           A_nso(9) => SHIFT_n_8_9_port, A_nso(8) => 
                           SHIFT_n_8_8_port, A_nso(7) => SHIFT_n_8_7_port, 
                           A_nso(6) => SHIFT_n_8_6_port, A_nso(5) => 
                           SHIFT_n_8_5_port, A_nso(4) => SHIFT_n_8_4_port, 
                           A_nso(3) => SHIFT_n_8_3_port, A_nso(2) => 
                           SHIFT_n_8_2_port, A_nso(1) => n_1115, A_nso(0) => 
                           n_1116);
   ENC_8 : BOOTHENC_NBIT50_i16 port map( A_s(49) => SHIFT_8_47_port, A_s(48) =>
                           SHIFT_8_47_port, A_s(47) => SHIFT_8_47_port, A_s(46)
                           => SHIFT_8_46_port, A_s(45) => SHIFT_8_45_port, 
                           A_s(44) => SHIFT_8_44_port, A_s(43) => 
                           SHIFT_8_43_port, A_s(42) => SHIFT_8_42_port, A_s(41)
                           => SHIFT_8_41_port, A_s(40) => SHIFT_8_40_port, 
                           A_s(39) => SHIFT_8_39_port, A_s(38) => 
                           SHIFT_8_38_port, A_s(37) => SHIFT_8_37_port, A_s(36)
                           => SHIFT_8_36_port, A_s(35) => SHIFT_8_35_port, 
                           A_s(34) => SHIFT_8_34_port, A_s(33) => 
                           SHIFT_8_33_port, A_s(32) => SHIFT_8_32_port, A_s(31)
                           => SHIFT_8_31_port, A_s(30) => SHIFT_8_30_port, 
                           A_s(29) => SHIFT_8_29_port, A_s(28) => 
                           SHIFT_8_28_port, A_s(27) => SHIFT_8_27_port, A_s(26)
                           => SHIFT_8_26_port, A_s(25) => SHIFT_8_25_port, 
                           A_s(24) => SHIFT_8_24_port, A_s(23) => 
                           SHIFT_8_23_port, A_s(22) => SHIFT_8_22_port, A_s(21)
                           => SHIFT_8_21_port, A_s(20) => SHIFT_8_20_port, 
                           A_s(19) => SHIFT_8_19_port, A_s(18) => 
                           SHIFT_8_18_port, A_s(17) => SHIFT_8_17_port, A_s(16)
                           => SHIFT_8_16_port, A_s(15) => SHIFT_8_15_port, 
                           A_s(14) => SHIFT_8_14_port, A_s(13) => 
                           SHIFT_8_13_port, A_s(12) => SHIFT_8_12_port, A_s(11)
                           => SHIFT_8_11_port, A_s(10) => SHIFT_8_10_port, 
                           A_s(9) => SHIFT_8_9_port, A_s(8) => SHIFT_8_8_port, 
                           A_s(7) => SHIFT_8_7_port, A_s(6) => SHIFT_8_6_port, 
                           A_s(5) => SHIFT_8_5_port, A_s(4) => SHIFT_8_4_port, 
                           A_s(3) => SHIFT_8_3_port, A_s(2) => SHIFT_8_2_port, 
                           A_s(1) => SHIFT_8_1_port, A_s(0) => SHIFT_8_0_port, 
                           A_ns(49) => SHIFT_n_8_47_port, A_ns(48) => 
                           SHIFT_n_8_47_port, A_ns(47) => SHIFT_n_8_47_port, 
                           A_ns(46) => SHIFT_n_8_46_port, A_ns(45) => 
                           SHIFT_n_8_45_port, A_ns(44) => SHIFT_n_8_44_port, 
                           A_ns(43) => SHIFT_n_8_43_port, A_ns(42) => 
                           SHIFT_n_8_42_port, A_ns(41) => SHIFT_n_8_41_port, 
                           A_ns(40) => SHIFT_n_8_40_port, A_ns(39) => 
                           SHIFT_n_8_39_port, A_ns(38) => SHIFT_n_8_38_port, 
                           A_ns(37) => SHIFT_n_8_37_port, A_ns(36) => 
                           SHIFT_n_8_36_port, A_ns(35) => SHIFT_n_8_35_port, 
                           A_ns(34) => SHIFT_n_8_34_port, A_ns(33) => 
                           SHIFT_n_8_33_port, A_ns(32) => SHIFT_n_8_32_port, 
                           A_ns(31) => SHIFT_n_8_31_port, A_ns(30) => 
                           SHIFT_n_8_30_port, A_ns(29) => SHIFT_n_8_29_port, 
                           A_ns(28) => SHIFT_n_8_28_port, A_ns(27) => 
                           SHIFT_n_8_27_port, A_ns(26) => SHIFT_n_8_26_port, 
                           A_ns(25) => SHIFT_n_8_25_port, A_ns(24) => 
                           SHIFT_n_8_24_port, A_ns(23) => SHIFT_n_8_23_port, 
                           A_ns(22) => SHIFT_n_8_22_port, A_ns(21) => 
                           SHIFT_n_8_21_port, A_ns(20) => SHIFT_n_8_20_port, 
                           A_ns(19) => SHIFT_n_8_19_port, A_ns(18) => 
                           SHIFT_n_8_18_port, A_ns(17) => SHIFT_n_8_17_port, 
                           A_ns(16) => SHIFT_n_8_16_port, A_ns(15) => 
                           SHIFT_n_8_15_port, A_ns(14) => SHIFT_n_8_14_port, 
                           A_ns(13) => SHIFT_n_8_13_port, A_ns(12) => 
                           SHIFT_n_8_12_port, A_ns(11) => SHIFT_n_8_11_port, 
                           A_ns(10) => SHIFT_n_8_10_port, A_ns(9) => 
                           SHIFT_n_8_9_port, A_ns(8) => SHIFT_n_8_8_port, 
                           A_ns(7) => SHIFT_n_8_7_port, A_ns(6) => 
                           SHIFT_n_8_6_port, A_ns(5) => SHIFT_n_8_5_port, 
                           A_ns(4) => SHIFT_n_8_4_port, A_ns(3) => 
                           SHIFT_n_8_3_port, A_ns(2) => SHIFT_n_8_2_port, 
                           A_ns(1) => SHIFT_n_8_1_port, A_ns(0) => 
                           SHIFT_n_8_0_port, B(49) => B(31), B(48) => B(31), 
                           B(47) => B(31), B(46) => B(31), B(45) => B(31), 
                           B(44) => B(31), B(43) => B(31), B(42) => B(31), 
                           B(41) => B(31), B(40) => B(31), B(39) => B(31), 
                           B(38) => B(31), B(37) => B(31), B(36) => B(31), 
                           B(35) => B(31), B(34) => B(31), B(33) => B(31), 
                           B(32) => B(31), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), O(49) => OTMP_8_49_port, O(48) 
                           => OTMP_8_48_port, O(47) => OTMP_8_47_port, O(46) =>
                           OTMP_8_46_port, O(45) => OTMP_8_45_port, O(44) => 
                           OTMP_8_44_port, O(43) => OTMP_8_43_port, O(42) => 
                           OTMP_8_42_port, O(41) => OTMP_8_41_port, O(40) => 
                           OTMP_8_40_port, O(39) => OTMP_8_39_port, O(38) => 
                           OTMP_8_38_port, O(37) => OTMP_8_37_port, O(36) => 
                           OTMP_8_36_port, O(35) => OTMP_8_35_port, O(34) => 
                           OTMP_8_34_port, O(33) => OTMP_8_33_port, O(32) => 
                           OTMP_8_32_port, O(31) => OTMP_8_31_port, O(30) => 
                           OTMP_8_30_port, O(29) => OTMP_8_29_port, O(28) => 
                           OTMP_8_28_port, O(27) => OTMP_8_27_port, O(26) => 
                           OTMP_8_26_port, O(25) => OTMP_8_25_port, O(24) => 
                           OTMP_8_24_port, O(23) => OTMP_8_23_port, O(22) => 
                           OTMP_8_22_port, O(21) => OTMP_8_21_port, O(20) => 
                           OTMP_8_20_port, O(19) => OTMP_8_19_port, O(18) => 
                           OTMP_8_18_port, O(17) => OTMP_8_17_port, O(16) => 
                           OTMP_8_16_port, O(15) => OTMP_8_15_port, O(14) => 
                           OTMP_8_14_port, O(13) => OTMP_8_13_port, O(12) => 
                           OTMP_8_12_port, O(11) => OTMP_8_11_port, O(10) => 
                           OTMP_8_10_port, O(9) => OTMP_8_9_port, O(8) => 
                           OTMP_8_8_port, O(7) => OTMP_8_7_port, O(6) => 
                           OTMP_8_6_port, O(5) => OTMP_8_5_port, O(4) => 
                           OTMP_8_4_port, O(3) => OTMP_8_3_port, O(2) => 
                           OTMP_8_2_port, O(1) => OTMP_8_1_port, O(0) => n_1117
                           , A_so(49) => SHIFT_9_49_port, A_so(48) => 
                           SHIFT_9_48_port, A_so(47) => SHIFT_9_47_port, 
                           A_so(46) => SHIFT_9_46_port, A_so(45) => 
                           SHIFT_9_45_port, A_so(44) => SHIFT_9_44_port, 
                           A_so(43) => SHIFT_9_43_port, A_so(42) => 
                           SHIFT_9_42_port, A_so(41) => SHIFT_9_41_port, 
                           A_so(40) => SHIFT_9_40_port, A_so(39) => 
                           SHIFT_9_39_port, A_so(38) => SHIFT_9_38_port, 
                           A_so(37) => SHIFT_9_37_port, A_so(36) => 
                           SHIFT_9_36_port, A_so(35) => SHIFT_9_35_port, 
                           A_so(34) => SHIFT_9_34_port, A_so(33) => 
                           SHIFT_9_33_port, A_so(32) => SHIFT_9_32_port, 
                           A_so(31) => SHIFT_9_31_port, A_so(30) => 
                           SHIFT_9_30_port, A_so(29) => SHIFT_9_29_port, 
                           A_so(28) => SHIFT_9_28_port, A_so(27) => 
                           SHIFT_9_27_port, A_so(26) => SHIFT_9_26_port, 
                           A_so(25) => SHIFT_9_25_port, A_so(24) => 
                           SHIFT_9_24_port, A_so(23) => SHIFT_9_23_port, 
                           A_so(22) => SHIFT_9_22_port, A_so(21) => 
                           SHIFT_9_21_port, A_so(20) => SHIFT_9_20_port, 
                           A_so(19) => SHIFT_9_19_port, A_so(18) => 
                           SHIFT_9_18_port, A_so(17) => SHIFT_9_17_port, 
                           A_so(16) => SHIFT_9_16_port, A_so(15) => 
                           SHIFT_9_15_port, A_so(14) => SHIFT_9_14_port, 
                           A_so(13) => SHIFT_9_13_port, A_so(12) => 
                           SHIFT_9_12_port, A_so(11) => SHIFT_9_11_port, 
                           A_so(10) => SHIFT_9_10_port, A_so(9) => 
                           SHIFT_9_9_port, A_so(8) => SHIFT_9_8_port, A_so(7) 
                           => SHIFT_9_7_port, A_so(6) => SHIFT_9_6_port, 
                           A_so(5) => SHIFT_9_5_port, A_so(4) => SHIFT_9_4_port
                           , A_so(3) => SHIFT_9_3_port, A_so(2) => 
                           SHIFT_9_2_port, A_so(1) => n_1118, A_so(0) => n_1119
                           , A_nso(49) => SHIFT_n_9_49_port, A_nso(48) => 
                           SHIFT_n_9_48_port, A_nso(47) => SHIFT_n_9_47_port, 
                           A_nso(46) => SHIFT_n_9_46_port, A_nso(45) => 
                           SHIFT_n_9_45_port, A_nso(44) => SHIFT_n_9_44_port, 
                           A_nso(43) => SHIFT_n_9_43_port, A_nso(42) => 
                           SHIFT_n_9_42_port, A_nso(41) => SHIFT_n_9_41_port, 
                           A_nso(40) => SHIFT_n_9_40_port, A_nso(39) => 
                           SHIFT_n_9_39_port, A_nso(38) => SHIFT_n_9_38_port, 
                           A_nso(37) => SHIFT_n_9_37_port, A_nso(36) => 
                           SHIFT_n_9_36_port, A_nso(35) => SHIFT_n_9_35_port, 
                           A_nso(34) => SHIFT_n_9_34_port, A_nso(33) => 
                           SHIFT_n_9_33_port, A_nso(32) => SHIFT_n_9_32_port, 
                           A_nso(31) => SHIFT_n_9_31_port, A_nso(30) => 
                           SHIFT_n_9_30_port, A_nso(29) => SHIFT_n_9_29_port, 
                           A_nso(28) => SHIFT_n_9_28_port, A_nso(27) => 
                           SHIFT_n_9_27_port, A_nso(26) => SHIFT_n_9_26_port, 
                           A_nso(25) => SHIFT_n_9_25_port, A_nso(24) => 
                           SHIFT_n_9_24_port, A_nso(23) => SHIFT_n_9_23_port, 
                           A_nso(22) => SHIFT_n_9_22_port, A_nso(21) => 
                           SHIFT_n_9_21_port, A_nso(20) => SHIFT_n_9_20_port, 
                           A_nso(19) => SHIFT_n_9_19_port, A_nso(18) => 
                           SHIFT_n_9_18_port, A_nso(17) => SHIFT_n_9_17_port, 
                           A_nso(16) => SHIFT_n_9_16_port, A_nso(15) => 
                           SHIFT_n_9_15_port, A_nso(14) => SHIFT_n_9_14_port, 
                           A_nso(13) => SHIFT_n_9_13_port, A_nso(12) => 
                           SHIFT_n_9_12_port, A_nso(11) => SHIFT_n_9_11_port, 
                           A_nso(10) => SHIFT_n_9_10_port, A_nso(9) => 
                           SHIFT_n_9_9_port, A_nso(8) => SHIFT_n_9_8_port, 
                           A_nso(7) => SHIFT_n_9_7_port, A_nso(6) => 
                           SHIFT_n_9_6_port, A_nso(5) => SHIFT_n_9_5_port, 
                           A_nso(4) => SHIFT_n_9_4_port, A_nso(3) => 
                           SHIFT_n_9_3_port, A_nso(2) => SHIFT_n_9_2_port, 
                           A_nso(1) => n_1120, A_nso(0) => n_1121);
   ENC_9 : BOOTHENC_NBIT52_i18 port map( A_s(51) => SHIFT_9_49_port, A_s(50) =>
                           SHIFT_9_49_port, A_s(49) => SHIFT_9_49_port, A_s(48)
                           => SHIFT_9_48_port, A_s(47) => SHIFT_9_47_port, 
                           A_s(46) => SHIFT_9_46_port, A_s(45) => 
                           SHIFT_9_45_port, A_s(44) => SHIFT_9_44_port, A_s(43)
                           => SHIFT_9_43_port, A_s(42) => SHIFT_9_42_port, 
                           A_s(41) => SHIFT_9_41_port, A_s(40) => 
                           SHIFT_9_40_port, A_s(39) => SHIFT_9_39_port, A_s(38)
                           => SHIFT_9_38_port, A_s(37) => SHIFT_9_37_port, 
                           A_s(36) => SHIFT_9_36_port, A_s(35) => 
                           SHIFT_9_35_port, A_s(34) => SHIFT_9_34_port, A_s(33)
                           => SHIFT_9_33_port, A_s(32) => SHIFT_9_32_port, 
                           A_s(31) => SHIFT_9_31_port, A_s(30) => 
                           SHIFT_9_30_port, A_s(29) => SHIFT_9_29_port, A_s(28)
                           => SHIFT_9_28_port, A_s(27) => SHIFT_9_27_port, 
                           A_s(26) => SHIFT_9_26_port, A_s(25) => 
                           SHIFT_9_25_port, A_s(24) => SHIFT_9_24_port, A_s(23)
                           => SHIFT_9_23_port, A_s(22) => SHIFT_9_22_port, 
                           A_s(21) => SHIFT_9_21_port, A_s(20) => 
                           SHIFT_9_20_port, A_s(19) => SHIFT_9_19_port, A_s(18)
                           => SHIFT_9_18_port, A_s(17) => SHIFT_9_17_port, 
                           A_s(16) => SHIFT_9_16_port, A_s(15) => 
                           SHIFT_9_15_port, A_s(14) => SHIFT_9_14_port, A_s(13)
                           => SHIFT_9_13_port, A_s(12) => SHIFT_9_12_port, 
                           A_s(11) => SHIFT_9_11_port, A_s(10) => 
                           SHIFT_9_10_port, A_s(9) => SHIFT_9_9_port, A_s(8) =>
                           SHIFT_9_8_port, A_s(7) => SHIFT_9_7_port, A_s(6) => 
                           SHIFT_9_6_port, A_s(5) => SHIFT_9_5_port, A_s(4) => 
                           SHIFT_9_4_port, A_s(3) => SHIFT_9_3_port, A_s(2) => 
                           SHIFT_9_2_port, A_s(1) => SHIFT_9_1_port, A_s(0) => 
                           SHIFT_9_0_port, A_ns(51) => SHIFT_n_9_49_port, 
                           A_ns(50) => SHIFT_n_9_49_port, A_ns(49) => 
                           SHIFT_n_9_49_port, A_ns(48) => SHIFT_n_9_48_port, 
                           A_ns(47) => SHIFT_n_9_47_port, A_ns(46) => 
                           SHIFT_n_9_46_port, A_ns(45) => SHIFT_n_9_45_port, 
                           A_ns(44) => SHIFT_n_9_44_port, A_ns(43) => 
                           SHIFT_n_9_43_port, A_ns(42) => SHIFT_n_9_42_port, 
                           A_ns(41) => SHIFT_n_9_41_port, A_ns(40) => 
                           SHIFT_n_9_40_port, A_ns(39) => SHIFT_n_9_39_port, 
                           A_ns(38) => SHIFT_n_9_38_port, A_ns(37) => 
                           SHIFT_n_9_37_port, A_ns(36) => SHIFT_n_9_36_port, 
                           A_ns(35) => SHIFT_n_9_35_port, A_ns(34) => 
                           SHIFT_n_9_34_port, A_ns(33) => SHIFT_n_9_33_port, 
                           A_ns(32) => SHIFT_n_9_32_port, A_ns(31) => 
                           SHIFT_n_9_31_port, A_ns(30) => SHIFT_n_9_30_port, 
                           A_ns(29) => SHIFT_n_9_29_port, A_ns(28) => 
                           SHIFT_n_9_28_port, A_ns(27) => SHIFT_n_9_27_port, 
                           A_ns(26) => SHIFT_n_9_26_port, A_ns(25) => 
                           SHIFT_n_9_25_port, A_ns(24) => SHIFT_n_9_24_port, 
                           A_ns(23) => SHIFT_n_9_23_port, A_ns(22) => 
                           SHIFT_n_9_22_port, A_ns(21) => SHIFT_n_9_21_port, 
                           A_ns(20) => SHIFT_n_9_20_port, A_ns(19) => 
                           SHIFT_n_9_19_port, A_ns(18) => SHIFT_n_9_18_port, 
                           A_ns(17) => SHIFT_n_9_17_port, A_ns(16) => 
                           SHIFT_n_9_16_port, A_ns(15) => SHIFT_n_9_15_port, 
                           A_ns(14) => SHIFT_n_9_14_port, A_ns(13) => 
                           SHIFT_n_9_13_port, A_ns(12) => SHIFT_n_9_12_port, 
                           A_ns(11) => SHIFT_n_9_11_port, A_ns(10) => 
                           SHIFT_n_9_10_port, A_ns(9) => SHIFT_n_9_9_port, 
                           A_ns(8) => SHIFT_n_9_8_port, A_ns(7) => 
                           SHIFT_n_9_7_port, A_ns(6) => SHIFT_n_9_6_port, 
                           A_ns(5) => SHIFT_n_9_5_port, A_ns(4) => 
                           SHIFT_n_9_4_port, A_ns(3) => SHIFT_n_9_3_port, 
                           A_ns(2) => SHIFT_n_9_2_port, A_ns(1) => 
                           SHIFT_n_9_1_port, A_ns(0) => SHIFT_n_9_0_port, B(51)
                           => B(31), B(50) => B(31), B(49) => B(31), B(48) => 
                           B(31), B(47) => B(31), B(46) => B(31), B(45) => 
                           B(31), B(44) => B(31), B(43) => B(31), B(42) => 
                           B(31), B(41) => B(31), B(40) => B(31), B(39) => 
                           B(31), B(38) => B(31), B(37) => B(31), B(36) => 
                           B(31), B(35) => B(31), B(34) => B(31), B(33) => 
                           B(31), B(32) => B(31), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), O(51) => OTMP_9_51_port, 
                           O(50) => OTMP_9_50_port, O(49) => OTMP_9_49_port, 
                           O(48) => OTMP_9_48_port, O(47) => OTMP_9_47_port, 
                           O(46) => OTMP_9_46_port, O(45) => OTMP_9_45_port, 
                           O(44) => OTMP_9_44_port, O(43) => OTMP_9_43_port, 
                           O(42) => OTMP_9_42_port, O(41) => OTMP_9_41_port, 
                           O(40) => OTMP_9_40_port, O(39) => OTMP_9_39_port, 
                           O(38) => OTMP_9_38_port, O(37) => OTMP_9_37_port, 
                           O(36) => OTMP_9_36_port, O(35) => OTMP_9_35_port, 
                           O(34) => OTMP_9_34_port, O(33) => OTMP_9_33_port, 
                           O(32) => OTMP_9_32_port, O(31) => OTMP_9_31_port, 
                           O(30) => OTMP_9_30_port, O(29) => OTMP_9_29_port, 
                           O(28) => OTMP_9_28_port, O(27) => OTMP_9_27_port, 
                           O(26) => OTMP_9_26_port, O(25) => OTMP_9_25_port, 
                           O(24) => OTMP_9_24_port, O(23) => OTMP_9_23_port, 
                           O(22) => OTMP_9_22_port, O(21) => OTMP_9_21_port, 
                           O(20) => OTMP_9_20_port, O(19) => OTMP_9_19_port, 
                           O(18) => OTMP_9_18_port, O(17) => OTMP_9_17_port, 
                           O(16) => OTMP_9_16_port, O(15) => OTMP_9_15_port, 
                           O(14) => OTMP_9_14_port, O(13) => OTMP_9_13_port, 
                           O(12) => OTMP_9_12_port, O(11) => OTMP_9_11_port, 
                           O(10) => OTMP_9_10_port, O(9) => OTMP_9_9_port, O(8)
                           => OTMP_9_8_port, O(7) => OTMP_9_7_port, O(6) => 
                           OTMP_9_6_port, O(5) => OTMP_9_5_port, O(4) => 
                           OTMP_9_4_port, O(3) => OTMP_9_3_port, O(2) => 
                           OTMP_9_2_port, O(1) => OTMP_9_1_port, O(0) => n_1122
                           , A_so(51) => SHIFT_10_51_port, A_so(50) => 
                           SHIFT_10_50_port, A_so(49) => SHIFT_10_49_port, 
                           A_so(48) => SHIFT_10_48_port, A_so(47) => 
                           SHIFT_10_47_port, A_so(46) => SHIFT_10_46_port, 
                           A_so(45) => SHIFT_10_45_port, A_so(44) => 
                           SHIFT_10_44_port, A_so(43) => SHIFT_10_43_port, 
                           A_so(42) => SHIFT_10_42_port, A_so(41) => 
                           SHIFT_10_41_port, A_so(40) => SHIFT_10_40_port, 
                           A_so(39) => SHIFT_10_39_port, A_so(38) => 
                           SHIFT_10_38_port, A_so(37) => SHIFT_10_37_port, 
                           A_so(36) => SHIFT_10_36_port, A_so(35) => 
                           SHIFT_10_35_port, A_so(34) => SHIFT_10_34_port, 
                           A_so(33) => SHIFT_10_33_port, A_so(32) => 
                           SHIFT_10_32_port, A_so(31) => SHIFT_10_31_port, 
                           A_so(30) => SHIFT_10_30_port, A_so(29) => 
                           SHIFT_10_29_port, A_so(28) => SHIFT_10_28_port, 
                           A_so(27) => SHIFT_10_27_port, A_so(26) => 
                           SHIFT_10_26_port, A_so(25) => SHIFT_10_25_port, 
                           A_so(24) => SHIFT_10_24_port, A_so(23) => 
                           SHIFT_10_23_port, A_so(22) => SHIFT_10_22_port, 
                           A_so(21) => SHIFT_10_21_port, A_so(20) => 
                           SHIFT_10_20_port, A_so(19) => SHIFT_10_19_port, 
                           A_so(18) => SHIFT_10_18_port, A_so(17) => 
                           SHIFT_10_17_port, A_so(16) => SHIFT_10_16_port, 
                           A_so(15) => SHIFT_10_15_port, A_so(14) => 
                           SHIFT_10_14_port, A_so(13) => SHIFT_10_13_port, 
                           A_so(12) => SHIFT_10_12_port, A_so(11) => 
                           SHIFT_10_11_port, A_so(10) => SHIFT_10_10_port, 
                           A_so(9) => SHIFT_10_9_port, A_so(8) => 
                           SHIFT_10_8_port, A_so(7) => SHIFT_10_7_port, A_so(6)
                           => SHIFT_10_6_port, A_so(5) => SHIFT_10_5_port, 
                           A_so(4) => SHIFT_10_4_port, A_so(3) => 
                           SHIFT_10_3_port, A_so(2) => SHIFT_10_2_port, A_so(1)
                           => n_1123, A_so(0) => n_1124, A_nso(51) => 
                           SHIFT_n_10_51_port, A_nso(50) => SHIFT_n_10_50_port,
                           A_nso(49) => SHIFT_n_10_49_port, A_nso(48) => 
                           SHIFT_n_10_48_port, A_nso(47) => SHIFT_n_10_47_port,
                           A_nso(46) => SHIFT_n_10_46_port, A_nso(45) => 
                           SHIFT_n_10_45_port, A_nso(44) => SHIFT_n_10_44_port,
                           A_nso(43) => SHIFT_n_10_43_port, A_nso(42) => 
                           SHIFT_n_10_42_port, A_nso(41) => SHIFT_n_10_41_port,
                           A_nso(40) => SHIFT_n_10_40_port, A_nso(39) => 
                           SHIFT_n_10_39_port, A_nso(38) => SHIFT_n_10_38_port,
                           A_nso(37) => SHIFT_n_10_37_port, A_nso(36) => 
                           SHIFT_n_10_36_port, A_nso(35) => SHIFT_n_10_35_port,
                           A_nso(34) => SHIFT_n_10_34_port, A_nso(33) => 
                           SHIFT_n_10_33_port, A_nso(32) => SHIFT_n_10_32_port,
                           A_nso(31) => SHIFT_n_10_31_port, A_nso(30) => 
                           SHIFT_n_10_30_port, A_nso(29) => SHIFT_n_10_29_port,
                           A_nso(28) => SHIFT_n_10_28_port, A_nso(27) => 
                           SHIFT_n_10_27_port, A_nso(26) => SHIFT_n_10_26_port,
                           A_nso(25) => SHIFT_n_10_25_port, A_nso(24) => 
                           SHIFT_n_10_24_port, A_nso(23) => SHIFT_n_10_23_port,
                           A_nso(22) => SHIFT_n_10_22_port, A_nso(21) => 
                           SHIFT_n_10_21_port, A_nso(20) => SHIFT_n_10_20_port,
                           A_nso(19) => SHIFT_n_10_19_port, A_nso(18) => 
                           SHIFT_n_10_18_port, A_nso(17) => SHIFT_n_10_17_port,
                           A_nso(16) => SHIFT_n_10_16_port, A_nso(15) => 
                           SHIFT_n_10_15_port, A_nso(14) => SHIFT_n_10_14_port,
                           A_nso(13) => SHIFT_n_10_13_port, A_nso(12) => 
                           SHIFT_n_10_12_port, A_nso(11) => SHIFT_n_10_11_port,
                           A_nso(10) => SHIFT_n_10_10_port, A_nso(9) => 
                           SHIFT_n_10_9_port, A_nso(8) => SHIFT_n_10_8_port, 
                           A_nso(7) => SHIFT_n_10_7_port, A_nso(6) => 
                           SHIFT_n_10_6_port, A_nso(5) => SHIFT_n_10_5_port, 
                           A_nso(4) => SHIFT_n_10_4_port, A_nso(3) => 
                           SHIFT_n_10_3_port, A_nso(2) => SHIFT_n_10_2_port, 
                           A_nso(1) => n_1125, A_nso(0) => n_1126);
   ENC_10 : BOOTHENC_NBIT54_i20 port map( A_s(53) => SHIFT_10_51_port, A_s(52) 
                           => SHIFT_10_51_port, A_s(51) => SHIFT_10_51_port, 
                           A_s(50) => SHIFT_10_50_port, A_s(49) => 
                           SHIFT_10_49_port, A_s(48) => SHIFT_10_48_port, 
                           A_s(47) => SHIFT_10_47_port, A_s(46) => 
                           SHIFT_10_46_port, A_s(45) => SHIFT_10_45_port, 
                           A_s(44) => SHIFT_10_44_port, A_s(43) => 
                           SHIFT_10_43_port, A_s(42) => SHIFT_10_42_port, 
                           A_s(41) => SHIFT_10_41_port, A_s(40) => 
                           SHIFT_10_40_port, A_s(39) => SHIFT_10_39_port, 
                           A_s(38) => SHIFT_10_38_port, A_s(37) => 
                           SHIFT_10_37_port, A_s(36) => SHIFT_10_36_port, 
                           A_s(35) => SHIFT_10_35_port, A_s(34) => 
                           SHIFT_10_34_port, A_s(33) => SHIFT_10_33_port, 
                           A_s(32) => SHIFT_10_32_port, A_s(31) => 
                           SHIFT_10_31_port, A_s(30) => SHIFT_10_30_port, 
                           A_s(29) => SHIFT_10_29_port, A_s(28) => 
                           SHIFT_10_28_port, A_s(27) => SHIFT_10_27_port, 
                           A_s(26) => SHIFT_10_26_port, A_s(25) => 
                           SHIFT_10_25_port, A_s(24) => SHIFT_10_24_port, 
                           A_s(23) => SHIFT_10_23_port, A_s(22) => 
                           SHIFT_10_22_port, A_s(21) => SHIFT_10_21_port, 
                           A_s(20) => SHIFT_10_20_port, A_s(19) => 
                           SHIFT_10_19_port, A_s(18) => SHIFT_10_18_port, 
                           A_s(17) => SHIFT_10_17_port, A_s(16) => 
                           SHIFT_10_16_port, A_s(15) => SHIFT_10_15_port, 
                           A_s(14) => SHIFT_10_14_port, A_s(13) => 
                           SHIFT_10_13_port, A_s(12) => SHIFT_10_12_port, 
                           A_s(11) => SHIFT_10_11_port, A_s(10) => 
                           SHIFT_10_10_port, A_s(9) => SHIFT_10_9_port, A_s(8) 
                           => SHIFT_10_8_port, A_s(7) => SHIFT_10_7_port, 
                           A_s(6) => SHIFT_10_6_port, A_s(5) => SHIFT_10_5_port
                           , A_s(4) => SHIFT_10_4_port, A_s(3) => 
                           SHIFT_10_3_port, A_s(2) => SHIFT_10_2_port, A_s(1) 
                           => SHIFT_10_1_port, A_s(0) => SHIFT_10_0_port, 
                           A_ns(53) => SHIFT_n_10_51_port, A_ns(52) => 
                           SHIFT_n_10_51_port, A_ns(51) => SHIFT_n_10_51_port, 
                           A_ns(50) => SHIFT_n_10_50_port, A_ns(49) => 
                           SHIFT_n_10_49_port, A_ns(48) => SHIFT_n_10_48_port, 
                           A_ns(47) => SHIFT_n_10_47_port, A_ns(46) => 
                           SHIFT_n_10_46_port, A_ns(45) => SHIFT_n_10_45_port, 
                           A_ns(44) => SHIFT_n_10_44_port, A_ns(43) => 
                           SHIFT_n_10_43_port, A_ns(42) => SHIFT_n_10_42_port, 
                           A_ns(41) => SHIFT_n_10_41_port, A_ns(40) => 
                           SHIFT_n_10_40_port, A_ns(39) => SHIFT_n_10_39_port, 
                           A_ns(38) => SHIFT_n_10_38_port, A_ns(37) => 
                           SHIFT_n_10_37_port, A_ns(36) => SHIFT_n_10_36_port, 
                           A_ns(35) => SHIFT_n_10_35_port, A_ns(34) => 
                           SHIFT_n_10_34_port, A_ns(33) => SHIFT_n_10_33_port, 
                           A_ns(32) => SHIFT_n_10_32_port, A_ns(31) => 
                           SHIFT_n_10_31_port, A_ns(30) => SHIFT_n_10_30_port, 
                           A_ns(29) => SHIFT_n_10_29_port, A_ns(28) => 
                           SHIFT_n_10_28_port, A_ns(27) => SHIFT_n_10_27_port, 
                           A_ns(26) => SHIFT_n_10_26_port, A_ns(25) => 
                           SHIFT_n_10_25_port, A_ns(24) => SHIFT_n_10_24_port, 
                           A_ns(23) => SHIFT_n_10_23_port, A_ns(22) => 
                           SHIFT_n_10_22_port, A_ns(21) => SHIFT_n_10_21_port, 
                           A_ns(20) => SHIFT_n_10_20_port, A_ns(19) => 
                           SHIFT_n_10_19_port, A_ns(18) => SHIFT_n_10_18_port, 
                           A_ns(17) => SHIFT_n_10_17_port, A_ns(16) => 
                           SHIFT_n_10_16_port, A_ns(15) => SHIFT_n_10_15_port, 
                           A_ns(14) => SHIFT_n_10_14_port, A_ns(13) => 
                           SHIFT_n_10_13_port, A_ns(12) => SHIFT_n_10_12_port, 
                           A_ns(11) => SHIFT_n_10_11_port, A_ns(10) => 
                           SHIFT_n_10_10_port, A_ns(9) => SHIFT_n_10_9_port, 
                           A_ns(8) => SHIFT_n_10_8_port, A_ns(7) => 
                           SHIFT_n_10_7_port, A_ns(6) => SHIFT_n_10_6_port, 
                           A_ns(5) => SHIFT_n_10_5_port, A_ns(4) => 
                           SHIFT_n_10_4_port, A_ns(3) => SHIFT_n_10_3_port, 
                           A_ns(2) => SHIFT_n_10_2_port, A_ns(1) => 
                           SHIFT_n_10_1_port, A_ns(0) => SHIFT_n_10_0_port, 
                           B(53) => B(31), B(52) => B(31), B(51) => B(31), 
                           B(50) => B(31), B(49) => B(31), B(48) => B(31), 
                           B(47) => B(31), B(46) => B(31), B(45) => B(31), 
                           B(44) => B(31), B(43) => B(31), B(42) => B(31), 
                           B(41) => B(31), B(40) => B(31), B(39) => B(31), 
                           B(38) => B(31), B(37) => B(31), B(36) => B(31), 
                           B(35) => B(31), B(34) => B(31), B(33) => B(31), 
                           B(32) => B(31), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), O(53) => OTMP_10_53_port, O(52) 
                           => OTMP_10_52_port, O(51) => OTMP_10_51_port, O(50) 
                           => OTMP_10_50_port, O(49) => OTMP_10_49_port, O(48) 
                           => OTMP_10_48_port, O(47) => OTMP_10_47_port, O(46) 
                           => OTMP_10_46_port, O(45) => OTMP_10_45_port, O(44) 
                           => OTMP_10_44_port, O(43) => OTMP_10_43_port, O(42) 
                           => OTMP_10_42_port, O(41) => OTMP_10_41_port, O(40) 
                           => OTMP_10_40_port, O(39) => OTMP_10_39_port, O(38) 
                           => OTMP_10_38_port, O(37) => OTMP_10_37_port, O(36) 
                           => OTMP_10_36_port, O(35) => OTMP_10_35_port, O(34) 
                           => OTMP_10_34_port, O(33) => OTMP_10_33_port, O(32) 
                           => OTMP_10_32_port, O(31) => OTMP_10_31_port, O(30) 
                           => OTMP_10_30_port, O(29) => OTMP_10_29_port, O(28) 
                           => OTMP_10_28_port, O(27) => OTMP_10_27_port, O(26) 
                           => OTMP_10_26_port, O(25) => OTMP_10_25_port, O(24) 
                           => OTMP_10_24_port, O(23) => OTMP_10_23_port, O(22) 
                           => OTMP_10_22_port, O(21) => OTMP_10_21_port, O(20) 
                           => OTMP_10_20_port, O(19) => OTMP_10_19_port, O(18) 
                           => OTMP_10_18_port, O(17) => OTMP_10_17_port, O(16) 
                           => OTMP_10_16_port, O(15) => OTMP_10_15_port, O(14) 
                           => OTMP_10_14_port, O(13) => OTMP_10_13_port, O(12) 
                           => OTMP_10_12_port, O(11) => OTMP_10_11_port, O(10) 
                           => OTMP_10_10_port, O(9) => OTMP_10_9_port, O(8) => 
                           OTMP_10_8_port, O(7) => OTMP_10_7_port, O(6) => 
                           OTMP_10_6_port, O(5) => OTMP_10_5_port, O(4) => 
                           OTMP_10_4_port, O(3) => OTMP_10_3_port, O(2) => 
                           OTMP_10_2_port, O(1) => OTMP_10_1_port, O(0) => 
                           n_1127, A_so(53) => SHIFT_11_53_port, A_so(52) => 
                           SHIFT_11_52_port, A_so(51) => SHIFT_11_51_port, 
                           A_so(50) => SHIFT_11_50_port, A_so(49) => 
                           SHIFT_11_49_port, A_so(48) => SHIFT_11_48_port, 
                           A_so(47) => SHIFT_11_47_port, A_so(46) => 
                           SHIFT_11_46_port, A_so(45) => SHIFT_11_45_port, 
                           A_so(44) => SHIFT_11_44_port, A_so(43) => 
                           SHIFT_11_43_port, A_so(42) => SHIFT_11_42_port, 
                           A_so(41) => SHIFT_11_41_port, A_so(40) => 
                           SHIFT_11_40_port, A_so(39) => SHIFT_11_39_port, 
                           A_so(38) => SHIFT_11_38_port, A_so(37) => 
                           SHIFT_11_37_port, A_so(36) => SHIFT_11_36_port, 
                           A_so(35) => SHIFT_11_35_port, A_so(34) => 
                           SHIFT_11_34_port, A_so(33) => SHIFT_11_33_port, 
                           A_so(32) => SHIFT_11_32_port, A_so(31) => 
                           SHIFT_11_31_port, A_so(30) => SHIFT_11_30_port, 
                           A_so(29) => SHIFT_11_29_port, A_so(28) => 
                           SHIFT_11_28_port, A_so(27) => SHIFT_11_27_port, 
                           A_so(26) => SHIFT_11_26_port, A_so(25) => 
                           SHIFT_11_25_port, A_so(24) => SHIFT_11_24_port, 
                           A_so(23) => SHIFT_11_23_port, A_so(22) => 
                           SHIFT_11_22_port, A_so(21) => SHIFT_11_21_port, 
                           A_so(20) => SHIFT_11_20_port, A_so(19) => 
                           SHIFT_11_19_port, A_so(18) => SHIFT_11_18_port, 
                           A_so(17) => SHIFT_11_17_port, A_so(16) => 
                           SHIFT_11_16_port, A_so(15) => SHIFT_11_15_port, 
                           A_so(14) => SHIFT_11_14_port, A_so(13) => 
                           SHIFT_11_13_port, A_so(12) => SHIFT_11_12_port, 
                           A_so(11) => SHIFT_11_11_port, A_so(10) => 
                           SHIFT_11_10_port, A_so(9) => SHIFT_11_9_port, 
                           A_so(8) => SHIFT_11_8_port, A_so(7) => 
                           SHIFT_11_7_port, A_so(6) => SHIFT_11_6_port, A_so(5)
                           => SHIFT_11_5_port, A_so(4) => SHIFT_11_4_port, 
                           A_so(3) => SHIFT_11_3_port, A_so(2) => 
                           SHIFT_11_2_port, A_so(1) => n_1128, A_so(0) => 
                           n_1129, A_nso(53) => SHIFT_n_11_53_port, A_nso(52) 
                           => SHIFT_n_11_52_port, A_nso(51) => 
                           SHIFT_n_11_51_port, A_nso(50) => SHIFT_n_11_50_port,
                           A_nso(49) => SHIFT_n_11_49_port, A_nso(48) => 
                           SHIFT_n_11_48_port, A_nso(47) => SHIFT_n_11_47_port,
                           A_nso(46) => SHIFT_n_11_46_port, A_nso(45) => 
                           SHIFT_n_11_45_port, A_nso(44) => SHIFT_n_11_44_port,
                           A_nso(43) => SHIFT_n_11_43_port, A_nso(42) => 
                           SHIFT_n_11_42_port, A_nso(41) => SHIFT_n_11_41_port,
                           A_nso(40) => SHIFT_n_11_40_port, A_nso(39) => 
                           SHIFT_n_11_39_port, A_nso(38) => SHIFT_n_11_38_port,
                           A_nso(37) => SHIFT_n_11_37_port, A_nso(36) => 
                           SHIFT_n_11_36_port, A_nso(35) => SHIFT_n_11_35_port,
                           A_nso(34) => SHIFT_n_11_34_port, A_nso(33) => 
                           SHIFT_n_11_33_port, A_nso(32) => SHIFT_n_11_32_port,
                           A_nso(31) => SHIFT_n_11_31_port, A_nso(30) => 
                           SHIFT_n_11_30_port, A_nso(29) => SHIFT_n_11_29_port,
                           A_nso(28) => SHIFT_n_11_28_port, A_nso(27) => 
                           SHIFT_n_11_27_port, A_nso(26) => SHIFT_n_11_26_port,
                           A_nso(25) => SHIFT_n_11_25_port, A_nso(24) => 
                           SHIFT_n_11_24_port, A_nso(23) => SHIFT_n_11_23_port,
                           A_nso(22) => SHIFT_n_11_22_port, A_nso(21) => 
                           SHIFT_n_11_21_port, A_nso(20) => SHIFT_n_11_20_port,
                           A_nso(19) => SHIFT_n_11_19_port, A_nso(18) => 
                           SHIFT_n_11_18_port, A_nso(17) => SHIFT_n_11_17_port,
                           A_nso(16) => SHIFT_n_11_16_port, A_nso(15) => 
                           SHIFT_n_11_15_port, A_nso(14) => SHIFT_n_11_14_port,
                           A_nso(13) => SHIFT_n_11_13_port, A_nso(12) => 
                           SHIFT_n_11_12_port, A_nso(11) => SHIFT_n_11_11_port,
                           A_nso(10) => SHIFT_n_11_10_port, A_nso(9) => 
                           SHIFT_n_11_9_port, A_nso(8) => SHIFT_n_11_8_port, 
                           A_nso(7) => SHIFT_n_11_7_port, A_nso(6) => 
                           SHIFT_n_11_6_port, A_nso(5) => SHIFT_n_11_5_port, 
                           A_nso(4) => SHIFT_n_11_4_port, A_nso(3) => 
                           SHIFT_n_11_3_port, A_nso(2) => SHIFT_n_11_2_port, 
                           A_nso(1) => n_1130, A_nso(0) => n_1131);
   ENC_11 : BOOTHENC_NBIT56_i22 port map( A_s(55) => SHIFT_11_53_port, A_s(54) 
                           => SHIFT_11_53_port, A_s(53) => SHIFT_11_53_port, 
                           A_s(52) => SHIFT_11_52_port, A_s(51) => 
                           SHIFT_11_51_port, A_s(50) => SHIFT_11_50_port, 
                           A_s(49) => SHIFT_11_49_port, A_s(48) => 
                           SHIFT_11_48_port, A_s(47) => SHIFT_11_47_port, 
                           A_s(46) => SHIFT_11_46_port, A_s(45) => 
                           SHIFT_11_45_port, A_s(44) => SHIFT_11_44_port, 
                           A_s(43) => SHIFT_11_43_port, A_s(42) => 
                           SHIFT_11_42_port, A_s(41) => SHIFT_11_41_port, 
                           A_s(40) => SHIFT_11_40_port, A_s(39) => 
                           SHIFT_11_39_port, A_s(38) => SHIFT_11_38_port, 
                           A_s(37) => SHIFT_11_37_port, A_s(36) => 
                           SHIFT_11_36_port, A_s(35) => SHIFT_11_35_port, 
                           A_s(34) => SHIFT_11_34_port, A_s(33) => 
                           SHIFT_11_33_port, A_s(32) => SHIFT_11_32_port, 
                           A_s(31) => SHIFT_11_31_port, A_s(30) => 
                           SHIFT_11_30_port, A_s(29) => SHIFT_11_29_port, 
                           A_s(28) => SHIFT_11_28_port, A_s(27) => 
                           SHIFT_11_27_port, A_s(26) => SHIFT_11_26_port, 
                           A_s(25) => SHIFT_11_25_port, A_s(24) => 
                           SHIFT_11_24_port, A_s(23) => SHIFT_11_23_port, 
                           A_s(22) => SHIFT_11_22_port, A_s(21) => 
                           SHIFT_11_21_port, A_s(20) => SHIFT_11_20_port, 
                           A_s(19) => SHIFT_11_19_port, A_s(18) => 
                           SHIFT_11_18_port, A_s(17) => SHIFT_11_17_port, 
                           A_s(16) => SHIFT_11_16_port, A_s(15) => 
                           SHIFT_11_15_port, A_s(14) => SHIFT_11_14_port, 
                           A_s(13) => SHIFT_11_13_port, A_s(12) => 
                           SHIFT_11_12_port, A_s(11) => SHIFT_11_11_port, 
                           A_s(10) => SHIFT_11_10_port, A_s(9) => 
                           SHIFT_11_9_port, A_s(8) => SHIFT_11_8_port, A_s(7) 
                           => SHIFT_11_7_port, A_s(6) => SHIFT_11_6_port, 
                           A_s(5) => SHIFT_11_5_port, A_s(4) => SHIFT_11_4_port
                           , A_s(3) => SHIFT_11_3_port, A_s(2) => 
                           SHIFT_11_2_port, A_s(1) => SHIFT_11_1_port, A_s(0) 
                           => SHIFT_11_0_port, A_ns(55) => SHIFT_n_11_53_port, 
                           A_ns(54) => SHIFT_n_11_53_port, A_ns(53) => 
                           SHIFT_n_11_53_port, A_ns(52) => SHIFT_n_11_52_port, 
                           A_ns(51) => SHIFT_n_11_51_port, A_ns(50) => 
                           SHIFT_n_11_50_port, A_ns(49) => SHIFT_n_11_49_port, 
                           A_ns(48) => SHIFT_n_11_48_port, A_ns(47) => 
                           SHIFT_n_11_47_port, A_ns(46) => SHIFT_n_11_46_port, 
                           A_ns(45) => SHIFT_n_11_45_port, A_ns(44) => 
                           SHIFT_n_11_44_port, A_ns(43) => SHIFT_n_11_43_port, 
                           A_ns(42) => SHIFT_n_11_42_port, A_ns(41) => 
                           SHIFT_n_11_41_port, A_ns(40) => SHIFT_n_11_40_port, 
                           A_ns(39) => SHIFT_n_11_39_port, A_ns(38) => 
                           SHIFT_n_11_38_port, A_ns(37) => SHIFT_n_11_37_port, 
                           A_ns(36) => SHIFT_n_11_36_port, A_ns(35) => 
                           SHIFT_n_11_35_port, A_ns(34) => SHIFT_n_11_34_port, 
                           A_ns(33) => SHIFT_n_11_33_port, A_ns(32) => 
                           SHIFT_n_11_32_port, A_ns(31) => SHIFT_n_11_31_port, 
                           A_ns(30) => SHIFT_n_11_30_port, A_ns(29) => 
                           SHIFT_n_11_29_port, A_ns(28) => SHIFT_n_11_28_port, 
                           A_ns(27) => SHIFT_n_11_27_port, A_ns(26) => 
                           SHIFT_n_11_26_port, A_ns(25) => SHIFT_n_11_25_port, 
                           A_ns(24) => SHIFT_n_11_24_port, A_ns(23) => 
                           SHIFT_n_11_23_port, A_ns(22) => SHIFT_n_11_22_port, 
                           A_ns(21) => SHIFT_n_11_21_port, A_ns(20) => 
                           SHIFT_n_11_20_port, A_ns(19) => SHIFT_n_11_19_port, 
                           A_ns(18) => SHIFT_n_11_18_port, A_ns(17) => 
                           SHIFT_n_11_17_port, A_ns(16) => SHIFT_n_11_16_port, 
                           A_ns(15) => SHIFT_n_11_15_port, A_ns(14) => 
                           SHIFT_n_11_14_port, A_ns(13) => SHIFT_n_11_13_port, 
                           A_ns(12) => SHIFT_n_11_12_port, A_ns(11) => 
                           SHIFT_n_11_11_port, A_ns(10) => SHIFT_n_11_10_port, 
                           A_ns(9) => SHIFT_n_11_9_port, A_ns(8) => 
                           SHIFT_n_11_8_port, A_ns(7) => SHIFT_n_11_7_port, 
                           A_ns(6) => SHIFT_n_11_6_port, A_ns(5) => 
                           SHIFT_n_11_5_port, A_ns(4) => SHIFT_n_11_4_port, 
                           A_ns(3) => SHIFT_n_11_3_port, A_ns(2) => 
                           SHIFT_n_11_2_port, A_ns(1) => SHIFT_n_11_1_port, 
                           A_ns(0) => SHIFT_n_11_0_port, B(55) => B(31), B(54) 
                           => B(31), B(53) => B(31), B(52) => B(31), B(51) => 
                           B(31), B(50) => B(31), B(49) => B(31), B(48) => 
                           B(31), B(47) => B(31), B(46) => B(31), B(45) => 
                           B(31), B(44) => B(31), B(43) => B(31), B(42) => 
                           B(31), B(41) => B(31), B(40) => B(31), B(39) => 
                           B(31), B(38) => B(31), B(37) => B(31), B(36) => 
                           B(31), B(35) => B(31), B(34) => B(31), B(33) => 
                           B(31), B(32) => B(31), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), O(55) => OTMP_11_55_port, 
                           O(54) => OTMP_11_54_port, O(53) => OTMP_11_53_port, 
                           O(52) => OTMP_11_52_port, O(51) => OTMP_11_51_port, 
                           O(50) => OTMP_11_50_port, O(49) => OTMP_11_49_port, 
                           O(48) => OTMP_11_48_port, O(47) => OTMP_11_47_port, 
                           O(46) => OTMP_11_46_port, O(45) => OTMP_11_45_port, 
                           O(44) => OTMP_11_44_port, O(43) => OTMP_11_43_port, 
                           O(42) => OTMP_11_42_port, O(41) => OTMP_11_41_port, 
                           O(40) => OTMP_11_40_port, O(39) => OTMP_11_39_port, 
                           O(38) => OTMP_11_38_port, O(37) => OTMP_11_37_port, 
                           O(36) => OTMP_11_36_port, O(35) => OTMP_11_35_port, 
                           O(34) => OTMP_11_34_port, O(33) => OTMP_11_33_port, 
                           O(32) => OTMP_11_32_port, O(31) => OTMP_11_31_port, 
                           O(30) => OTMP_11_30_port, O(29) => OTMP_11_29_port, 
                           O(28) => OTMP_11_28_port, O(27) => OTMP_11_27_port, 
                           O(26) => OTMP_11_26_port, O(25) => OTMP_11_25_port, 
                           O(24) => OTMP_11_24_port, O(23) => OTMP_11_23_port, 
                           O(22) => OTMP_11_22_port, O(21) => OTMP_11_21_port, 
                           O(20) => OTMP_11_20_port, O(19) => OTMP_11_19_port, 
                           O(18) => OTMP_11_18_port, O(17) => OTMP_11_17_port, 
                           O(16) => OTMP_11_16_port, O(15) => OTMP_11_15_port, 
                           O(14) => OTMP_11_14_port, O(13) => OTMP_11_13_port, 
                           O(12) => OTMP_11_12_port, O(11) => OTMP_11_11_port, 
                           O(10) => OTMP_11_10_port, O(9) => OTMP_11_9_port, 
                           O(8) => OTMP_11_8_port, O(7) => OTMP_11_7_port, O(6)
                           => OTMP_11_6_port, O(5) => OTMP_11_5_port, O(4) => 
                           OTMP_11_4_port, O(3) => OTMP_11_3_port, O(2) => 
                           OTMP_11_2_port, O(1) => OTMP_11_1_port, O(0) => 
                           n_1132, A_so(55) => SHIFT_12_55_port, A_so(54) => 
                           SHIFT_12_54_port, A_so(53) => SHIFT_12_53_port, 
                           A_so(52) => SHIFT_12_52_port, A_so(51) => 
                           SHIFT_12_51_port, A_so(50) => SHIFT_12_50_port, 
                           A_so(49) => SHIFT_12_49_port, A_so(48) => 
                           SHIFT_12_48_port, A_so(47) => SHIFT_12_47_port, 
                           A_so(46) => SHIFT_12_46_port, A_so(45) => 
                           SHIFT_12_45_port, A_so(44) => SHIFT_12_44_port, 
                           A_so(43) => SHIFT_12_43_port, A_so(42) => 
                           SHIFT_12_42_port, A_so(41) => SHIFT_12_41_port, 
                           A_so(40) => SHIFT_12_40_port, A_so(39) => 
                           SHIFT_12_39_port, A_so(38) => SHIFT_12_38_port, 
                           A_so(37) => SHIFT_12_37_port, A_so(36) => 
                           SHIFT_12_36_port, A_so(35) => SHIFT_12_35_port, 
                           A_so(34) => SHIFT_12_34_port, A_so(33) => 
                           SHIFT_12_33_port, A_so(32) => SHIFT_12_32_port, 
                           A_so(31) => SHIFT_12_31_port, A_so(30) => 
                           SHIFT_12_30_port, A_so(29) => SHIFT_12_29_port, 
                           A_so(28) => SHIFT_12_28_port, A_so(27) => 
                           SHIFT_12_27_port, A_so(26) => SHIFT_12_26_port, 
                           A_so(25) => SHIFT_12_25_port, A_so(24) => 
                           SHIFT_12_24_port, A_so(23) => SHIFT_12_23_port, 
                           A_so(22) => SHIFT_12_22_port, A_so(21) => 
                           SHIFT_12_21_port, A_so(20) => SHIFT_12_20_port, 
                           A_so(19) => SHIFT_12_19_port, A_so(18) => 
                           SHIFT_12_18_port, A_so(17) => SHIFT_12_17_port, 
                           A_so(16) => SHIFT_12_16_port, A_so(15) => 
                           SHIFT_12_15_port, A_so(14) => SHIFT_12_14_port, 
                           A_so(13) => SHIFT_12_13_port, A_so(12) => 
                           SHIFT_12_12_port, A_so(11) => SHIFT_12_11_port, 
                           A_so(10) => SHIFT_12_10_port, A_so(9) => 
                           SHIFT_12_9_port, A_so(8) => SHIFT_12_8_port, A_so(7)
                           => SHIFT_12_7_port, A_so(6) => SHIFT_12_6_port, 
                           A_so(5) => SHIFT_12_5_port, A_so(4) => 
                           SHIFT_12_4_port, A_so(3) => SHIFT_12_3_port, A_so(2)
                           => SHIFT_12_2_port, A_so(1) => n_1133, A_so(0) => 
                           n_1134, A_nso(55) => SHIFT_n_12_55_port, A_nso(54) 
                           => SHIFT_n_12_54_port, A_nso(53) => 
                           SHIFT_n_12_53_port, A_nso(52) => SHIFT_n_12_52_port,
                           A_nso(51) => SHIFT_n_12_51_port, A_nso(50) => 
                           SHIFT_n_12_50_port, A_nso(49) => SHIFT_n_12_49_port,
                           A_nso(48) => SHIFT_n_12_48_port, A_nso(47) => 
                           SHIFT_n_12_47_port, A_nso(46) => SHIFT_n_12_46_port,
                           A_nso(45) => SHIFT_n_12_45_port, A_nso(44) => 
                           SHIFT_n_12_44_port, A_nso(43) => SHIFT_n_12_43_port,
                           A_nso(42) => SHIFT_n_12_42_port, A_nso(41) => 
                           SHIFT_n_12_41_port, A_nso(40) => SHIFT_n_12_40_port,
                           A_nso(39) => SHIFT_n_12_39_port, A_nso(38) => 
                           SHIFT_n_12_38_port, A_nso(37) => SHIFT_n_12_37_port,
                           A_nso(36) => SHIFT_n_12_36_port, A_nso(35) => 
                           SHIFT_n_12_35_port, A_nso(34) => SHIFT_n_12_34_port,
                           A_nso(33) => SHIFT_n_12_33_port, A_nso(32) => 
                           SHIFT_n_12_32_port, A_nso(31) => SHIFT_n_12_31_port,
                           A_nso(30) => SHIFT_n_12_30_port, A_nso(29) => 
                           SHIFT_n_12_29_port, A_nso(28) => SHIFT_n_12_28_port,
                           A_nso(27) => SHIFT_n_12_27_port, A_nso(26) => 
                           SHIFT_n_12_26_port, A_nso(25) => SHIFT_n_12_25_port,
                           A_nso(24) => SHIFT_n_12_24_port, A_nso(23) => 
                           SHIFT_n_12_23_port, A_nso(22) => SHIFT_n_12_22_port,
                           A_nso(21) => SHIFT_n_12_21_port, A_nso(20) => 
                           SHIFT_n_12_20_port, A_nso(19) => SHIFT_n_12_19_port,
                           A_nso(18) => SHIFT_n_12_18_port, A_nso(17) => 
                           SHIFT_n_12_17_port, A_nso(16) => SHIFT_n_12_16_port,
                           A_nso(15) => SHIFT_n_12_15_port, A_nso(14) => 
                           SHIFT_n_12_14_port, A_nso(13) => SHIFT_n_12_13_port,
                           A_nso(12) => SHIFT_n_12_12_port, A_nso(11) => 
                           SHIFT_n_12_11_port, A_nso(10) => SHIFT_n_12_10_port,
                           A_nso(9) => SHIFT_n_12_9_port, A_nso(8) => 
                           SHIFT_n_12_8_port, A_nso(7) => SHIFT_n_12_7_port, 
                           A_nso(6) => SHIFT_n_12_6_port, A_nso(5) => 
                           SHIFT_n_12_5_port, A_nso(4) => SHIFT_n_12_4_port, 
                           A_nso(3) => SHIFT_n_12_3_port, A_nso(2) => 
                           SHIFT_n_12_2_port, A_nso(1) => n_1135, A_nso(0) => 
                           n_1136);
   ENC_12 : BOOTHENC_NBIT58_i24 port map( A_s(57) => SHIFT_12_55_port, A_s(56) 
                           => SHIFT_12_55_port, A_s(55) => SHIFT_12_55_port, 
                           A_s(54) => SHIFT_12_54_port, A_s(53) => 
                           SHIFT_12_53_port, A_s(52) => SHIFT_12_52_port, 
                           A_s(51) => SHIFT_12_51_port, A_s(50) => 
                           SHIFT_12_50_port, A_s(49) => SHIFT_12_49_port, 
                           A_s(48) => SHIFT_12_48_port, A_s(47) => 
                           SHIFT_12_47_port, A_s(46) => SHIFT_12_46_port, 
                           A_s(45) => SHIFT_12_45_port, A_s(44) => 
                           SHIFT_12_44_port, A_s(43) => SHIFT_12_43_port, 
                           A_s(42) => SHIFT_12_42_port, A_s(41) => 
                           SHIFT_12_41_port, A_s(40) => SHIFT_12_40_port, 
                           A_s(39) => SHIFT_12_39_port, A_s(38) => 
                           SHIFT_12_38_port, A_s(37) => SHIFT_12_37_port, 
                           A_s(36) => SHIFT_12_36_port, A_s(35) => 
                           SHIFT_12_35_port, A_s(34) => SHIFT_12_34_port, 
                           A_s(33) => SHIFT_12_33_port, A_s(32) => 
                           SHIFT_12_32_port, A_s(31) => SHIFT_12_31_port, 
                           A_s(30) => SHIFT_12_30_port, A_s(29) => 
                           SHIFT_12_29_port, A_s(28) => SHIFT_12_28_port, 
                           A_s(27) => SHIFT_12_27_port, A_s(26) => 
                           SHIFT_12_26_port, A_s(25) => SHIFT_12_25_port, 
                           A_s(24) => SHIFT_12_24_port, A_s(23) => 
                           SHIFT_12_23_port, A_s(22) => SHIFT_12_22_port, 
                           A_s(21) => SHIFT_12_21_port, A_s(20) => 
                           SHIFT_12_20_port, A_s(19) => SHIFT_12_19_port, 
                           A_s(18) => SHIFT_12_18_port, A_s(17) => 
                           SHIFT_12_17_port, A_s(16) => SHIFT_12_16_port, 
                           A_s(15) => SHIFT_12_15_port, A_s(14) => 
                           SHIFT_12_14_port, A_s(13) => SHIFT_12_13_port, 
                           A_s(12) => SHIFT_12_12_port, A_s(11) => 
                           SHIFT_12_11_port, A_s(10) => SHIFT_12_10_port, 
                           A_s(9) => SHIFT_12_9_port, A_s(8) => SHIFT_12_8_port
                           , A_s(7) => SHIFT_12_7_port, A_s(6) => 
                           SHIFT_12_6_port, A_s(5) => SHIFT_12_5_port, A_s(4) 
                           => SHIFT_12_4_port, A_s(3) => SHIFT_12_3_port, 
                           A_s(2) => SHIFT_12_2_port, A_s(1) => SHIFT_12_1_port
                           , A_s(0) => SHIFT_12_0_port, A_ns(57) => 
                           SHIFT_n_12_55_port, A_ns(56) => SHIFT_n_12_55_port, 
                           A_ns(55) => SHIFT_n_12_55_port, A_ns(54) => 
                           SHIFT_n_12_54_port, A_ns(53) => SHIFT_n_12_53_port, 
                           A_ns(52) => SHIFT_n_12_52_port, A_ns(51) => 
                           SHIFT_n_12_51_port, A_ns(50) => SHIFT_n_12_50_port, 
                           A_ns(49) => SHIFT_n_12_49_port, A_ns(48) => 
                           SHIFT_n_12_48_port, A_ns(47) => SHIFT_n_12_47_port, 
                           A_ns(46) => SHIFT_n_12_46_port, A_ns(45) => 
                           SHIFT_n_12_45_port, A_ns(44) => SHIFT_n_12_44_port, 
                           A_ns(43) => SHIFT_n_12_43_port, A_ns(42) => 
                           SHIFT_n_12_42_port, A_ns(41) => SHIFT_n_12_41_port, 
                           A_ns(40) => SHIFT_n_12_40_port, A_ns(39) => 
                           SHIFT_n_12_39_port, A_ns(38) => SHIFT_n_12_38_port, 
                           A_ns(37) => SHIFT_n_12_37_port, A_ns(36) => 
                           SHIFT_n_12_36_port, A_ns(35) => SHIFT_n_12_35_port, 
                           A_ns(34) => SHIFT_n_12_34_port, A_ns(33) => 
                           SHIFT_n_12_33_port, A_ns(32) => SHIFT_n_12_32_port, 
                           A_ns(31) => SHIFT_n_12_31_port, A_ns(30) => 
                           SHIFT_n_12_30_port, A_ns(29) => SHIFT_n_12_29_port, 
                           A_ns(28) => SHIFT_n_12_28_port, A_ns(27) => 
                           SHIFT_n_12_27_port, A_ns(26) => SHIFT_n_12_26_port, 
                           A_ns(25) => SHIFT_n_12_25_port, A_ns(24) => 
                           SHIFT_n_12_24_port, A_ns(23) => SHIFT_n_12_23_port, 
                           A_ns(22) => SHIFT_n_12_22_port, A_ns(21) => 
                           SHIFT_n_12_21_port, A_ns(20) => SHIFT_n_12_20_port, 
                           A_ns(19) => SHIFT_n_12_19_port, A_ns(18) => 
                           SHIFT_n_12_18_port, A_ns(17) => SHIFT_n_12_17_port, 
                           A_ns(16) => SHIFT_n_12_16_port, A_ns(15) => 
                           SHIFT_n_12_15_port, A_ns(14) => SHIFT_n_12_14_port, 
                           A_ns(13) => SHIFT_n_12_13_port, A_ns(12) => 
                           SHIFT_n_12_12_port, A_ns(11) => SHIFT_n_12_11_port, 
                           A_ns(10) => SHIFT_n_12_10_port, A_ns(9) => 
                           SHIFT_n_12_9_port, A_ns(8) => SHIFT_n_12_8_port, 
                           A_ns(7) => SHIFT_n_12_7_port, A_ns(6) => 
                           SHIFT_n_12_6_port, A_ns(5) => SHIFT_n_12_5_port, 
                           A_ns(4) => SHIFT_n_12_4_port, A_ns(3) => 
                           SHIFT_n_12_3_port, A_ns(2) => SHIFT_n_12_2_port, 
                           A_ns(1) => SHIFT_n_12_1_port, A_ns(0) => 
                           SHIFT_n_12_0_port, B(57) => B(31), B(56) => B(31), 
                           B(55) => B(31), B(54) => B(31), B(53) => B(31), 
                           B(52) => B(31), B(51) => B(31), B(50) => B(31), 
                           B(49) => B(31), B(48) => B(31), B(47) => B(31), 
                           B(46) => B(31), B(45) => B(31), B(44) => B(31), 
                           B(43) => B(31), B(42) => B(31), B(41) => B(31), 
                           B(40) => B(31), B(39) => B(31), B(38) => B(31), 
                           B(37) => B(31), B(36) => B(31), B(35) => B(31), 
                           B(34) => B(31), B(33) => B(31), B(32) => B(31), 
                           B(31) => B(31), B(30) => B(30), B(29) => B(29), 
                           B(28) => B(28), B(27) => B(27), B(26) => B(26), 
                           B(25) => B(25), B(24) => B(24), B(23) => B(23), 
                           B(22) => B(22), B(21) => B(21), B(20) => B(20), 
                           B(19) => B(19), B(18) => B(18), B(17) => B(17), 
                           B(16) => B(16), B(15) => B(15), B(14) => B(14), 
                           B(13) => B(13), B(12) => B(12), B(11) => B(11), 
                           B(10) => B(10), B(9) => B(9), B(8) => B(8), B(7) => 
                           B(7), B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3)
                           => B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), 
                           O(57) => OTMP_12_57_port, O(56) => OTMP_12_56_port, 
                           O(55) => OTMP_12_55_port, O(54) => OTMP_12_54_port, 
                           O(53) => OTMP_12_53_port, O(52) => OTMP_12_52_port, 
                           O(51) => OTMP_12_51_port, O(50) => OTMP_12_50_port, 
                           O(49) => OTMP_12_49_port, O(48) => OTMP_12_48_port, 
                           O(47) => OTMP_12_47_port, O(46) => OTMP_12_46_port, 
                           O(45) => OTMP_12_45_port, O(44) => OTMP_12_44_port, 
                           O(43) => OTMP_12_43_port, O(42) => OTMP_12_42_port, 
                           O(41) => OTMP_12_41_port, O(40) => OTMP_12_40_port, 
                           O(39) => OTMP_12_39_port, O(38) => OTMP_12_38_port, 
                           O(37) => OTMP_12_37_port, O(36) => OTMP_12_36_port, 
                           O(35) => OTMP_12_35_port, O(34) => OTMP_12_34_port, 
                           O(33) => OTMP_12_33_port, O(32) => OTMP_12_32_port, 
                           O(31) => OTMP_12_31_port, O(30) => OTMP_12_30_port, 
                           O(29) => OTMP_12_29_port, O(28) => OTMP_12_28_port, 
                           O(27) => OTMP_12_27_port, O(26) => OTMP_12_26_port, 
                           O(25) => OTMP_12_25_port, O(24) => OTMP_12_24_port, 
                           O(23) => OTMP_12_23_port, O(22) => OTMP_12_22_port, 
                           O(21) => OTMP_12_21_port, O(20) => OTMP_12_20_port, 
                           O(19) => OTMP_12_19_port, O(18) => OTMP_12_18_port, 
                           O(17) => OTMP_12_17_port, O(16) => OTMP_12_16_port, 
                           O(15) => OTMP_12_15_port, O(14) => OTMP_12_14_port, 
                           O(13) => OTMP_12_13_port, O(12) => OTMP_12_12_port, 
                           O(11) => OTMP_12_11_port, O(10) => OTMP_12_10_port, 
                           O(9) => OTMP_12_9_port, O(8) => OTMP_12_8_port, O(7)
                           => OTMP_12_7_port, O(6) => OTMP_12_6_port, O(5) => 
                           OTMP_12_5_port, O(4) => OTMP_12_4_port, O(3) => 
                           OTMP_12_3_port, O(2) => OTMP_12_2_port, O(1) => 
                           OTMP_12_1_port, O(0) => n_1137, A_so(57) => 
                           SHIFT_13_57_port, A_so(56) => SHIFT_13_56_port, 
                           A_so(55) => SHIFT_13_55_port, A_so(54) => 
                           SHIFT_13_54_port, A_so(53) => SHIFT_13_53_port, 
                           A_so(52) => SHIFT_13_52_port, A_so(51) => 
                           SHIFT_13_51_port, A_so(50) => SHIFT_13_50_port, 
                           A_so(49) => SHIFT_13_49_port, A_so(48) => 
                           SHIFT_13_48_port, A_so(47) => SHIFT_13_47_port, 
                           A_so(46) => SHIFT_13_46_port, A_so(45) => 
                           SHIFT_13_45_port, A_so(44) => SHIFT_13_44_port, 
                           A_so(43) => SHIFT_13_43_port, A_so(42) => 
                           SHIFT_13_42_port, A_so(41) => SHIFT_13_41_port, 
                           A_so(40) => SHIFT_13_40_port, A_so(39) => 
                           SHIFT_13_39_port, A_so(38) => SHIFT_13_38_port, 
                           A_so(37) => SHIFT_13_37_port, A_so(36) => 
                           SHIFT_13_36_port, A_so(35) => SHIFT_13_35_port, 
                           A_so(34) => SHIFT_13_34_port, A_so(33) => 
                           SHIFT_13_33_port, A_so(32) => SHIFT_13_32_port, 
                           A_so(31) => SHIFT_13_31_port, A_so(30) => 
                           SHIFT_13_30_port, A_so(29) => SHIFT_13_29_port, 
                           A_so(28) => SHIFT_13_28_port, A_so(27) => 
                           SHIFT_13_27_port, A_so(26) => SHIFT_13_26_port, 
                           A_so(25) => SHIFT_13_25_port, A_so(24) => 
                           SHIFT_13_24_port, A_so(23) => SHIFT_13_23_port, 
                           A_so(22) => SHIFT_13_22_port, A_so(21) => 
                           SHIFT_13_21_port, A_so(20) => SHIFT_13_20_port, 
                           A_so(19) => SHIFT_13_19_port, A_so(18) => 
                           SHIFT_13_18_port, A_so(17) => SHIFT_13_17_port, 
                           A_so(16) => SHIFT_13_16_port, A_so(15) => 
                           SHIFT_13_15_port, A_so(14) => SHIFT_13_14_port, 
                           A_so(13) => SHIFT_13_13_port, A_so(12) => 
                           SHIFT_13_12_port, A_so(11) => SHIFT_13_11_port, 
                           A_so(10) => SHIFT_13_10_port, A_so(9) => 
                           SHIFT_13_9_port, A_so(8) => SHIFT_13_8_port, A_so(7)
                           => SHIFT_13_7_port, A_so(6) => SHIFT_13_6_port, 
                           A_so(5) => SHIFT_13_5_port, A_so(4) => 
                           SHIFT_13_4_port, A_so(3) => SHIFT_13_3_port, A_so(2)
                           => SHIFT_13_2_port, A_so(1) => n_1138, A_so(0) => 
                           n_1139, A_nso(57) => SHIFT_n_13_57_port, A_nso(56) 
                           => SHIFT_n_13_56_port, A_nso(55) => 
                           SHIFT_n_13_55_port, A_nso(54) => SHIFT_n_13_54_port,
                           A_nso(53) => SHIFT_n_13_53_port, A_nso(52) => 
                           SHIFT_n_13_52_port, A_nso(51) => SHIFT_n_13_51_port,
                           A_nso(50) => SHIFT_n_13_50_port, A_nso(49) => 
                           SHIFT_n_13_49_port, A_nso(48) => SHIFT_n_13_48_port,
                           A_nso(47) => SHIFT_n_13_47_port, A_nso(46) => 
                           SHIFT_n_13_46_port, A_nso(45) => SHIFT_n_13_45_port,
                           A_nso(44) => SHIFT_n_13_44_port, A_nso(43) => 
                           SHIFT_n_13_43_port, A_nso(42) => SHIFT_n_13_42_port,
                           A_nso(41) => SHIFT_n_13_41_port, A_nso(40) => 
                           SHIFT_n_13_40_port, A_nso(39) => SHIFT_n_13_39_port,
                           A_nso(38) => SHIFT_n_13_38_port, A_nso(37) => 
                           SHIFT_n_13_37_port, A_nso(36) => SHIFT_n_13_36_port,
                           A_nso(35) => SHIFT_n_13_35_port, A_nso(34) => 
                           SHIFT_n_13_34_port, A_nso(33) => SHIFT_n_13_33_port,
                           A_nso(32) => SHIFT_n_13_32_port, A_nso(31) => 
                           SHIFT_n_13_31_port, A_nso(30) => SHIFT_n_13_30_port,
                           A_nso(29) => SHIFT_n_13_29_port, A_nso(28) => 
                           SHIFT_n_13_28_port, A_nso(27) => SHIFT_n_13_27_port,
                           A_nso(26) => SHIFT_n_13_26_port, A_nso(25) => 
                           SHIFT_n_13_25_port, A_nso(24) => SHIFT_n_13_24_port,
                           A_nso(23) => SHIFT_n_13_23_port, A_nso(22) => 
                           SHIFT_n_13_22_port, A_nso(21) => SHIFT_n_13_21_port,
                           A_nso(20) => SHIFT_n_13_20_port, A_nso(19) => 
                           SHIFT_n_13_19_port, A_nso(18) => SHIFT_n_13_18_port,
                           A_nso(17) => SHIFT_n_13_17_port, A_nso(16) => 
                           SHIFT_n_13_16_port, A_nso(15) => SHIFT_n_13_15_port,
                           A_nso(14) => SHIFT_n_13_14_port, A_nso(13) => 
                           SHIFT_n_13_13_port, A_nso(12) => SHIFT_n_13_12_port,
                           A_nso(11) => SHIFT_n_13_11_port, A_nso(10) => 
                           SHIFT_n_13_10_port, A_nso(9) => SHIFT_n_13_9_port, 
                           A_nso(8) => SHIFT_n_13_8_port, A_nso(7) => 
                           SHIFT_n_13_7_port, A_nso(6) => SHIFT_n_13_6_port, 
                           A_nso(5) => SHIFT_n_13_5_port, A_nso(4) => 
                           SHIFT_n_13_4_port, A_nso(3) => SHIFT_n_13_3_port, 
                           A_nso(2) => SHIFT_n_13_2_port, A_nso(1) => n_1140, 
                           A_nso(0) => n_1141);
   ENC_13 : BOOTHENC_NBIT60_i26 port map( A_s(59) => SHIFT_13_57_port, A_s(58) 
                           => SHIFT_13_57_port, A_s(57) => SHIFT_13_57_port, 
                           A_s(56) => SHIFT_13_56_port, A_s(55) => 
                           SHIFT_13_55_port, A_s(54) => SHIFT_13_54_port, 
                           A_s(53) => SHIFT_13_53_port, A_s(52) => 
                           SHIFT_13_52_port, A_s(51) => SHIFT_13_51_port, 
                           A_s(50) => SHIFT_13_50_port, A_s(49) => 
                           SHIFT_13_49_port, A_s(48) => SHIFT_13_48_port, 
                           A_s(47) => SHIFT_13_47_port, A_s(46) => 
                           SHIFT_13_46_port, A_s(45) => SHIFT_13_45_port, 
                           A_s(44) => SHIFT_13_44_port, A_s(43) => 
                           SHIFT_13_43_port, A_s(42) => SHIFT_13_42_port, 
                           A_s(41) => SHIFT_13_41_port, A_s(40) => 
                           SHIFT_13_40_port, A_s(39) => SHIFT_13_39_port, 
                           A_s(38) => SHIFT_13_38_port, A_s(37) => 
                           SHIFT_13_37_port, A_s(36) => SHIFT_13_36_port, 
                           A_s(35) => SHIFT_13_35_port, A_s(34) => 
                           SHIFT_13_34_port, A_s(33) => SHIFT_13_33_port, 
                           A_s(32) => SHIFT_13_32_port, A_s(31) => 
                           SHIFT_13_31_port, A_s(30) => SHIFT_13_30_port, 
                           A_s(29) => SHIFT_13_29_port, A_s(28) => 
                           SHIFT_13_28_port, A_s(27) => SHIFT_13_27_port, 
                           A_s(26) => SHIFT_13_26_port, A_s(25) => 
                           SHIFT_13_25_port, A_s(24) => SHIFT_13_24_port, 
                           A_s(23) => SHIFT_13_23_port, A_s(22) => 
                           SHIFT_13_22_port, A_s(21) => SHIFT_13_21_port, 
                           A_s(20) => SHIFT_13_20_port, A_s(19) => 
                           SHIFT_13_19_port, A_s(18) => SHIFT_13_18_port, 
                           A_s(17) => SHIFT_13_17_port, A_s(16) => 
                           SHIFT_13_16_port, A_s(15) => SHIFT_13_15_port, 
                           A_s(14) => SHIFT_13_14_port, A_s(13) => 
                           SHIFT_13_13_port, A_s(12) => SHIFT_13_12_port, 
                           A_s(11) => SHIFT_13_11_port, A_s(10) => 
                           SHIFT_13_10_port, A_s(9) => SHIFT_13_9_port, A_s(8) 
                           => SHIFT_13_8_port, A_s(7) => SHIFT_13_7_port, 
                           A_s(6) => SHIFT_13_6_port, A_s(5) => SHIFT_13_5_port
                           , A_s(4) => SHIFT_13_4_port, A_s(3) => 
                           SHIFT_13_3_port, A_s(2) => SHIFT_13_2_port, A_s(1) 
                           => SHIFT_13_1_port, A_s(0) => SHIFT_13_0_port, 
                           A_ns(59) => SHIFT_n_13_57_port, A_ns(58) => 
                           SHIFT_n_13_57_port, A_ns(57) => SHIFT_n_13_57_port, 
                           A_ns(56) => SHIFT_n_13_56_port, A_ns(55) => 
                           SHIFT_n_13_55_port, A_ns(54) => SHIFT_n_13_54_port, 
                           A_ns(53) => SHIFT_n_13_53_port, A_ns(52) => 
                           SHIFT_n_13_52_port, A_ns(51) => SHIFT_n_13_51_port, 
                           A_ns(50) => SHIFT_n_13_50_port, A_ns(49) => 
                           SHIFT_n_13_49_port, A_ns(48) => SHIFT_n_13_48_port, 
                           A_ns(47) => SHIFT_n_13_47_port, A_ns(46) => 
                           SHIFT_n_13_46_port, A_ns(45) => SHIFT_n_13_45_port, 
                           A_ns(44) => SHIFT_n_13_44_port, A_ns(43) => 
                           SHIFT_n_13_43_port, A_ns(42) => SHIFT_n_13_42_port, 
                           A_ns(41) => SHIFT_n_13_41_port, A_ns(40) => 
                           SHIFT_n_13_40_port, A_ns(39) => SHIFT_n_13_39_port, 
                           A_ns(38) => SHIFT_n_13_38_port, A_ns(37) => 
                           SHIFT_n_13_37_port, A_ns(36) => SHIFT_n_13_36_port, 
                           A_ns(35) => SHIFT_n_13_35_port, A_ns(34) => 
                           SHIFT_n_13_34_port, A_ns(33) => SHIFT_n_13_33_port, 
                           A_ns(32) => SHIFT_n_13_32_port, A_ns(31) => 
                           SHIFT_n_13_31_port, A_ns(30) => SHIFT_n_13_30_port, 
                           A_ns(29) => SHIFT_n_13_29_port, A_ns(28) => 
                           SHIFT_n_13_28_port, A_ns(27) => SHIFT_n_13_27_port, 
                           A_ns(26) => SHIFT_n_13_26_port, A_ns(25) => 
                           SHIFT_n_13_25_port, A_ns(24) => SHIFT_n_13_24_port, 
                           A_ns(23) => SHIFT_n_13_23_port, A_ns(22) => 
                           SHIFT_n_13_22_port, A_ns(21) => SHIFT_n_13_21_port, 
                           A_ns(20) => SHIFT_n_13_20_port, A_ns(19) => 
                           SHIFT_n_13_19_port, A_ns(18) => SHIFT_n_13_18_port, 
                           A_ns(17) => SHIFT_n_13_17_port, A_ns(16) => 
                           SHIFT_n_13_16_port, A_ns(15) => SHIFT_n_13_15_port, 
                           A_ns(14) => SHIFT_n_13_14_port, A_ns(13) => 
                           SHIFT_n_13_13_port, A_ns(12) => SHIFT_n_13_12_port, 
                           A_ns(11) => SHIFT_n_13_11_port, A_ns(10) => 
                           SHIFT_n_13_10_port, A_ns(9) => SHIFT_n_13_9_port, 
                           A_ns(8) => SHIFT_n_13_8_port, A_ns(7) => 
                           SHIFT_n_13_7_port, A_ns(6) => SHIFT_n_13_6_port, 
                           A_ns(5) => SHIFT_n_13_5_port, A_ns(4) => 
                           SHIFT_n_13_4_port, A_ns(3) => SHIFT_n_13_3_port, 
                           A_ns(2) => SHIFT_n_13_2_port, A_ns(1) => 
                           SHIFT_n_13_1_port, A_ns(0) => SHIFT_n_13_0_port, 
                           B(59) => B(31), B(58) => B(31), B(57) => B(31), 
                           B(56) => B(31), B(55) => B(31), B(54) => B(31), 
                           B(53) => B(31), B(52) => B(31), B(51) => B(31), 
                           B(50) => B(31), B(49) => B(31), B(48) => B(31), 
                           B(47) => B(31), B(46) => B(31), B(45) => B(31), 
                           B(44) => B(31), B(43) => B(31), B(42) => B(31), 
                           B(41) => B(31), B(40) => B(31), B(39) => B(31), 
                           B(38) => B(31), B(37) => B(31), B(36) => B(31), 
                           B(35) => B(31), B(34) => B(31), B(33) => B(31), 
                           B(32) => B(31), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), O(59) => OTMP_13_59_port, O(58) 
                           => OTMP_13_58_port, O(57) => OTMP_13_57_port, O(56) 
                           => OTMP_13_56_port, O(55) => OTMP_13_55_port, O(54) 
                           => OTMP_13_54_port, O(53) => OTMP_13_53_port, O(52) 
                           => OTMP_13_52_port, O(51) => OTMP_13_51_port, O(50) 
                           => OTMP_13_50_port, O(49) => OTMP_13_49_port, O(48) 
                           => OTMP_13_48_port, O(47) => OTMP_13_47_port, O(46) 
                           => OTMP_13_46_port, O(45) => OTMP_13_45_port, O(44) 
                           => OTMP_13_44_port, O(43) => OTMP_13_43_port, O(42) 
                           => OTMP_13_42_port, O(41) => OTMP_13_41_port, O(40) 
                           => OTMP_13_40_port, O(39) => OTMP_13_39_port, O(38) 
                           => OTMP_13_38_port, O(37) => OTMP_13_37_port, O(36) 
                           => OTMP_13_36_port, O(35) => OTMP_13_35_port, O(34) 
                           => OTMP_13_34_port, O(33) => OTMP_13_33_port, O(32) 
                           => OTMP_13_32_port, O(31) => OTMP_13_31_port, O(30) 
                           => OTMP_13_30_port, O(29) => OTMP_13_29_port, O(28) 
                           => OTMP_13_28_port, O(27) => OTMP_13_27_port, O(26) 
                           => OTMP_13_26_port, O(25) => OTMP_13_25_port, O(24) 
                           => OTMP_13_24_port, O(23) => OTMP_13_23_port, O(22) 
                           => OTMP_13_22_port, O(21) => OTMP_13_21_port, O(20) 
                           => OTMP_13_20_port, O(19) => OTMP_13_19_port, O(18) 
                           => OTMP_13_18_port, O(17) => OTMP_13_17_port, O(16) 
                           => OTMP_13_16_port, O(15) => OTMP_13_15_port, O(14) 
                           => OTMP_13_14_port, O(13) => OTMP_13_13_port, O(12) 
                           => OTMP_13_12_port, O(11) => OTMP_13_11_port, O(10) 
                           => OTMP_13_10_port, O(9) => OTMP_13_9_port, O(8) => 
                           OTMP_13_8_port, O(7) => OTMP_13_7_port, O(6) => 
                           OTMP_13_6_port, O(5) => OTMP_13_5_port, O(4) => 
                           OTMP_13_4_port, O(3) => OTMP_13_3_port, O(2) => 
                           OTMP_13_2_port, O(1) => OTMP_13_1_port, O(0) => 
                           n_1142, A_so(59) => SHIFT_14_59_port, A_so(58) => 
                           SHIFT_14_58_port, A_so(57) => SHIFT_14_57_port, 
                           A_so(56) => SHIFT_14_56_port, A_so(55) => 
                           SHIFT_14_55_port, A_so(54) => SHIFT_14_54_port, 
                           A_so(53) => SHIFT_14_53_port, A_so(52) => 
                           SHIFT_14_52_port, A_so(51) => SHIFT_14_51_port, 
                           A_so(50) => SHIFT_14_50_port, A_so(49) => 
                           SHIFT_14_49_port, A_so(48) => SHIFT_14_48_port, 
                           A_so(47) => SHIFT_14_47_port, A_so(46) => 
                           SHIFT_14_46_port, A_so(45) => SHIFT_14_45_port, 
                           A_so(44) => SHIFT_14_44_port, A_so(43) => 
                           SHIFT_14_43_port, A_so(42) => SHIFT_14_42_port, 
                           A_so(41) => SHIFT_14_41_port, A_so(40) => 
                           SHIFT_14_40_port, A_so(39) => SHIFT_14_39_port, 
                           A_so(38) => SHIFT_14_38_port, A_so(37) => 
                           SHIFT_14_37_port, A_so(36) => SHIFT_14_36_port, 
                           A_so(35) => SHIFT_14_35_port, A_so(34) => 
                           SHIFT_14_34_port, A_so(33) => SHIFT_14_33_port, 
                           A_so(32) => SHIFT_14_32_port, A_so(31) => 
                           SHIFT_14_31_port, A_so(30) => SHIFT_14_30_port, 
                           A_so(29) => SHIFT_14_29_port, A_so(28) => 
                           SHIFT_14_28_port, A_so(27) => SHIFT_14_27_port, 
                           A_so(26) => SHIFT_14_26_port, A_so(25) => 
                           SHIFT_14_25_port, A_so(24) => SHIFT_14_24_port, 
                           A_so(23) => SHIFT_14_23_port, A_so(22) => 
                           SHIFT_14_22_port, A_so(21) => SHIFT_14_21_port, 
                           A_so(20) => SHIFT_14_20_port, A_so(19) => 
                           SHIFT_14_19_port, A_so(18) => SHIFT_14_18_port, 
                           A_so(17) => SHIFT_14_17_port, A_so(16) => 
                           SHIFT_14_16_port, A_so(15) => SHIFT_14_15_port, 
                           A_so(14) => SHIFT_14_14_port, A_so(13) => 
                           SHIFT_14_13_port, A_so(12) => SHIFT_14_12_port, 
                           A_so(11) => SHIFT_14_11_port, A_so(10) => 
                           SHIFT_14_10_port, A_so(9) => SHIFT_14_9_port, 
                           A_so(8) => SHIFT_14_8_port, A_so(7) => 
                           SHIFT_14_7_port, A_so(6) => SHIFT_14_6_port, A_so(5)
                           => SHIFT_14_5_port, A_so(4) => SHIFT_14_4_port, 
                           A_so(3) => SHIFT_14_3_port, A_so(2) => 
                           SHIFT_14_2_port, A_so(1) => n_1143, A_so(0) => 
                           n_1144, A_nso(59) => SHIFT_n_14_59_port, A_nso(58) 
                           => SHIFT_n_14_58_port, A_nso(57) => 
                           SHIFT_n_14_57_port, A_nso(56) => SHIFT_n_14_56_port,
                           A_nso(55) => SHIFT_n_14_55_port, A_nso(54) => 
                           SHIFT_n_14_54_port, A_nso(53) => SHIFT_n_14_53_port,
                           A_nso(52) => SHIFT_n_14_52_port, A_nso(51) => 
                           SHIFT_n_14_51_port, A_nso(50) => SHIFT_n_14_50_port,
                           A_nso(49) => SHIFT_n_14_49_port, A_nso(48) => 
                           SHIFT_n_14_48_port, A_nso(47) => SHIFT_n_14_47_port,
                           A_nso(46) => SHIFT_n_14_46_port, A_nso(45) => 
                           SHIFT_n_14_45_port, A_nso(44) => SHIFT_n_14_44_port,
                           A_nso(43) => SHIFT_n_14_43_port, A_nso(42) => 
                           SHIFT_n_14_42_port, A_nso(41) => SHIFT_n_14_41_port,
                           A_nso(40) => SHIFT_n_14_40_port, A_nso(39) => 
                           SHIFT_n_14_39_port, A_nso(38) => SHIFT_n_14_38_port,
                           A_nso(37) => SHIFT_n_14_37_port, A_nso(36) => 
                           SHIFT_n_14_36_port, A_nso(35) => SHIFT_n_14_35_port,
                           A_nso(34) => SHIFT_n_14_34_port, A_nso(33) => 
                           SHIFT_n_14_33_port, A_nso(32) => SHIFT_n_14_32_port,
                           A_nso(31) => SHIFT_n_14_31_port, A_nso(30) => 
                           SHIFT_n_14_30_port, A_nso(29) => SHIFT_n_14_29_port,
                           A_nso(28) => SHIFT_n_14_28_port, A_nso(27) => 
                           SHIFT_n_14_27_port, A_nso(26) => SHIFT_n_14_26_port,
                           A_nso(25) => SHIFT_n_14_25_port, A_nso(24) => 
                           SHIFT_n_14_24_port, A_nso(23) => SHIFT_n_14_23_port,
                           A_nso(22) => SHIFT_n_14_22_port, A_nso(21) => 
                           SHIFT_n_14_21_port, A_nso(20) => SHIFT_n_14_20_port,
                           A_nso(19) => SHIFT_n_14_19_port, A_nso(18) => 
                           SHIFT_n_14_18_port, A_nso(17) => SHIFT_n_14_17_port,
                           A_nso(16) => SHIFT_n_14_16_port, A_nso(15) => 
                           SHIFT_n_14_15_port, A_nso(14) => SHIFT_n_14_14_port,
                           A_nso(13) => SHIFT_n_14_13_port, A_nso(12) => 
                           SHIFT_n_14_12_port, A_nso(11) => SHIFT_n_14_11_port,
                           A_nso(10) => SHIFT_n_14_10_port, A_nso(9) => 
                           SHIFT_n_14_9_port, A_nso(8) => SHIFT_n_14_8_port, 
                           A_nso(7) => SHIFT_n_14_7_port, A_nso(6) => 
                           SHIFT_n_14_6_port, A_nso(5) => SHIFT_n_14_5_port, 
                           A_nso(4) => SHIFT_n_14_4_port, A_nso(3) => 
                           SHIFT_n_14_3_port, A_nso(2) => SHIFT_n_14_2_port, 
                           A_nso(1) => n_1145, A_nso(0) => n_1146);
   ENC_14 : BOOTHENC_NBIT62_i28 port map( A_s(61) => SHIFT_14_59_port, A_s(60) 
                           => SHIFT_14_59_port, A_s(59) => SHIFT_14_59_port, 
                           A_s(58) => SHIFT_14_58_port, A_s(57) => 
                           SHIFT_14_57_port, A_s(56) => SHIFT_14_56_port, 
                           A_s(55) => SHIFT_14_55_port, A_s(54) => 
                           SHIFT_14_54_port, A_s(53) => SHIFT_14_53_port, 
                           A_s(52) => SHIFT_14_52_port, A_s(51) => 
                           SHIFT_14_51_port, A_s(50) => SHIFT_14_50_port, 
                           A_s(49) => SHIFT_14_49_port, A_s(48) => 
                           SHIFT_14_48_port, A_s(47) => SHIFT_14_47_port, 
                           A_s(46) => SHIFT_14_46_port, A_s(45) => 
                           SHIFT_14_45_port, A_s(44) => SHIFT_14_44_port, 
                           A_s(43) => SHIFT_14_43_port, A_s(42) => 
                           SHIFT_14_42_port, A_s(41) => SHIFT_14_41_port, 
                           A_s(40) => SHIFT_14_40_port, A_s(39) => 
                           SHIFT_14_39_port, A_s(38) => SHIFT_14_38_port, 
                           A_s(37) => SHIFT_14_37_port, A_s(36) => 
                           SHIFT_14_36_port, A_s(35) => SHIFT_14_35_port, 
                           A_s(34) => SHIFT_14_34_port, A_s(33) => 
                           SHIFT_14_33_port, A_s(32) => SHIFT_14_32_port, 
                           A_s(31) => SHIFT_14_31_port, A_s(30) => 
                           SHIFT_14_30_port, A_s(29) => SHIFT_14_29_port, 
                           A_s(28) => SHIFT_14_28_port, A_s(27) => 
                           SHIFT_14_27_port, A_s(26) => SHIFT_14_26_port, 
                           A_s(25) => SHIFT_14_25_port, A_s(24) => 
                           SHIFT_14_24_port, A_s(23) => SHIFT_14_23_port, 
                           A_s(22) => SHIFT_14_22_port, A_s(21) => 
                           SHIFT_14_21_port, A_s(20) => SHIFT_14_20_port, 
                           A_s(19) => SHIFT_14_19_port, A_s(18) => 
                           SHIFT_14_18_port, A_s(17) => SHIFT_14_17_port, 
                           A_s(16) => SHIFT_14_16_port, A_s(15) => 
                           SHIFT_14_15_port, A_s(14) => SHIFT_14_14_port, 
                           A_s(13) => SHIFT_14_13_port, A_s(12) => 
                           SHIFT_14_12_port, A_s(11) => SHIFT_14_11_port, 
                           A_s(10) => SHIFT_14_10_port, A_s(9) => 
                           SHIFT_14_9_port, A_s(8) => SHIFT_14_8_port, A_s(7) 
                           => SHIFT_14_7_port, A_s(6) => SHIFT_14_6_port, 
                           A_s(5) => SHIFT_14_5_port, A_s(4) => SHIFT_14_4_port
                           , A_s(3) => SHIFT_14_3_port, A_s(2) => 
                           SHIFT_14_2_port, A_s(1) => SHIFT_14_1_port, A_s(0) 
                           => SHIFT_14_0_port, A_ns(61) => SHIFT_n_14_59_port, 
                           A_ns(60) => SHIFT_n_14_59_port, A_ns(59) => 
                           SHIFT_n_14_59_port, A_ns(58) => SHIFT_n_14_58_port, 
                           A_ns(57) => SHIFT_n_14_57_port, A_ns(56) => 
                           SHIFT_n_14_56_port, A_ns(55) => SHIFT_n_14_55_port, 
                           A_ns(54) => SHIFT_n_14_54_port, A_ns(53) => 
                           SHIFT_n_14_53_port, A_ns(52) => SHIFT_n_14_52_port, 
                           A_ns(51) => SHIFT_n_14_51_port, A_ns(50) => 
                           SHIFT_n_14_50_port, A_ns(49) => SHIFT_n_14_49_port, 
                           A_ns(48) => SHIFT_n_14_48_port, A_ns(47) => 
                           SHIFT_n_14_47_port, A_ns(46) => SHIFT_n_14_46_port, 
                           A_ns(45) => SHIFT_n_14_45_port, A_ns(44) => 
                           SHIFT_n_14_44_port, A_ns(43) => SHIFT_n_14_43_port, 
                           A_ns(42) => SHIFT_n_14_42_port, A_ns(41) => 
                           SHIFT_n_14_41_port, A_ns(40) => SHIFT_n_14_40_port, 
                           A_ns(39) => SHIFT_n_14_39_port, A_ns(38) => 
                           SHIFT_n_14_38_port, A_ns(37) => SHIFT_n_14_37_port, 
                           A_ns(36) => SHIFT_n_14_36_port, A_ns(35) => 
                           SHIFT_n_14_35_port, A_ns(34) => SHIFT_n_14_34_port, 
                           A_ns(33) => SHIFT_n_14_33_port, A_ns(32) => 
                           SHIFT_n_14_32_port, A_ns(31) => SHIFT_n_14_31_port, 
                           A_ns(30) => SHIFT_n_14_30_port, A_ns(29) => 
                           SHIFT_n_14_29_port, A_ns(28) => SHIFT_n_14_28_port, 
                           A_ns(27) => SHIFT_n_14_27_port, A_ns(26) => 
                           SHIFT_n_14_26_port, A_ns(25) => SHIFT_n_14_25_port, 
                           A_ns(24) => SHIFT_n_14_24_port, A_ns(23) => 
                           SHIFT_n_14_23_port, A_ns(22) => SHIFT_n_14_22_port, 
                           A_ns(21) => SHIFT_n_14_21_port, A_ns(20) => 
                           SHIFT_n_14_20_port, A_ns(19) => SHIFT_n_14_19_port, 
                           A_ns(18) => SHIFT_n_14_18_port, A_ns(17) => 
                           SHIFT_n_14_17_port, A_ns(16) => SHIFT_n_14_16_port, 
                           A_ns(15) => SHIFT_n_14_15_port, A_ns(14) => 
                           SHIFT_n_14_14_port, A_ns(13) => SHIFT_n_14_13_port, 
                           A_ns(12) => SHIFT_n_14_12_port, A_ns(11) => 
                           SHIFT_n_14_11_port, A_ns(10) => SHIFT_n_14_10_port, 
                           A_ns(9) => SHIFT_n_14_9_port, A_ns(8) => 
                           SHIFT_n_14_8_port, A_ns(7) => SHIFT_n_14_7_port, 
                           A_ns(6) => SHIFT_n_14_6_port, A_ns(5) => 
                           SHIFT_n_14_5_port, A_ns(4) => SHIFT_n_14_4_port, 
                           A_ns(3) => SHIFT_n_14_3_port, A_ns(2) => 
                           SHIFT_n_14_2_port, A_ns(1) => SHIFT_n_14_1_port, 
                           A_ns(0) => SHIFT_n_14_0_port, B(61) => B(31), B(60) 
                           => B(31), B(59) => B(31), B(58) => B(31), B(57) => 
                           B(31), B(56) => B(31), B(55) => B(31), B(54) => 
                           B(31), B(53) => B(31), B(52) => B(31), B(51) => 
                           B(31), B(50) => B(31), B(49) => B(31), B(48) => 
                           B(31), B(47) => B(31), B(46) => B(31), B(45) => 
                           B(31), B(44) => B(31), B(43) => B(31), B(42) => 
                           B(31), B(41) => B(31), B(40) => B(31), B(39) => 
                           B(31), B(38) => B(31), B(37) => B(31), B(36) => 
                           B(31), B(35) => B(31), B(34) => B(31), B(33) => 
                           B(31), B(32) => B(31), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), O(61) => OTMP_14_61_port, 
                           O(60) => OTMP_14_60_port, O(59) => OTMP_14_59_port, 
                           O(58) => OTMP_14_58_port, O(57) => OTMP_14_57_port, 
                           O(56) => OTMP_14_56_port, O(55) => OTMP_14_55_port, 
                           O(54) => OTMP_14_54_port, O(53) => OTMP_14_53_port, 
                           O(52) => OTMP_14_52_port, O(51) => OTMP_14_51_port, 
                           O(50) => OTMP_14_50_port, O(49) => OTMP_14_49_port, 
                           O(48) => OTMP_14_48_port, O(47) => OTMP_14_47_port, 
                           O(46) => OTMP_14_46_port, O(45) => OTMP_14_45_port, 
                           O(44) => OTMP_14_44_port, O(43) => OTMP_14_43_port, 
                           O(42) => OTMP_14_42_port, O(41) => OTMP_14_41_port, 
                           O(40) => OTMP_14_40_port, O(39) => OTMP_14_39_port, 
                           O(38) => OTMP_14_38_port, O(37) => OTMP_14_37_port, 
                           O(36) => OTMP_14_36_port, O(35) => OTMP_14_35_port, 
                           O(34) => OTMP_14_34_port, O(33) => OTMP_14_33_port, 
                           O(32) => OTMP_14_32_port, O(31) => OTMP_14_31_port, 
                           O(30) => OTMP_14_30_port, O(29) => OTMP_14_29_port, 
                           O(28) => OTMP_14_28_port, O(27) => OTMP_14_27_port, 
                           O(26) => OTMP_14_26_port, O(25) => OTMP_14_25_port, 
                           O(24) => OTMP_14_24_port, O(23) => OTMP_14_23_port, 
                           O(22) => OTMP_14_22_port, O(21) => OTMP_14_21_port, 
                           O(20) => OTMP_14_20_port, O(19) => OTMP_14_19_port, 
                           O(18) => OTMP_14_18_port, O(17) => OTMP_14_17_port, 
                           O(16) => OTMP_14_16_port, O(15) => OTMP_14_15_port, 
                           O(14) => OTMP_14_14_port, O(13) => OTMP_14_13_port, 
                           O(12) => OTMP_14_12_port, O(11) => OTMP_14_11_port, 
                           O(10) => OTMP_14_10_port, O(9) => OTMP_14_9_port, 
                           O(8) => OTMP_14_8_port, O(7) => OTMP_14_7_port, O(6)
                           => OTMP_14_6_port, O(5) => OTMP_14_5_port, O(4) => 
                           OTMP_14_4_port, O(3) => OTMP_14_3_port, O(2) => 
                           OTMP_14_2_port, O(1) => OTMP_14_1_port, O(0) => 
                           n_1147, A_so(61) => SHIFT_15_61_port, A_so(60) => 
                           SHIFT_15_60_port, A_so(59) => SHIFT_15_59_port, 
                           A_so(58) => SHIFT_15_58_port, A_so(57) => 
                           SHIFT_15_57_port, A_so(56) => SHIFT_15_56_port, 
                           A_so(55) => SHIFT_15_55_port, A_so(54) => 
                           SHIFT_15_54_port, A_so(53) => SHIFT_15_53_port, 
                           A_so(52) => SHIFT_15_52_port, A_so(51) => 
                           SHIFT_15_51_port, A_so(50) => SHIFT_15_50_port, 
                           A_so(49) => SHIFT_15_49_port, A_so(48) => 
                           SHIFT_15_48_port, A_so(47) => SHIFT_15_47_port, 
                           A_so(46) => SHIFT_15_46_port, A_so(45) => 
                           SHIFT_15_45_port, A_so(44) => SHIFT_15_44_port, 
                           A_so(43) => SHIFT_15_43_port, A_so(42) => 
                           SHIFT_15_42_port, A_so(41) => SHIFT_15_41_port, 
                           A_so(40) => SHIFT_15_40_port, A_so(39) => 
                           SHIFT_15_39_port, A_so(38) => SHIFT_15_38_port, 
                           A_so(37) => SHIFT_15_37_port, A_so(36) => 
                           SHIFT_15_36_port, A_so(35) => SHIFT_15_35_port, 
                           A_so(34) => SHIFT_15_34_port, A_so(33) => 
                           SHIFT_15_33_port, A_so(32) => SHIFT_15_32_port, 
                           A_so(31) => SHIFT_15_31_port, A_so(30) => 
                           SHIFT_15_30_port, A_so(29) => SHIFT_15_29_port, 
                           A_so(28) => SHIFT_15_28_port, A_so(27) => 
                           SHIFT_15_27_port, A_so(26) => SHIFT_15_26_port, 
                           A_so(25) => SHIFT_15_25_port, A_so(24) => 
                           SHIFT_15_24_port, A_so(23) => SHIFT_15_23_port, 
                           A_so(22) => SHIFT_15_22_port, A_so(21) => 
                           SHIFT_15_21_port, A_so(20) => SHIFT_15_20_port, 
                           A_so(19) => SHIFT_15_19_port, A_so(18) => 
                           SHIFT_15_18_port, A_so(17) => SHIFT_15_17_port, 
                           A_so(16) => SHIFT_15_16_port, A_so(15) => 
                           SHIFT_15_15_port, A_so(14) => SHIFT_15_14_port, 
                           A_so(13) => SHIFT_15_13_port, A_so(12) => 
                           SHIFT_15_12_port, A_so(11) => SHIFT_15_11_port, 
                           A_so(10) => SHIFT_15_10_port, A_so(9) => 
                           SHIFT_15_9_port, A_so(8) => SHIFT_15_8_port, A_so(7)
                           => SHIFT_15_7_port, A_so(6) => SHIFT_15_6_port, 
                           A_so(5) => SHIFT_15_5_port, A_so(4) => 
                           SHIFT_15_4_port, A_so(3) => SHIFT_15_3_port, A_so(2)
                           => SHIFT_15_2_port, A_so(1) => n_1148, A_so(0) => 
                           n_1149, A_nso(61) => SHIFT_n_15_61_port, A_nso(60) 
                           => SHIFT_n_15_60_port, A_nso(59) => 
                           SHIFT_n_15_59_port, A_nso(58) => SHIFT_n_15_58_port,
                           A_nso(57) => SHIFT_n_15_57_port, A_nso(56) => 
                           SHIFT_n_15_56_port, A_nso(55) => SHIFT_n_15_55_port,
                           A_nso(54) => SHIFT_n_15_54_port, A_nso(53) => 
                           SHIFT_n_15_53_port, A_nso(52) => SHIFT_n_15_52_port,
                           A_nso(51) => SHIFT_n_15_51_port, A_nso(50) => 
                           SHIFT_n_15_50_port, A_nso(49) => SHIFT_n_15_49_port,
                           A_nso(48) => SHIFT_n_15_48_port, A_nso(47) => 
                           SHIFT_n_15_47_port, A_nso(46) => SHIFT_n_15_46_port,
                           A_nso(45) => SHIFT_n_15_45_port, A_nso(44) => 
                           SHIFT_n_15_44_port, A_nso(43) => SHIFT_n_15_43_port,
                           A_nso(42) => SHIFT_n_15_42_port, A_nso(41) => 
                           SHIFT_n_15_41_port, A_nso(40) => SHIFT_n_15_40_port,
                           A_nso(39) => SHIFT_n_15_39_port, A_nso(38) => 
                           SHIFT_n_15_38_port, A_nso(37) => SHIFT_n_15_37_port,
                           A_nso(36) => SHIFT_n_15_36_port, A_nso(35) => 
                           SHIFT_n_15_35_port, A_nso(34) => SHIFT_n_15_34_port,
                           A_nso(33) => SHIFT_n_15_33_port, A_nso(32) => 
                           SHIFT_n_15_32_port, A_nso(31) => SHIFT_n_15_31_port,
                           A_nso(30) => SHIFT_n_15_30_port, A_nso(29) => 
                           SHIFT_n_15_29_port, A_nso(28) => SHIFT_n_15_28_port,
                           A_nso(27) => SHIFT_n_15_27_port, A_nso(26) => 
                           SHIFT_n_15_26_port, A_nso(25) => SHIFT_n_15_25_port,
                           A_nso(24) => SHIFT_n_15_24_port, A_nso(23) => 
                           SHIFT_n_15_23_port, A_nso(22) => SHIFT_n_15_22_port,
                           A_nso(21) => SHIFT_n_15_21_port, A_nso(20) => 
                           SHIFT_n_15_20_port, A_nso(19) => SHIFT_n_15_19_port,
                           A_nso(18) => SHIFT_n_15_18_port, A_nso(17) => 
                           SHIFT_n_15_17_port, A_nso(16) => SHIFT_n_15_16_port,
                           A_nso(15) => SHIFT_n_15_15_port, A_nso(14) => 
                           SHIFT_n_15_14_port, A_nso(13) => SHIFT_n_15_13_port,
                           A_nso(12) => SHIFT_n_15_12_port, A_nso(11) => 
                           SHIFT_n_15_11_port, A_nso(10) => SHIFT_n_15_10_port,
                           A_nso(9) => SHIFT_n_15_9_port, A_nso(8) => 
                           SHIFT_n_15_8_port, A_nso(7) => SHIFT_n_15_7_port, 
                           A_nso(6) => SHIFT_n_15_6_port, A_nso(5) => 
                           SHIFT_n_15_5_port, A_nso(4) => SHIFT_n_15_4_port, 
                           A_nso(3) => SHIFT_n_15_3_port, A_nso(2) => 
                           SHIFT_n_15_2_port, A_nso(1) => n_1150, A_nso(0) => 
                           n_1151);
   ENC_15 : BOOTHENC_NBIT64_i30 port map( A_s(63) => SHIFT_15_61_port, A_s(62) 
                           => SHIFT_15_61_port, A_s(61) => SHIFT_15_61_port, 
                           A_s(60) => SHIFT_15_60_port, A_s(59) => 
                           SHIFT_15_59_port, A_s(58) => SHIFT_15_58_port, 
                           A_s(57) => SHIFT_15_57_port, A_s(56) => 
                           SHIFT_15_56_port, A_s(55) => SHIFT_15_55_port, 
                           A_s(54) => SHIFT_15_54_port, A_s(53) => 
                           SHIFT_15_53_port, A_s(52) => SHIFT_15_52_port, 
                           A_s(51) => SHIFT_15_51_port, A_s(50) => 
                           SHIFT_15_50_port, A_s(49) => SHIFT_15_49_port, 
                           A_s(48) => SHIFT_15_48_port, A_s(47) => 
                           SHIFT_15_47_port, A_s(46) => SHIFT_15_46_port, 
                           A_s(45) => SHIFT_15_45_port, A_s(44) => 
                           SHIFT_15_44_port, A_s(43) => SHIFT_15_43_port, 
                           A_s(42) => SHIFT_15_42_port, A_s(41) => 
                           SHIFT_15_41_port, A_s(40) => SHIFT_15_40_port, 
                           A_s(39) => SHIFT_15_39_port, A_s(38) => 
                           SHIFT_15_38_port, A_s(37) => SHIFT_15_37_port, 
                           A_s(36) => SHIFT_15_36_port, A_s(35) => 
                           SHIFT_15_35_port, A_s(34) => SHIFT_15_34_port, 
                           A_s(33) => SHIFT_15_33_port, A_s(32) => 
                           SHIFT_15_32_port, A_s(31) => SHIFT_15_31_port, 
                           A_s(30) => SHIFT_15_30_port, A_s(29) => 
                           SHIFT_15_29_port, A_s(28) => SHIFT_15_28_port, 
                           A_s(27) => SHIFT_15_27_port, A_s(26) => 
                           SHIFT_15_26_port, A_s(25) => SHIFT_15_25_port, 
                           A_s(24) => SHIFT_15_24_port, A_s(23) => 
                           SHIFT_15_23_port, A_s(22) => SHIFT_15_22_port, 
                           A_s(21) => SHIFT_15_21_port, A_s(20) => 
                           SHIFT_15_20_port, A_s(19) => SHIFT_15_19_port, 
                           A_s(18) => SHIFT_15_18_port, A_s(17) => 
                           SHIFT_15_17_port, A_s(16) => SHIFT_15_16_port, 
                           A_s(15) => SHIFT_15_15_port, A_s(14) => 
                           SHIFT_15_14_port, A_s(13) => SHIFT_15_13_port, 
                           A_s(12) => SHIFT_15_12_port, A_s(11) => 
                           SHIFT_15_11_port, A_s(10) => SHIFT_15_10_port, 
                           A_s(9) => SHIFT_15_9_port, A_s(8) => SHIFT_15_8_port
                           , A_s(7) => SHIFT_15_7_port, A_s(6) => 
                           SHIFT_15_6_port, A_s(5) => SHIFT_15_5_port, A_s(4) 
                           => SHIFT_15_4_port, A_s(3) => SHIFT_15_3_port, 
                           A_s(2) => SHIFT_15_2_port, A_s(1) => SHIFT_15_1_port
                           , A_s(0) => SHIFT_15_0_port, A_ns(63) => 
                           SHIFT_n_15_61_port, A_ns(62) => SHIFT_n_15_61_port, 
                           A_ns(61) => SHIFT_n_15_61_port, A_ns(60) => 
                           SHIFT_n_15_60_port, A_ns(59) => SHIFT_n_15_59_port, 
                           A_ns(58) => SHIFT_n_15_58_port, A_ns(57) => 
                           SHIFT_n_15_57_port, A_ns(56) => SHIFT_n_15_56_port, 
                           A_ns(55) => SHIFT_n_15_55_port, A_ns(54) => 
                           SHIFT_n_15_54_port, A_ns(53) => SHIFT_n_15_53_port, 
                           A_ns(52) => SHIFT_n_15_52_port, A_ns(51) => 
                           SHIFT_n_15_51_port, A_ns(50) => SHIFT_n_15_50_port, 
                           A_ns(49) => SHIFT_n_15_49_port, A_ns(48) => 
                           SHIFT_n_15_48_port, A_ns(47) => SHIFT_n_15_47_port, 
                           A_ns(46) => SHIFT_n_15_46_port, A_ns(45) => 
                           SHIFT_n_15_45_port, A_ns(44) => SHIFT_n_15_44_port, 
                           A_ns(43) => SHIFT_n_15_43_port, A_ns(42) => 
                           SHIFT_n_15_42_port, A_ns(41) => SHIFT_n_15_41_port, 
                           A_ns(40) => SHIFT_n_15_40_port, A_ns(39) => 
                           SHIFT_n_15_39_port, A_ns(38) => SHIFT_n_15_38_port, 
                           A_ns(37) => SHIFT_n_15_37_port, A_ns(36) => 
                           SHIFT_n_15_36_port, A_ns(35) => SHIFT_n_15_35_port, 
                           A_ns(34) => SHIFT_n_15_34_port, A_ns(33) => 
                           SHIFT_n_15_33_port, A_ns(32) => SHIFT_n_15_32_port, 
                           A_ns(31) => SHIFT_n_15_31_port, A_ns(30) => 
                           SHIFT_n_15_30_port, A_ns(29) => SHIFT_n_15_29_port, 
                           A_ns(28) => SHIFT_n_15_28_port, A_ns(27) => 
                           SHIFT_n_15_27_port, A_ns(26) => SHIFT_n_15_26_port, 
                           A_ns(25) => SHIFT_n_15_25_port, A_ns(24) => 
                           SHIFT_n_15_24_port, A_ns(23) => SHIFT_n_15_23_port, 
                           A_ns(22) => SHIFT_n_15_22_port, A_ns(21) => 
                           SHIFT_n_15_21_port, A_ns(20) => SHIFT_n_15_20_port, 
                           A_ns(19) => SHIFT_n_15_19_port, A_ns(18) => 
                           SHIFT_n_15_18_port, A_ns(17) => SHIFT_n_15_17_port, 
                           A_ns(16) => SHIFT_n_15_16_port, A_ns(15) => 
                           SHIFT_n_15_15_port, A_ns(14) => SHIFT_n_15_14_port, 
                           A_ns(13) => SHIFT_n_15_13_port, A_ns(12) => 
                           SHIFT_n_15_12_port, A_ns(11) => SHIFT_n_15_11_port, 
                           A_ns(10) => SHIFT_n_15_10_port, A_ns(9) => 
                           SHIFT_n_15_9_port, A_ns(8) => SHIFT_n_15_8_port, 
                           A_ns(7) => SHIFT_n_15_7_port, A_ns(6) => 
                           SHIFT_n_15_6_port, A_ns(5) => SHIFT_n_15_5_port, 
                           A_ns(4) => SHIFT_n_15_4_port, A_ns(3) => 
                           SHIFT_n_15_3_port, A_ns(2) => SHIFT_n_15_2_port, 
                           A_ns(1) => SHIFT_n_15_1_port, A_ns(0) => 
                           SHIFT_n_15_0_port, B(63) => B(31), B(62) => B(31), 
                           B(61) => B(31), B(60) => B(31), B(59) => B(31), 
                           B(58) => B(31), B(57) => B(31), B(56) => B(31), 
                           B(55) => B(31), B(54) => B(31), B(53) => B(31), 
                           B(52) => B(31), B(51) => B(31), B(50) => B(31), 
                           B(49) => B(31), B(48) => B(31), B(47) => B(31), 
                           B(46) => B(31), B(45) => B(31), B(44) => B(31), 
                           B(43) => B(31), B(42) => B(31), B(41) => B(31), 
                           B(40) => B(31), B(39) => B(31), B(38) => B(31), 
                           B(37) => B(31), B(36) => B(31), B(35) => B(31), 
                           B(34) => B(31), B(33) => B(31), B(32) => B(31), 
                           B(31) => B(31), B(30) => B(30), B(29) => B(29), 
                           B(28) => B(28), B(27) => B(27), B(26) => B(26), 
                           B(25) => B(25), B(24) => B(24), B(23) => B(23), 
                           B(22) => B(22), B(21) => B(21), B(20) => B(20), 
                           B(19) => B(19), B(18) => B(18), B(17) => B(17), 
                           B(16) => B(16), B(15) => B(15), B(14) => B(14), 
                           B(13) => B(13), B(12) => B(12), B(11) => B(11), 
                           B(10) => B(10), B(9) => B(9), B(8) => B(8), B(7) => 
                           B(7), B(6) => B(6), B(5) => B(5), B(4) => B(4), B(3)
                           => B(3), B(2) => B(2), B(1) => B(1), B(0) => B(0), 
                           O(63) => OTMP_15_63_port, O(62) => OTMP_15_62_port, 
                           O(61) => OTMP_15_61_port, O(60) => OTMP_15_60_port, 
                           O(59) => OTMP_15_59_port, O(58) => OTMP_15_58_port, 
                           O(57) => OTMP_15_57_port, O(56) => OTMP_15_56_port, 
                           O(55) => OTMP_15_55_port, O(54) => OTMP_15_54_port, 
                           O(53) => OTMP_15_53_port, O(52) => OTMP_15_52_port, 
                           O(51) => OTMP_15_51_port, O(50) => OTMP_15_50_port, 
                           O(49) => OTMP_15_49_port, O(48) => OTMP_15_48_port, 
                           O(47) => OTMP_15_47_port, O(46) => OTMP_15_46_port, 
                           O(45) => OTMP_15_45_port, O(44) => OTMP_15_44_port, 
                           O(43) => OTMP_15_43_port, O(42) => OTMP_15_42_port, 
                           O(41) => OTMP_15_41_port, O(40) => OTMP_15_40_port, 
                           O(39) => OTMP_15_39_port, O(38) => OTMP_15_38_port, 
                           O(37) => OTMP_15_37_port, O(36) => OTMP_15_36_port, 
                           O(35) => OTMP_15_35_port, O(34) => OTMP_15_34_port, 
                           O(33) => OTMP_15_33_port, O(32) => OTMP_15_32_port, 
                           O(31) => OTMP_15_31_port, O(30) => OTMP_15_30_port, 
                           O(29) => OTMP_15_29_port, O(28) => OTMP_15_28_port, 
                           O(27) => OTMP_15_27_port, O(26) => OTMP_15_26_port, 
                           O(25) => OTMP_15_25_port, O(24) => OTMP_15_24_port, 
                           O(23) => OTMP_15_23_port, O(22) => OTMP_15_22_port, 
                           O(21) => OTMP_15_21_port, O(20) => OTMP_15_20_port, 
                           O(19) => OTMP_15_19_port, O(18) => OTMP_15_18_port, 
                           O(17) => OTMP_15_17_port, O(16) => OTMP_15_16_port, 
                           O(15) => OTMP_15_15_port, O(14) => OTMP_15_14_port, 
                           O(13) => OTMP_15_13_port, O(12) => OTMP_15_12_port, 
                           O(11) => OTMP_15_11_port, O(10) => OTMP_15_10_port, 
                           O(9) => OTMP_15_9_port, O(8) => OTMP_15_8_port, O(7)
                           => OTMP_15_7_port, O(6) => OTMP_15_6_port, O(5) => 
                           OTMP_15_5_port, O(4) => OTMP_15_4_port, O(3) => 
                           OTMP_15_3_port, O(2) => OTMP_15_2_port, O(1) => 
                           OTMP_15_1_port, O(0) => n_1152, A_so(63) => n_1153, 
                           A_so(62) => n_1154, A_so(61) => n_1155, A_so(60) => 
                           n_1156, A_so(59) => n_1157, A_so(58) => n_1158, 
                           A_so(57) => n_1159, A_so(56) => n_1160, A_so(55) => 
                           n_1161, A_so(54) => n_1162, A_so(53) => n_1163, 
                           A_so(52) => n_1164, A_so(51) => n_1165, A_so(50) => 
                           n_1166, A_so(49) => n_1167, A_so(48) => n_1168, 
                           A_so(47) => n_1169, A_so(46) => n_1170, A_so(45) => 
                           n_1171, A_so(44) => n_1172, A_so(43) => n_1173, 
                           A_so(42) => n_1174, A_so(41) => n_1175, A_so(40) => 
                           n_1176, A_so(39) => n_1177, A_so(38) => n_1178, 
                           A_so(37) => n_1179, A_so(36) => n_1180, A_so(35) => 
                           n_1181, A_so(34) => n_1182, A_so(33) => n_1183, 
                           A_so(32) => n_1184, A_so(31) => n_1185, A_so(30) => 
                           n_1186, A_so(29) => n_1187, A_so(28) => n_1188, 
                           A_so(27) => n_1189, A_so(26) => n_1190, A_so(25) => 
                           n_1191, A_so(24) => n_1192, A_so(23) => n_1193, 
                           A_so(22) => n_1194, A_so(21) => n_1195, A_so(20) => 
                           n_1196, A_so(19) => n_1197, A_so(18) => n_1198, 
                           A_so(17) => n_1199, A_so(16) => n_1200, A_so(15) => 
                           n_1201, A_so(14) => n_1202, A_so(13) => n_1203, 
                           A_so(12) => n_1204, A_so(11) => n_1205, A_so(10) => 
                           n_1206, A_so(9) => n_1207, A_so(8) => n_1208, 
                           A_so(7) => n_1209, A_so(6) => n_1210, A_so(5) => 
                           n_1211, A_so(4) => n_1212, A_so(3) => n_1213, 
                           A_so(2) => n_1214, A_so(1) => n_1215, A_so(0) => 
                           n_1216, A_nso(63) => n_1217, A_nso(62) => n_1218, 
                           A_nso(61) => n_1219, A_nso(60) => n_1220, A_nso(59) 
                           => n_1221, A_nso(58) => n_1222, A_nso(57) => n_1223,
                           A_nso(56) => n_1224, A_nso(55) => n_1225, A_nso(54) 
                           => n_1226, A_nso(53) => n_1227, A_nso(52) => n_1228,
                           A_nso(51) => n_1229, A_nso(50) => n_1230, A_nso(49) 
                           => n_1231, A_nso(48) => n_1232, A_nso(47) => n_1233,
                           A_nso(46) => n_1234, A_nso(45) => n_1235, A_nso(44) 
                           => n_1236, A_nso(43) => n_1237, A_nso(42) => n_1238,
                           A_nso(41) => n_1239, A_nso(40) => n_1240, A_nso(39) 
                           => n_1241, A_nso(38) => n_1242, A_nso(37) => n_1243,
                           A_nso(36) => n_1244, A_nso(35) => n_1245, A_nso(34) 
                           => n_1246, A_nso(33) => n_1247, A_nso(32) => n_1248,
                           A_nso(31) => n_1249, A_nso(30) => n_1250, A_nso(29) 
                           => n_1251, A_nso(28) => n_1252, A_nso(27) => n_1253,
                           A_nso(26) => n_1254, A_nso(25) => n_1255, A_nso(24) 
                           => n_1256, A_nso(23) => n_1257, A_nso(22) => n_1258,
                           A_nso(21) => n_1259, A_nso(20) => n_1260, A_nso(19) 
                           => n_1261, A_nso(18) => n_1262, A_nso(17) => n_1263,
                           A_nso(16) => n_1264, A_nso(15) => n_1265, A_nso(14) 
                           => n_1266, A_nso(13) => n_1267, A_nso(12) => n_1268,
                           A_nso(11) => n_1269, A_nso(10) => n_1270, A_nso(9) 
                           => n_1271, A_nso(8) => n_1272, A_nso(7) => n_1273, 
                           A_nso(6) => n_1274, A_nso(5) => n_1275, A_nso(4) => 
                           n_1276, A_nso(3) => n_1277, A_nso(2) => n_1278, 
                           A_nso(1) => n_1279, A_nso(0) => n_1280);
   ADDER1 : RCA_NBIT36 port map( A(35) => OTMP_0_34_port, A(34) => 
                           OTMP_0_34_port, A(33) => OTMP_0_34_port, A(32) => 
                           OTMP_0_32_port, A(31) => OTMP_0_31_port, A(30) => 
                           OTMP_0_30_port, A(29) => OTMP_0_29_port, A(28) => 
                           OTMP_0_28_port, A(27) => OTMP_0_27_port, A(26) => 
                           OTMP_0_26_port, A(25) => OTMP_0_25_port, A(24) => 
                           OTMP_0_24_port, A(23) => OTMP_0_23_port, A(22) => 
                           OTMP_0_22_port, A(21) => OTMP_0_21_port, A(20) => 
                           OTMP_0_20_port, A(19) => OTMP_0_19_port, A(18) => 
                           OTMP_0_18_port, A(17) => OTMP_0_17_port, A(16) => 
                           OTMP_0_16_port, A(15) => OTMP_0_15_port, A(14) => 
                           OTMP_0_14_port, A(13) => OTMP_0_13_port, A(12) => 
                           OTMP_0_12_port, A(11) => OTMP_0_11_port, A(10) => 
                           OTMP_0_10_port, A(9) => OTMP_0_9_port, A(8) => 
                           OTMP_0_8_port, A(7) => OTMP_0_7_port, A(6) => 
                           OTMP_0_6_port, A(5) => OTMP_0_5_port, A(4) => 
                           OTMP_0_4_port, A(3) => OTMP_0_3_port, A(2) => 
                           OTMP_0_2_port, A(1) => OTMP_0_1_port, A(0) => 
                           OTMP_0_0_port, B(35) => OTMP_1_35_port, B(34) => 
                           OTMP_1_34_port, B(33) => OTMP_1_33_port, B(32) => 
                           OTMP_1_32_port, B(31) => OTMP_1_31_port, B(30) => 
                           OTMP_1_30_port, B(29) => OTMP_1_29_port, B(28) => 
                           OTMP_1_28_port, B(27) => OTMP_1_27_port, B(26) => 
                           OTMP_1_26_port, B(25) => OTMP_1_25_port, B(24) => 
                           OTMP_1_24_port, B(23) => OTMP_1_23_port, B(22) => 
                           OTMP_1_22_port, B(21) => OTMP_1_21_port, B(20) => 
                           OTMP_1_20_port, B(19) => OTMP_1_19_port, B(18) => 
                           OTMP_1_18_port, B(17) => OTMP_1_17_port, B(16) => 
                           OTMP_1_16_port, B(15) => OTMP_1_15_port, B(14) => 
                           OTMP_1_14_port, B(13) => OTMP_1_13_port, B(12) => 
                           OTMP_1_12_port, B(11) => OTMP_1_11_port, B(10) => 
                           OTMP_1_10_port, B(9) => OTMP_1_9_port, B(8) => 
                           OTMP_1_8_port, B(7) => OTMP_1_7_port, B(6) => 
                           OTMP_1_6_port, B(5) => OTMP_1_5_port, B(4) => 
                           OTMP_1_4_port, B(3) => OTMP_1_3_port, B(2) => 
                           OTMP_1_2_port, B(1) => OTMP_1_1_port, B(0) => 
                           OTMP_1_0_port, Ci => X_Logic0_port, S(35) => 
                           PTMP_0_36_port, S(34) => PTMP_0_34_port, S(33) => 
                           PTMP_0_33_port, S(32) => PTMP_0_32_port, S(31) => 
                           PTMP_0_31_port, S(30) => PTMP_0_30_port, S(29) => 
                           PTMP_0_29_port, S(28) => PTMP_0_28_port, S(27) => 
                           PTMP_0_27_port, S(26) => PTMP_0_26_port, S(25) => 
                           PTMP_0_25_port, S(24) => PTMP_0_24_port, S(23) => 
                           PTMP_0_23_port, S(22) => PTMP_0_22_port, S(21) => 
                           PTMP_0_21_port, S(20) => PTMP_0_20_port, S(19) => 
                           PTMP_0_19_port, S(18) => PTMP_0_18_port, S(17) => 
                           PTMP_0_17_port, S(16) => PTMP_0_16_port, S(15) => 
                           PTMP_0_15_port, S(14) => PTMP_0_14_port, S(13) => 
                           PTMP_0_13_port, S(12) => PTMP_0_12_port, S(11) => 
                           PTMP_0_11_port, S(10) => PTMP_0_10_port, S(9) => 
                           PTMP_0_9_port, S(8) => PTMP_0_8_port, S(7) => 
                           PTMP_0_7_port, S(6) => PTMP_0_6_port, S(5) => 
                           PTMP_0_5_port, S(4) => PTMP_0_4_port, S(3) => 
                           PTMP_0_3_port, S(2) => PTMP_0_2_port, S(1) => 
                           PTMP_0_1_port, S(0) => PTMP_0_0_port, Co => n_1281);
   ADDER_2 : RCA_NBIT38 port map( A(37) => PTMP_0_36_port, A(36) => 
                           PTMP_0_36_port, A(35) => PTMP_0_36_port, A(34) => 
                           PTMP_0_34_port, A(33) => PTMP_0_33_port, A(32) => 
                           PTMP_0_32_port, A(31) => PTMP_0_31_port, A(30) => 
                           PTMP_0_30_port, A(29) => PTMP_0_29_port, A(28) => 
                           PTMP_0_28_port, A(27) => PTMP_0_27_port, A(26) => 
                           PTMP_0_26_port, A(25) => PTMP_0_25_port, A(24) => 
                           PTMP_0_24_port, A(23) => PTMP_0_23_port, A(22) => 
                           PTMP_0_22_port, A(21) => PTMP_0_21_port, A(20) => 
                           PTMP_0_20_port, A(19) => PTMP_0_19_port, A(18) => 
                           PTMP_0_18_port, A(17) => PTMP_0_17_port, A(16) => 
                           PTMP_0_16_port, A(15) => PTMP_0_15_port, A(14) => 
                           PTMP_0_14_port, A(13) => PTMP_0_13_port, A(12) => 
                           PTMP_0_12_port, A(11) => PTMP_0_11_port, A(10) => 
                           PTMP_0_10_port, A(9) => PTMP_0_9_port, A(8) => 
                           PTMP_0_8_port, A(7) => PTMP_0_7_port, A(6) => 
                           PTMP_0_6_port, A(5) => PTMP_0_5_port, A(4) => 
                           PTMP_0_4_port, A(3) => PTMP_0_3_port, A(2) => 
                           PTMP_0_2_port, A(1) => PTMP_0_1_port, A(0) => 
                           PTMP_0_0_port, B(37) => OTMP_2_37_port, B(36) => 
                           OTMP_2_36_port, B(35) => OTMP_2_35_port, B(34) => 
                           OTMP_2_34_port, B(33) => OTMP_2_33_port, B(32) => 
                           OTMP_2_32_port, B(31) => OTMP_2_31_port, B(30) => 
                           OTMP_2_30_port, B(29) => OTMP_2_29_port, B(28) => 
                           OTMP_2_28_port, B(27) => OTMP_2_27_port, B(26) => 
                           OTMP_2_26_port, B(25) => OTMP_2_25_port, B(24) => 
                           OTMP_2_24_port, B(23) => OTMP_2_23_port, B(22) => 
                           OTMP_2_22_port, B(21) => OTMP_2_21_port, B(20) => 
                           OTMP_2_20_port, B(19) => OTMP_2_19_port, B(18) => 
                           OTMP_2_18_port, B(17) => OTMP_2_17_port, B(16) => 
                           OTMP_2_16_port, B(15) => OTMP_2_15_port, B(14) => 
                           OTMP_2_14_port, B(13) => OTMP_2_13_port, B(12) => 
                           OTMP_2_12_port, B(11) => OTMP_2_11_port, B(10) => 
                           OTMP_2_10_port, B(9) => OTMP_2_9_port, B(8) => 
                           OTMP_2_8_port, B(7) => OTMP_2_7_port, B(6) => 
                           OTMP_2_6_port, B(5) => OTMP_2_5_port, B(4) => 
                           OTMP_2_4_port, B(3) => OTMP_2_3_port, B(2) => 
                           OTMP_2_2_port, B(1) => OTMP_2_1_port, B(0) => 
                           OTMP_2_0_port, Ci => X_Logic0_port, S(37) => 
                           PTMP_1_37_port, S(36) => PTMP_1_36_port, S(35) => 
                           PTMP_1_35_port, S(34) => PTMP_1_34_port, S(33) => 
                           PTMP_1_33_port, S(32) => PTMP_1_32_port, S(31) => 
                           PTMP_1_31_port, S(30) => PTMP_1_30_port, S(29) => 
                           PTMP_1_29_port, S(28) => PTMP_1_28_port, S(27) => 
                           PTMP_1_27_port, S(26) => PTMP_1_26_port, S(25) => 
                           PTMP_1_25_port, S(24) => PTMP_1_24_port, S(23) => 
                           PTMP_1_23_port, S(22) => PTMP_1_22_port, S(21) => 
                           PTMP_1_21_port, S(20) => PTMP_1_20_port, S(19) => 
                           PTMP_1_19_port, S(18) => PTMP_1_18_port, S(17) => 
                           PTMP_1_17_port, S(16) => PTMP_1_16_port, S(15) => 
                           PTMP_1_15_port, S(14) => PTMP_1_14_port, S(13) => 
                           PTMP_1_13_port, S(12) => PTMP_1_12_port, S(11) => 
                           PTMP_1_11_port, S(10) => PTMP_1_10_port, S(9) => 
                           PTMP_1_9_port, S(8) => PTMP_1_8_port, S(7) => 
                           PTMP_1_7_port, S(6) => PTMP_1_6_port, S(5) => 
                           PTMP_1_5_port, S(4) => PTMP_1_4_port, S(3) => 
                           PTMP_1_3_port, S(2) => PTMP_1_2_port, S(1) => 
                           PTMP_1_1_port, S(0) => PTMP_1_0_port, Co => n_1282);
   ADDER_3 : RCA_NBIT40 port map( A(39) => PTMP_1_37_port, A(38) => 
                           PTMP_1_37_port, A(37) => PTMP_1_37_port, A(36) => 
                           PTMP_1_36_port, A(35) => PTMP_1_35_port, A(34) => 
                           PTMP_1_34_port, A(33) => PTMP_1_33_port, A(32) => 
                           PTMP_1_32_port, A(31) => PTMP_1_31_port, A(30) => 
                           PTMP_1_30_port, A(29) => PTMP_1_29_port, A(28) => 
                           PTMP_1_28_port, A(27) => PTMP_1_27_port, A(26) => 
                           PTMP_1_26_port, A(25) => PTMP_1_25_port, A(24) => 
                           PTMP_1_24_port, A(23) => PTMP_1_23_port, A(22) => 
                           PTMP_1_22_port, A(21) => PTMP_1_21_port, A(20) => 
                           PTMP_1_20_port, A(19) => PTMP_1_19_port, A(18) => 
                           PTMP_1_18_port, A(17) => PTMP_1_17_port, A(16) => 
                           PTMP_1_16_port, A(15) => PTMP_1_15_port, A(14) => 
                           PTMP_1_14_port, A(13) => PTMP_1_13_port, A(12) => 
                           PTMP_1_12_port, A(11) => PTMP_1_11_port, A(10) => 
                           PTMP_1_10_port, A(9) => PTMP_1_9_port, A(8) => 
                           PTMP_1_8_port, A(7) => PTMP_1_7_port, A(6) => 
                           PTMP_1_6_port, A(5) => PTMP_1_5_port, A(4) => 
                           PTMP_1_4_port, A(3) => PTMP_1_3_port, A(2) => 
                           PTMP_1_2_port, A(1) => PTMP_1_1_port, A(0) => 
                           PTMP_1_0_port, B(39) => OTMP_3_39_port, B(38) => 
                           OTMP_3_38_port, B(37) => OTMP_3_37_port, B(36) => 
                           OTMP_3_36_port, B(35) => OTMP_3_35_port, B(34) => 
                           OTMP_3_34_port, B(33) => OTMP_3_33_port, B(32) => 
                           OTMP_3_32_port, B(31) => OTMP_3_31_port, B(30) => 
                           OTMP_3_30_port, B(29) => OTMP_3_29_port, B(28) => 
                           OTMP_3_28_port, B(27) => OTMP_3_27_port, B(26) => 
                           OTMP_3_26_port, B(25) => OTMP_3_25_port, B(24) => 
                           OTMP_3_24_port, B(23) => OTMP_3_23_port, B(22) => 
                           OTMP_3_22_port, B(21) => OTMP_3_21_port, B(20) => 
                           OTMP_3_20_port, B(19) => OTMP_3_19_port, B(18) => 
                           OTMP_3_18_port, B(17) => OTMP_3_17_port, B(16) => 
                           OTMP_3_16_port, B(15) => OTMP_3_15_port, B(14) => 
                           OTMP_3_14_port, B(13) => OTMP_3_13_port, B(12) => 
                           OTMP_3_12_port, B(11) => OTMP_3_11_port, B(10) => 
                           OTMP_3_10_port, B(9) => OTMP_3_9_port, B(8) => 
                           OTMP_3_8_port, B(7) => OTMP_3_7_port, B(6) => 
                           OTMP_3_6_port, B(5) => OTMP_3_5_port, B(4) => 
                           OTMP_3_4_port, B(3) => OTMP_3_3_port, B(2) => 
                           OTMP_3_2_port, B(1) => OTMP_3_1_port, B(0) => 
                           OTMP_3_0_port, Ci => X_Logic0_port, S(39) => 
                           PTMP_2_39_port, S(38) => PTMP_2_38_port, S(37) => 
                           PTMP_2_37_port, S(36) => PTMP_2_36_port, S(35) => 
                           PTMP_2_35_port, S(34) => PTMP_2_34_port, S(33) => 
                           PTMP_2_33_port, S(32) => PTMP_2_32_port, S(31) => 
                           PTMP_2_31_port, S(30) => PTMP_2_30_port, S(29) => 
                           PTMP_2_29_port, S(28) => PTMP_2_28_port, S(27) => 
                           PTMP_2_27_port, S(26) => PTMP_2_26_port, S(25) => 
                           PTMP_2_25_port, S(24) => PTMP_2_24_port, S(23) => 
                           PTMP_2_23_port, S(22) => PTMP_2_22_port, S(21) => 
                           PTMP_2_21_port, S(20) => PTMP_2_20_port, S(19) => 
                           PTMP_2_19_port, S(18) => PTMP_2_18_port, S(17) => 
                           PTMP_2_17_port, S(16) => PTMP_2_16_port, S(15) => 
                           PTMP_2_15_port, S(14) => PTMP_2_14_port, S(13) => 
                           PTMP_2_13_port, S(12) => PTMP_2_12_port, S(11) => 
                           PTMP_2_11_port, S(10) => PTMP_2_10_port, S(9) => 
                           PTMP_2_9_port, S(8) => PTMP_2_8_port, S(7) => 
                           PTMP_2_7_port, S(6) => PTMP_2_6_port, S(5) => 
                           PTMP_2_5_port, S(4) => PTMP_2_4_port, S(3) => 
                           PTMP_2_3_port, S(2) => PTMP_2_2_port, S(1) => 
                           PTMP_2_1_port, S(0) => PTMP_2_0_port, Co => n_1283);
   ADDER_4 : RCA_NBIT42 port map( A(41) => PTMP_2_39_port, A(40) => 
                           PTMP_2_39_port, A(39) => PTMP_2_39_port, A(38) => 
                           PTMP_2_38_port, A(37) => PTMP_2_37_port, A(36) => 
                           PTMP_2_36_port, A(35) => PTMP_2_35_port, A(34) => 
                           PTMP_2_34_port, A(33) => PTMP_2_33_port, A(32) => 
                           PTMP_2_32_port, A(31) => PTMP_2_31_port, A(30) => 
                           PTMP_2_30_port, A(29) => PTMP_2_29_port, A(28) => 
                           PTMP_2_28_port, A(27) => PTMP_2_27_port, A(26) => 
                           PTMP_2_26_port, A(25) => PTMP_2_25_port, A(24) => 
                           PTMP_2_24_port, A(23) => PTMP_2_23_port, A(22) => 
                           PTMP_2_22_port, A(21) => PTMP_2_21_port, A(20) => 
                           PTMP_2_20_port, A(19) => PTMP_2_19_port, A(18) => 
                           PTMP_2_18_port, A(17) => PTMP_2_17_port, A(16) => 
                           PTMP_2_16_port, A(15) => PTMP_2_15_port, A(14) => 
                           PTMP_2_14_port, A(13) => PTMP_2_13_port, A(12) => 
                           PTMP_2_12_port, A(11) => PTMP_2_11_port, A(10) => 
                           PTMP_2_10_port, A(9) => PTMP_2_9_port, A(8) => 
                           PTMP_2_8_port, A(7) => PTMP_2_7_port, A(6) => 
                           PTMP_2_6_port, A(5) => PTMP_2_5_port, A(4) => 
                           PTMP_2_4_port, A(3) => PTMP_2_3_port, A(2) => 
                           PTMP_2_2_port, A(1) => PTMP_2_1_port, A(0) => 
                           PTMP_2_0_port, B(41) => OTMP_4_41_port, B(40) => 
                           OTMP_4_40_port, B(39) => OTMP_4_39_port, B(38) => 
                           OTMP_4_38_port, B(37) => OTMP_4_37_port, B(36) => 
                           OTMP_4_36_port, B(35) => OTMP_4_35_port, B(34) => 
                           OTMP_4_34_port, B(33) => OTMP_4_33_port, B(32) => 
                           OTMP_4_32_port, B(31) => OTMP_4_31_port, B(30) => 
                           OTMP_4_30_port, B(29) => OTMP_4_29_port, B(28) => 
                           OTMP_4_28_port, B(27) => OTMP_4_27_port, B(26) => 
                           OTMP_4_26_port, B(25) => OTMP_4_25_port, B(24) => 
                           OTMP_4_24_port, B(23) => OTMP_4_23_port, B(22) => 
                           OTMP_4_22_port, B(21) => OTMP_4_21_port, B(20) => 
                           OTMP_4_20_port, B(19) => OTMP_4_19_port, B(18) => 
                           OTMP_4_18_port, B(17) => OTMP_4_17_port, B(16) => 
                           OTMP_4_16_port, B(15) => OTMP_4_15_port, B(14) => 
                           OTMP_4_14_port, B(13) => OTMP_4_13_port, B(12) => 
                           OTMP_4_12_port, B(11) => OTMP_4_11_port, B(10) => 
                           OTMP_4_10_port, B(9) => OTMP_4_9_port, B(8) => 
                           OTMP_4_8_port, B(7) => OTMP_4_7_port, B(6) => 
                           OTMP_4_6_port, B(5) => OTMP_4_5_port, B(4) => 
                           OTMP_4_4_port, B(3) => OTMP_4_3_port, B(2) => 
                           OTMP_4_2_port, B(1) => OTMP_4_1_port, B(0) => 
                           OTMP_4_0_port, Ci => X_Logic0_port, S(41) => 
                           PTMP_3_41_port, S(40) => PTMP_3_40_port, S(39) => 
                           PTMP_3_39_port, S(38) => PTMP_3_38_port, S(37) => 
                           PTMP_3_37_port, S(36) => PTMP_3_36_port, S(35) => 
                           PTMP_3_35_port, S(34) => PTMP_3_34_port, S(33) => 
                           PTMP_3_33_port, S(32) => PTMP_3_32_port, S(31) => 
                           PTMP_3_31_port, S(30) => PTMP_3_30_port, S(29) => 
                           PTMP_3_29_port, S(28) => PTMP_3_28_port, S(27) => 
                           PTMP_3_27_port, S(26) => PTMP_3_26_port, S(25) => 
                           PTMP_3_25_port, S(24) => PTMP_3_24_port, S(23) => 
                           PTMP_3_23_port, S(22) => PTMP_3_22_port, S(21) => 
                           PTMP_3_21_port, S(20) => PTMP_3_20_port, S(19) => 
                           PTMP_3_19_port, S(18) => PTMP_3_18_port, S(17) => 
                           PTMP_3_17_port, S(16) => PTMP_3_16_port, S(15) => 
                           PTMP_3_15_port, S(14) => PTMP_3_14_port, S(13) => 
                           PTMP_3_13_port, S(12) => PTMP_3_12_port, S(11) => 
                           PTMP_3_11_port, S(10) => PTMP_3_10_port, S(9) => 
                           PTMP_3_9_port, S(8) => PTMP_3_8_port, S(7) => 
                           PTMP_3_7_port, S(6) => PTMP_3_6_port, S(5) => 
                           PTMP_3_5_port, S(4) => PTMP_3_4_port, S(3) => 
                           PTMP_3_3_port, S(2) => PTMP_3_2_port, S(1) => 
                           PTMP_3_1_port, S(0) => PTMP_3_0_port, Co => n_1284);
   ADDER_5 : RCA_NBIT44 port map( A(43) => PTMP_3_41_port, A(42) => 
                           PTMP_3_41_port, A(41) => PTMP_3_41_port, A(40) => 
                           PTMP_3_40_port, A(39) => PTMP_3_39_port, A(38) => 
                           PTMP_3_38_port, A(37) => PTMP_3_37_port, A(36) => 
                           PTMP_3_36_port, A(35) => PTMP_3_35_port, A(34) => 
                           PTMP_3_34_port, A(33) => PTMP_3_33_port, A(32) => 
                           PTMP_3_32_port, A(31) => PTMP_3_31_port, A(30) => 
                           PTMP_3_30_port, A(29) => PTMP_3_29_port, A(28) => 
                           PTMP_3_28_port, A(27) => PTMP_3_27_port, A(26) => 
                           PTMP_3_26_port, A(25) => PTMP_3_25_port, A(24) => 
                           PTMP_3_24_port, A(23) => PTMP_3_23_port, A(22) => 
                           PTMP_3_22_port, A(21) => PTMP_3_21_port, A(20) => 
                           PTMP_3_20_port, A(19) => PTMP_3_19_port, A(18) => 
                           PTMP_3_18_port, A(17) => PTMP_3_17_port, A(16) => 
                           PTMP_3_16_port, A(15) => PTMP_3_15_port, A(14) => 
                           PTMP_3_14_port, A(13) => PTMP_3_13_port, A(12) => 
                           PTMP_3_12_port, A(11) => PTMP_3_11_port, A(10) => 
                           PTMP_3_10_port, A(9) => PTMP_3_9_port, A(8) => 
                           PTMP_3_8_port, A(7) => PTMP_3_7_port, A(6) => 
                           PTMP_3_6_port, A(5) => PTMP_3_5_port, A(4) => 
                           PTMP_3_4_port, A(3) => PTMP_3_3_port, A(2) => 
                           PTMP_3_2_port, A(1) => PTMP_3_1_port, A(0) => 
                           PTMP_3_0_port, B(43) => OTMP_5_43_port, B(42) => 
                           OTMP_5_42_port, B(41) => OTMP_5_41_port, B(40) => 
                           OTMP_5_40_port, B(39) => OTMP_5_39_port, B(38) => 
                           OTMP_5_38_port, B(37) => OTMP_5_37_port, B(36) => 
                           OTMP_5_36_port, B(35) => OTMP_5_35_port, B(34) => 
                           OTMP_5_34_port, B(33) => OTMP_5_33_port, B(32) => 
                           OTMP_5_32_port, B(31) => OTMP_5_31_port, B(30) => 
                           OTMP_5_30_port, B(29) => OTMP_5_29_port, B(28) => 
                           OTMP_5_28_port, B(27) => OTMP_5_27_port, B(26) => 
                           OTMP_5_26_port, B(25) => OTMP_5_25_port, B(24) => 
                           OTMP_5_24_port, B(23) => OTMP_5_23_port, B(22) => 
                           OTMP_5_22_port, B(21) => OTMP_5_21_port, B(20) => 
                           OTMP_5_20_port, B(19) => OTMP_5_19_port, B(18) => 
                           OTMP_5_18_port, B(17) => OTMP_5_17_port, B(16) => 
                           OTMP_5_16_port, B(15) => OTMP_5_15_port, B(14) => 
                           OTMP_5_14_port, B(13) => OTMP_5_13_port, B(12) => 
                           OTMP_5_12_port, B(11) => OTMP_5_11_port, B(10) => 
                           OTMP_5_10_port, B(9) => OTMP_5_9_port, B(8) => 
                           OTMP_5_8_port, B(7) => OTMP_5_7_port, B(6) => 
                           OTMP_5_6_port, B(5) => OTMP_5_5_port, B(4) => 
                           OTMP_5_4_port, B(3) => OTMP_5_3_port, B(2) => 
                           OTMP_5_2_port, B(1) => OTMP_5_1_port, B(0) => 
                           OTMP_5_0_port, Ci => X_Logic0_port, S(43) => 
                           PTMP_4_43_port, S(42) => PTMP_4_42_port, S(41) => 
                           PTMP_4_41_port, S(40) => PTMP_4_40_port, S(39) => 
                           PTMP_4_39_port, S(38) => PTMP_4_38_port, S(37) => 
                           PTMP_4_37_port, S(36) => PTMP_4_36_port, S(35) => 
                           PTMP_4_35_port, S(34) => PTMP_4_34_port, S(33) => 
                           PTMP_4_33_port, S(32) => PTMP_4_32_port, S(31) => 
                           PTMP_4_31_port, S(30) => PTMP_4_30_port, S(29) => 
                           PTMP_4_29_port, S(28) => PTMP_4_28_port, S(27) => 
                           PTMP_4_27_port, S(26) => PTMP_4_26_port, S(25) => 
                           PTMP_4_25_port, S(24) => PTMP_4_24_port, S(23) => 
                           PTMP_4_23_port, S(22) => PTMP_4_22_port, S(21) => 
                           PTMP_4_21_port, S(20) => PTMP_4_20_port, S(19) => 
                           PTMP_4_19_port, S(18) => PTMP_4_18_port, S(17) => 
                           PTMP_4_17_port, S(16) => PTMP_4_16_port, S(15) => 
                           PTMP_4_15_port, S(14) => PTMP_4_14_port, S(13) => 
                           PTMP_4_13_port, S(12) => PTMP_4_12_port, S(11) => 
                           PTMP_4_11_port, S(10) => PTMP_4_10_port, S(9) => 
                           PTMP_4_9_port, S(8) => PTMP_4_8_port, S(7) => 
                           PTMP_4_7_port, S(6) => PTMP_4_6_port, S(5) => 
                           PTMP_4_5_port, S(4) => PTMP_4_4_port, S(3) => 
                           PTMP_4_3_port, S(2) => PTMP_4_2_port, S(1) => 
                           PTMP_4_1_port, S(0) => PTMP_4_0_port, Co => n_1285);
   ADDER_6 : RCA_NBIT46 port map( A(45) => PTMP_4_43_port, A(44) => 
                           PTMP_4_43_port, A(43) => PTMP_4_43_port, A(42) => 
                           PTMP_4_42_port, A(41) => PTMP_4_41_port, A(40) => 
                           PTMP_4_40_port, A(39) => PTMP_4_39_port, A(38) => 
                           PTMP_4_38_port, A(37) => PTMP_4_37_port, A(36) => 
                           PTMP_4_36_port, A(35) => PTMP_4_35_port, A(34) => 
                           PTMP_4_34_port, A(33) => PTMP_4_33_port, A(32) => 
                           PTMP_4_32_port, A(31) => PTMP_4_31_port, A(30) => 
                           PTMP_4_30_port, A(29) => PTMP_4_29_port, A(28) => 
                           PTMP_4_28_port, A(27) => PTMP_4_27_port, A(26) => 
                           PTMP_4_26_port, A(25) => PTMP_4_25_port, A(24) => 
                           PTMP_4_24_port, A(23) => PTMP_4_23_port, A(22) => 
                           PTMP_4_22_port, A(21) => PTMP_4_21_port, A(20) => 
                           PTMP_4_20_port, A(19) => PTMP_4_19_port, A(18) => 
                           PTMP_4_18_port, A(17) => PTMP_4_17_port, A(16) => 
                           PTMP_4_16_port, A(15) => PTMP_4_15_port, A(14) => 
                           PTMP_4_14_port, A(13) => PTMP_4_13_port, A(12) => 
                           PTMP_4_12_port, A(11) => PTMP_4_11_port, A(10) => 
                           PTMP_4_10_port, A(9) => PTMP_4_9_port, A(8) => 
                           PTMP_4_8_port, A(7) => PTMP_4_7_port, A(6) => 
                           PTMP_4_6_port, A(5) => PTMP_4_5_port, A(4) => 
                           PTMP_4_4_port, A(3) => PTMP_4_3_port, A(2) => 
                           PTMP_4_2_port, A(1) => PTMP_4_1_port, A(0) => 
                           PTMP_4_0_port, B(45) => OTMP_6_45_port, B(44) => 
                           OTMP_6_44_port, B(43) => OTMP_6_43_port, B(42) => 
                           OTMP_6_42_port, B(41) => OTMP_6_41_port, B(40) => 
                           OTMP_6_40_port, B(39) => OTMP_6_39_port, B(38) => 
                           OTMP_6_38_port, B(37) => OTMP_6_37_port, B(36) => 
                           OTMP_6_36_port, B(35) => OTMP_6_35_port, B(34) => 
                           OTMP_6_34_port, B(33) => OTMP_6_33_port, B(32) => 
                           OTMP_6_32_port, B(31) => OTMP_6_31_port, B(30) => 
                           OTMP_6_30_port, B(29) => OTMP_6_29_port, B(28) => 
                           OTMP_6_28_port, B(27) => OTMP_6_27_port, B(26) => 
                           OTMP_6_26_port, B(25) => OTMP_6_25_port, B(24) => 
                           OTMP_6_24_port, B(23) => OTMP_6_23_port, B(22) => 
                           OTMP_6_22_port, B(21) => OTMP_6_21_port, B(20) => 
                           OTMP_6_20_port, B(19) => OTMP_6_19_port, B(18) => 
                           OTMP_6_18_port, B(17) => OTMP_6_17_port, B(16) => 
                           OTMP_6_16_port, B(15) => OTMP_6_15_port, B(14) => 
                           OTMP_6_14_port, B(13) => OTMP_6_13_port, B(12) => 
                           OTMP_6_12_port, B(11) => OTMP_6_11_port, B(10) => 
                           OTMP_6_10_port, B(9) => OTMP_6_9_port, B(8) => 
                           OTMP_6_8_port, B(7) => OTMP_6_7_port, B(6) => 
                           OTMP_6_6_port, B(5) => OTMP_6_5_port, B(4) => 
                           OTMP_6_4_port, B(3) => OTMP_6_3_port, B(2) => 
                           OTMP_6_2_port, B(1) => OTMP_6_1_port, B(0) => 
                           OTMP_6_0_port, Ci => X_Logic0_port, S(45) => 
                           PTMP_5_45_port, S(44) => PTMP_5_44_port, S(43) => 
                           PTMP_5_43_port, S(42) => PTMP_5_42_port, S(41) => 
                           PTMP_5_41_port, S(40) => PTMP_5_40_port, S(39) => 
                           PTMP_5_39_port, S(38) => PTMP_5_38_port, S(37) => 
                           PTMP_5_37_port, S(36) => PTMP_5_36_port, S(35) => 
                           PTMP_5_35_port, S(34) => PTMP_5_34_port, S(33) => 
                           PTMP_5_33_port, S(32) => PTMP_5_32_port, S(31) => 
                           PTMP_5_31_port, S(30) => PTMP_5_30_port, S(29) => 
                           PTMP_5_29_port, S(28) => PTMP_5_28_port, S(27) => 
                           PTMP_5_27_port, S(26) => PTMP_5_26_port, S(25) => 
                           PTMP_5_25_port, S(24) => PTMP_5_24_port, S(23) => 
                           PTMP_5_23_port, S(22) => PTMP_5_22_port, S(21) => 
                           PTMP_5_21_port, S(20) => PTMP_5_20_port, S(19) => 
                           PTMP_5_19_port, S(18) => PTMP_5_18_port, S(17) => 
                           PTMP_5_17_port, S(16) => PTMP_5_16_port, S(15) => 
                           PTMP_5_15_port, S(14) => PTMP_5_14_port, S(13) => 
                           PTMP_5_13_port, S(12) => PTMP_5_12_port, S(11) => 
                           PTMP_5_11_port, S(10) => PTMP_5_10_port, S(9) => 
                           PTMP_5_9_port, S(8) => PTMP_5_8_port, S(7) => 
                           PTMP_5_7_port, S(6) => PTMP_5_6_port, S(5) => 
                           PTMP_5_5_port, S(4) => PTMP_5_4_port, S(3) => 
                           PTMP_5_3_port, S(2) => PTMP_5_2_port, S(1) => 
                           PTMP_5_1_port, S(0) => PTMP_5_0_port, Co => n_1286);
   ADDER_7 : RCA_NBIT48 port map( A(47) => PTMP_5_45_port, A(46) => 
                           PTMP_5_45_port, A(45) => PTMP_5_45_port, A(44) => 
                           PTMP_5_44_port, A(43) => PTMP_5_43_port, A(42) => 
                           PTMP_5_42_port, A(41) => PTMP_5_41_port, A(40) => 
                           PTMP_5_40_port, A(39) => PTMP_5_39_port, A(38) => 
                           PTMP_5_38_port, A(37) => PTMP_5_37_port, A(36) => 
                           PTMP_5_36_port, A(35) => PTMP_5_35_port, A(34) => 
                           PTMP_5_34_port, A(33) => PTMP_5_33_port, A(32) => 
                           PTMP_5_32_port, A(31) => PTMP_5_31_port, A(30) => 
                           PTMP_5_30_port, A(29) => PTMP_5_29_port, A(28) => 
                           PTMP_5_28_port, A(27) => PTMP_5_27_port, A(26) => 
                           PTMP_5_26_port, A(25) => PTMP_5_25_port, A(24) => 
                           PTMP_5_24_port, A(23) => PTMP_5_23_port, A(22) => 
                           PTMP_5_22_port, A(21) => PTMP_5_21_port, A(20) => 
                           PTMP_5_20_port, A(19) => PTMP_5_19_port, A(18) => 
                           PTMP_5_18_port, A(17) => PTMP_5_17_port, A(16) => 
                           PTMP_5_16_port, A(15) => PTMP_5_15_port, A(14) => 
                           PTMP_5_14_port, A(13) => PTMP_5_13_port, A(12) => 
                           PTMP_5_12_port, A(11) => PTMP_5_11_port, A(10) => 
                           PTMP_5_10_port, A(9) => PTMP_5_9_port, A(8) => 
                           PTMP_5_8_port, A(7) => PTMP_5_7_port, A(6) => 
                           PTMP_5_6_port, A(5) => PTMP_5_5_port, A(4) => 
                           PTMP_5_4_port, A(3) => PTMP_5_3_port, A(2) => 
                           PTMP_5_2_port, A(1) => PTMP_5_1_port, A(0) => 
                           PTMP_5_0_port, B(47) => OTMP_7_47_port, B(46) => 
                           OTMP_7_46_port, B(45) => OTMP_7_45_port, B(44) => 
                           OTMP_7_44_port, B(43) => OTMP_7_43_port, B(42) => 
                           OTMP_7_42_port, B(41) => OTMP_7_41_port, B(40) => 
                           OTMP_7_40_port, B(39) => OTMP_7_39_port, B(38) => 
                           OTMP_7_38_port, B(37) => OTMP_7_37_port, B(36) => 
                           OTMP_7_36_port, B(35) => OTMP_7_35_port, B(34) => 
                           OTMP_7_34_port, B(33) => OTMP_7_33_port, B(32) => 
                           OTMP_7_32_port, B(31) => OTMP_7_31_port, B(30) => 
                           OTMP_7_30_port, B(29) => OTMP_7_29_port, B(28) => 
                           OTMP_7_28_port, B(27) => OTMP_7_27_port, B(26) => 
                           OTMP_7_26_port, B(25) => OTMP_7_25_port, B(24) => 
                           OTMP_7_24_port, B(23) => OTMP_7_23_port, B(22) => 
                           OTMP_7_22_port, B(21) => OTMP_7_21_port, B(20) => 
                           OTMP_7_20_port, B(19) => OTMP_7_19_port, B(18) => 
                           OTMP_7_18_port, B(17) => OTMP_7_17_port, B(16) => 
                           OTMP_7_16_port, B(15) => OTMP_7_15_port, B(14) => 
                           OTMP_7_14_port, B(13) => OTMP_7_13_port, B(12) => 
                           OTMP_7_12_port, B(11) => OTMP_7_11_port, B(10) => 
                           OTMP_7_10_port, B(9) => OTMP_7_9_port, B(8) => 
                           OTMP_7_8_port, B(7) => OTMP_7_7_port, B(6) => 
                           OTMP_7_6_port, B(5) => OTMP_7_5_port, B(4) => 
                           OTMP_7_4_port, B(3) => OTMP_7_3_port, B(2) => 
                           OTMP_7_2_port, B(1) => OTMP_7_1_port, B(0) => 
                           OTMP_7_0_port, Ci => X_Logic0_port, S(47) => 
                           PTMP_6_47_port, S(46) => PTMP_6_46_port, S(45) => 
                           PTMP_6_45_port, S(44) => PTMP_6_44_port, S(43) => 
                           PTMP_6_43_port, S(42) => PTMP_6_42_port, S(41) => 
                           PTMP_6_41_port, S(40) => PTMP_6_40_port, S(39) => 
                           PTMP_6_39_port, S(38) => PTMP_6_38_port, S(37) => 
                           PTMP_6_37_port, S(36) => PTMP_6_36_port, S(35) => 
                           PTMP_6_35_port, S(34) => PTMP_6_34_port, S(33) => 
                           PTMP_6_33_port, S(32) => PTMP_6_32_port, S(31) => 
                           PTMP_6_31_port, S(30) => PTMP_6_30_port, S(29) => 
                           PTMP_6_29_port, S(28) => PTMP_6_28_port, S(27) => 
                           PTMP_6_27_port, S(26) => PTMP_6_26_port, S(25) => 
                           PTMP_6_25_port, S(24) => PTMP_6_24_port, S(23) => 
                           PTMP_6_23_port, S(22) => PTMP_6_22_port, S(21) => 
                           PTMP_6_21_port, S(20) => PTMP_6_20_port, S(19) => 
                           PTMP_6_19_port, S(18) => PTMP_6_18_port, S(17) => 
                           PTMP_6_17_port, S(16) => PTMP_6_16_port, S(15) => 
                           PTMP_6_15_port, S(14) => PTMP_6_14_port, S(13) => 
                           PTMP_6_13_port, S(12) => PTMP_6_12_port, S(11) => 
                           PTMP_6_11_port, S(10) => PTMP_6_10_port, S(9) => 
                           PTMP_6_9_port, S(8) => PTMP_6_8_port, S(7) => 
                           PTMP_6_7_port, S(6) => PTMP_6_6_port, S(5) => 
                           PTMP_6_5_port, S(4) => PTMP_6_4_port, S(3) => 
                           PTMP_6_3_port, S(2) => PTMP_6_2_port, S(1) => 
                           PTMP_6_1_port, S(0) => PTMP_6_0_port, Co => n_1287);
   ADDER_8 : RCA_NBIT50 port map( A(49) => PTMP_6_47_port, A(48) => 
                           PTMP_6_47_port, A(47) => PTMP_6_47_port, A(46) => 
                           PTMP_6_46_port, A(45) => PTMP_6_45_port, A(44) => 
                           PTMP_6_44_port, A(43) => PTMP_6_43_port, A(42) => 
                           PTMP_6_42_port, A(41) => PTMP_6_41_port, A(40) => 
                           PTMP_6_40_port, A(39) => PTMP_6_39_port, A(38) => 
                           PTMP_6_38_port, A(37) => PTMP_6_37_port, A(36) => 
                           PTMP_6_36_port, A(35) => PTMP_6_35_port, A(34) => 
                           PTMP_6_34_port, A(33) => PTMP_6_33_port, A(32) => 
                           PTMP_6_32_port, A(31) => PTMP_6_31_port, A(30) => 
                           PTMP_6_30_port, A(29) => PTMP_6_29_port, A(28) => 
                           PTMP_6_28_port, A(27) => PTMP_6_27_port, A(26) => 
                           PTMP_6_26_port, A(25) => PTMP_6_25_port, A(24) => 
                           PTMP_6_24_port, A(23) => PTMP_6_23_port, A(22) => 
                           PTMP_6_22_port, A(21) => PTMP_6_21_port, A(20) => 
                           PTMP_6_20_port, A(19) => PTMP_6_19_port, A(18) => 
                           PTMP_6_18_port, A(17) => PTMP_6_17_port, A(16) => 
                           PTMP_6_16_port, A(15) => PTMP_6_15_port, A(14) => 
                           PTMP_6_14_port, A(13) => PTMP_6_13_port, A(12) => 
                           PTMP_6_12_port, A(11) => PTMP_6_11_port, A(10) => 
                           PTMP_6_10_port, A(9) => PTMP_6_9_port, A(8) => 
                           PTMP_6_8_port, A(7) => PTMP_6_7_port, A(6) => 
                           PTMP_6_6_port, A(5) => PTMP_6_5_port, A(4) => 
                           PTMP_6_4_port, A(3) => PTMP_6_3_port, A(2) => 
                           PTMP_6_2_port, A(1) => PTMP_6_1_port, A(0) => 
                           PTMP_6_0_port, B(49) => OTMP_8_49_port, B(48) => 
                           OTMP_8_48_port, B(47) => OTMP_8_47_port, B(46) => 
                           OTMP_8_46_port, B(45) => OTMP_8_45_port, B(44) => 
                           OTMP_8_44_port, B(43) => OTMP_8_43_port, B(42) => 
                           OTMP_8_42_port, B(41) => OTMP_8_41_port, B(40) => 
                           OTMP_8_40_port, B(39) => OTMP_8_39_port, B(38) => 
                           OTMP_8_38_port, B(37) => OTMP_8_37_port, B(36) => 
                           OTMP_8_36_port, B(35) => OTMP_8_35_port, B(34) => 
                           OTMP_8_34_port, B(33) => OTMP_8_33_port, B(32) => 
                           OTMP_8_32_port, B(31) => OTMP_8_31_port, B(30) => 
                           OTMP_8_30_port, B(29) => OTMP_8_29_port, B(28) => 
                           OTMP_8_28_port, B(27) => OTMP_8_27_port, B(26) => 
                           OTMP_8_26_port, B(25) => OTMP_8_25_port, B(24) => 
                           OTMP_8_24_port, B(23) => OTMP_8_23_port, B(22) => 
                           OTMP_8_22_port, B(21) => OTMP_8_21_port, B(20) => 
                           OTMP_8_20_port, B(19) => OTMP_8_19_port, B(18) => 
                           OTMP_8_18_port, B(17) => OTMP_8_17_port, B(16) => 
                           OTMP_8_16_port, B(15) => OTMP_8_15_port, B(14) => 
                           OTMP_8_14_port, B(13) => OTMP_8_13_port, B(12) => 
                           OTMP_8_12_port, B(11) => OTMP_8_11_port, B(10) => 
                           OTMP_8_10_port, B(9) => OTMP_8_9_port, B(8) => 
                           OTMP_8_8_port, B(7) => OTMP_8_7_port, B(6) => 
                           OTMP_8_6_port, B(5) => OTMP_8_5_port, B(4) => 
                           OTMP_8_4_port, B(3) => OTMP_8_3_port, B(2) => 
                           OTMP_8_2_port, B(1) => OTMP_8_1_port, B(0) => 
                           OTMP_8_0_port, Ci => X_Logic0_port, S(49) => 
                           PTMP_7_49_port, S(48) => PTMP_7_48_port, S(47) => 
                           PTMP_7_47_port, S(46) => PTMP_7_46_port, S(45) => 
                           PTMP_7_45_port, S(44) => PTMP_7_44_port, S(43) => 
                           PTMP_7_43_port, S(42) => PTMP_7_42_port, S(41) => 
                           PTMP_7_41_port, S(40) => PTMP_7_40_port, S(39) => 
                           PTMP_7_39_port, S(38) => PTMP_7_38_port, S(37) => 
                           PTMP_7_37_port, S(36) => PTMP_7_36_port, S(35) => 
                           PTMP_7_35_port, S(34) => PTMP_7_34_port, S(33) => 
                           PTMP_7_33_port, S(32) => PTMP_7_32_port, S(31) => 
                           PTMP_7_31_port, S(30) => PTMP_7_30_port, S(29) => 
                           PTMP_7_29_port, S(28) => PTMP_7_28_port, S(27) => 
                           PTMP_7_27_port, S(26) => PTMP_7_26_port, S(25) => 
                           PTMP_7_25_port, S(24) => PTMP_7_24_port, S(23) => 
                           PTMP_7_23_port, S(22) => PTMP_7_22_port, S(21) => 
                           PTMP_7_21_port, S(20) => PTMP_7_20_port, S(19) => 
                           PTMP_7_19_port, S(18) => PTMP_7_18_port, S(17) => 
                           PTMP_7_17_port, S(16) => PTMP_7_16_port, S(15) => 
                           PTMP_7_15_port, S(14) => PTMP_7_14_port, S(13) => 
                           PTMP_7_13_port, S(12) => PTMP_7_12_port, S(11) => 
                           PTMP_7_11_port, S(10) => PTMP_7_10_port, S(9) => 
                           PTMP_7_9_port, S(8) => PTMP_7_8_port, S(7) => 
                           PTMP_7_7_port, S(6) => PTMP_7_6_port, S(5) => 
                           PTMP_7_5_port, S(4) => PTMP_7_4_port, S(3) => 
                           PTMP_7_3_port, S(2) => PTMP_7_2_port, S(1) => 
                           PTMP_7_1_port, S(0) => PTMP_7_0_port, Co => n_1288);
   ADDER_9 : RCA_NBIT52 port map( A(51) => PTMP_7_49_port, A(50) => 
                           PTMP_7_49_port, A(49) => PTMP_7_49_port, A(48) => 
                           PTMP_7_48_port, A(47) => PTMP_7_47_port, A(46) => 
                           PTMP_7_46_port, A(45) => PTMP_7_45_port, A(44) => 
                           PTMP_7_44_port, A(43) => PTMP_7_43_port, A(42) => 
                           PTMP_7_42_port, A(41) => PTMP_7_41_port, A(40) => 
                           PTMP_7_40_port, A(39) => PTMP_7_39_port, A(38) => 
                           PTMP_7_38_port, A(37) => PTMP_7_37_port, A(36) => 
                           PTMP_7_36_port, A(35) => PTMP_7_35_port, A(34) => 
                           PTMP_7_34_port, A(33) => PTMP_7_33_port, A(32) => 
                           PTMP_7_32_port, A(31) => PTMP_7_31_port, A(30) => 
                           PTMP_7_30_port, A(29) => PTMP_7_29_port, A(28) => 
                           PTMP_7_28_port, A(27) => PTMP_7_27_port, A(26) => 
                           PTMP_7_26_port, A(25) => PTMP_7_25_port, A(24) => 
                           PTMP_7_24_port, A(23) => PTMP_7_23_port, A(22) => 
                           PTMP_7_22_port, A(21) => PTMP_7_21_port, A(20) => 
                           PTMP_7_20_port, A(19) => PTMP_7_19_port, A(18) => 
                           PTMP_7_18_port, A(17) => PTMP_7_17_port, A(16) => 
                           PTMP_7_16_port, A(15) => PTMP_7_15_port, A(14) => 
                           PTMP_7_14_port, A(13) => PTMP_7_13_port, A(12) => 
                           PTMP_7_12_port, A(11) => PTMP_7_11_port, A(10) => 
                           PTMP_7_10_port, A(9) => PTMP_7_9_port, A(8) => 
                           PTMP_7_8_port, A(7) => PTMP_7_7_port, A(6) => 
                           PTMP_7_6_port, A(5) => PTMP_7_5_port, A(4) => 
                           PTMP_7_4_port, A(3) => PTMP_7_3_port, A(2) => 
                           PTMP_7_2_port, A(1) => PTMP_7_1_port, A(0) => 
                           PTMP_7_0_port, B(51) => OTMP_9_51_port, B(50) => 
                           OTMP_9_50_port, B(49) => OTMP_9_49_port, B(48) => 
                           OTMP_9_48_port, B(47) => OTMP_9_47_port, B(46) => 
                           OTMP_9_46_port, B(45) => OTMP_9_45_port, B(44) => 
                           OTMP_9_44_port, B(43) => OTMP_9_43_port, B(42) => 
                           OTMP_9_42_port, B(41) => OTMP_9_41_port, B(40) => 
                           OTMP_9_40_port, B(39) => OTMP_9_39_port, B(38) => 
                           OTMP_9_38_port, B(37) => OTMP_9_37_port, B(36) => 
                           OTMP_9_36_port, B(35) => OTMP_9_35_port, B(34) => 
                           OTMP_9_34_port, B(33) => OTMP_9_33_port, B(32) => 
                           OTMP_9_32_port, B(31) => OTMP_9_31_port, B(30) => 
                           OTMP_9_30_port, B(29) => OTMP_9_29_port, B(28) => 
                           OTMP_9_28_port, B(27) => OTMP_9_27_port, B(26) => 
                           OTMP_9_26_port, B(25) => OTMP_9_25_port, B(24) => 
                           OTMP_9_24_port, B(23) => OTMP_9_23_port, B(22) => 
                           OTMP_9_22_port, B(21) => OTMP_9_21_port, B(20) => 
                           OTMP_9_20_port, B(19) => OTMP_9_19_port, B(18) => 
                           OTMP_9_18_port, B(17) => OTMP_9_17_port, B(16) => 
                           OTMP_9_16_port, B(15) => OTMP_9_15_port, B(14) => 
                           OTMP_9_14_port, B(13) => OTMP_9_13_port, B(12) => 
                           OTMP_9_12_port, B(11) => OTMP_9_11_port, B(10) => 
                           OTMP_9_10_port, B(9) => OTMP_9_9_port, B(8) => 
                           OTMP_9_8_port, B(7) => OTMP_9_7_port, B(6) => 
                           OTMP_9_6_port, B(5) => OTMP_9_5_port, B(4) => 
                           OTMP_9_4_port, B(3) => OTMP_9_3_port, B(2) => 
                           OTMP_9_2_port, B(1) => OTMP_9_1_port, B(0) => 
                           OTMP_9_0_port, Ci => X_Logic0_port, S(51) => 
                           PTMP_8_51_port, S(50) => PTMP_8_50_port, S(49) => 
                           PTMP_8_49_port, S(48) => PTMP_8_48_port, S(47) => 
                           PTMP_8_47_port, S(46) => PTMP_8_46_port, S(45) => 
                           PTMP_8_45_port, S(44) => PTMP_8_44_port, S(43) => 
                           PTMP_8_43_port, S(42) => PTMP_8_42_port, S(41) => 
                           PTMP_8_41_port, S(40) => PTMP_8_40_port, S(39) => 
                           PTMP_8_39_port, S(38) => PTMP_8_38_port, S(37) => 
                           PTMP_8_37_port, S(36) => PTMP_8_36_port, S(35) => 
                           PTMP_8_35_port, S(34) => PTMP_8_34_port, S(33) => 
                           PTMP_8_33_port, S(32) => PTMP_8_32_port, S(31) => 
                           PTMP_8_31_port, S(30) => PTMP_8_30_port, S(29) => 
                           PTMP_8_29_port, S(28) => PTMP_8_28_port, S(27) => 
                           PTMP_8_27_port, S(26) => PTMP_8_26_port, S(25) => 
                           PTMP_8_25_port, S(24) => PTMP_8_24_port, S(23) => 
                           PTMP_8_23_port, S(22) => PTMP_8_22_port, S(21) => 
                           PTMP_8_21_port, S(20) => PTMP_8_20_port, S(19) => 
                           PTMP_8_19_port, S(18) => PTMP_8_18_port, S(17) => 
                           PTMP_8_17_port, S(16) => PTMP_8_16_port, S(15) => 
                           PTMP_8_15_port, S(14) => PTMP_8_14_port, S(13) => 
                           PTMP_8_13_port, S(12) => PTMP_8_12_port, S(11) => 
                           PTMP_8_11_port, S(10) => PTMP_8_10_port, S(9) => 
                           PTMP_8_9_port, S(8) => PTMP_8_8_port, S(7) => 
                           PTMP_8_7_port, S(6) => PTMP_8_6_port, S(5) => 
                           PTMP_8_5_port, S(4) => PTMP_8_4_port, S(3) => 
                           PTMP_8_3_port, S(2) => PTMP_8_2_port, S(1) => 
                           PTMP_8_1_port, S(0) => PTMP_8_0_port, Co => n_1289);
   ADDER_10 : RCA_NBIT54 port map( A(53) => PTMP_8_51_port, A(52) => 
                           PTMP_8_51_port, A(51) => PTMP_8_51_port, A(50) => 
                           PTMP_8_50_port, A(49) => PTMP_8_49_port, A(48) => 
                           PTMP_8_48_port, A(47) => PTMP_8_47_port, A(46) => 
                           PTMP_8_46_port, A(45) => PTMP_8_45_port, A(44) => 
                           PTMP_8_44_port, A(43) => PTMP_8_43_port, A(42) => 
                           PTMP_8_42_port, A(41) => PTMP_8_41_port, A(40) => 
                           PTMP_8_40_port, A(39) => PTMP_8_39_port, A(38) => 
                           PTMP_8_38_port, A(37) => PTMP_8_37_port, A(36) => 
                           PTMP_8_36_port, A(35) => PTMP_8_35_port, A(34) => 
                           PTMP_8_34_port, A(33) => PTMP_8_33_port, A(32) => 
                           PTMP_8_32_port, A(31) => PTMP_8_31_port, A(30) => 
                           PTMP_8_30_port, A(29) => PTMP_8_29_port, A(28) => 
                           PTMP_8_28_port, A(27) => PTMP_8_27_port, A(26) => 
                           PTMP_8_26_port, A(25) => PTMP_8_25_port, A(24) => 
                           PTMP_8_24_port, A(23) => PTMP_8_23_port, A(22) => 
                           PTMP_8_22_port, A(21) => PTMP_8_21_port, A(20) => 
                           PTMP_8_20_port, A(19) => PTMP_8_19_port, A(18) => 
                           PTMP_8_18_port, A(17) => PTMP_8_17_port, A(16) => 
                           PTMP_8_16_port, A(15) => PTMP_8_15_port, A(14) => 
                           PTMP_8_14_port, A(13) => PTMP_8_13_port, A(12) => 
                           PTMP_8_12_port, A(11) => PTMP_8_11_port, A(10) => 
                           PTMP_8_10_port, A(9) => PTMP_8_9_port, A(8) => 
                           PTMP_8_8_port, A(7) => PTMP_8_7_port, A(6) => 
                           PTMP_8_6_port, A(5) => PTMP_8_5_port, A(4) => 
                           PTMP_8_4_port, A(3) => PTMP_8_3_port, A(2) => 
                           PTMP_8_2_port, A(1) => PTMP_8_1_port, A(0) => 
                           PTMP_8_0_port, B(53) => OTMP_10_53_port, B(52) => 
                           OTMP_10_52_port, B(51) => OTMP_10_51_port, B(50) => 
                           OTMP_10_50_port, B(49) => OTMP_10_49_port, B(48) => 
                           OTMP_10_48_port, B(47) => OTMP_10_47_port, B(46) => 
                           OTMP_10_46_port, B(45) => OTMP_10_45_port, B(44) => 
                           OTMP_10_44_port, B(43) => OTMP_10_43_port, B(42) => 
                           OTMP_10_42_port, B(41) => OTMP_10_41_port, B(40) => 
                           OTMP_10_40_port, B(39) => OTMP_10_39_port, B(38) => 
                           OTMP_10_38_port, B(37) => OTMP_10_37_port, B(36) => 
                           OTMP_10_36_port, B(35) => OTMP_10_35_port, B(34) => 
                           OTMP_10_34_port, B(33) => OTMP_10_33_port, B(32) => 
                           OTMP_10_32_port, B(31) => OTMP_10_31_port, B(30) => 
                           OTMP_10_30_port, B(29) => OTMP_10_29_port, B(28) => 
                           OTMP_10_28_port, B(27) => OTMP_10_27_port, B(26) => 
                           OTMP_10_26_port, B(25) => OTMP_10_25_port, B(24) => 
                           OTMP_10_24_port, B(23) => OTMP_10_23_port, B(22) => 
                           OTMP_10_22_port, B(21) => OTMP_10_21_port, B(20) => 
                           OTMP_10_20_port, B(19) => OTMP_10_19_port, B(18) => 
                           OTMP_10_18_port, B(17) => OTMP_10_17_port, B(16) => 
                           OTMP_10_16_port, B(15) => OTMP_10_15_port, B(14) => 
                           OTMP_10_14_port, B(13) => OTMP_10_13_port, B(12) => 
                           OTMP_10_12_port, B(11) => OTMP_10_11_port, B(10) => 
                           OTMP_10_10_port, B(9) => OTMP_10_9_port, B(8) => 
                           OTMP_10_8_port, B(7) => OTMP_10_7_port, B(6) => 
                           OTMP_10_6_port, B(5) => OTMP_10_5_port, B(4) => 
                           OTMP_10_4_port, B(3) => OTMP_10_3_port, B(2) => 
                           OTMP_10_2_port, B(1) => OTMP_10_1_port, B(0) => 
                           OTMP_10_0_port, Ci => X_Logic0_port, S(53) => 
                           PTMP_9_53_port, S(52) => PTMP_9_52_port, S(51) => 
                           PTMP_9_51_port, S(50) => PTMP_9_50_port, S(49) => 
                           PTMP_9_49_port, S(48) => PTMP_9_48_port, S(47) => 
                           PTMP_9_47_port, S(46) => PTMP_9_46_port, S(45) => 
                           PTMP_9_45_port, S(44) => PTMP_9_44_port, S(43) => 
                           PTMP_9_43_port, S(42) => PTMP_9_42_port, S(41) => 
                           PTMP_9_41_port, S(40) => PTMP_9_40_port, S(39) => 
                           PTMP_9_39_port, S(38) => PTMP_9_38_port, S(37) => 
                           PTMP_9_37_port, S(36) => PTMP_9_36_port, S(35) => 
                           PTMP_9_35_port, S(34) => PTMP_9_34_port, S(33) => 
                           PTMP_9_33_port, S(32) => PTMP_9_32_port, S(31) => 
                           PTMP_9_31_port, S(30) => PTMP_9_30_port, S(29) => 
                           PTMP_9_29_port, S(28) => PTMP_9_28_port, S(27) => 
                           PTMP_9_27_port, S(26) => PTMP_9_26_port, S(25) => 
                           PTMP_9_25_port, S(24) => PTMP_9_24_port, S(23) => 
                           PTMP_9_23_port, S(22) => PTMP_9_22_port, S(21) => 
                           PTMP_9_21_port, S(20) => PTMP_9_20_port, S(19) => 
                           PTMP_9_19_port, S(18) => PTMP_9_18_port, S(17) => 
                           PTMP_9_17_port, S(16) => PTMP_9_16_port, S(15) => 
                           PTMP_9_15_port, S(14) => PTMP_9_14_port, S(13) => 
                           PTMP_9_13_port, S(12) => PTMP_9_12_port, S(11) => 
                           PTMP_9_11_port, S(10) => PTMP_9_10_port, S(9) => 
                           PTMP_9_9_port, S(8) => PTMP_9_8_port, S(7) => 
                           PTMP_9_7_port, S(6) => PTMP_9_6_port, S(5) => 
                           PTMP_9_5_port, S(4) => PTMP_9_4_port, S(3) => 
                           PTMP_9_3_port, S(2) => PTMP_9_2_port, S(1) => 
                           PTMP_9_1_port, S(0) => PTMP_9_0_port, Co => n_1290);
   ADDER_11 : RCA_NBIT56 port map( A(55) => PTMP_9_53_port, A(54) => 
                           PTMP_9_53_port, A(53) => PTMP_9_53_port, A(52) => 
                           PTMP_9_52_port, A(51) => PTMP_9_51_port, A(50) => 
                           PTMP_9_50_port, A(49) => PTMP_9_49_port, A(48) => 
                           PTMP_9_48_port, A(47) => PTMP_9_47_port, A(46) => 
                           PTMP_9_46_port, A(45) => PTMP_9_45_port, A(44) => 
                           PTMP_9_44_port, A(43) => PTMP_9_43_port, A(42) => 
                           PTMP_9_42_port, A(41) => PTMP_9_41_port, A(40) => 
                           PTMP_9_40_port, A(39) => PTMP_9_39_port, A(38) => 
                           PTMP_9_38_port, A(37) => PTMP_9_37_port, A(36) => 
                           PTMP_9_36_port, A(35) => PTMP_9_35_port, A(34) => 
                           PTMP_9_34_port, A(33) => PTMP_9_33_port, A(32) => 
                           PTMP_9_32_port, A(31) => PTMP_9_31_port, A(30) => 
                           PTMP_9_30_port, A(29) => PTMP_9_29_port, A(28) => 
                           PTMP_9_28_port, A(27) => PTMP_9_27_port, A(26) => 
                           PTMP_9_26_port, A(25) => PTMP_9_25_port, A(24) => 
                           PTMP_9_24_port, A(23) => PTMP_9_23_port, A(22) => 
                           PTMP_9_22_port, A(21) => PTMP_9_21_port, A(20) => 
                           PTMP_9_20_port, A(19) => PTMP_9_19_port, A(18) => 
                           PTMP_9_18_port, A(17) => PTMP_9_17_port, A(16) => 
                           PTMP_9_16_port, A(15) => PTMP_9_15_port, A(14) => 
                           PTMP_9_14_port, A(13) => PTMP_9_13_port, A(12) => 
                           PTMP_9_12_port, A(11) => PTMP_9_11_port, A(10) => 
                           PTMP_9_10_port, A(9) => PTMP_9_9_port, A(8) => 
                           PTMP_9_8_port, A(7) => PTMP_9_7_port, A(6) => 
                           PTMP_9_6_port, A(5) => PTMP_9_5_port, A(4) => 
                           PTMP_9_4_port, A(3) => PTMP_9_3_port, A(2) => 
                           PTMP_9_2_port, A(1) => PTMP_9_1_port, A(0) => 
                           PTMP_9_0_port, B(55) => OTMP_11_55_port, B(54) => 
                           OTMP_11_54_port, B(53) => OTMP_11_53_port, B(52) => 
                           OTMP_11_52_port, B(51) => OTMP_11_51_port, B(50) => 
                           OTMP_11_50_port, B(49) => OTMP_11_49_port, B(48) => 
                           OTMP_11_48_port, B(47) => OTMP_11_47_port, B(46) => 
                           OTMP_11_46_port, B(45) => OTMP_11_45_port, B(44) => 
                           OTMP_11_44_port, B(43) => OTMP_11_43_port, B(42) => 
                           OTMP_11_42_port, B(41) => OTMP_11_41_port, B(40) => 
                           OTMP_11_40_port, B(39) => OTMP_11_39_port, B(38) => 
                           OTMP_11_38_port, B(37) => OTMP_11_37_port, B(36) => 
                           OTMP_11_36_port, B(35) => OTMP_11_35_port, B(34) => 
                           OTMP_11_34_port, B(33) => OTMP_11_33_port, B(32) => 
                           OTMP_11_32_port, B(31) => OTMP_11_31_port, B(30) => 
                           OTMP_11_30_port, B(29) => OTMP_11_29_port, B(28) => 
                           OTMP_11_28_port, B(27) => OTMP_11_27_port, B(26) => 
                           OTMP_11_26_port, B(25) => OTMP_11_25_port, B(24) => 
                           OTMP_11_24_port, B(23) => OTMP_11_23_port, B(22) => 
                           OTMP_11_22_port, B(21) => OTMP_11_21_port, B(20) => 
                           OTMP_11_20_port, B(19) => OTMP_11_19_port, B(18) => 
                           OTMP_11_18_port, B(17) => OTMP_11_17_port, B(16) => 
                           OTMP_11_16_port, B(15) => OTMP_11_15_port, B(14) => 
                           OTMP_11_14_port, B(13) => OTMP_11_13_port, B(12) => 
                           OTMP_11_12_port, B(11) => OTMP_11_11_port, B(10) => 
                           OTMP_11_10_port, B(9) => OTMP_11_9_port, B(8) => 
                           OTMP_11_8_port, B(7) => OTMP_11_7_port, B(6) => 
                           OTMP_11_6_port, B(5) => OTMP_11_5_port, B(4) => 
                           OTMP_11_4_port, B(3) => OTMP_11_3_port, B(2) => 
                           OTMP_11_2_port, B(1) => OTMP_11_1_port, B(0) => 
                           OTMP_11_0_port, Ci => X_Logic0_port, S(55) => 
                           PTMP_10_55_port, S(54) => PTMP_10_54_port, S(53) => 
                           PTMP_10_53_port, S(52) => PTMP_10_52_port, S(51) => 
                           PTMP_10_51_port, S(50) => PTMP_10_50_port, S(49) => 
                           PTMP_10_49_port, S(48) => PTMP_10_48_port, S(47) => 
                           PTMP_10_47_port, S(46) => PTMP_10_46_port, S(45) => 
                           PTMP_10_45_port, S(44) => PTMP_10_44_port, S(43) => 
                           PTMP_10_43_port, S(42) => PTMP_10_42_port, S(41) => 
                           PTMP_10_41_port, S(40) => PTMP_10_40_port, S(39) => 
                           PTMP_10_39_port, S(38) => PTMP_10_38_port, S(37) => 
                           PTMP_10_37_port, S(36) => PTMP_10_36_port, S(35) => 
                           PTMP_10_35_port, S(34) => PTMP_10_34_port, S(33) => 
                           PTMP_10_33_port, S(32) => PTMP_10_32_port, S(31) => 
                           PTMP_10_31_port, S(30) => PTMP_10_30_port, S(29) => 
                           PTMP_10_29_port, S(28) => PTMP_10_28_port, S(27) => 
                           PTMP_10_27_port, S(26) => PTMP_10_26_port, S(25) => 
                           PTMP_10_25_port, S(24) => PTMP_10_24_port, S(23) => 
                           PTMP_10_23_port, S(22) => PTMP_10_22_port, S(21) => 
                           PTMP_10_21_port, S(20) => PTMP_10_20_port, S(19) => 
                           PTMP_10_19_port, S(18) => PTMP_10_18_port, S(17) => 
                           PTMP_10_17_port, S(16) => PTMP_10_16_port, S(15) => 
                           PTMP_10_15_port, S(14) => PTMP_10_14_port, S(13) => 
                           PTMP_10_13_port, S(12) => PTMP_10_12_port, S(11) => 
                           PTMP_10_11_port, S(10) => PTMP_10_10_port, S(9) => 
                           PTMP_10_9_port, S(8) => PTMP_10_8_port, S(7) => 
                           PTMP_10_7_port, S(6) => PTMP_10_6_port, S(5) => 
                           PTMP_10_5_port, S(4) => PTMP_10_4_port, S(3) => 
                           PTMP_10_3_port, S(2) => PTMP_10_2_port, S(1) => 
                           PTMP_10_1_port, S(0) => PTMP_10_0_port, Co => n_1291
                           );
   ADDER_12 : RCA_NBIT58 port map( A(57) => PTMP_10_55_port, A(56) => 
                           PTMP_10_55_port, A(55) => PTMP_10_55_port, A(54) => 
                           PTMP_10_54_port, A(53) => PTMP_10_53_port, A(52) => 
                           PTMP_10_52_port, A(51) => PTMP_10_51_port, A(50) => 
                           PTMP_10_50_port, A(49) => PTMP_10_49_port, A(48) => 
                           PTMP_10_48_port, A(47) => PTMP_10_47_port, A(46) => 
                           PTMP_10_46_port, A(45) => PTMP_10_45_port, A(44) => 
                           PTMP_10_44_port, A(43) => PTMP_10_43_port, A(42) => 
                           PTMP_10_42_port, A(41) => PTMP_10_41_port, A(40) => 
                           PTMP_10_40_port, A(39) => PTMP_10_39_port, A(38) => 
                           PTMP_10_38_port, A(37) => PTMP_10_37_port, A(36) => 
                           PTMP_10_36_port, A(35) => PTMP_10_35_port, A(34) => 
                           PTMP_10_34_port, A(33) => PTMP_10_33_port, A(32) => 
                           PTMP_10_32_port, A(31) => PTMP_10_31_port, A(30) => 
                           PTMP_10_30_port, A(29) => PTMP_10_29_port, A(28) => 
                           PTMP_10_28_port, A(27) => PTMP_10_27_port, A(26) => 
                           PTMP_10_26_port, A(25) => PTMP_10_25_port, A(24) => 
                           PTMP_10_24_port, A(23) => PTMP_10_23_port, A(22) => 
                           PTMP_10_22_port, A(21) => PTMP_10_21_port, A(20) => 
                           PTMP_10_20_port, A(19) => PTMP_10_19_port, A(18) => 
                           PTMP_10_18_port, A(17) => PTMP_10_17_port, A(16) => 
                           PTMP_10_16_port, A(15) => PTMP_10_15_port, A(14) => 
                           PTMP_10_14_port, A(13) => PTMP_10_13_port, A(12) => 
                           PTMP_10_12_port, A(11) => PTMP_10_11_port, A(10) => 
                           PTMP_10_10_port, A(9) => PTMP_10_9_port, A(8) => 
                           PTMP_10_8_port, A(7) => PTMP_10_7_port, A(6) => 
                           PTMP_10_6_port, A(5) => PTMP_10_5_port, A(4) => 
                           PTMP_10_4_port, A(3) => PTMP_10_3_port, A(2) => 
                           PTMP_10_2_port, A(1) => PTMP_10_1_port, A(0) => 
                           PTMP_10_0_port, B(57) => OTMP_12_57_port, B(56) => 
                           OTMP_12_56_port, B(55) => OTMP_12_55_port, B(54) => 
                           OTMP_12_54_port, B(53) => OTMP_12_53_port, B(52) => 
                           OTMP_12_52_port, B(51) => OTMP_12_51_port, B(50) => 
                           OTMP_12_50_port, B(49) => OTMP_12_49_port, B(48) => 
                           OTMP_12_48_port, B(47) => OTMP_12_47_port, B(46) => 
                           OTMP_12_46_port, B(45) => OTMP_12_45_port, B(44) => 
                           OTMP_12_44_port, B(43) => OTMP_12_43_port, B(42) => 
                           OTMP_12_42_port, B(41) => OTMP_12_41_port, B(40) => 
                           OTMP_12_40_port, B(39) => OTMP_12_39_port, B(38) => 
                           OTMP_12_38_port, B(37) => OTMP_12_37_port, B(36) => 
                           OTMP_12_36_port, B(35) => OTMP_12_35_port, B(34) => 
                           OTMP_12_34_port, B(33) => OTMP_12_33_port, B(32) => 
                           OTMP_12_32_port, B(31) => OTMP_12_31_port, B(30) => 
                           OTMP_12_30_port, B(29) => OTMP_12_29_port, B(28) => 
                           OTMP_12_28_port, B(27) => OTMP_12_27_port, B(26) => 
                           OTMP_12_26_port, B(25) => OTMP_12_25_port, B(24) => 
                           OTMP_12_24_port, B(23) => OTMP_12_23_port, B(22) => 
                           OTMP_12_22_port, B(21) => OTMP_12_21_port, B(20) => 
                           OTMP_12_20_port, B(19) => OTMP_12_19_port, B(18) => 
                           OTMP_12_18_port, B(17) => OTMP_12_17_port, B(16) => 
                           OTMP_12_16_port, B(15) => OTMP_12_15_port, B(14) => 
                           OTMP_12_14_port, B(13) => OTMP_12_13_port, B(12) => 
                           OTMP_12_12_port, B(11) => OTMP_12_11_port, B(10) => 
                           OTMP_12_10_port, B(9) => OTMP_12_9_port, B(8) => 
                           OTMP_12_8_port, B(7) => OTMP_12_7_port, B(6) => 
                           OTMP_12_6_port, B(5) => OTMP_12_5_port, B(4) => 
                           OTMP_12_4_port, B(3) => OTMP_12_3_port, B(2) => 
                           OTMP_12_2_port, B(1) => OTMP_12_1_port, B(0) => 
                           OTMP_12_0_port, Ci => X_Logic0_port, S(57) => 
                           PTMP_11_57_port, S(56) => PTMP_11_56_port, S(55) => 
                           PTMP_11_55_port, S(54) => PTMP_11_54_port, S(53) => 
                           PTMP_11_53_port, S(52) => PTMP_11_52_port, S(51) => 
                           PTMP_11_51_port, S(50) => PTMP_11_50_port, S(49) => 
                           PTMP_11_49_port, S(48) => PTMP_11_48_port, S(47) => 
                           PTMP_11_47_port, S(46) => PTMP_11_46_port, S(45) => 
                           PTMP_11_45_port, S(44) => PTMP_11_44_port, S(43) => 
                           PTMP_11_43_port, S(42) => PTMP_11_42_port, S(41) => 
                           PTMP_11_41_port, S(40) => PTMP_11_40_port, S(39) => 
                           PTMP_11_39_port, S(38) => PTMP_11_38_port, S(37) => 
                           PTMP_11_37_port, S(36) => PTMP_11_36_port, S(35) => 
                           PTMP_11_35_port, S(34) => PTMP_11_34_port, S(33) => 
                           PTMP_11_33_port, S(32) => PTMP_11_32_port, S(31) => 
                           PTMP_11_31_port, S(30) => PTMP_11_30_port, S(29) => 
                           PTMP_11_29_port, S(28) => PTMP_11_28_port, S(27) => 
                           PTMP_11_27_port, S(26) => PTMP_11_26_port, S(25) => 
                           PTMP_11_25_port, S(24) => PTMP_11_24_port, S(23) => 
                           PTMP_11_23_port, S(22) => PTMP_11_22_port, S(21) => 
                           PTMP_11_21_port, S(20) => PTMP_11_20_port, S(19) => 
                           PTMP_11_19_port, S(18) => PTMP_11_18_port, S(17) => 
                           PTMP_11_17_port, S(16) => PTMP_11_16_port, S(15) => 
                           PTMP_11_15_port, S(14) => PTMP_11_14_port, S(13) => 
                           PTMP_11_13_port, S(12) => PTMP_11_12_port, S(11) => 
                           PTMP_11_11_port, S(10) => PTMP_11_10_port, S(9) => 
                           PTMP_11_9_port, S(8) => PTMP_11_8_port, S(7) => 
                           PTMP_11_7_port, S(6) => PTMP_11_6_port, S(5) => 
                           PTMP_11_5_port, S(4) => PTMP_11_4_port, S(3) => 
                           PTMP_11_3_port, S(2) => PTMP_11_2_port, S(1) => 
                           PTMP_11_1_port, S(0) => PTMP_11_0_port, Co => n_1292
                           );
   ADDER_13 : RCA_NBIT60 port map( A(59) => PTMP_11_57_port, A(58) => 
                           PTMP_11_57_port, A(57) => PTMP_11_57_port, A(56) => 
                           PTMP_11_56_port, A(55) => PTMP_11_55_port, A(54) => 
                           PTMP_11_54_port, A(53) => PTMP_11_53_port, A(52) => 
                           PTMP_11_52_port, A(51) => PTMP_11_51_port, A(50) => 
                           PTMP_11_50_port, A(49) => PTMP_11_49_port, A(48) => 
                           PTMP_11_48_port, A(47) => PTMP_11_47_port, A(46) => 
                           PTMP_11_46_port, A(45) => PTMP_11_45_port, A(44) => 
                           PTMP_11_44_port, A(43) => PTMP_11_43_port, A(42) => 
                           PTMP_11_42_port, A(41) => PTMP_11_41_port, A(40) => 
                           PTMP_11_40_port, A(39) => PTMP_11_39_port, A(38) => 
                           PTMP_11_38_port, A(37) => PTMP_11_37_port, A(36) => 
                           PTMP_11_36_port, A(35) => PTMP_11_35_port, A(34) => 
                           PTMP_11_34_port, A(33) => PTMP_11_33_port, A(32) => 
                           PTMP_11_32_port, A(31) => PTMP_11_31_port, A(30) => 
                           PTMP_11_30_port, A(29) => PTMP_11_29_port, A(28) => 
                           PTMP_11_28_port, A(27) => PTMP_11_27_port, A(26) => 
                           PTMP_11_26_port, A(25) => PTMP_11_25_port, A(24) => 
                           PTMP_11_24_port, A(23) => PTMP_11_23_port, A(22) => 
                           PTMP_11_22_port, A(21) => PTMP_11_21_port, A(20) => 
                           PTMP_11_20_port, A(19) => PTMP_11_19_port, A(18) => 
                           PTMP_11_18_port, A(17) => PTMP_11_17_port, A(16) => 
                           PTMP_11_16_port, A(15) => PTMP_11_15_port, A(14) => 
                           PTMP_11_14_port, A(13) => PTMP_11_13_port, A(12) => 
                           PTMP_11_12_port, A(11) => PTMP_11_11_port, A(10) => 
                           PTMP_11_10_port, A(9) => PTMP_11_9_port, A(8) => 
                           PTMP_11_8_port, A(7) => PTMP_11_7_port, A(6) => 
                           PTMP_11_6_port, A(5) => PTMP_11_5_port, A(4) => 
                           PTMP_11_4_port, A(3) => PTMP_11_3_port, A(2) => 
                           PTMP_11_2_port, A(1) => PTMP_11_1_port, A(0) => 
                           PTMP_11_0_port, B(59) => OTMP_13_59_port, B(58) => 
                           OTMP_13_58_port, B(57) => OTMP_13_57_port, B(56) => 
                           OTMP_13_56_port, B(55) => OTMP_13_55_port, B(54) => 
                           OTMP_13_54_port, B(53) => OTMP_13_53_port, B(52) => 
                           OTMP_13_52_port, B(51) => OTMP_13_51_port, B(50) => 
                           OTMP_13_50_port, B(49) => OTMP_13_49_port, B(48) => 
                           OTMP_13_48_port, B(47) => OTMP_13_47_port, B(46) => 
                           OTMP_13_46_port, B(45) => OTMP_13_45_port, B(44) => 
                           OTMP_13_44_port, B(43) => OTMP_13_43_port, B(42) => 
                           OTMP_13_42_port, B(41) => OTMP_13_41_port, B(40) => 
                           OTMP_13_40_port, B(39) => OTMP_13_39_port, B(38) => 
                           OTMP_13_38_port, B(37) => OTMP_13_37_port, B(36) => 
                           OTMP_13_36_port, B(35) => OTMP_13_35_port, B(34) => 
                           OTMP_13_34_port, B(33) => OTMP_13_33_port, B(32) => 
                           OTMP_13_32_port, B(31) => OTMP_13_31_port, B(30) => 
                           OTMP_13_30_port, B(29) => OTMP_13_29_port, B(28) => 
                           OTMP_13_28_port, B(27) => OTMP_13_27_port, B(26) => 
                           OTMP_13_26_port, B(25) => OTMP_13_25_port, B(24) => 
                           OTMP_13_24_port, B(23) => OTMP_13_23_port, B(22) => 
                           OTMP_13_22_port, B(21) => OTMP_13_21_port, B(20) => 
                           OTMP_13_20_port, B(19) => OTMP_13_19_port, B(18) => 
                           OTMP_13_18_port, B(17) => OTMP_13_17_port, B(16) => 
                           OTMP_13_16_port, B(15) => OTMP_13_15_port, B(14) => 
                           OTMP_13_14_port, B(13) => OTMP_13_13_port, B(12) => 
                           OTMP_13_12_port, B(11) => OTMP_13_11_port, B(10) => 
                           OTMP_13_10_port, B(9) => OTMP_13_9_port, B(8) => 
                           OTMP_13_8_port, B(7) => OTMP_13_7_port, B(6) => 
                           OTMP_13_6_port, B(5) => OTMP_13_5_port, B(4) => 
                           OTMP_13_4_port, B(3) => OTMP_13_3_port, B(2) => 
                           OTMP_13_2_port, B(1) => OTMP_13_1_port, B(0) => 
                           OTMP_13_0_port, Ci => X_Logic0_port, S(59) => 
                           PTMP_12_59_port, S(58) => PTMP_12_58_port, S(57) => 
                           PTMP_12_57_port, S(56) => PTMP_12_56_port, S(55) => 
                           PTMP_12_55_port, S(54) => PTMP_12_54_port, S(53) => 
                           PTMP_12_53_port, S(52) => PTMP_12_52_port, S(51) => 
                           PTMP_12_51_port, S(50) => PTMP_12_50_port, S(49) => 
                           PTMP_12_49_port, S(48) => PTMP_12_48_port, S(47) => 
                           PTMP_12_47_port, S(46) => PTMP_12_46_port, S(45) => 
                           PTMP_12_45_port, S(44) => PTMP_12_44_port, S(43) => 
                           PTMP_12_43_port, S(42) => PTMP_12_42_port, S(41) => 
                           PTMP_12_41_port, S(40) => PTMP_12_40_port, S(39) => 
                           PTMP_12_39_port, S(38) => PTMP_12_38_port, S(37) => 
                           PTMP_12_37_port, S(36) => PTMP_12_36_port, S(35) => 
                           PTMP_12_35_port, S(34) => PTMP_12_34_port, S(33) => 
                           PTMP_12_33_port, S(32) => PTMP_12_32_port, S(31) => 
                           PTMP_12_31_port, S(30) => PTMP_12_30_port, S(29) => 
                           PTMP_12_29_port, S(28) => PTMP_12_28_port, S(27) => 
                           PTMP_12_27_port, S(26) => PTMP_12_26_port, S(25) => 
                           PTMP_12_25_port, S(24) => PTMP_12_24_port, S(23) => 
                           PTMP_12_23_port, S(22) => PTMP_12_22_port, S(21) => 
                           PTMP_12_21_port, S(20) => PTMP_12_20_port, S(19) => 
                           PTMP_12_19_port, S(18) => PTMP_12_18_port, S(17) => 
                           PTMP_12_17_port, S(16) => PTMP_12_16_port, S(15) => 
                           PTMP_12_15_port, S(14) => PTMP_12_14_port, S(13) => 
                           PTMP_12_13_port, S(12) => PTMP_12_12_port, S(11) => 
                           PTMP_12_11_port, S(10) => PTMP_12_10_port, S(9) => 
                           PTMP_12_9_port, S(8) => PTMP_12_8_port, S(7) => 
                           PTMP_12_7_port, S(6) => PTMP_12_6_port, S(5) => 
                           PTMP_12_5_port, S(4) => PTMP_12_4_port, S(3) => 
                           PTMP_12_3_port, S(2) => PTMP_12_2_port, S(1) => 
                           PTMP_12_1_port, S(0) => PTMP_12_0_port, Co => n_1293
                           );
   ADDER_14 : RCA_NBIT62 port map( A(61) => PTMP_12_59_port, A(60) => 
                           PTMP_12_59_port, A(59) => PTMP_12_59_port, A(58) => 
                           PTMP_12_58_port, A(57) => PTMP_12_57_port, A(56) => 
                           PTMP_12_56_port, A(55) => PTMP_12_55_port, A(54) => 
                           PTMP_12_54_port, A(53) => PTMP_12_53_port, A(52) => 
                           PTMP_12_52_port, A(51) => PTMP_12_51_port, A(50) => 
                           PTMP_12_50_port, A(49) => PTMP_12_49_port, A(48) => 
                           PTMP_12_48_port, A(47) => PTMP_12_47_port, A(46) => 
                           PTMP_12_46_port, A(45) => PTMP_12_45_port, A(44) => 
                           PTMP_12_44_port, A(43) => PTMP_12_43_port, A(42) => 
                           PTMP_12_42_port, A(41) => PTMP_12_41_port, A(40) => 
                           PTMP_12_40_port, A(39) => PTMP_12_39_port, A(38) => 
                           PTMP_12_38_port, A(37) => PTMP_12_37_port, A(36) => 
                           PTMP_12_36_port, A(35) => PTMP_12_35_port, A(34) => 
                           PTMP_12_34_port, A(33) => PTMP_12_33_port, A(32) => 
                           PTMP_12_32_port, A(31) => PTMP_12_31_port, A(30) => 
                           PTMP_12_30_port, A(29) => PTMP_12_29_port, A(28) => 
                           PTMP_12_28_port, A(27) => PTMP_12_27_port, A(26) => 
                           PTMP_12_26_port, A(25) => PTMP_12_25_port, A(24) => 
                           PTMP_12_24_port, A(23) => PTMP_12_23_port, A(22) => 
                           PTMP_12_22_port, A(21) => PTMP_12_21_port, A(20) => 
                           PTMP_12_20_port, A(19) => PTMP_12_19_port, A(18) => 
                           PTMP_12_18_port, A(17) => PTMP_12_17_port, A(16) => 
                           PTMP_12_16_port, A(15) => PTMP_12_15_port, A(14) => 
                           PTMP_12_14_port, A(13) => PTMP_12_13_port, A(12) => 
                           PTMP_12_12_port, A(11) => PTMP_12_11_port, A(10) => 
                           PTMP_12_10_port, A(9) => PTMP_12_9_port, A(8) => 
                           PTMP_12_8_port, A(7) => PTMP_12_7_port, A(6) => 
                           PTMP_12_6_port, A(5) => PTMP_12_5_port, A(4) => 
                           PTMP_12_4_port, A(3) => PTMP_12_3_port, A(2) => 
                           PTMP_12_2_port, A(1) => PTMP_12_1_port, A(0) => 
                           PTMP_12_0_port, B(61) => OTMP_14_61_port, B(60) => 
                           OTMP_14_60_port, B(59) => OTMP_14_59_port, B(58) => 
                           OTMP_14_58_port, B(57) => OTMP_14_57_port, B(56) => 
                           OTMP_14_56_port, B(55) => OTMP_14_55_port, B(54) => 
                           OTMP_14_54_port, B(53) => OTMP_14_53_port, B(52) => 
                           OTMP_14_52_port, B(51) => OTMP_14_51_port, B(50) => 
                           OTMP_14_50_port, B(49) => OTMP_14_49_port, B(48) => 
                           OTMP_14_48_port, B(47) => OTMP_14_47_port, B(46) => 
                           OTMP_14_46_port, B(45) => OTMP_14_45_port, B(44) => 
                           OTMP_14_44_port, B(43) => OTMP_14_43_port, B(42) => 
                           OTMP_14_42_port, B(41) => OTMP_14_41_port, B(40) => 
                           OTMP_14_40_port, B(39) => OTMP_14_39_port, B(38) => 
                           OTMP_14_38_port, B(37) => OTMP_14_37_port, B(36) => 
                           OTMP_14_36_port, B(35) => OTMP_14_35_port, B(34) => 
                           OTMP_14_34_port, B(33) => OTMP_14_33_port, B(32) => 
                           OTMP_14_32_port, B(31) => OTMP_14_31_port, B(30) => 
                           OTMP_14_30_port, B(29) => OTMP_14_29_port, B(28) => 
                           OTMP_14_28_port, B(27) => OTMP_14_27_port, B(26) => 
                           OTMP_14_26_port, B(25) => OTMP_14_25_port, B(24) => 
                           OTMP_14_24_port, B(23) => OTMP_14_23_port, B(22) => 
                           OTMP_14_22_port, B(21) => OTMP_14_21_port, B(20) => 
                           OTMP_14_20_port, B(19) => OTMP_14_19_port, B(18) => 
                           OTMP_14_18_port, B(17) => OTMP_14_17_port, B(16) => 
                           OTMP_14_16_port, B(15) => OTMP_14_15_port, B(14) => 
                           OTMP_14_14_port, B(13) => OTMP_14_13_port, B(12) => 
                           OTMP_14_12_port, B(11) => OTMP_14_11_port, B(10) => 
                           OTMP_14_10_port, B(9) => OTMP_14_9_port, B(8) => 
                           OTMP_14_8_port, B(7) => OTMP_14_7_port, B(6) => 
                           OTMP_14_6_port, B(5) => OTMP_14_5_port, B(4) => 
                           OTMP_14_4_port, B(3) => OTMP_14_3_port, B(2) => 
                           OTMP_14_2_port, B(1) => OTMP_14_1_port, B(0) => 
                           OTMP_14_0_port, Ci => X_Logic0_port, S(61) => 
                           PTMP_13_61_port, S(60) => PTMP_13_60_port, S(59) => 
                           PTMP_13_59_port, S(58) => PTMP_13_58_port, S(57) => 
                           PTMP_13_57_port, S(56) => PTMP_13_56_port, S(55) => 
                           PTMP_13_55_port, S(54) => PTMP_13_54_port, S(53) => 
                           PTMP_13_53_port, S(52) => PTMP_13_52_port, S(51) => 
                           PTMP_13_51_port, S(50) => PTMP_13_50_port, S(49) => 
                           PTMP_13_49_port, S(48) => PTMP_13_48_port, S(47) => 
                           PTMP_13_47_port, S(46) => PTMP_13_46_port, S(45) => 
                           PTMP_13_45_port, S(44) => PTMP_13_44_port, S(43) => 
                           PTMP_13_43_port, S(42) => PTMP_13_42_port, S(41) => 
                           PTMP_13_41_port, S(40) => PTMP_13_40_port, S(39) => 
                           PTMP_13_39_port, S(38) => PTMP_13_38_port, S(37) => 
                           PTMP_13_37_port, S(36) => PTMP_13_36_port, S(35) => 
                           PTMP_13_35_port, S(34) => PTMP_13_34_port, S(33) => 
                           PTMP_13_33_port, S(32) => PTMP_13_32_port, S(31) => 
                           PTMP_13_31_port, S(30) => PTMP_13_30_port, S(29) => 
                           PTMP_13_29_port, S(28) => PTMP_13_28_port, S(27) => 
                           PTMP_13_27_port, S(26) => PTMP_13_26_port, S(25) => 
                           PTMP_13_25_port, S(24) => PTMP_13_24_port, S(23) => 
                           PTMP_13_23_port, S(22) => PTMP_13_22_port, S(21) => 
                           PTMP_13_21_port, S(20) => PTMP_13_20_port, S(19) => 
                           PTMP_13_19_port, S(18) => PTMP_13_18_port, S(17) => 
                           PTMP_13_17_port, S(16) => PTMP_13_16_port, S(15) => 
                           PTMP_13_15_port, S(14) => PTMP_13_14_port, S(13) => 
                           PTMP_13_13_port, S(12) => PTMP_13_12_port, S(11) => 
                           PTMP_13_11_port, S(10) => PTMP_13_10_port, S(9) => 
                           PTMP_13_9_port, S(8) => PTMP_13_8_port, S(7) => 
                           PTMP_13_7_port, S(6) => PTMP_13_6_port, S(5) => 
                           PTMP_13_5_port, S(4) => PTMP_13_4_port, S(3) => 
                           PTMP_13_3_port, S(2) => PTMP_13_2_port, S(1) => 
                           PTMP_13_1_port, S(0) => PTMP_13_0_port, Co => n_1294
                           );
   ADDER_15 : RCA_NBIT64 port map( A(63) => PTMP_13_61_port, A(62) => 
                           PTMP_13_61_port, A(61) => PTMP_13_61_port, A(60) => 
                           PTMP_13_60_port, A(59) => PTMP_13_59_port, A(58) => 
                           PTMP_13_58_port, A(57) => PTMP_13_57_port, A(56) => 
                           PTMP_13_56_port, A(55) => PTMP_13_55_port, A(54) => 
                           PTMP_13_54_port, A(53) => PTMP_13_53_port, A(52) => 
                           PTMP_13_52_port, A(51) => PTMP_13_51_port, A(50) => 
                           PTMP_13_50_port, A(49) => PTMP_13_49_port, A(48) => 
                           PTMP_13_48_port, A(47) => PTMP_13_47_port, A(46) => 
                           PTMP_13_46_port, A(45) => PTMP_13_45_port, A(44) => 
                           PTMP_13_44_port, A(43) => PTMP_13_43_port, A(42) => 
                           PTMP_13_42_port, A(41) => PTMP_13_41_port, A(40) => 
                           PTMP_13_40_port, A(39) => PTMP_13_39_port, A(38) => 
                           PTMP_13_38_port, A(37) => PTMP_13_37_port, A(36) => 
                           PTMP_13_36_port, A(35) => PTMP_13_35_port, A(34) => 
                           PTMP_13_34_port, A(33) => PTMP_13_33_port, A(32) => 
                           PTMP_13_32_port, A(31) => PTMP_13_31_port, A(30) => 
                           PTMP_13_30_port, A(29) => PTMP_13_29_port, A(28) => 
                           PTMP_13_28_port, A(27) => PTMP_13_27_port, A(26) => 
                           PTMP_13_26_port, A(25) => PTMP_13_25_port, A(24) => 
                           PTMP_13_24_port, A(23) => PTMP_13_23_port, A(22) => 
                           PTMP_13_22_port, A(21) => PTMP_13_21_port, A(20) => 
                           PTMP_13_20_port, A(19) => PTMP_13_19_port, A(18) => 
                           PTMP_13_18_port, A(17) => PTMP_13_17_port, A(16) => 
                           PTMP_13_16_port, A(15) => PTMP_13_15_port, A(14) => 
                           PTMP_13_14_port, A(13) => PTMP_13_13_port, A(12) => 
                           PTMP_13_12_port, A(11) => PTMP_13_11_port, A(10) => 
                           PTMP_13_10_port, A(9) => PTMP_13_9_port, A(8) => 
                           PTMP_13_8_port, A(7) => PTMP_13_7_port, A(6) => 
                           PTMP_13_6_port, A(5) => PTMP_13_5_port, A(4) => 
                           PTMP_13_4_port, A(3) => PTMP_13_3_port, A(2) => 
                           PTMP_13_2_port, A(1) => PTMP_13_1_port, A(0) => 
                           PTMP_13_0_port, B(63) => OTMP_15_63_port, B(62) => 
                           OTMP_15_62_port, B(61) => OTMP_15_61_port, B(60) => 
                           OTMP_15_60_port, B(59) => OTMP_15_59_port, B(58) => 
                           OTMP_15_58_port, B(57) => OTMP_15_57_port, B(56) => 
                           OTMP_15_56_port, B(55) => OTMP_15_55_port, B(54) => 
                           OTMP_15_54_port, B(53) => OTMP_15_53_port, B(52) => 
                           OTMP_15_52_port, B(51) => OTMP_15_51_port, B(50) => 
                           OTMP_15_50_port, B(49) => OTMP_15_49_port, B(48) => 
                           OTMP_15_48_port, B(47) => OTMP_15_47_port, B(46) => 
                           OTMP_15_46_port, B(45) => OTMP_15_45_port, B(44) => 
                           OTMP_15_44_port, B(43) => OTMP_15_43_port, B(42) => 
                           OTMP_15_42_port, B(41) => OTMP_15_41_port, B(40) => 
                           OTMP_15_40_port, B(39) => OTMP_15_39_port, B(38) => 
                           OTMP_15_38_port, B(37) => OTMP_15_37_port, B(36) => 
                           OTMP_15_36_port, B(35) => OTMP_15_35_port, B(34) => 
                           OTMP_15_34_port, B(33) => OTMP_15_33_port, B(32) => 
                           OTMP_15_32_port, B(31) => OTMP_15_31_port, B(30) => 
                           OTMP_15_30_port, B(29) => OTMP_15_29_port, B(28) => 
                           OTMP_15_28_port, B(27) => OTMP_15_27_port, B(26) => 
                           OTMP_15_26_port, B(25) => OTMP_15_25_port, B(24) => 
                           OTMP_15_24_port, B(23) => OTMP_15_23_port, B(22) => 
                           OTMP_15_22_port, B(21) => OTMP_15_21_port, B(20) => 
                           OTMP_15_20_port, B(19) => OTMP_15_19_port, B(18) => 
                           OTMP_15_18_port, B(17) => OTMP_15_17_port, B(16) => 
                           OTMP_15_16_port, B(15) => OTMP_15_15_port, B(14) => 
                           OTMP_15_14_port, B(13) => OTMP_15_13_port, B(12) => 
                           OTMP_15_12_port, B(11) => OTMP_15_11_port, B(10) => 
                           OTMP_15_10_port, B(9) => OTMP_15_9_port, B(8) => 
                           OTMP_15_8_port, B(7) => OTMP_15_7_port, B(6) => 
                           OTMP_15_6_port, B(5) => OTMP_15_5_port, B(4) => 
                           OTMP_15_4_port, B(3) => OTMP_15_3_port, B(2) => 
                           OTMP_15_2_port, B(1) => OTMP_15_1_port, B(0) => 
                           OTMP_15_0_port, Ci => X_Logic0_port, S(63) => S(63),
                           S(62) => S(62), S(61) => S(61), S(60) => S(60), 
                           S(59) => S(59), S(58) => S(58), S(57) => S(57), 
                           S(56) => S(56), S(55) => S(55), S(54) => S(54), 
                           S(53) => S(53), S(52) => S(52), S(51) => S(51), 
                           S(50) => S(50), S(49) => S(49), S(48) => S(48), 
                           S(47) => S(47), S(46) => S(46), S(45) => S(45), 
                           S(44) => S(44), S(43) => S(43), S(42) => S(42), 
                           S(41) => S(41), S(40) => S(40), S(39) => S(39), 
                           S(38) => S(38), S(37) => S(37), S(36) => S(36), 
                           S(35) => S(35), S(34) => S(34), S(33) => S(33), 
                           S(32) => S(32), S(31) => S(31), S(30) => S(30), 
                           S(29) => S(29), S(28) => S(28), S(27) => S(27), 
                           S(26) => S(26), S(25) => S(25), S(24) => S(24), 
                           S(23) => S(23), S(22) => S(22), S(21) => S(21), 
                           S(20) => S(20), S(19) => S(19), S(18) => S(18), 
                           S(17) => S(17), S(16) => S(16), S(15) => S(15), 
                           S(14) => S(14), S(13) => S(13), S(12) => S(12), 
                           S(11) => S(11), S(10) => S(10), S(9) => S(9), S(8) 
                           => S(8), S(7) => S(7), S(6) => S(6), S(5) => S(5), 
                           S(4) => S(4), S(3) => S(3), S(2) => S(2), S(1) => 
                           S(1), S(0) => S(0), Co => n_1295);
   sub_101 : BOOTHMUL_NBIT32_DW01_sub_0 port map( A(31) => n1, A(30) => n1, 
                           A(29) => n1, A(28) => n1, A(27) => n1, A(26) => n1, 
                           A(25) => n1, A(24) => n1, A(23) => n1, A(22) => n1, 
                           A(21) => n1, A(20) => n1, A(19) => n1, A(18) => n1, 
                           A(17) => n1, A(16) => n1, A(15) => n1, A(14) => n1, 
                           A(13) => n1, A(12) => n1, A(11) => n1, A(10) => n1, 
                           A(9) => n1, A(8) => n1, A(7) => n1, A(6) => n1, A(5)
                           => n1, A(4) => n1, A(3) => n1, A(2) => n1, A(1) => 
                           n1, A(0) => n1, B(31) => A(31), B(30) => A(30), 
                           B(29) => A(29), B(28) => A(28), B(27) => A(27), 
                           B(26) => A(26), B(25) => A(25), B(24) => A(24), 
                           B(23) => A(23), B(22) => A(22), B(21) => A(21), 
                           B(20) => A(20), B(19) => A(19), B(18) => A(18), 
                           B(17) => A(17), B(16) => A(16), B(15) => A(15), 
                           B(14) => A(14), B(13) => A(13), B(12) => A(12), 
                           B(11) => A(11), B(10) => A(10), B(9) => A(9), B(8) 
                           => A(8), B(7) => A(7), B(6) => A(6), B(5) => A(5), 
                           B(4) => A(4), B(3) => A(3), B(2) => A(2), B(1) => 
                           A(1), B(0) => A(0), CI => n2, DIFF(31) => A_n_65, 
                           DIFF(30) => A_n_30_port, DIFF(29) => A_n_29_port, 
                           DIFF(28) => A_n_28_port, DIFF(27) => A_n_27_port, 
                           DIFF(26) => A_n_26_port, DIFF(25) => A_n_25_port, 
                           DIFF(24) => A_n_24_port, DIFF(23) => A_n_23_port, 
                           DIFF(22) => A_n_22_port, DIFF(21) => A_n_21_port, 
                           DIFF(20) => A_n_20_port, DIFF(19) => A_n_19_port, 
                           DIFF(18) => A_n_18_port, DIFF(17) => A_n_17_port, 
                           DIFF(16) => A_n_16_port, DIFF(15) => A_n_15_port, 
                           DIFF(14) => A_n_14_port, DIFF(13) => A_n_13_port, 
                           DIFF(12) => A_n_12_port, DIFF(11) => A_n_11_port, 
                           DIFF(10) => A_n_10_port, DIFF(9) => A_n_9_port, 
                           DIFF(8) => A_n_8_port, DIFF(7) => A_n_7_port, 
                           DIFF(6) => A_n_6_port, DIFF(5) => A_n_5_port, 
                           DIFF(4) => A_n_4_port, DIFF(3) => A_n_3_port, 
                           DIFF(2) => A_n_2_port, DIFF(1) => A_n_1_port, 
                           DIFF(0) => A_n_0_port, CO => n_1296);
   OTMP_15_0_port <= '0';
   SHIFT_n_15_0_port <= '0';
   SHIFT_n_15_1_port <= '0';
   SHIFT_15_0_port <= '0';
   SHIFT_15_1_port <= '0';
   OTMP_14_0_port <= '0';
   SHIFT_n_14_0_port <= '0';
   SHIFT_n_14_1_port <= '0';
   SHIFT_14_0_port <= '0';
   SHIFT_14_1_port <= '0';
   OTMP_13_0_port <= '0';
   SHIFT_n_13_0_port <= '0';
   SHIFT_n_13_1_port <= '0';
   SHIFT_13_0_port <= '0';
   SHIFT_13_1_port <= '0';
   OTMP_12_0_port <= '0';
   SHIFT_n_12_0_port <= '0';
   SHIFT_n_12_1_port <= '0';
   SHIFT_12_0_port <= '0';
   SHIFT_12_1_port <= '0';
   OTMP_11_0_port <= '0';
   SHIFT_n_11_0_port <= '0';
   SHIFT_n_11_1_port <= '0';
   SHIFT_11_0_port <= '0';
   SHIFT_11_1_port <= '0';
   OTMP_10_0_port <= '0';
   SHIFT_n_10_0_port <= '0';
   SHIFT_n_10_1_port <= '0';
   SHIFT_10_0_port <= '0';
   SHIFT_10_1_port <= '0';
   OTMP_9_0_port <= '0';
   SHIFT_n_9_0_port <= '0';
   SHIFT_n_9_1_port <= '0';
   SHIFT_9_0_port <= '0';
   SHIFT_9_1_port <= '0';
   OTMP_8_0_port <= '0';
   SHIFT_n_8_0_port <= '0';
   SHIFT_n_8_1_port <= '0';
   SHIFT_8_0_port <= '0';
   SHIFT_8_1_port <= '0';
   OTMP_7_0_port <= '0';
   SHIFT_n_7_0_port <= '0';
   SHIFT_n_7_1_port <= '0';
   SHIFT_7_0_port <= '0';
   SHIFT_7_1_port <= '0';
   OTMP_6_0_port <= '0';
   SHIFT_n_6_0_port <= '0';
   SHIFT_n_6_1_port <= '0';
   SHIFT_6_0_port <= '0';
   SHIFT_6_1_port <= '0';
   OTMP_5_0_port <= '0';
   SHIFT_n_5_0_port <= '0';
   SHIFT_n_5_1_port <= '0';
   SHIFT_5_0_port <= '0';
   SHIFT_5_1_port <= '0';
   OTMP_4_0_port <= '0';
   SHIFT_n_4_0_port <= '0';
   SHIFT_n_4_1_port <= '0';
   SHIFT_4_0_port <= '0';
   SHIFT_4_1_port <= '0';
   OTMP_3_0_port <= '0';
   SHIFT_n_3_0_port <= '0';
   SHIFT_n_3_1_port <= '0';
   SHIFT_3_0_port <= '0';
   SHIFT_3_1_port <= '0';
   OTMP_2_0_port <= '0';
   SHIFT_n_2_0_port <= '0';
   SHIFT_n_2_1_port <= '0';
   SHIFT_2_0_port <= '0';
   SHIFT_2_1_port <= '0';
   OTMP_1_0_port <= '0';
   SHIFT_n_1_0_port <= '0';
   SHIFT_1_0_port <= '0';

end SYN_BEHAVIOURAL;
