PACKAGE CONSTANTS IS
   CONSTANT NumBit : INTEGER := 64;
END CONSTANTS;