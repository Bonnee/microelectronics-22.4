LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL; --  libreria IEEE con definizione tipi standard logic
USE WORK.constants.ALL; -- libreria WORK user-defined

ENTITY IV IS
	PORT (
		A : IN STD_LOGIC;
		Y : OUT STD_LOGIC);
END IV;
ARCHITECTURE BEHAVIORAL OF IV IS

BEGIN
	Y <= NOT(A);

END BEHAVIORAL;

CONFIGURATION CFG_IV_BEHAVIORAL OF IV IS
	FOR BEHAVIORAL
	END FOR;
END CFG_IV_BEHAVIORAL;
