PACKAGE CONSTANTS IS
   CONSTANT NumBit : INTEGER := 6;
   CONSTANT TP_MUX : TIME := 0.5 ns;
END CONSTANTS;