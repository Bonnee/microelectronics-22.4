/home/ms22.4/cap1/vhdlsim/constants.vhd