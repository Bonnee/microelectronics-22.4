PACKAGE CONSTANTS IS
   CONSTANT NumBit : INTEGER := 6;
END CONSTANTS;