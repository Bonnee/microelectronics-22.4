
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_RF_ADDR_W5_DATA_W32 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_RF_ADDR_W5_DATA_W32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_RF_ADDR_W5_DATA_W32.all;

entity RF_ADDR_W5_DATA_W32 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end RF_ADDR_W5_DATA_W32;

architecture SYN_Behavioural of RF_ADDR_W5_DATA_W32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X4
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal OUT1_31_port, OUT1_30_port, OUT1_29_port, OUT1_28_port, OUT1_27_port,
      OUT1_26_port, OUT1_25_port, OUT1_24_port, OUT1_23_port, OUT1_22_port, 
      OUT1_21_port, OUT1_20_port, OUT1_19_port, OUT1_18_port, OUT1_17_port, 
      OUT1_16_port, OUT1_15_port, OUT1_14_port, OUT1_13_port, OUT1_12_port, 
      OUT1_11_port, OUT1_10_port, OUT1_9_port, OUT1_8_port, OUT1_7_port, 
      OUT1_6_port, OUT1_5_port, OUT1_4_port, OUT1_3_port, OUT1_2_port, 
      OUT1_1_port, OUT1_0_port, OUT2_31_port, OUT2_30_port, OUT2_29_port, 
      OUT2_28_port, OUT2_27_port, OUT2_26_port, OUT2_25_port, OUT2_24_port, 
      OUT2_23_port, OUT2_22_port, OUT2_21_port, OUT2_20_port, OUT2_19_port, 
      OUT2_18_port, OUT2_17_port, OUT2_16_port, OUT2_15_port, OUT2_14_port, 
      OUT2_13_port, OUT2_12_port, OUT2_11_port, OUT2_10_port, OUT2_9_port, 
      OUT2_8_port, OUT2_7_port, OUT2_6_port, OUT2_5_port, OUT2_4_port, 
      OUT2_3_port, OUT2_2_port, OUT2_1_port, OUT2_0_port, n1, n2, n3, n4, n5, 
      n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, 
      n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35
      , n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, 
      n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64
      , n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
      n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, 
      n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, 
      n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, 
      n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, 
      n189, n190, n191, n192, n257, n258, n259, n260, n261, n262, n263, n264, 
      n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, 
      n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, 
      n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, 
      n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, 
      n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, 
      n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, 
      n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, 
      n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, 
      n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, 
      n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, 
      n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, 
      n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, 
      n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, 
      n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, 
      n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, 
      n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, 
      n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, 
      n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, 
      n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, 
      n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, 
      n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, 
      n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, 
      n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, 
      n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, 
      n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, 
      n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, 
      n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, 
      n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, 
      n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, 
      n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, 
      n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, 
      n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, 
      n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, 
      n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, 
      n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, 
      n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, 
      n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, 
      n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, 
      n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, 
      n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, 
      n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, 
      n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, 
      n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, 
      n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, 
      n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, 
      n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, 
      n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, 
      n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, 
      n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, 
      n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, 
      n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, 
      n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, 
      n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, 
      n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, 
      n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, 
      n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, 
      n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, 
      n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, 
      n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, 
      n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, 
      n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, 
      n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, 
      n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, 
      n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, 
      n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, 
      n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, 
      n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, 
      n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, 
      n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, 
      n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, 
      n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, 
      n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, 
      n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, 
      n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, 
      n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, 
      n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, 
      n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, 
      n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, 
      n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, 
      n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, 
      n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, 
      n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, 
      n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, 
      n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, 
      n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, 
      n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, 
      n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, 
      n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, 
      n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, 
      n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, 
      n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, 
      n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, 
      n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, 
      n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, 
      n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, 
      n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, 
      n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, 
      n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, 
      n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, 
      n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, 
      n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, 
      n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, 
      n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, 
      n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, 
      n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, 
      n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, 
      n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, 
      n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, 
      n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, 
      n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, 
      n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, 
      n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, 
      n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, 
      n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, 
      n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, 
      n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, 
      n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, 
      n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, 
      n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, 
      n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, 
      n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, 
      n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, 
      n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, 
      n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, 
      n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, 
      n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, 
      n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, 
      n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, 
      n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, 
      n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, 
      n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, 
      n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, 
      n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, 
      n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, 
      n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, 
      n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, 
      n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, 
      n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, 
      n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, 
      n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, 
      n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, 
      n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, 
      n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, 
      n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, 
      n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, 
      n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, 
      n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, 
      n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, 
      n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, 
      n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, 
      n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, 
      n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, 
      n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, 
      n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, 
      n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, 
      n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, 
      n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, 
      n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, 
      n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, 
      n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, 
      n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, 
      n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, 
      n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, 
      n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, 
      n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, 
      n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, 
      n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, 
      n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, 
      n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, 
      n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, 
      n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, 
      n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, 
      n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, 
      n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, 
      n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, 
      n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, 
      n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, 
      n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, 
      n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, 
      n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, 
      n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, 
      n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, 
      n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, 
      n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, 
      n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, 
      n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, 
      n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, 
      n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, 
      n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, 
      n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, 
      n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, 
      n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, 
      n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, 
      n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, 
      n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, 
      n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, 
      n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, 
      n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, 
      n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, 
      n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, 
      n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, 
      n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, 
      n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, 
      n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, 
      n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, 
      n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, 
      n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, 
      n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, 
      n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, 
      n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, 
      n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, 
      n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, 
      n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, 
      n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, 
      n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, 
      n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, 
      n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, 
      n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, 
      n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, 
      n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, 
      n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, 
      n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, 
      n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, 
      n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, 
      n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, 
      n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, 
      n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, 
      n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, 
      n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, 
      n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, 
      n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, 
      n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, 
      n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, 
      n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, 
      n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, 
      n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, 
      n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, 
      n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, 
      n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, 
      n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, 
      n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, 
      n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, 
      n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, 
      n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, 
      n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, 
      n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, 
      n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, 
      n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, 
      n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, 
      n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, 
      n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, 
      n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, 
      n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, 
      n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, 
      n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, 
      n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, 
      n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, 
      n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, 
      n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, 
      n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, 
      n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, 
      n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, 
      n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, 
      n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, 
      n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, 
      n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, 
      n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, 
      n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, 
      n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, 
      n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, 
      n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, 
      n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, 
      n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, 
      n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, 
      n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, 
      n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, 
      n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, 
      n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, 
      n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, 
      n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, 
      n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, 
      n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, 
      n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, 
      n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, 
      n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, 
      n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, 
      n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, 
      n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, 
      n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, 
      n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, 
      n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, 
      n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, 
      n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, 
      n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, 
      n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, 
      n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, 
      n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, 
      n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, 
      n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, 
      n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, 
      n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, 
      n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, 
      n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, 
      n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, 
      n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, 
      n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, 
      n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, 
      n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, 
      n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, 
      n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, 
      n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, 
      n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, 
      n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, 
      n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, 
      n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, 
      n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, 
      n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, 
      n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, 
      n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, 
      n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, 
      n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, 
      n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, 
      n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, 
      n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, 
      n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, 
      n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, 
      n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, 
      n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, 
      n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, 
      n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, 
      n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, 
      n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, 
      n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, 
      n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, 
      n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, 
      n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, 
      n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, 
      n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, 
      n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, 
      n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, 
      n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, 
      n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, 
      n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, 
      n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, 
      n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, 
      n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, 
      n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, 
      n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, 
      n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, 
      n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, 
      n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, 
      n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, 
      n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, 
      n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, 
      n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, 
      n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, 
      n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, 
      n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, 
      n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, 
      n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, 
      n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, 
      n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, 
      n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, 
      n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, 
      n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, 
      n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, 
      n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, 
      n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, 
      n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, 
      n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, 
      n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, 
      n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, 
      n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, 
      n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, 
      n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, 
      n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, 
      n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, 
      n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, 
      n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, 
      n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, 
      n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, 
      n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, 
      n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, 
      n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, 
      n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, 
      n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, 
      n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, 
      n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, 
      n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, 
      n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, 
      n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, 
      n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, 
      n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, 
      n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, 
      n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, 
      n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, 
      n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, 
      n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, 
      n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, 
      n6416, n6417, n6418, n_1000, n_1001, n_1002, n_1003, n_1004, n_1005, 
      n_1006, n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, 
      n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, 
      n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, 
      n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, 
      n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, 
      n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, 
      n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, 
      n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, 
      n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, 
      n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, 
      n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, 
      n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, 
      n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, 
      n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, 
      n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, 
      n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, 
      n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, 
      n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, 
      n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, 
      n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, 
      n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, 
      n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, 
      n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, 
      n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, 
      n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, 
      n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, 
      n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, 
      n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, 
      n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, 
      n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, 
      n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, 
      n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, 
      n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, 
      n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, 
      n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, 
      n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, 
      n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, 
      n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, 
      n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, 
      n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, 
      n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, 
      n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, 
      n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, 
      n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, 
      n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, 
      n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, 
      n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, 
      n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, 
      n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, 
      n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, 
      n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, 
      n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, 
      n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, 
      n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, 
      n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, 
      n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, n_1509, 
      n_1510, n_1511 : std_logic;

begin
   OUT1 <= ( OUT1_31_port, OUT1_30_port, OUT1_29_port, OUT1_28_port, 
      OUT1_27_port, OUT1_26_port, OUT1_25_port, OUT1_24_port, OUT1_23_port, 
      OUT1_22_port, OUT1_21_port, OUT1_20_port, OUT1_19_port, OUT1_18_port, 
      OUT1_17_port, OUT1_16_port, OUT1_15_port, OUT1_14_port, OUT1_13_port, 
      OUT1_12_port, OUT1_11_port, OUT1_10_port, OUT1_9_port, OUT1_8_port, 
      OUT1_7_port, OUT1_6_port, OUT1_5_port, OUT1_4_port, OUT1_3_port, 
      OUT1_2_port, OUT1_1_port, OUT1_0_port );
   OUT2 <= ( OUT2_31_port, OUT2_30_port, OUT2_29_port, OUT2_28_port, 
      OUT2_27_port, OUT2_26_port, OUT2_25_port, OUT2_24_port, OUT2_23_port, 
      OUT2_22_port, OUT2_21_port, OUT2_20_port, OUT2_19_port, OUT2_18_port, 
      OUT2_17_port, OUT2_16_port, OUT2_15_port, OUT2_14_port, OUT2_13_port, 
      OUT2_12_port, OUT2_11_port, OUT2_10_port, OUT2_9_port, OUT2_8_port, 
      OUT2_7_port, OUT2_6_port, OUT2_5_port, OUT2_4_port, OUT2_3_port, 
      OUT2_2_port, OUT2_1_port, OUT2_0_port );
   
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n3613, CK => CLK, Q => n4382
                           , QN => n1);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n3612, CK => CLK, Q => n4383
                           , QN => n2);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n3611, CK => CLK, Q => n4384
                           , QN => n3);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n3610, CK => CLK, Q => n4385
                           , QN => n4);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n3609, CK => CLK, Q => n4386
                           , QN => n5);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n3608, CK => CLK, Q => n4387
                           , QN => n6);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n3607, CK => CLK, Q => n4388
                           , QN => n7);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n3606, CK => CLK, Q => n4389
                           , QN => n8);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n3605, CK => CLK, Q => n4390
                           , QN => n9);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n3604, CK => CLK, Q => n4391
                           , QN => n10);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n3603, CK => CLK, Q => n4392
                           , QN => n11);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n3602, CK => CLK, Q => n4393
                           , QN => n12);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n3601, CK => CLK, Q => n4394
                           , QN => n13);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n3600, CK => CLK, Q => n4395
                           , QN => n14);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n3599, CK => CLK, Q => n4396
                           , QN => n15);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n3598, CK => CLK, Q => n4397
                           , QN => n16);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n3597, CK => CLK, Q => n4398
                           , QN => n17);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n3596, CK => CLK, Q => n4399
                           , QN => n18);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n3595, CK => CLK, Q => n4400
                           , QN => n19);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n3594, CK => CLK, Q => n4401
                           , QN => n20);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n3593, CK => CLK, Q => n4402
                           , QN => n21);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n3592, CK => CLK, Q => n4403
                           , QN => n22);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n3591, CK => CLK, Q => n4404,
                           QN => n23);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n3590, CK => CLK, Q => n4405,
                           QN => n24);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n3589, CK => CLK, Q => n4406,
                           QN => n25);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n3588, CK => CLK, Q => n4407,
                           QN => n26);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n3587, CK => CLK, Q => n4408,
                           QN => n27);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n3586, CK => CLK, Q => n4409,
                           QN => n28);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n3585, CK => CLK, Q => n4410,
                           QN => n29);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n3584, CK => CLK, Q => n4411,
                           QN => n30);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n3583, CK => CLK, Q => n4412,
                           QN => n31);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n3582, CK => CLK, Q => n4413,
                           QN => n32);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n3581, CK => CLK, Q => n4446
                           , QN => n33);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n3580, CK => CLK, Q => n4447
                           , QN => n34);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n3579, CK => CLK, Q => n4448
                           , QN => n35);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n3578, CK => CLK, Q => n4449
                           , QN => n36);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n3577, CK => CLK, Q => n4450
                           , QN => n37);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n3576, CK => CLK, Q => n4451
                           , QN => n38);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n3575, CK => CLK, Q => n4452
                           , QN => n39);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n3574, CK => CLK, Q => n4453
                           , QN => n40);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n3573, CK => CLK, Q => n4454
                           , QN => n41);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n3572, CK => CLK, Q => n4455
                           , QN => n42);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n3571, CK => CLK, Q => n4456
                           , QN => n43);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n3570, CK => CLK, Q => n4457
                           , QN => n44);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n3569, CK => CLK, Q => n4458
                           , QN => n45);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n3568, CK => CLK, Q => n4459
                           , QN => n46);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n3567, CK => CLK, Q => n4460
                           , QN => n47);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n3566, CK => CLK, Q => n4461
                           , QN => n48);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n3565, CK => CLK, Q => n4462
                           , QN => n49);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n3564, CK => CLK, Q => n4463
                           , QN => n50);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n3563, CK => CLK, Q => n4464
                           , QN => n51);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n3562, CK => CLK, Q => n4465
                           , QN => n52);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n3561, CK => CLK, Q => n4466
                           , QN => n53);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n3560, CK => CLK, Q => n4467
                           , QN => n54);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n3559, CK => CLK, Q => n4468,
                           QN => n55);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n3558, CK => CLK, Q => n4469,
                           QN => n56);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n3557, CK => CLK, Q => n4470,
                           QN => n57);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n3556, CK => CLK, Q => n4471,
                           QN => n58);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n3555, CK => CLK, Q => n4472,
                           QN => n59);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n3554, CK => CLK, Q => n4473,
                           QN => n60);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n3553, CK => CLK, Q => n4474,
                           QN => n61);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n3552, CK => CLK, Q => n4475,
                           QN => n62);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n3551, CK => CLK, Q => n4476,
                           QN => n63);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n3550, CK => CLK, Q => n4477,
                           QN => n64);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n3549, CK => CLK, Q => n6098
                           , QN => n_1000);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n3548, CK => CLK, Q => n6094
                           , QN => n_1001);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n3547, CK => CLK, Q => n6090
                           , QN => n_1002);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n3546, CK => CLK, Q => n6086
                           , QN => n_1003);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n3545, CK => CLK, Q => n6082
                           , QN => n_1004);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n3544, CK => CLK, Q => n6078
                           , QN => n_1005);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n3543, CK => CLK, Q => n6074
                           , QN => n_1006);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n3542, CK => CLK, Q => n6070
                           , QN => n_1007);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n3541, CK => CLK, Q => n6066
                           , QN => n_1008);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n3540, CK => CLK, Q => n6062
                           , QN => n_1009);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n3539, CK => CLK, Q => n6058
                           , QN => n_1010);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n3538, CK => CLK, Q => n6054
                           , QN => n_1011);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n3537, CK => CLK, Q => n6050
                           , QN => n_1012);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n3536, CK => CLK, Q => n6046
                           , QN => n_1013);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n3535, CK => CLK, Q => n6042
                           , QN => n_1014);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n3534, CK => CLK, Q => n6038
                           , QN => n_1015);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n3533, CK => CLK, Q => n6034
                           , QN => n_1016);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n3532, CK => CLK, Q => n6030
                           , QN => n_1017);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n3531, CK => CLK, Q => n6026
                           , QN => n_1018);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n3530, CK => CLK, Q => n6022
                           , QN => n_1019);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n3529, CK => CLK, Q => n6018
                           , QN => n_1020);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n3528, CK => CLK, Q => n6014
                           , QN => n_1021);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n3527, CK => CLK, Q => n6010,
                           QN => n_1022);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n3526, CK => CLK, Q => n6006,
                           QN => n_1023);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n3525, CK => CLK, Q => n6002,
                           QN => n_1024);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n3524, CK => CLK, Q => n5998,
                           QN => n_1025);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n3523, CK => CLK, Q => n5994,
                           QN => n_1026);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n3522, CK => CLK, Q => n5990,
                           QN => n_1027);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n3521, CK => CLK, Q => n5986,
                           QN => n_1028);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n3520, CK => CLK, Q => n5982,
                           QN => n_1029);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n3519, CK => CLK, Q => n5978,
                           QN => n_1030);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n3518, CK => CLK, Q => n5974,
                           QN => n_1031);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n3517, CK => CLK, Q => n6097
                           , QN => n_1032);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n3516, CK => CLK, Q => n6093
                           , QN => n_1033);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n3515, CK => CLK, Q => n6089
                           , QN => n_1034);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n3514, CK => CLK, Q => n6085
                           , QN => n_1035);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n3513, CK => CLK, Q => n6081
                           , QN => n_1036);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n3512, CK => CLK, Q => n6077
                           , QN => n_1037);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n3511, CK => CLK, Q => n6073
                           , QN => n_1038);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n3510, CK => CLK, Q => n6069
                           , QN => n_1039);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n3509, CK => CLK, Q => n6065
                           , QN => n_1040);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n3508, CK => CLK, Q => n6061
                           , QN => n_1041);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n3507, CK => CLK, Q => n6057
                           , QN => n_1042);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n3506, CK => CLK, Q => n6053
                           , QN => n_1043);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n3505, CK => CLK, Q => n6049
                           , QN => n_1044);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n3504, CK => CLK, Q => n6045
                           , QN => n_1045);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n3503, CK => CLK, Q => n6041
                           , QN => n_1046);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n3502, CK => CLK, Q => n6037
                           , QN => n_1047);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n3501, CK => CLK, Q => n6033
                           , QN => n_1048);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n3500, CK => CLK, Q => n6029
                           , QN => n_1049);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n3499, CK => CLK, Q => n6025
                           , QN => n_1050);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n3498, CK => CLK, Q => n6021
                           , QN => n_1051);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n3497, CK => CLK, Q => n6017
                           , QN => n_1052);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n3496, CK => CLK, Q => n6013
                           , QN => n_1053);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n3495, CK => CLK, Q => n6009,
                           QN => n_1054);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n3494, CK => CLK, Q => n6005,
                           QN => n_1055);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n3493, CK => CLK, Q => n6001,
                           QN => n_1056);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n3492, CK => CLK, Q => n5997,
                           QN => n_1057);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n3491, CK => CLK, Q => n5993,
                           QN => n_1058);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n3490, CK => CLK, Q => n5989,
                           QN => n_1059);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n3489, CK => CLK, Q => n5985,
                           QN => n_1060);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n3488, CK => CLK, Q => n5981,
                           QN => n_1061);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n3487, CK => CLK, Q => n5977,
                           QN => n_1062);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n3486, CK => CLK, Q => n5973,
                           QN => n_1063);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n3485, CK => CLK, Q => n4414
                           , QN => n129);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n3484, CK => CLK, Q => n4415
                           , QN => n130);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n3483, CK => CLK, Q => n4416
                           , QN => n131);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n3482, CK => CLK, Q => n4417
                           , QN => n132);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n3481, CK => CLK, Q => n4418
                           , QN => n133);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n3480, CK => CLK, Q => n4419
                           , QN => n134);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n3479, CK => CLK, Q => n4420
                           , QN => n135);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n3478, CK => CLK, Q => n4421
                           , QN => n136);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n3477, CK => CLK, Q => n4422
                           , QN => n137);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n3476, CK => CLK, Q => n4423
                           , QN => n138);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n3475, CK => CLK, Q => n4424
                           , QN => n139);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n3474, CK => CLK, Q => n4425
                           , QN => n140);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n3473, CK => CLK, Q => n4426
                           , QN => n141);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n3472, CK => CLK, Q => n4427
                           , QN => n142);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n3471, CK => CLK, Q => n4428
                           , QN => n143);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n3470, CK => CLK, Q => n4429
                           , QN => n144);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n3469, CK => CLK, Q => n4430
                           , QN => n145);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n3468, CK => CLK, Q => n4431
                           , QN => n146);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n3467, CK => CLK, Q => n4432
                           , QN => n147);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n3466, CK => CLK, Q => n4433
                           , QN => n148);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n3465, CK => CLK, Q => n4434
                           , QN => n149);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n3464, CK => CLK, Q => n4435
                           , QN => n150);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n3463, CK => CLK, Q => n4436,
                           QN => n151);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n3462, CK => CLK, Q => n4437,
                           QN => n152);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n3461, CK => CLK, Q => n4438,
                           QN => n153);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n3460, CK => CLK, Q => n4439,
                           QN => n154);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n3459, CK => CLK, Q => n4440,
                           QN => n155);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n3458, CK => CLK, Q => n4441,
                           QN => n156);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n3457, CK => CLK, Q => n4442,
                           QN => n157);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n3456, CK => CLK, Q => n4443,
                           QN => n158);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n3455, CK => CLK, Q => n4444,
                           QN => n159);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n3454, CK => CLK, Q => n4445,
                           QN => n160);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n3453, CK => CLK, Q => n4478
                           , QN => n161);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n3452, CK => CLK, Q => n4479
                           , QN => n162);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n3451, CK => CLK, Q => n4480
                           , QN => n163);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n3450, CK => CLK, Q => n4481
                           , QN => n164);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n3449, CK => CLK, Q => n4482
                           , QN => n165);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n3448, CK => CLK, Q => n4483
                           , QN => n166);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n3447, CK => CLK, Q => n4484
                           , QN => n167);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n3446, CK => CLK, Q => n4485
                           , QN => n168);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n3445, CK => CLK, Q => n4486
                           , QN => n169);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n3444, CK => CLK, Q => n4487
                           , QN => n170);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n3443, CK => CLK, Q => n4488
                           , QN => n171);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n3442, CK => CLK, Q => n4489
                           , QN => n172);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n3441, CK => CLK, Q => n4490
                           , QN => n173);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n3440, CK => CLK, Q => n4491
                           , QN => n174);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n3439, CK => CLK, Q => n4492
                           , QN => n175);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n3438, CK => CLK, Q => n4493
                           , QN => n176);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n3437, CK => CLK, Q => n4494
                           , QN => n177);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n3436, CK => CLK, Q => n4495
                           , QN => n178);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n3435, CK => CLK, Q => n4496
                           , QN => n179);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n3434, CK => CLK, Q => n4497
                           , QN => n180);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n3433, CK => CLK, Q => n4498
                           , QN => n181);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n3432, CK => CLK, Q => n4499
                           , QN => n182);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n3431, CK => CLK, Q => n4500,
                           QN => n183);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n3430, CK => CLK, Q => n4501,
                           QN => n184);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n3429, CK => CLK, Q => n4502,
                           QN => n185);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n3428, CK => CLK, Q => n4503,
                           QN => n186);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n3427, CK => CLK, Q => n4504,
                           QN => n187);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n3426, CK => CLK, Q => n4505,
                           QN => n188);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n3425, CK => CLK, Q => n4506,
                           QN => n189);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n3424, CK => CLK, Q => n4507,
                           QN => n190);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n3423, CK => CLK, Q => n4508,
                           QN => n191);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n3422, CK => CLK, Q => n4509,
                           QN => n192);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n3421, CK => CLK, Q => n6096
                           , QN => n_1064);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n3420, CK => CLK, Q => n6092
                           , QN => n_1065);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n3419, CK => CLK, Q => n6088
                           , QN => n_1066);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n3418, CK => CLK, Q => n6084
                           , QN => n_1067);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n3417, CK => CLK, Q => n6080
                           , QN => n_1068);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n3416, CK => CLK, Q => n6076
                           , QN => n_1069);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n3415, CK => CLK, Q => n6072
                           , QN => n_1070);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n3414, CK => CLK, Q => n6068
                           , QN => n_1071);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n3413, CK => CLK, Q => n6064
                           , QN => n_1072);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n3412, CK => CLK, Q => n6060
                           , QN => n_1073);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n3411, CK => CLK, Q => n6056
                           , QN => n_1074);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n3410, CK => CLK, Q => n6052
                           , QN => n_1075);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n3409, CK => CLK, Q => n6048
                           , QN => n_1076);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n3408, CK => CLK, Q => n6044
                           , QN => n_1077);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n3407, CK => CLK, Q => n6040
                           , QN => n_1078);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n3406, CK => CLK, Q => n6036
                           , QN => n_1079);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n3405, CK => CLK, Q => n6032
                           , QN => n_1080);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n3404, CK => CLK, Q => n6028
                           , QN => n_1081);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n3403, CK => CLK, Q => n6024
                           , QN => n_1082);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n3402, CK => CLK, Q => n6020
                           , QN => n_1083);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n3401, CK => CLK, Q => n6016
                           , QN => n_1084);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n3400, CK => CLK, Q => n6012
                           , QN => n_1085);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n3399, CK => CLK, Q => n6008,
                           QN => n_1086);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n3398, CK => CLK, Q => n6004,
                           QN => n_1087);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n3397, CK => CLK, Q => n6000,
                           QN => n_1088);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n3396, CK => CLK, Q => n5996,
                           QN => n_1089);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n3395, CK => CLK, Q => n5992,
                           QN => n_1090);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n3394, CK => CLK, Q => n5988,
                           QN => n_1091);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n3393, CK => CLK, Q => n5984,
                           QN => n_1092);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n3392, CK => CLK, Q => n5980,
                           QN => n_1093);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n3391, CK => CLK, Q => n5976,
                           QN => n_1094);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n3390, CK => CLK, Q => n5972,
                           QN => n_1095);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n3389, CK => CLK, Q => n6095
                           , QN => n_1096);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n3388, CK => CLK, Q => n6091
                           , QN => n_1097);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n3387, CK => CLK, Q => n6087
                           , QN => n_1098);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n3386, CK => CLK, Q => n6083
                           , QN => n_1099);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n3385, CK => CLK, Q => n6079
                           , QN => n_1100);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n3384, CK => CLK, Q => n6075
                           , QN => n_1101);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n3383, CK => CLK, Q => n6071
                           , QN => n_1102);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n3382, CK => CLK, Q => n6067
                           , QN => n_1103);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n3381, CK => CLK, Q => n6063
                           , QN => n_1104);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n3380, CK => CLK, Q => n6059
                           , QN => n_1105);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n3379, CK => CLK, Q => n6055
                           , QN => n_1106);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n3378, CK => CLK, Q => n6051
                           , QN => n_1107);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n3377, CK => CLK, Q => n6047
                           , QN => n_1108);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n3376, CK => CLK, Q => n6043
                           , QN => n_1109);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n3375, CK => CLK, Q => n6039
                           , QN => n_1110);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n3374, CK => CLK, Q => n6035
                           , QN => n_1111);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n3373, CK => CLK, Q => n6031
                           , QN => n_1112);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n3372, CK => CLK, Q => n6027
                           , QN => n_1113);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n3371, CK => CLK, Q => n6023
                           , QN => n_1114);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n3370, CK => CLK, Q => n6019
                           , QN => n_1115);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n3369, CK => CLK, Q => n6015
                           , QN => n_1116);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n3368, CK => CLK, Q => n6011
                           , QN => n_1117);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n3367, CK => CLK, Q => n6007,
                           QN => n_1118);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n3366, CK => CLK, Q => n6003,
                           QN => n_1119);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n3365, CK => CLK, Q => n5999,
                           QN => n_1120);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n3364, CK => CLK, Q => n5995,
                           QN => n_1121);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n3363, CK => CLK, Q => n5991,
                           QN => n_1122);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n3362, CK => CLK, Q => n5987,
                           QN => n_1123);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n3361, CK => CLK, Q => n5983,
                           QN => n_1124);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n3360, CK => CLK, Q => n5979,
                           QN => n_1125);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n3359, CK => CLK, Q => n5975,
                           QN => n_1126);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n3358, CK => CLK, Q => n5971,
                           QN => n_1127);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n3357, CK => CLK, Q => n3934
                           , QN => n257);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n3356, CK => CLK, Q => n3935
                           , QN => n258);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n3355, CK => CLK, Q => n3936
                           , QN => n259);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n3354, CK => CLK, Q => n3937
                           , QN => n260);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n3353, CK => CLK, Q => n3938
                           , QN => n261);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n3352, CK => CLK, Q => n3939
                           , QN => n262);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n3351, CK => CLK, Q => n3940
                           , QN => n263);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n3350, CK => CLK, Q => n3941
                           , QN => n264);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n3349, CK => CLK, Q => n3942
                           , QN => n265);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n3348, CK => CLK, Q => n3943
                           , QN => n266);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n3347, CK => CLK, Q => n3944
                           , QN => n267);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n3346, CK => CLK, Q => n3945
                           , QN => n268);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n3345, CK => CLK, Q => n3946
                           , QN => n269);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n3344, CK => CLK, Q => n3947
                           , QN => n270);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n3343, CK => CLK, Q => n3948
                           , QN => n271);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n3342, CK => CLK, Q => n3949
                           , QN => n272);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n3341, CK => CLK, Q => n3950
                           , QN => n273);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n3340, CK => CLK, Q => n3951
                           , QN => n274);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n3339, CK => CLK, Q => n3952
                           , QN => n275);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n3338, CK => CLK, Q => n3953
                           , QN => n276);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n3337, CK => CLK, Q => n3954
                           , QN => n277);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n3336, CK => CLK, Q => n3955
                           , QN => n278);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n3335, CK => CLK, Q => n3956,
                           QN => n279);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n3334, CK => CLK, Q => n3957,
                           QN => n280);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n3333, CK => CLK, Q => n3958,
                           QN => n281);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n3332, CK => CLK, Q => n3959,
                           QN => n282);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n3331, CK => CLK, Q => n3960,
                           QN => n283);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n3330, CK => CLK, Q => n3961,
                           QN => n284);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n3329, CK => CLK, Q => n3962,
                           QN => n285);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n3328, CK => CLK, Q => n3963,
                           QN => n286);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n3327, CK => CLK, Q => n3964,
                           QN => n287);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n3326, CK => CLK, Q => n3965,
                           QN => n288);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n3325, CK => CLK, Q => n4318
                           , QN => n289);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n3324, CK => CLK, Q => n4319
                           , QN => n290);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n3323, CK => CLK, Q => n4320
                           , QN => n291);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n3322, CK => CLK, Q => n4321
                           , QN => n292);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n3321, CK => CLK, Q => n4322
                           , QN => n293);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n3320, CK => CLK, Q => n4323
                           , QN => n294);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n3319, CK => CLK, Q => n4324
                           , QN => n295);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n3318, CK => CLK, Q => n4325
                           , QN => n296);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n3317, CK => CLK, Q => n4326
                           , QN => n297);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n3316, CK => CLK, Q => n4327
                           , QN => n298);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n3315, CK => CLK, Q => n4328
                           , QN => n299);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n3314, CK => CLK, Q => n4329
                           , QN => n300);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n3313, CK => CLK, Q => n4330
                           , QN => n301);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n3312, CK => CLK, Q => n4331
                           , QN => n302);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n3311, CK => CLK, Q => n4332
                           , QN => n303);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n3310, CK => CLK, Q => n4333
                           , QN => n304);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n3309, CK => CLK, Q => n4334
                           , QN => n305);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n3308, CK => CLK, Q => n4335
                           , QN => n306);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n3307, CK => CLK, Q => n4336
                           , QN => n307);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n3306, CK => CLK, Q => n4337
                           , QN => n308);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n3305, CK => CLK, Q => n4338
                           , QN => n309);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n3304, CK => CLK, Q => n4339
                           , QN => n310);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n3303, CK => CLK, Q => n4340,
                           QN => n311);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n3302, CK => CLK, Q => n4341,
                           QN => n312);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n3301, CK => CLK, Q => n4342,
                           QN => n313);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n3300, CK => CLK, Q => n4343,
                           QN => n314);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n3299, CK => CLK, Q => n4344,
                           QN => n315);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n3298, CK => CLK, Q => n4345,
                           QN => n316);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n3297, CK => CLK, Q => n4346,
                           QN => n317);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n3296, CK => CLK, Q => n4347,
                           QN => n318);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n3295, CK => CLK, Q => n4348,
                           QN => n319);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n3294, CK => CLK, Q => n4349,
                           QN => n320);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n3293, CK => CLK, Q => 
                           n3966, QN => n321);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n3292, CK => CLK, Q => 
                           n3967, QN => n322);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n3291, CK => CLK, Q => 
                           n3968, QN => n323);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n3290, CK => CLK, Q => 
                           n3969, QN => n324);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n3289, CK => CLK, Q => 
                           n3970, QN => n325);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n3288, CK => CLK, Q => 
                           n3971, QN => n326);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n3287, CK => CLK, Q => 
                           n3972, QN => n327);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n3286, CK => CLK, Q => 
                           n3973, QN => n328);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n3285, CK => CLK, Q => 
                           n3974, QN => n329);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n3284, CK => CLK, Q => 
                           n3975, QN => n330);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n3283, CK => CLK, Q => 
                           n3976, QN => n331);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n3282, CK => CLK, Q => 
                           n3977, QN => n332);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n3281, CK => CLK, Q => 
                           n3978, QN => n333);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n3280, CK => CLK, Q => 
                           n3979, QN => n334);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n3279, CK => CLK, Q => 
                           n3980, QN => n335);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n3278, CK => CLK, Q => 
                           n3981, QN => n336);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n3277, CK => CLK, Q => 
                           n3982, QN => n337);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n3276, CK => CLK, Q => 
                           n3983, QN => n338);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n3275, CK => CLK, Q => 
                           n3984, QN => n339);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n3274, CK => CLK, Q => 
                           n3985, QN => n340);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n3273, CK => CLK, Q => 
                           n3986, QN => n341);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n3272, CK => CLK, Q => 
                           n3987, QN => n342);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n3271, CK => CLK, Q => n3988
                           , QN => n343);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n3270, CK => CLK, Q => n3989
                           , QN => n344);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n3269, CK => CLK, Q => n3990
                           , QN => n345);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n3268, CK => CLK, Q => n3991
                           , QN => n346);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n3267, CK => CLK, Q => n3992
                           , QN => n347);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n3266, CK => CLK, Q => n3993
                           , QN => n348);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n3265, CK => CLK, Q => n3994
                           , QN => n349);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n3264, CK => CLK, Q => n3995
                           , QN => n350);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n3263, CK => CLK, Q => n3996
                           , QN => n351);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n3262, CK => CLK, Q => n3997
                           , QN => n352);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n3261, CK => CLK, Q => 
                           n4350, QN => n353);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n3260, CK => CLK, Q => 
                           n4351, QN => n354);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n3259, CK => CLK, Q => 
                           n4352, QN => n355);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n3258, CK => CLK, Q => 
                           n4353, QN => n356);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n3257, CK => CLK, Q => 
                           n4354, QN => n357);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n3256, CK => CLK, Q => 
                           n4355, QN => n358);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n3255, CK => CLK, Q => 
                           n4356, QN => n359);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n3254, CK => CLK, Q => 
                           n4357, QN => n360);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n3253, CK => CLK, Q => 
                           n4358, QN => n361);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n3252, CK => CLK, Q => 
                           n4359, QN => n362);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n3251, CK => CLK, Q => 
                           n4360, QN => n363);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n3250, CK => CLK, Q => 
                           n4361, QN => n364);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n3249, CK => CLK, Q => 
                           n4362, QN => n365);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n3248, CK => CLK, Q => 
                           n4363, QN => n366);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n3247, CK => CLK, Q => 
                           n4364, QN => n367);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n3246, CK => CLK, Q => 
                           n4365, QN => n368);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n3245, CK => CLK, Q => 
                           n4366, QN => n369);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n3244, CK => CLK, Q => 
                           n4367, QN => n370);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n3243, CK => CLK, Q => 
                           n4368, QN => n371);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n3242, CK => CLK, Q => 
                           n4369, QN => n372);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n3241, CK => CLK, Q => 
                           n4370, QN => n373);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n3240, CK => CLK, Q => 
                           n4371, QN => n374);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n3239, CK => CLK, Q => n4372
                           , QN => n375);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n3238, CK => CLK, Q => n4373
                           , QN => n376);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n3237, CK => CLK, Q => n4374
                           , QN => n377);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n3236, CK => CLK, Q => n4375
                           , QN => n378);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n3235, CK => CLK, Q => n4376
                           , QN => n379);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n3234, CK => CLK, Q => n4377
                           , QN => n380);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n3233, CK => CLK, Q => n4378
                           , QN => n381);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n3232, CK => CLK, Q => n4379
                           , QN => n382);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n3231, CK => CLK, Q => n4380
                           , QN => n383);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n3230, CK => CLK, Q => n4381
                           , QN => n384);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n3229, CK => CLK, Q => 
                           n3614, QN => n_1128);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n3228, CK => CLK, Q => 
                           n3619, QN => n_1129);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n3227, CK => CLK, Q => 
                           n3624, QN => n_1130);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n3226, CK => CLK, Q => 
                           n3629, QN => n_1131);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n3225, CK => CLK, Q => 
                           n3634, QN => n_1132);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n3224, CK => CLK, Q => 
                           n3639, QN => n_1133);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n3223, CK => CLK, Q => 
                           n3644, QN => n_1134);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n3222, CK => CLK, Q => 
                           n3649, QN => n_1135);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n3221, CK => CLK, Q => 
                           n3654, QN => n_1136);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n3220, CK => CLK, Q => 
                           n3659, QN => n_1137);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n3219, CK => CLK, Q => 
                           n3664, QN => n_1138);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n3218, CK => CLK, Q => 
                           n3669, QN => n_1139);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n3217, CK => CLK, Q => 
                           n3674, QN => n_1140);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n3216, CK => CLK, Q => 
                           n3679, QN => n_1141);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n3215, CK => CLK, Q => 
                           n3684, QN => n_1142);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n3214, CK => CLK, Q => 
                           n3689, QN => n_1143);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n3213, CK => CLK, Q => 
                           n3694, QN => n_1144);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n3212, CK => CLK, Q => 
                           n3699, QN => n_1145);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n3211, CK => CLK, Q => 
                           n3704, QN => n_1146);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n3210, CK => CLK, Q => 
                           n3709, QN => n_1147);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n3209, CK => CLK, Q => 
                           n3714, QN => n_1148);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n3208, CK => CLK, Q => 
                           n3719, QN => n_1149);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n3207, CK => CLK, Q => n3724
                           , QN => n_1150);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n3206, CK => CLK, Q => n3729
                           , QN => n_1151);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n3205, CK => CLK, Q => n3734
                           , QN => n_1152);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n3204, CK => CLK, Q => n3739
                           , QN => n_1153);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n3203, CK => CLK, Q => n3744
                           , QN => n_1154);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n3202, CK => CLK, Q => n3749
                           , QN => n_1155);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n3201, CK => CLK, Q => n3754
                           , QN => n_1156);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n3200, CK => CLK, Q => n3759
                           , QN => n_1157);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n3199, CK => CLK, Q => n3764
                           , QN => n_1158);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n3198, CK => CLK, Q => n3769
                           , QN => n_1159);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n3197, CK => CLK, Q => 
                           n3998, QN => n_1160);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n3196, CK => CLK, Q => 
                           n4003, QN => n_1161);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n3195, CK => CLK, Q => 
                           n4008, QN => n_1162);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n3194, CK => CLK, Q => 
                           n4013, QN => n_1163);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n3193, CK => CLK, Q => 
                           n4018, QN => n_1164);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n3192, CK => CLK, Q => 
                           n4023, QN => n_1165);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n3191, CK => CLK, Q => 
                           n4028, QN => n_1166);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n3190, CK => CLK, Q => 
                           n4033, QN => n_1167);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n3189, CK => CLK, Q => 
                           n4038, QN => n_1168);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n3188, CK => CLK, Q => 
                           n4043, QN => n_1169);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n3187, CK => CLK, Q => 
                           n4048, QN => n_1170);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n3186, CK => CLK, Q => 
                           n4053, QN => n_1171);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n3185, CK => CLK, Q => 
                           n4058, QN => n_1172);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n3184, CK => CLK, Q => 
                           n4063, QN => n_1173);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n3183, CK => CLK, Q => 
                           n4068, QN => n_1174);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n3182, CK => CLK, Q => 
                           n4073, QN => n_1175);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n3181, CK => CLK, Q => 
                           n4078, QN => n_1176);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n3180, CK => CLK, Q => 
                           n4083, QN => n_1177);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n3179, CK => CLK, Q => 
                           n4088, QN => n_1178);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n3178, CK => CLK, Q => 
                           n4093, QN => n_1179);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n3177, CK => CLK, Q => 
                           n4098, QN => n_1180);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n3176, CK => CLK, Q => 
                           n4103, QN => n_1181);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n3175, CK => CLK, Q => n4108
                           , QN => n_1182);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n3174, CK => CLK, Q => n4113
                           , QN => n_1183);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n3173, CK => CLK, Q => n4118
                           , QN => n_1184);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n3172, CK => CLK, Q => n4123
                           , QN => n_1185);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n3171, CK => CLK, Q => n4128
                           , QN => n_1186);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n3170, CK => CLK, Q => n4133
                           , QN => n_1187);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n3169, CK => CLK, Q => n4138
                           , QN => n_1188);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n3168, CK => CLK, Q => n4143
                           , QN => n_1189);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n3167, CK => CLK, Q => n4148
                           , QN => n_1190);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n3166, CK => CLK, Q => n4153
                           , QN => n_1191);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n3165, CK => CLK, Q => 
                           n6418, QN => n4158);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n3164, CK => CLK, Q => 
                           n6417, QN => n4163);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n3163, CK => CLK, Q => 
                           n6416, QN => n4168);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n3162, CK => CLK, Q => 
                           n6415, QN => n4173);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n3161, CK => CLK, Q => 
                           n6414, QN => n4178);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n3160, CK => CLK, Q => 
                           n6413, QN => n4183);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n3159, CK => CLK, Q => 
                           n6412, QN => n4188);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n3158, CK => CLK, Q => 
                           n6411, QN => n4193);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n3157, CK => CLK, Q => 
                           n6410, QN => n4198);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n3156, CK => CLK, Q => 
                           n6409, QN => n4203);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n3155, CK => CLK, Q => 
                           n6408, QN => n4208);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n3154, CK => CLK, Q => 
                           n6407, QN => n4213);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n3153, CK => CLK, Q => 
                           n6406, QN => n4218);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n3152, CK => CLK, Q => 
                           n6405, QN => n4223);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n3151, CK => CLK, Q => 
                           n6404, QN => n4228);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n3150, CK => CLK, Q => 
                           n6403, QN => n4233);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n3149, CK => CLK, Q => 
                           n6402, QN => n4238);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n3148, CK => CLK, Q => 
                           n6401, QN => n4243);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n3147, CK => CLK, Q => 
                           n6400, QN => n4248);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n3146, CK => CLK, Q => 
                           n6399, QN => n4253);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n3145, CK => CLK, Q => 
                           n6398, QN => n4258);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n3144, CK => CLK, Q => 
                           n6397, QN => n4263);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n3143, CK => CLK, Q => n6396
                           , QN => n4268);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n3142, CK => CLK, Q => n6395
                           , QN => n4273);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n3141, CK => CLK, Q => n6394
                           , QN => n4278);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n3140, CK => CLK, Q => n6393
                           , QN => n4283);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n3139, CK => CLK, Q => n6392
                           , QN => n4288);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n3138, CK => CLK, Q => n6391
                           , QN => n4293);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n3137, CK => CLK, Q => n6390
                           , QN => n4298);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n3136, CK => CLK, Q => n6389
                           , QN => n4303);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n3135, CK => CLK, Q => n6388
                           , QN => n4308);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n3134, CK => CLK, Q => n6387
                           , QN => n4313);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n3133, CK => CLK, Q => 
                           n6386, QN => n3774);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n3132, CK => CLK, Q => 
                           n6385, QN => n3779);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n3131, CK => CLK, Q => 
                           n6384, QN => n3784);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n3130, CK => CLK, Q => 
                           n6383, QN => n3789);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n3129, CK => CLK, Q => 
                           n6382, QN => n3794);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n3128, CK => CLK, Q => 
                           n6381, QN => n3799);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n3127, CK => CLK, Q => 
                           n6380, QN => n3804);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n3126, CK => CLK, Q => 
                           n6379, QN => n3809);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n3125, CK => CLK, Q => 
                           n6378, QN => n3814);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n3124, CK => CLK, Q => 
                           n6377, QN => n3819);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n3123, CK => CLK, Q => 
                           n6376, QN => n3824);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n3122, CK => CLK, Q => 
                           n6375, QN => n3829);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n3121, CK => CLK, Q => 
                           n6374, QN => n3834);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n3120, CK => CLK, Q => 
                           n6373, QN => n3839);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n3119, CK => CLK, Q => 
                           n6372, QN => n3844);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n3118, CK => CLK, Q => 
                           n6371, QN => n3849);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n3117, CK => CLK, Q => 
                           n6370, QN => n3854);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n3116, CK => CLK, Q => 
                           n6369, QN => n3859);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n3115, CK => CLK, Q => 
                           n6368, QN => n3864);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n3114, CK => CLK, Q => 
                           n6367, QN => n3869);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n3113, CK => CLK, Q => 
                           n6366, QN => n3874);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n3112, CK => CLK, Q => 
                           n6365, QN => n3879);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n3111, CK => CLK, Q => n6364
                           , QN => n3884);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n3110, CK => CLK, Q => n6363
                           , QN => n3889);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n3109, CK => CLK, Q => n6362
                           , QN => n3894);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n3108, CK => CLK, Q => n6361
                           , QN => n3899);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n3107, CK => CLK, Q => n6360
                           , QN => n3904);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n3106, CK => CLK, Q => n6359
                           , QN => n3909);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n3105, CK => CLK, Q => n6358
                           , QN => n3914);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n3104, CK => CLK, Q => n6357
                           , QN => n3919);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n3103, CK => CLK, Q => n6356
                           , QN => n3924);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n3102, CK => CLK, Q => n6355
                           , QN => n3929);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n3101, CK => CLK, Q => 
                           n3615, QN => n_1192);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n3100, CK => CLK, Q => 
                           n3620, QN => n_1193);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n3099, CK => CLK, Q => 
                           n3625, QN => n_1194);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n3098, CK => CLK, Q => 
                           n3630, QN => n_1195);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n3097, CK => CLK, Q => 
                           n3635, QN => n_1196);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n3096, CK => CLK, Q => 
                           n3640, QN => n_1197);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n3095, CK => CLK, Q => 
                           n3645, QN => n_1198);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n3094, CK => CLK, Q => 
                           n3650, QN => n_1199);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n3093, CK => CLK, Q => 
                           n3655, QN => n_1200);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n3092, CK => CLK, Q => 
                           n3660, QN => n_1201);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n3091, CK => CLK, Q => 
                           n3665, QN => n_1202);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n3090, CK => CLK, Q => 
                           n3670, QN => n_1203);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n3089, CK => CLK, Q => 
                           n3675, QN => n_1204);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n3088, CK => CLK, Q => 
                           n3680, QN => n_1205);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n3087, CK => CLK, Q => 
                           n3685, QN => n_1206);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n3086, CK => CLK, Q => 
                           n3690, QN => n_1207);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n3085, CK => CLK, Q => 
                           n3695, QN => n_1208);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n3084, CK => CLK, Q => 
                           n3700, QN => n_1209);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n3083, CK => CLK, Q => 
                           n3705, QN => n_1210);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n3082, CK => CLK, Q => 
                           n3710, QN => n_1211);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n3081, CK => CLK, Q => 
                           n3715, QN => n_1212);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n3080, CK => CLK, Q => 
                           n3720, QN => n_1213);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n3079, CK => CLK, Q => n3725
                           , QN => n_1214);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n3078, CK => CLK, Q => n3730
                           , QN => n_1215);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n3077, CK => CLK, Q => n3735
                           , QN => n_1216);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n3076, CK => CLK, Q => n3740
                           , QN => n_1217);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n3075, CK => CLK, Q => n3745
                           , QN => n_1218);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n3074, CK => CLK, Q => n3750
                           , QN => n_1219);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n3073, CK => CLK, Q => n3755
                           , QN => n_1220);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n3072, CK => CLK, Q => n3760
                           , QN => n_1221);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n3071, CK => CLK, Q => n3765
                           , QN => n_1222);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n3070, CK => CLK, Q => n3770
                           , QN => n_1223);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n3069, CK => CLK, Q => 
                           n3999, QN => n_1224);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n3068, CK => CLK, Q => 
                           n4004, QN => n_1225);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n3067, CK => CLK, Q => 
                           n4009, QN => n_1226);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n3066, CK => CLK, Q => 
                           n4014, QN => n_1227);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n3065, CK => CLK, Q => 
                           n4019, QN => n_1228);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n3064, CK => CLK, Q => 
                           n4024, QN => n_1229);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n3063, CK => CLK, Q => 
                           n4029, QN => n_1230);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n3062, CK => CLK, Q => 
                           n4034, QN => n_1231);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n3061, CK => CLK, Q => 
                           n4039, QN => n_1232);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n3060, CK => CLK, Q => 
                           n4044, QN => n_1233);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n3059, CK => CLK, Q => 
                           n4049, QN => n_1234);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n3058, CK => CLK, Q => 
                           n4054, QN => n_1235);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n3057, CK => CLK, Q => 
                           n4059, QN => n_1236);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n3056, CK => CLK, Q => 
                           n4064, QN => n_1237);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n3055, CK => CLK, Q => 
                           n4069, QN => n_1238);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n3054, CK => CLK, Q => 
                           n4074, QN => n_1239);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n3053, CK => CLK, Q => 
                           n4079, QN => n_1240);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n3052, CK => CLK, Q => 
                           n4084, QN => n_1241);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n3051, CK => CLK, Q => 
                           n4089, QN => n_1242);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n3050, CK => CLK, Q => 
                           n4094, QN => n_1243);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n3049, CK => CLK, Q => 
                           n4099, QN => n_1244);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n3048, CK => CLK, Q => 
                           n4104, QN => n_1245);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n3047, CK => CLK, Q => n4109
                           , QN => n_1246);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n3046, CK => CLK, Q => n4114
                           , QN => n_1247);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n3045, CK => CLK, Q => n4119
                           , QN => n_1248);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n3044, CK => CLK, Q => n4124
                           , QN => n_1249);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n3043, CK => CLK, Q => n4129
                           , QN => n_1250);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n3042, CK => CLK, Q => n4134
                           , QN => n_1251);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n3041, CK => CLK, Q => n4139
                           , QN => n_1252);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n3040, CK => CLK, Q => n4144
                           , QN => n_1253);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n3039, CK => CLK, Q => n4149
                           , QN => n_1254);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n3038, CK => CLK, Q => n4154
                           , QN => n_1255);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n3037, CK => CLK, Q => 
                           n6354, QN => n4159);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n3036, CK => CLK, Q => 
                           n6353, QN => n4164);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n3035, CK => CLK, Q => 
                           n6352, QN => n4169);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n3034, CK => CLK, Q => 
                           n6351, QN => n4174);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n3033, CK => CLK, Q => 
                           n6350, QN => n4179);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n3032, CK => CLK, Q => 
                           n6349, QN => n4184);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n3031, CK => CLK, Q => 
                           n6348, QN => n4189);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n3030, CK => CLK, Q => 
                           n6347, QN => n4194);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n3029, CK => CLK, Q => 
                           n6346, QN => n4199);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n3028, CK => CLK, Q => 
                           n6345, QN => n4204);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n3027, CK => CLK, Q => 
                           n6344, QN => n4209);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n3026, CK => CLK, Q => 
                           n6343, QN => n4214);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n3025, CK => CLK, Q => 
                           n6342, QN => n4219);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n3024, CK => CLK, Q => 
                           n6341, QN => n4224);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n3023, CK => CLK, Q => 
                           n6340, QN => n4229);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n3022, CK => CLK, Q => 
                           n6339, QN => n4234);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n3021, CK => CLK, Q => 
                           n6338, QN => n4239);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n3020, CK => CLK, Q => 
                           n6337, QN => n4244);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n3019, CK => CLK, Q => 
                           n6336, QN => n4249);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n3018, CK => CLK, Q => 
                           n6335, QN => n4254);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n3017, CK => CLK, Q => 
                           n6334, QN => n4259);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n3016, CK => CLK, Q => 
                           n6333, QN => n4264);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n3015, CK => CLK, Q => n6332
                           , QN => n4269);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n3014, CK => CLK, Q => n6331
                           , QN => n4274);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n3013, CK => CLK, Q => n6330
                           , QN => n4279);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n3012, CK => CLK, Q => n6329
                           , QN => n4284);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n3011, CK => CLK, Q => n6328
                           , QN => n4289);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n3010, CK => CLK, Q => n6327
                           , QN => n4294);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n3009, CK => CLK, Q => n6326
                           , QN => n4299);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n3008, CK => CLK, Q => n6325
                           , QN => n4304);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n3007, CK => CLK, Q => n6324
                           , QN => n4309);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n3006, CK => CLK, Q => n6323
                           , QN => n4314);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n3005, CK => CLK, Q => 
                           n6322, QN => n3775);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n3004, CK => CLK, Q => 
                           n6321, QN => n3780);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n3003, CK => CLK, Q => 
                           n6320, QN => n3785);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n3002, CK => CLK, Q => 
                           n6319, QN => n3790);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n3001, CK => CLK, Q => 
                           n6318, QN => n3795);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n3000, CK => CLK, Q => 
                           n6317, QN => n3800);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n2999, CK => CLK, Q => 
                           n6316, QN => n3805);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n2998, CK => CLK, Q => 
                           n6315, QN => n3810);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n2997, CK => CLK, Q => 
                           n6314, QN => n3815);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n2996, CK => CLK, Q => 
                           n6313, QN => n3820);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n2995, CK => CLK, Q => 
                           n6312, QN => n3825);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n2994, CK => CLK, Q => 
                           n6311, QN => n3830);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n2993, CK => CLK, Q => 
                           n6310, QN => n3835);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n2992, CK => CLK, Q => 
                           n6309, QN => n3840);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n2991, CK => CLK, Q => 
                           n6308, QN => n3845);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n2990, CK => CLK, Q => 
                           n6307, QN => n3850);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n2989, CK => CLK, Q => 
                           n6306, QN => n3855);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n2988, CK => CLK, Q => 
                           n6305, QN => n3860);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n2987, CK => CLK, Q => 
                           n6304, QN => n3865);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n2986, CK => CLK, Q => 
                           n6303, QN => n3870);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n2985, CK => CLK, Q => 
                           n6302, QN => n3875);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n2984, CK => CLK, Q => 
                           n6301, QN => n3880);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n2983, CK => CLK, Q => n6300
                           , QN => n3885);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n2982, CK => CLK, Q => n6299
                           , QN => n3890);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n2981, CK => CLK, Q => n6298
                           , QN => n3895);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n2980, CK => CLK, Q => n6297
                           , QN => n3900);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n2979, CK => CLK, Q => n6296
                           , QN => n3905);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n2978, CK => CLK, Q => n6295
                           , QN => n3910);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n2977, CK => CLK, Q => n6294
                           , QN => n3915);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n2976, CK => CLK, Q => n6293
                           , QN => n3920);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n2975, CK => CLK, Q => n6292
                           , QN => n3925);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n2974, CK => CLK, Q => n6291
                           , QN => n3930);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n2973, CK => CLK, Q => 
                           n3616, QN => n_1256);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n2972, CK => CLK, Q => 
                           n3621, QN => n_1257);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n2971, CK => CLK, Q => 
                           n3626, QN => n_1258);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n2970, CK => CLK, Q => 
                           n3631, QN => n_1259);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n2969, CK => CLK, Q => 
                           n3636, QN => n_1260);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n2968, CK => CLK, Q => 
                           n3641, QN => n_1261);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n2967, CK => CLK, Q => 
                           n3646, QN => n_1262);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n2966, CK => CLK, Q => 
                           n3651, QN => n_1263);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n2965, CK => CLK, Q => 
                           n3656, QN => n_1264);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n2964, CK => CLK, Q => 
                           n3661, QN => n_1265);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n2963, CK => CLK, Q => 
                           n3666, QN => n_1266);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n2962, CK => CLK, Q => 
                           n3671, QN => n_1267);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n2961, CK => CLK, Q => 
                           n3676, QN => n_1268);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n2960, CK => CLK, Q => 
                           n3681, QN => n_1269);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n2959, CK => CLK, Q => 
                           n3686, QN => n_1270);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n2958, CK => CLK, Q => 
                           n3691, QN => n_1271);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n2957, CK => CLK, Q => 
                           n3696, QN => n_1272);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n2956, CK => CLK, Q => 
                           n3701, QN => n_1273);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n2955, CK => CLK, Q => 
                           n3706, QN => n_1274);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n2954, CK => CLK, Q => 
                           n3711, QN => n_1275);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n2953, CK => CLK, Q => 
                           n3716, QN => n_1276);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n2952, CK => CLK, Q => 
                           n3721, QN => n_1277);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n2951, CK => CLK, Q => n3726
                           , QN => n_1278);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n2950, CK => CLK, Q => n3731
                           , QN => n_1279);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n2949, CK => CLK, Q => n3736
                           , QN => n_1280);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n2948, CK => CLK, Q => n3741
                           , QN => n_1281);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n2947, CK => CLK, Q => n3746
                           , QN => n_1282);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n2946, CK => CLK, Q => n3751
                           , QN => n_1283);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n2945, CK => CLK, Q => n3756
                           , QN => n_1284);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n2944, CK => CLK, Q => n3761
                           , QN => n_1285);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n2943, CK => CLK, Q => n3766
                           , QN => n_1286);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n2942, CK => CLK, Q => n3771
                           , QN => n_1287);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n2941, CK => CLK, Q => 
                           n4000, QN => n_1288);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n2940, CK => CLK, Q => 
                           n4005, QN => n_1289);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n2939, CK => CLK, Q => 
                           n4010, QN => n_1290);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n2938, CK => CLK, Q => 
                           n4015, QN => n_1291);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n2937, CK => CLK, Q => 
                           n4020, QN => n_1292);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n2936, CK => CLK, Q => 
                           n4025, QN => n_1293);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n2935, CK => CLK, Q => 
                           n4030, QN => n_1294);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n2934, CK => CLK, Q => 
                           n4035, QN => n_1295);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n2933, CK => CLK, Q => 
                           n4040, QN => n_1296);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n2932, CK => CLK, Q => 
                           n4045, QN => n_1297);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n2931, CK => CLK, Q => 
                           n4050, QN => n_1298);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n2930, CK => CLK, Q => 
                           n4055, QN => n_1299);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n2929, CK => CLK, Q => 
                           n4060, QN => n_1300);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n2928, CK => CLK, Q => 
                           n4065, QN => n_1301);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n2927, CK => CLK, Q => 
                           n4070, QN => n_1302);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n2926, CK => CLK, Q => 
                           n4075, QN => n_1303);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n2925, CK => CLK, Q => 
                           n4080, QN => n_1304);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n2924, CK => CLK, Q => 
                           n4085, QN => n_1305);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n2923, CK => CLK, Q => 
                           n4090, QN => n_1306);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n2922, CK => CLK, Q => 
                           n4095, QN => n_1307);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n2921, CK => CLK, Q => 
                           n4100, QN => n_1308);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n2920, CK => CLK, Q => 
                           n4105, QN => n_1309);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n2919, CK => CLK, Q => n4110
                           , QN => n_1310);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n2918, CK => CLK, Q => n4115
                           , QN => n_1311);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n2917, CK => CLK, Q => n4120
                           , QN => n_1312);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n2916, CK => CLK, Q => n4125
                           , QN => n_1313);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n2915, CK => CLK, Q => n4130
                           , QN => n_1314);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n2914, CK => CLK, Q => n4135
                           , QN => n_1315);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n2913, CK => CLK, Q => n4140
                           , QN => n_1316);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n2912, CK => CLK, Q => n4145
                           , QN => n_1317);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n2911, CK => CLK, Q => n4150
                           , QN => n_1318);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n2910, CK => CLK, Q => n4155
                           , QN => n_1319);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n2909, CK => CLK, Q => 
                           n6290, QN => n4160);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n2908, CK => CLK, Q => 
                           n6289, QN => n4165);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n2907, CK => CLK, Q => 
                           n6288, QN => n4170);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n2906, CK => CLK, Q => 
                           n6287, QN => n4175);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n2905, CK => CLK, Q => 
                           n6286, QN => n4180);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n2904, CK => CLK, Q => 
                           n6285, QN => n4185);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n2903, CK => CLK, Q => 
                           n6284, QN => n4190);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n2902, CK => CLK, Q => 
                           n6283, QN => n4195);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n2901, CK => CLK, Q => 
                           n6282, QN => n4200);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n2900, CK => CLK, Q => 
                           n6281, QN => n4205);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n2899, CK => CLK, Q => 
                           n6280, QN => n4210);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n2898, CK => CLK, Q => 
                           n6279, QN => n4215);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n2897, CK => CLK, Q => 
                           n6278, QN => n4220);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n2896, CK => CLK, Q => 
                           n6277, QN => n4225);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n2895, CK => CLK, Q => 
                           n6276, QN => n4230);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n2894, CK => CLK, Q => 
                           n6275, QN => n4235);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n2893, CK => CLK, Q => 
                           n6274, QN => n4240);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n2892, CK => CLK, Q => 
                           n6273, QN => n4245);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n2891, CK => CLK, Q => 
                           n6272, QN => n4250);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n2890, CK => CLK, Q => 
                           n6271, QN => n4255);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n2889, CK => CLK, Q => 
                           n6270, QN => n4260);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n2888, CK => CLK, Q => 
                           n6269, QN => n4265);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n2887, CK => CLK, Q => n6268
                           , QN => n4270);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n2886, CK => CLK, Q => n6267
                           , QN => n4275);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n2885, CK => CLK, Q => n6266
                           , QN => n4280);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n2884, CK => CLK, Q => n6265
                           , QN => n4285);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n2883, CK => CLK, Q => n6264
                           , QN => n4290);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n2882, CK => CLK, Q => n6263
                           , QN => n4295);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n2881, CK => CLK, Q => n6262
                           , QN => n4300);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n2880, CK => CLK, Q => n6261
                           , QN => n4305);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n2879, CK => CLK, Q => n6260
                           , QN => n4310);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n2878, CK => CLK, Q => n6259
                           , QN => n4315);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n2877, CK => CLK, Q => 
                           n6258, QN => n3776);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n2876, CK => CLK, Q => 
                           n6257, QN => n3781);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n2875, CK => CLK, Q => 
                           n6256, QN => n3786);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n2874, CK => CLK, Q => 
                           n6255, QN => n3791);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n2873, CK => CLK, Q => 
                           n6254, QN => n3796);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n2872, CK => CLK, Q => 
                           n6253, QN => n3801);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n2871, CK => CLK, Q => 
                           n6252, QN => n3806);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n2870, CK => CLK, Q => 
                           n6251, QN => n3811);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n2869, CK => CLK, Q => 
                           n6250, QN => n3816);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n2868, CK => CLK, Q => 
                           n6249, QN => n3821);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n2867, CK => CLK, Q => 
                           n6248, QN => n3826);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n2866, CK => CLK, Q => 
                           n6247, QN => n3831);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n2865, CK => CLK, Q => 
                           n6246, QN => n3836);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n2864, CK => CLK, Q => 
                           n6245, QN => n3841);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n2863, CK => CLK, Q => 
                           n6244, QN => n3846);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n2862, CK => CLK, Q => 
                           n6243, QN => n3851);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n2861, CK => CLK, Q => 
                           n6242, QN => n3856);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n2860, CK => CLK, Q => 
                           n6241, QN => n3861);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n2859, CK => CLK, Q => 
                           n6240, QN => n3866);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n2858, CK => CLK, Q => 
                           n6239, QN => n3871);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n2857, CK => CLK, Q => 
                           n6238, QN => n3876);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n2856, CK => CLK, Q => 
                           n6237, QN => n3881);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n2855, CK => CLK, Q => n6236
                           , QN => n3886);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n2854, CK => CLK, Q => n6235
                           , QN => n3891);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n2853, CK => CLK, Q => n6234
                           , QN => n3896);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n2852, CK => CLK, Q => n6233
                           , QN => n3901);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n2851, CK => CLK, Q => n6232
                           , QN => n3906);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n2850, CK => CLK, Q => n6231
                           , QN => n3911);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n2849, CK => CLK, Q => n6230
                           , QN => n3916);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n2848, CK => CLK, Q => n6229
                           , QN => n3921);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n2847, CK => CLK, Q => n6228
                           , QN => n3926);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n2846, CK => CLK, Q => n6227
                           , QN => n3931);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n2845, CK => CLK, Q => 
                           n6226, QN => n4161);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n2844, CK => CLK, Q => 
                           n6225, QN => n4166);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n2843, CK => CLK, Q => 
                           n6224, QN => n4171);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n2842, CK => CLK, Q => 
                           n6223, QN => n4176);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n2841, CK => CLK, Q => 
                           n6222, QN => n4181);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n2840, CK => CLK, Q => 
                           n6221, QN => n4186);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n2839, CK => CLK, Q => 
                           n6220, QN => n4191);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n2838, CK => CLK, Q => 
                           n6219, QN => n4196);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n2837, CK => CLK, Q => 
                           n6218, QN => n4201);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n2836, CK => CLK, Q => 
                           n6217, QN => n4206);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n2835, CK => CLK, Q => 
                           n6216, QN => n4211);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n2834, CK => CLK, Q => 
                           n6215, QN => n4216);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n2833, CK => CLK, Q => 
                           n6214, QN => n4221);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n2832, CK => CLK, Q => 
                           n6213, QN => n4226);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n2831, CK => CLK, Q => 
                           n6212, QN => n4231);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n2830, CK => CLK, Q => 
                           n6211, QN => n4236);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n2829, CK => CLK, Q => 
                           n6210, QN => n4241);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n2828, CK => CLK, Q => 
                           n6209, QN => n4246);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n2827, CK => CLK, Q => 
                           n6208, QN => n4251);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n2826, CK => CLK, Q => 
                           n6207, QN => n4256);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n2825, CK => CLK, Q => 
                           n6206, QN => n4261);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n2824, CK => CLK, Q => 
                           n6205, QN => n4266);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n2823, CK => CLK, Q => n6204
                           , QN => n4271);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n2822, CK => CLK, Q => n6203
                           , QN => n4276);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n2821, CK => CLK, Q => n6202
                           , QN => n4281);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n2820, CK => CLK, Q => n6201
                           , QN => n4286);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n2819, CK => CLK, Q => n6200
                           , QN => n4291);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n2818, CK => CLK, Q => n6199
                           , QN => n4296);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n2817, CK => CLK, Q => n6198
                           , QN => n4301);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n2816, CK => CLK, Q => n6197
                           , QN => n4306);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n2815, CK => CLK, Q => n6196
                           , QN => n4311);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n2814, CK => CLK, Q => n6195
                           , QN => n4316);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n2813, CK => CLK, Q => 
                           n6194, QN => n3777);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n2812, CK => CLK, Q => 
                           n6193, QN => n3782);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n2811, CK => CLK, Q => 
                           n6192, QN => n3787);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n2810, CK => CLK, Q => 
                           n6191, QN => n3792);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n2809, CK => CLK, Q => 
                           n6190, QN => n3797);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n2808, CK => CLK, Q => 
                           n6189, QN => n3802);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n2807, CK => CLK, Q => 
                           n6188, QN => n3807);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n2806, CK => CLK, Q => 
                           n6187, QN => n3812);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n2805, CK => CLK, Q => 
                           n6186, QN => n3817);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n2804, CK => CLK, Q => 
                           n6185, QN => n3822);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n2803, CK => CLK, Q => 
                           n6184, QN => n3827);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n2802, CK => CLK, Q => 
                           n6183, QN => n3832);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n2801, CK => CLK, Q => 
                           n6182, QN => n3837);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n2800, CK => CLK, Q => 
                           n6181, QN => n3842);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n2799, CK => CLK, Q => 
                           n6180, QN => n3847);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n2798, CK => CLK, Q => 
                           n6179, QN => n3852);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n2797, CK => CLK, Q => 
                           n6178, QN => n3857);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n2796, CK => CLK, Q => 
                           n6177, QN => n3862);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n2795, CK => CLK, Q => 
                           n6176, QN => n3867);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n2794, CK => CLK, Q => 
                           n6175, QN => n3872);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n2793, CK => CLK, Q => 
                           n6174, QN => n3877);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n2792, CK => CLK, Q => 
                           n6173, QN => n3882);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n2791, CK => CLK, Q => n6172
                           , QN => n3887);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n2790, CK => CLK, Q => n6171
                           , QN => n3892);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n2789, CK => CLK, Q => n6170
                           , QN => n3897);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n2788, CK => CLK, Q => n6169
                           , QN => n3902);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n2787, CK => CLK, Q => n6168
                           , QN => n3907);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n2786, CK => CLK, Q => n6167
                           , QN => n3912);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n2785, CK => CLK, Q => n6166
                           , QN => n3917);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n2784, CK => CLK, Q => n6165
                           , QN => n3922);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n2783, CK => CLK, Q => n6164
                           , QN => n3927);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n2782, CK => CLK, Q => n6163
                           , QN => n3932);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n2781, CK => CLK, Q => 
                           n3617, QN => n_1320);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n2780, CK => CLK, Q => 
                           n3622, QN => n_1321);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n2779, CK => CLK, Q => 
                           n3627, QN => n_1322);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n2778, CK => CLK, Q => 
                           n3632, QN => n_1323);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n2777, CK => CLK, Q => 
                           n3637, QN => n_1324);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n2776, CK => CLK, Q => 
                           n3642, QN => n_1325);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n2775, CK => CLK, Q => 
                           n3647, QN => n_1326);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n2774, CK => CLK, Q => 
                           n3652, QN => n_1327);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n2773, CK => CLK, Q => 
                           n3657, QN => n_1328);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n2772, CK => CLK, Q => 
                           n3662, QN => n_1329);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n2771, CK => CLK, Q => 
                           n3667, QN => n_1330);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n2770, CK => CLK, Q => 
                           n3672, QN => n_1331);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n2769, CK => CLK, Q => 
                           n3677, QN => n_1332);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n2768, CK => CLK, Q => 
                           n3682, QN => n_1333);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n2767, CK => CLK, Q => 
                           n3687, QN => n_1334);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n2766, CK => CLK, Q => 
                           n3692, QN => n_1335);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n2765, CK => CLK, Q => 
                           n3697, QN => n_1336);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n2764, CK => CLK, Q => 
                           n3702, QN => n_1337);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n2763, CK => CLK, Q => 
                           n3707, QN => n_1338);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n2762, CK => CLK, Q => 
                           n3712, QN => n_1339);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n2761, CK => CLK, Q => 
                           n3717, QN => n_1340);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n2760, CK => CLK, Q => 
                           n3722, QN => n_1341);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n2759, CK => CLK, Q => n3727
                           , QN => n_1342);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n2758, CK => CLK, Q => n3732
                           , QN => n_1343);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n2757, CK => CLK, Q => n3737
                           , QN => n_1344);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n2756, CK => CLK, Q => n3742
                           , QN => n_1345);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n2755, CK => CLK, Q => n3747
                           , QN => n_1346);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n2754, CK => CLK, Q => n3752
                           , QN => n_1347);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n2753, CK => CLK, Q => n3757
                           , QN => n_1348);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n2752, CK => CLK, Q => n3762
                           , QN => n_1349);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n2751, CK => CLK, Q => n3767
                           , QN => n_1350);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n2750, CK => CLK, Q => n3772
                           , QN => n_1351);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n2749, CK => CLK, Q => 
                           n4001, QN => n_1352);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n2748, CK => CLK, Q => 
                           n4006, QN => n_1353);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n2747, CK => CLK, Q => 
                           n4011, QN => n_1354);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n2746, CK => CLK, Q => 
                           n4016, QN => n_1355);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n2745, CK => CLK, Q => 
                           n4021, QN => n_1356);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n2744, CK => CLK, Q => 
                           n4026, QN => n_1357);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n2743, CK => CLK, Q => 
                           n4031, QN => n_1358);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n2742, CK => CLK, Q => 
                           n4036, QN => n_1359);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n2741, CK => CLK, Q => 
                           n4041, QN => n_1360);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n2740, CK => CLK, Q => 
                           n4046, QN => n_1361);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n2739, CK => CLK, Q => 
                           n4051, QN => n_1362);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n2738, CK => CLK, Q => 
                           n4056, QN => n_1363);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n2737, CK => CLK, Q => 
                           n4061, QN => n_1364);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n2736, CK => CLK, Q => 
                           n4066, QN => n_1365);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n2735, CK => CLK, Q => 
                           n4071, QN => n_1366);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n2734, CK => CLK, Q => 
                           n4076, QN => n_1367);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n2733, CK => CLK, Q => 
                           n4081, QN => n_1368);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n2732, CK => CLK, Q => 
                           n4086, QN => n_1369);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n2731, CK => CLK, Q => 
                           n4091, QN => n_1370);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n2730, CK => CLK, Q => 
                           n4096, QN => n_1371);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n2729, CK => CLK, Q => 
                           n4101, QN => n_1372);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n2728, CK => CLK, Q => 
                           n4106, QN => n_1373);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n2727, CK => CLK, Q => n4111
                           , QN => n_1374);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n2726, CK => CLK, Q => n4116
                           , QN => n_1375);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n2725, CK => CLK, Q => n4121
                           , QN => n_1376);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n2724, CK => CLK, Q => n4126
                           , QN => n_1377);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n2723, CK => CLK, Q => n4131
                           , QN => n_1378);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n2722, CK => CLK, Q => n4136
                           , QN => n_1379);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n2721, CK => CLK, Q => n4141
                           , QN => n_1380);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n2720, CK => CLK, Q => n4146
                           , QN => n_1381);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n2719, CK => CLK, Q => n4151
                           , QN => n_1382);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n2718, CK => CLK, Q => n4156
                           , QN => n_1383);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n2717, CK => CLK, Q => 
                           n6162, QN => n4162);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n2716, CK => CLK, Q => 
                           n6161, QN => n4167);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n2715, CK => CLK, Q => 
                           n6160, QN => n4172);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n2714, CK => CLK, Q => 
                           n6159, QN => n4177);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n2713, CK => CLK, Q => 
                           n6158, QN => n4182);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n2712, CK => CLK, Q => 
                           n6157, QN => n4187);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n2711, CK => CLK, Q => 
                           n6156, QN => n4192);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n2710, CK => CLK, Q => 
                           n6155, QN => n4197);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n2709, CK => CLK, Q => 
                           n6154, QN => n4202);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n2708, CK => CLK, Q => 
                           n6153, QN => n4207);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n2707, CK => CLK, Q => 
                           n6152, QN => n4212);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n2706, CK => CLK, Q => 
                           n6151, QN => n4217);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n2705, CK => CLK, Q => 
                           n6150, QN => n4222);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n2704, CK => CLK, Q => 
                           n6149, QN => n4227);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n2703, CK => CLK, Q => 
                           n6148, QN => n4232);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n2702, CK => CLK, Q => 
                           n6147, QN => n4237);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n2701, CK => CLK, Q => 
                           n6146, QN => n4242);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n2700, CK => CLK, Q => 
                           n6145, QN => n4247);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n2699, CK => CLK, Q => 
                           n6144, QN => n4252);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n2698, CK => CLK, Q => 
                           n6143, QN => n4257);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n2697, CK => CLK, Q => 
                           n6142, QN => n4262);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n2696, CK => CLK, Q => 
                           n6141, QN => n4267);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n2695, CK => CLK, Q => n6140
                           , QN => n4272);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n2694, CK => CLK, Q => n6139
                           , QN => n4277);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n2693, CK => CLK, Q => n6138
                           , QN => n4282);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n2692, CK => CLK, Q => n6137
                           , QN => n4287);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n2691, CK => CLK, Q => n6136
                           , QN => n4292);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n2690, CK => CLK, Q => n6135
                           , QN => n4297);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n2689, CK => CLK, Q => n6134
                           , QN => n4302);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n2688, CK => CLK, Q => n6133
                           , QN => n4307);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n2687, CK => CLK, Q => n6132
                           , QN => n4312);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n2686, CK => CLK, Q => n6131
                           , QN => n4317);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n2685, CK => CLK, Q => 
                           n6130, QN => n3778);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n2684, CK => CLK, Q => 
                           n6129, QN => n3783);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n2683, CK => CLK, Q => 
                           n6128, QN => n3788);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n2682, CK => CLK, Q => 
                           n6127, QN => n3793);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n2681, CK => CLK, Q => 
                           n6126, QN => n3798);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n2680, CK => CLK, Q => 
                           n6125, QN => n3803);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n2679, CK => CLK, Q => 
                           n6124, QN => n3808);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n2678, CK => CLK, Q => 
                           n6123, QN => n3813);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n2677, CK => CLK, Q => 
                           n6122, QN => n3818);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n2676, CK => CLK, Q => 
                           n6121, QN => n3823);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n2675, CK => CLK, Q => 
                           n6120, QN => n3828);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n2674, CK => CLK, Q => 
                           n6119, QN => n3833);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n2673, CK => CLK, Q => 
                           n6118, QN => n3838);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n2672, CK => CLK, Q => 
                           n6117, QN => n3843);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n2671, CK => CLK, Q => 
                           n6116, QN => n3848);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n2670, CK => CLK, Q => 
                           n6115, QN => n3853);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n2669, CK => CLK, Q => 
                           n6114, QN => n3858);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n2668, CK => CLK, Q => 
                           n6113, QN => n3863);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n2667, CK => CLK, Q => 
                           n6112, QN => n3868);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n2666, CK => CLK, Q => 
                           n6111, QN => n3873);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n2665, CK => CLK, Q => 
                           n6110, QN => n3878);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n2664, CK => CLK, Q => 
                           n6109, QN => n3883);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n2663, CK => CLK, Q => n6108
                           , QN => n3888);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n2662, CK => CLK, Q => n6107
                           , QN => n3893);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n2661, CK => CLK, Q => n6106
                           , QN => n3898);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n2660, CK => CLK, Q => n6105
                           , QN => n3903);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n2659, CK => CLK, Q => n6104
                           , QN => n3908);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n2658, CK => CLK, Q => n6103
                           , QN => n3913);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n2657, CK => CLK, Q => n6102
                           , QN => n3918);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n2656, CK => CLK, Q => n6101
                           , QN => n3923);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n2655, CK => CLK, Q => n6100
                           , QN => n3928);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n2654, CK => CLK, Q => n6099
                           , QN => n3933);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n2653, CK => CLK, Q => 
                           n3618, QN => n_1384);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n2652, CK => CLK, Q => 
                           n3623, QN => n_1385);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n2651, CK => CLK, Q => 
                           n3628, QN => n_1386);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n2650, CK => CLK, Q => 
                           n3633, QN => n_1387);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n2649, CK => CLK, Q => 
                           n3638, QN => n_1388);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n2648, CK => CLK, Q => 
                           n3643, QN => n_1389);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n2647, CK => CLK, Q => 
                           n3648, QN => n_1390);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n2646, CK => CLK, Q => 
                           n3653, QN => n_1391);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n2645, CK => CLK, Q => 
                           n3658, QN => n_1392);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n2644, CK => CLK, Q => 
                           n3663, QN => n_1393);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n2643, CK => CLK, Q => 
                           n3668, QN => n_1394);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n2642, CK => CLK, Q => 
                           n3673, QN => n_1395);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n2641, CK => CLK, Q => 
                           n3678, QN => n_1396);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n2640, CK => CLK, Q => 
                           n3683, QN => n_1397);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n2639, CK => CLK, Q => 
                           n3688, QN => n_1398);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n2638, CK => CLK, Q => 
                           n3693, QN => n_1399);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n2637, CK => CLK, Q => 
                           n3698, QN => n_1400);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n2636, CK => CLK, Q => 
                           n3703, QN => n_1401);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n2635, CK => CLK, Q => 
                           n3708, QN => n_1402);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n2634, CK => CLK, Q => 
                           n3713, QN => n_1403);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n2633, CK => CLK, Q => 
                           n3718, QN => n_1404);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n2632, CK => CLK, Q => 
                           n3723, QN => n_1405);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n2631, CK => CLK, Q => n3728
                           , QN => n_1406);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n2630, CK => CLK, Q => n3733
                           , QN => n_1407);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n2629, CK => CLK, Q => n3738
                           , QN => n_1408);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n2628, CK => CLK, Q => n3743
                           , QN => n_1409);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n2627, CK => CLK, Q => n3748
                           , QN => n_1410);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n2626, CK => CLK, Q => n3753
                           , QN => n_1411);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n2625, CK => CLK, Q => n3758
                           , QN => n_1412);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n2624, CK => CLK, Q => n3763
                           , QN => n_1413);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n2623, CK => CLK, Q => n3768
                           , QN => n_1414);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n2622, CK => CLK, Q => n3773
                           , QN => n_1415);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n2621, CK => CLK, Q => 
                           n4002, QN => n_1416);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n2620, CK => CLK, Q => 
                           n4007, QN => n_1417);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n2619, CK => CLK, Q => 
                           n4012, QN => n_1418);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n2618, CK => CLK, Q => 
                           n4017, QN => n_1419);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n2617, CK => CLK, Q => 
                           n4022, QN => n_1420);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n2616, CK => CLK, Q => 
                           n4027, QN => n_1421);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n2615, CK => CLK, Q => 
                           n4032, QN => n_1422);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n2614, CK => CLK, Q => 
                           n4037, QN => n_1423);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n2613, CK => CLK, Q => 
                           n4042, QN => n_1424);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n2612, CK => CLK, Q => 
                           n4047, QN => n_1425);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n2611, CK => CLK, Q => 
                           n4052, QN => n_1426);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n2610, CK => CLK, Q => 
                           n4057, QN => n_1427);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n2609, CK => CLK, Q => 
                           n4062, QN => n_1428);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n2608, CK => CLK, Q => 
                           n4067, QN => n_1429);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n2607, CK => CLK, Q => 
                           n4072, QN => n_1430);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n2606, CK => CLK, Q => 
                           n4077, QN => n_1431);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n2605, CK => CLK, Q => 
                           n4082, QN => n_1432);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n2604, CK => CLK, Q => 
                           n4087, QN => n_1433);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n2603, CK => CLK, Q => 
                           n4092, QN => n_1434);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n2602, CK => CLK, Q => 
                           n4097, QN => n_1435);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n2601, CK => CLK, Q => 
                           n4102, QN => n_1436);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n2600, CK => CLK, Q => 
                           n4107, QN => n_1437);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n2599, CK => CLK, Q => n4112
                           , QN => n_1438);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n2598, CK => CLK, Q => n4117
                           , QN => n_1439);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n2597, CK => CLK, Q => n4122
                           , QN => n_1440);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n2596, CK => CLK, Q => n4127
                           , QN => n_1441);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n2595, CK => CLK, Q => n4132
                           , QN => n_1442);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n2594, CK => CLK, Q => n4137
                           , QN => n_1443);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n2593, CK => CLK, Q => n4142
                           , QN => n_1444);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n2592, CK => CLK, Q => n4147
                           , QN => n_1445);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n2591, CK => CLK, Q => n4152
                           , QN => n_1446);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n2590, CK => CLK, Q => n4157
                           , QN => n_1447);
   OUT2_reg_31_inst : DFF_X1 port map( D => n2589, CK => CLK, Q => OUT2_31_port
                           , QN => n_1448);
   OUT2_reg_30_inst : DFF_X1 port map( D => n2588, CK => CLK, Q => OUT2_30_port
                           , QN => n_1449);
   OUT2_reg_29_inst : DFF_X1 port map( D => n2587, CK => CLK, Q => OUT2_29_port
                           , QN => n_1450);
   OUT2_reg_28_inst : DFF_X1 port map( D => n2586, CK => CLK, Q => OUT2_28_port
                           , QN => n_1451);
   OUT2_reg_27_inst : DFF_X1 port map( D => n2585, CK => CLK, Q => OUT2_27_port
                           , QN => n_1452);
   OUT2_reg_26_inst : DFF_X1 port map( D => n2584, CK => CLK, Q => OUT2_26_port
                           , QN => n_1453);
   OUT2_reg_25_inst : DFF_X1 port map( D => n2583, CK => CLK, Q => OUT2_25_port
                           , QN => n_1454);
   OUT2_reg_24_inst : DFF_X1 port map( D => n2582, CK => CLK, Q => OUT2_24_port
                           , QN => n_1455);
   OUT2_reg_23_inst : DFF_X1 port map( D => n2581, CK => CLK, Q => OUT2_23_port
                           , QN => n_1456);
   OUT2_reg_22_inst : DFF_X1 port map( D => n2580, CK => CLK, Q => OUT2_22_port
                           , QN => n_1457);
   OUT2_reg_21_inst : DFF_X1 port map( D => n2579, CK => CLK, Q => OUT2_21_port
                           , QN => n_1458);
   OUT2_reg_20_inst : DFF_X1 port map( D => n2578, CK => CLK, Q => OUT2_20_port
                           , QN => n_1459);
   OUT2_reg_19_inst : DFF_X1 port map( D => n2577, CK => CLK, Q => OUT2_19_port
                           , QN => n_1460);
   OUT2_reg_18_inst : DFF_X1 port map( D => n2576, CK => CLK, Q => OUT2_18_port
                           , QN => n_1461);
   OUT2_reg_17_inst : DFF_X1 port map( D => n2575, CK => CLK, Q => OUT2_17_port
                           , QN => n_1462);
   OUT2_reg_16_inst : DFF_X1 port map( D => n2574, CK => CLK, Q => OUT2_16_port
                           , QN => n_1463);
   OUT2_reg_15_inst : DFF_X1 port map( D => n2573, CK => CLK, Q => OUT2_15_port
                           , QN => n_1464);
   OUT2_reg_14_inst : DFF_X1 port map( D => n2572, CK => CLK, Q => OUT2_14_port
                           , QN => n_1465);
   OUT2_reg_13_inst : DFF_X1 port map( D => n2571, CK => CLK, Q => OUT2_13_port
                           , QN => n_1466);
   OUT2_reg_12_inst : DFF_X1 port map( D => n2570, CK => CLK, Q => OUT2_12_port
                           , QN => n_1467);
   OUT2_reg_11_inst : DFF_X1 port map( D => n2569, CK => CLK, Q => OUT2_11_port
                           , QN => n_1468);
   OUT2_reg_10_inst : DFF_X1 port map( D => n2568, CK => CLK, Q => OUT2_10_port
                           , QN => n_1469);
   OUT2_reg_9_inst : DFF_X1 port map( D => n2567, CK => CLK, Q => OUT2_9_port, 
                           QN => n_1470);
   OUT2_reg_8_inst : DFF_X1 port map( D => n2566, CK => CLK, Q => OUT2_8_port, 
                           QN => n_1471);
   OUT2_reg_7_inst : DFF_X1 port map( D => n2565, CK => CLK, Q => OUT2_7_port, 
                           QN => n_1472);
   OUT2_reg_6_inst : DFF_X1 port map( D => n2564, CK => CLK, Q => OUT2_6_port, 
                           QN => n_1473);
   OUT2_reg_5_inst : DFF_X1 port map( D => n2563, CK => CLK, Q => OUT2_5_port, 
                           QN => n_1474);
   OUT2_reg_4_inst : DFF_X1 port map( D => n2562, CK => CLK, Q => OUT2_4_port, 
                           QN => n_1475);
   OUT2_reg_3_inst : DFF_X1 port map( D => n2561, CK => CLK, Q => OUT2_3_port, 
                           QN => n_1476);
   OUT2_reg_2_inst : DFF_X1 port map( D => n2560, CK => CLK, Q => OUT2_2_port, 
                           QN => n_1477);
   OUT2_reg_1_inst : DFF_X1 port map( D => n2559, CK => CLK, Q => OUT2_1_port, 
                           QN => n_1478);
   OUT2_reg_0_inst : DFF_X1 port map( D => n2558, CK => CLK, Q => OUT2_0_port, 
                           QN => n_1479);
   OUT1_reg_31_inst : DFF_X1 port map( D => n2557, CK => CLK, Q => OUT1_31_port
                           , QN => n_1480);
   OUT1_reg_30_inst : DFF_X1 port map( D => n2556, CK => CLK, Q => OUT1_30_port
                           , QN => n_1481);
   OUT1_reg_29_inst : DFF_X1 port map( D => n2555, CK => CLK, Q => OUT1_29_port
                           , QN => n_1482);
   OUT1_reg_28_inst : DFF_X1 port map( D => n2554, CK => CLK, Q => OUT1_28_port
                           , QN => n_1483);
   OUT1_reg_27_inst : DFF_X1 port map( D => n2553, CK => CLK, Q => OUT1_27_port
                           , QN => n_1484);
   OUT1_reg_26_inst : DFF_X1 port map( D => n2552, CK => CLK, Q => OUT1_26_port
                           , QN => n_1485);
   OUT1_reg_25_inst : DFF_X1 port map( D => n2551, CK => CLK, Q => OUT1_25_port
                           , QN => n_1486);
   OUT1_reg_24_inst : DFF_X1 port map( D => n2550, CK => CLK, Q => OUT1_24_port
                           , QN => n_1487);
   OUT1_reg_23_inst : DFF_X1 port map( D => n2549, CK => CLK, Q => OUT1_23_port
                           , QN => n_1488);
   OUT1_reg_22_inst : DFF_X1 port map( D => n2548, CK => CLK, Q => OUT1_22_port
                           , QN => n_1489);
   OUT1_reg_21_inst : DFF_X1 port map( D => n2547, CK => CLK, Q => OUT1_21_port
                           , QN => n_1490);
   OUT1_reg_20_inst : DFF_X1 port map( D => n2546, CK => CLK, Q => OUT1_20_port
                           , QN => n_1491);
   OUT1_reg_19_inst : DFF_X1 port map( D => n2545, CK => CLK, Q => OUT1_19_port
                           , QN => n_1492);
   OUT1_reg_18_inst : DFF_X1 port map( D => n2544, CK => CLK, Q => OUT1_18_port
                           , QN => n_1493);
   OUT1_reg_17_inst : DFF_X1 port map( D => n2543, CK => CLK, Q => OUT1_17_port
                           , QN => n_1494);
   OUT1_reg_16_inst : DFF_X1 port map( D => n2542, CK => CLK, Q => OUT1_16_port
                           , QN => n_1495);
   OUT1_reg_15_inst : DFF_X1 port map( D => n2541, CK => CLK, Q => OUT1_15_port
                           , QN => n_1496);
   OUT1_reg_14_inst : DFF_X1 port map( D => n2540, CK => CLK, Q => OUT1_14_port
                           , QN => n_1497);
   OUT1_reg_13_inst : DFF_X1 port map( D => n2539, CK => CLK, Q => OUT1_13_port
                           , QN => n_1498);
   OUT1_reg_12_inst : DFF_X1 port map( D => n2538, CK => CLK, Q => OUT1_12_port
                           , QN => n_1499);
   OUT1_reg_11_inst : DFF_X1 port map( D => n2537, CK => CLK, Q => OUT1_11_port
                           , QN => n_1500);
   OUT1_reg_10_inst : DFF_X1 port map( D => n2536, CK => CLK, Q => OUT1_10_port
                           , QN => n_1501);
   OUT1_reg_9_inst : DFF_X1 port map( D => n2535, CK => CLK, Q => OUT1_9_port, 
                           QN => n_1502);
   OUT1_reg_8_inst : DFF_X1 port map( D => n2534, CK => CLK, Q => OUT1_8_port, 
                           QN => n_1503);
   OUT1_reg_7_inst : DFF_X1 port map( D => n2533, CK => CLK, Q => OUT1_7_port, 
                           QN => n_1504);
   OUT1_reg_6_inst : DFF_X1 port map( D => n2532, CK => CLK, Q => OUT1_6_port, 
                           QN => n_1505);
   OUT1_reg_5_inst : DFF_X1 port map( D => n2531, CK => CLK, Q => OUT1_5_port, 
                           QN => n_1506);
   OUT1_reg_4_inst : DFF_X1 port map( D => n2530, CK => CLK, Q => OUT1_4_port, 
                           QN => n_1507);
   OUT1_reg_3_inst : DFF_X1 port map( D => n2529, CK => CLK, Q => OUT1_3_port, 
                           QN => n_1508);
   OUT1_reg_2_inst : DFF_X1 port map( D => n2528, CK => CLK, Q => OUT1_2_port, 
                           QN => n_1509);
   OUT1_reg_1_inst : DFF_X1 port map( D => n2527, CK => CLK, Q => OUT1_1_port, 
                           QN => n_1510);
   OUT1_reg_0_inst : DFF_X1 port map( D => n2526, CK => CLK, Q => OUT1_0_port, 
                           QN => n_1511);
   U2528 : AND3_X2 port map( A1 => ENABLE, A2 => n4607, A3 => RD2, ZN => n4656)
                           ;
   U2529 : AND3_X2 port map( A1 => ENABLE, A2 => n4607, A3 => RD1, ZN => n5314)
                           ;
   U2530 : INV_X1 port map( A => n4642, ZN => n4510);
   U2531 : INV_X2 port map( A => n4510, ZN => n4511);
   U2532 : INV_X1 port map( A => n4643, ZN => n4512);
   U2533 : INV_X2 port map( A => n4512, ZN => n4513);
   U2534 : INV_X1 port map( A => n4648, ZN => n4514);
   U2535 : INV_X2 port map( A => n4514, ZN => n4515);
   U2536 : INV_X1 port map( A => n4649, ZN => n4516);
   U2537 : INV_X2 port map( A => n4516, ZN => n4517);
   U2538 : INV_X1 port map( A => n4650, ZN => n4518);
   U2539 : INV_X2 port map( A => n4518, ZN => n4519);
   U2540 : INV_X1 port map( A => n4651, ZN => n4520);
   U2541 : INV_X2 port map( A => n4520, ZN => n4521);
   U2542 : INV_X1 port map( A => n4652, ZN => n4522);
   U2543 : INV_X2 port map( A => n4522, ZN => n4523);
   U2544 : INV_X1 port map( A => n4653, ZN => n4524);
   U2545 : INV_X2 port map( A => n4524, ZN => n4525);
   U2546 : INV_X1 port map( A => n4654, ZN => n4526);
   U2547 : INV_X2 port map( A => n4526, ZN => n4527);
   U2548 : INV_X1 port map( A => n4640, ZN => n4528);
   U2549 : INV_X2 port map( A => n4528, ZN => n4529);
   U2550 : INV_X1 port map( A => n4641, ZN => n4530);
   U2551 : INV_X2 port map( A => n4530, ZN => n4531);
   U2552 : INV_X1 port map( A => n4638, ZN => n4532);
   U2553 : INV_X2 port map( A => n4532, ZN => n4533);
   U2554 : INV_X1 port map( A => n4639, ZN => n4534);
   U2555 : INV_X2 port map( A => n4534, ZN => n4535);
   U2556 : INV_X1 port map( A => n4636, ZN => n4536);
   U2557 : INV_X2 port map( A => n4536, ZN => n4537);
   U2558 : INV_X1 port map( A => n4637, ZN => n4538);
   U2559 : INV_X2 port map( A => n4538, ZN => n4539);
   U2560 : INV_X1 port map( A => n4633, ZN => n4540);
   U2561 : INV_X2 port map( A => n4540, ZN => n4541);
   U2562 : INV_X1 port map( A => n4634, ZN => n4542);
   U2563 : INV_X2 port map( A => n4542, ZN => n4543);
   U2564 : INV_X1 port map( A => n4631, ZN => n4544);
   U2565 : INV_X2 port map( A => n4544, ZN => n4545);
   U2566 : INV_X1 port map( A => n4632, ZN => n4546);
   U2567 : INV_X2 port map( A => n4546, ZN => n4547);
   U2568 : INV_X1 port map( A => n4629, ZN => n4548);
   U2569 : INV_X2 port map( A => n4548, ZN => n4549);
   U2570 : INV_X1 port map( A => n4630, ZN => n4550);
   U2571 : INV_X2 port map( A => n4550, ZN => n4551);
   U2572 : INV_X1 port map( A => n4627, ZN => n4552);
   U2573 : INV_X2 port map( A => n4552, ZN => n4553);
   U2574 : INV_X1 port map( A => n4628, ZN => n4554);
   U2575 : INV_X2 port map( A => n4554, ZN => n4555);
   U2576 : INV_X1 port map( A => n4620, ZN => n4556);
   U2577 : INV_X2 port map( A => n4556, ZN => n4557);
   U2578 : INV_X1 port map( A => n4625, ZN => n4558);
   U2579 : INV_X2 port map( A => n4558, ZN => n4559);
   U2580 : INV_X1 port map( A => n4616, ZN => n4560);
   U2581 : INV_X2 port map( A => n4560, ZN => n4561);
   U2582 : INV_X1 port map( A => n4618, ZN => n4562);
   U2583 : INV_X2 port map( A => n4562, ZN => n4563);
   U2584 : INV_X1 port map( A => n4612, ZN => n4564);
   U2585 : INV_X2 port map( A => n4564, ZN => n4565);
   U2586 : INV_X1 port map( A => n4614, ZN => n4566);
   U2587 : INV_X2 port map( A => n4566, ZN => n4567);
   U2588 : INV_X1 port map( A => n4608, ZN => n4568);
   U2589 : INV_X2 port map( A => n4568, ZN => n4569);
   U2590 : INV_X1 port map( A => n4610, ZN => n4570);
   U2591 : INV_X2 port map( A => n4570, ZN => n4571);
   U2592 : OAI21_X4 port map( B1 => n4605, B2 => n4606, A => n4607, ZN => n4573
                           );
   U2593 : INV_X4 port map( A => RESET, ZN => n4607);
   U2594 : AND2_X2 port map( A1 => n5961, A2 => n5946, ZN => n5349);
   U2595 : NOR2_X2 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), ZN => n5946);
   U2596 : AND2_X2 port map( A1 => n5285, A2 => n5290, ZN => n4672);
   U2597 : AND2_X2 port map( A1 => n5288, A2 => n5294, ZN => n4677);
   U2598 : AND2_X2 port map( A1 => n5943, A2 => n5948, ZN => n5330);
   U2599 : AND2_X2 port map( A1 => n5944, A2 => n5952, ZN => n5335);
   U2600 : AND2_X2 port map( A1 => n5303, A2 => n5291, ZN => n4696);
   U2601 : AND2_X2 port map( A1 => n5308, A2 => n5286, ZN => n4701);
   U2602 : AND2_X2 port map( A1 => n5961, A2 => n5949, ZN => n5354);
   U2603 : AND2_X2 port map( A1 => n5285, A2 => n5286, ZN => n4667);
   U2604 : AND2_X2 port map( A1 => n5943, A2 => n5944, ZN => n5325);
   U2605 : AND2_X2 port map( A1 => n5303, A2 => n5288, ZN => n4691);
   U2606 : AND2_X2 port map( A1 => n5308, A2 => n5290, ZN => n4706);
   U2607 : AND2_X2 port map( A1 => n5291, A2 => n5294, ZN => n4682);
   U2608 : AND2_X2 port map( A1 => n5966, A2 => n5948, ZN => n5364);
   U2609 : AND2_X2 port map( A1 => n5949, A2 => n5952, ZN => n5340);
   U2610 : NAND2_X2 port map( A1 => n5946, A2 => n5953, ZN => n5332);
   U2611 : AND2_X2 port map( A1 => n5966, A2 => n5944, ZN => n5359);
   U2612 : NAND2_X2 port map( A1 => n5287, A2 => n5291, ZN => n4669);
   U2613 : NAND2_X2 port map( A1 => n5286, A2 => n5295, ZN => n4674);
   U2614 : NAND2_X2 port map( A1 => n5945, A2 => n5949, ZN => n5327);
   U2615 : NAND2_X2 port map( A1 => n5304, A2 => n5290, ZN => n4693);
   U2616 : NAND2_X2 port map( A1 => n5309, A2 => n5288, ZN => n4698);
   U2617 : NAND2_X2 port map( A1 => n5962, A2 => n5948, ZN => n5351);
   U2618 : NAND2_X2 port map( A1 => n5967, A2 => n5946, ZN => n5356);
   U2619 : NAND2_X2 port map( A1 => n5287, A2 => n5288, ZN => n4664);
   U2620 : NAND2_X2 port map( A1 => n5945, A2 => n5946, ZN => n5322);
   U2621 : NAND2_X2 port map( A1 => n5304, A2 => n5286, ZN => n4688);
   U2622 : NAND2_X2 port map( A1 => n5309, A2 => n5291, ZN => n4703);
   U2623 : NAND2_X2 port map( A1 => n5295, A2 => n5290, ZN => n4679);
   U2624 : NAND2_X2 port map( A1 => n5967, A2 => n5949, ZN => n5361);
   U2625 : NAND2_X2 port map( A1 => n5953, A2 => n5948, ZN => n5337);
   U2626 : NAND2_X2 port map( A1 => n5961, A2 => n5944, ZN => n5345);
   U2627 : NAND2_X2 port map( A1 => n5962, A2 => n5944, ZN => n5346);
   U2628 : NAND2_X2 port map( A1 => n5285, A2 => n5291, ZN => n4668);
   U2629 : NAND2_X2 port map( A1 => n5286, A2 => n5294, ZN => n4673);
   U2630 : NAND2_X2 port map( A1 => n5943, A2 => n5949, ZN => n5326);
   U2631 : NAND2_X2 port map( A1 => n5946, A2 => n5952, ZN => n5331);
   U2632 : NAND2_X2 port map( A1 => n5303, A2 => n5290, ZN => n4692);
   U2633 : NAND2_X2 port map( A1 => n5308, A2 => n5288, ZN => n4697);
   U2634 : NAND2_X2 port map( A1 => n5961, A2 => n5948, ZN => n5350);
   U2635 : NAND2_X2 port map( A1 => n5285, A2 => n5288, ZN => n4663);
   U2636 : NAND2_X2 port map( A1 => n5943, A2 => n5946, ZN => n5321);
   U2637 : NAND2_X2 port map( A1 => n5303, A2 => n5286, ZN => n4687);
   U2638 : NAND2_X2 port map( A1 => n5308, A2 => n5291, ZN => n4702);
   U2639 : NAND2_X2 port map( A1 => n5290, A2 => n5294, ZN => n4678);
   U2640 : NAND2_X2 port map( A1 => n5966, A2 => n5949, ZN => n5360);
   U2641 : NAND2_X2 port map( A1 => n5948, A2 => n5952, ZN => n5336);
   U2642 : AND2_X2 port map( A1 => n5944, A2 => n5953, ZN => n5334);
   U2643 : NAND2_X2 port map( A1 => n5966, A2 => n5946, ZN => n5355);
   U2644 : AND2_X2 port map( A1 => n5287, A2 => n5290, ZN => n4671);
   U2645 : AND2_X2 port map( A1 => n5288, A2 => n5295, ZN => n4676);
   U2646 : AND2_X2 port map( A1 => n5945, A2 => n5948, ZN => n5329);
   U2647 : AND2_X2 port map( A1 => n5304, A2 => n5291, ZN => n4695);
   U2648 : AND2_X2 port map( A1 => n5309, A2 => n5286, ZN => n4700);
   U2649 : AND2_X2 port map( A1 => n5962, A2 => n5949, ZN => n5353);
   U2650 : AND2_X2 port map( A1 => n5967, A2 => n5944, ZN => n5358);
   U2651 : AND2_X2 port map( A1 => n5287, A2 => n5286, ZN => n4666);
   U2652 : AND2_X2 port map( A1 => n5945, A2 => n5944, ZN => n5324);
   U2653 : AND2_X2 port map( A1 => n5304, A2 => n5288, ZN => n4690);
   U2654 : AND2_X2 port map( A1 => n5309, A2 => n5290, ZN => n4705);
   U2655 : AND2_X2 port map( A1 => n5291, A2 => n5295, ZN => n4681);
   U2656 : AND2_X2 port map( A1 => n5962, A2 => n5946, ZN => n5348);
   U2657 : AND2_X2 port map( A1 => n5967, A2 => n5948, ZN => n5363);
   U2658 : AND2_X2 port map( A1 => n5949, A2 => n5953, ZN => n5339);
   U2659 : MUX2_X1 port map( A => n4382, B => n4572, S => n4573, Z => n3613);
   U2660 : MUX2_X1 port map( A => n4383, B => n4574, S => n4573, Z => n3612);
   U2661 : MUX2_X1 port map( A => n4384, B => n4575, S => n4573, Z => n3611);
   U2662 : MUX2_X1 port map( A => n4385, B => n4576, S => n4573, Z => n3610);
   U2663 : MUX2_X1 port map( A => n4386, B => n4577, S => n4573, Z => n3609);
   U2664 : MUX2_X1 port map( A => n4387, B => n4578, S => n4573, Z => n3608);
   U2665 : MUX2_X1 port map( A => n4388, B => n4579, S => n4573, Z => n3607);
   U2666 : MUX2_X1 port map( A => n4389, B => n4580, S => n4573, Z => n3606);
   U2667 : MUX2_X1 port map( A => n4390, B => n4581, S => n4573, Z => n3605);
   U2668 : MUX2_X1 port map( A => n4391, B => n4582, S => n4573, Z => n3604);
   U2669 : MUX2_X1 port map( A => n4392, B => n4583, S => n4573, Z => n3603);
   U2670 : MUX2_X1 port map( A => n4393, B => n4584, S => n4573, Z => n3602);
   U2671 : MUX2_X1 port map( A => n4394, B => n4585, S => n4573, Z => n3601);
   U2672 : MUX2_X1 port map( A => n4395, B => n4586, S => n4573, Z => n3600);
   U2673 : MUX2_X1 port map( A => n4396, B => n4587, S => n4573, Z => n3599);
   U2674 : MUX2_X1 port map( A => n4397, B => n4588, S => n4573, Z => n3598);
   U2675 : MUX2_X1 port map( A => n4398, B => n4589, S => n4573, Z => n3597);
   U2676 : MUX2_X1 port map( A => n4399, B => n4590, S => n4573, Z => n3596);
   U2677 : MUX2_X1 port map( A => n4400, B => n4591, S => n4573, Z => n3595);
   U2678 : MUX2_X1 port map( A => n4401, B => n4592, S => n4573, Z => n3594);
   U2679 : MUX2_X1 port map( A => n4402, B => n4593, S => n4573, Z => n3593);
   U2680 : MUX2_X1 port map( A => n4403, B => n4594, S => n4573, Z => n3592);
   U2681 : MUX2_X1 port map( A => n4404, B => n4595, S => n4573, Z => n3591);
   U2682 : MUX2_X1 port map( A => n4405, B => n4596, S => n4573, Z => n3590);
   U2683 : MUX2_X1 port map( A => n4406, B => n4597, S => n4573, Z => n3589);
   U2684 : MUX2_X1 port map( A => n4407, B => n4598, S => n4573, Z => n3588);
   U2685 : MUX2_X1 port map( A => n4408, B => n4599, S => n4573, Z => n3587);
   U2686 : MUX2_X1 port map( A => n4409, B => n4600, S => n4573, Z => n3586);
   U2687 : MUX2_X1 port map( A => n4410, B => n4601, S => n4573, Z => n3585);
   U2688 : MUX2_X1 port map( A => n4411, B => n4602, S => n4573, Z => n3584);
   U2689 : MUX2_X1 port map( A => n4412, B => n4603, S => n4573, Z => n3583);
   U2690 : MUX2_X1 port map( A => n4413, B => n4604, S => n4573, Z => n3582);
   U2691 : MUX2_X1 port map( A => n4446, B => n4572, S => n4569, Z => n3581);
   U2692 : MUX2_X1 port map( A => n4447, B => n4574, S => n4569, Z => n3580);
   U2693 : MUX2_X1 port map( A => n4448, B => n4575, S => n4569, Z => n3579);
   U2694 : MUX2_X1 port map( A => n4449, B => n4576, S => n4569, Z => n3578);
   U2695 : MUX2_X1 port map( A => n4450, B => n4577, S => n4569, Z => n3577);
   U2696 : MUX2_X1 port map( A => n4451, B => n4578, S => n4569, Z => n3576);
   U2697 : MUX2_X1 port map( A => n4452, B => n4579, S => n4569, Z => n3575);
   U2698 : MUX2_X1 port map( A => n4453, B => n4580, S => n4569, Z => n3574);
   U2699 : MUX2_X1 port map( A => n4454, B => n4581, S => n4569, Z => n3573);
   U2700 : MUX2_X1 port map( A => n4455, B => n4582, S => n4569, Z => n3572);
   U2701 : MUX2_X1 port map( A => n4456, B => n4583, S => n4569, Z => n3571);
   U2702 : MUX2_X1 port map( A => n4457, B => n4584, S => n4569, Z => n3570);
   U2703 : MUX2_X1 port map( A => n4458, B => n4585, S => n4569, Z => n3569);
   U2704 : MUX2_X1 port map( A => n4459, B => n4586, S => n4569, Z => n3568);
   U2705 : MUX2_X1 port map( A => n4460, B => n4587, S => n4569, Z => n3567);
   U2706 : MUX2_X1 port map( A => n4461, B => n4588, S => n4569, Z => n3566);
   U2707 : MUX2_X1 port map( A => n4462, B => n4589, S => n4569, Z => n3565);
   U2708 : MUX2_X1 port map( A => n4463, B => n4590, S => n4569, Z => n3564);
   U2709 : MUX2_X1 port map( A => n4464, B => n4591, S => n4569, Z => n3563);
   U2710 : MUX2_X1 port map( A => n4465, B => n4592, S => n4569, Z => n3562);
   U2711 : MUX2_X1 port map( A => n4466, B => n4593, S => n4569, Z => n3561);
   U2712 : MUX2_X1 port map( A => n4467, B => n4594, S => n4569, Z => n3560);
   U2713 : MUX2_X1 port map( A => n4468, B => n4595, S => n4569, Z => n3559);
   U2714 : MUX2_X1 port map( A => n4469, B => n4596, S => n4569, Z => n3558);
   U2715 : MUX2_X1 port map( A => n4470, B => n4597, S => n4569, Z => n3557);
   U2716 : MUX2_X1 port map( A => n4471, B => n4598, S => n4569, Z => n3556);
   U2717 : MUX2_X1 port map( A => n4472, B => n4599, S => n4569, Z => n3555);
   U2718 : MUX2_X1 port map( A => n4473, B => n4600, S => n4569, Z => n3554);
   U2719 : MUX2_X1 port map( A => n4474, B => n4601, S => n4569, Z => n3553);
   U2720 : MUX2_X1 port map( A => n4475, B => n4602, S => n4569, Z => n3552);
   U2721 : MUX2_X1 port map( A => n4476, B => n4603, S => n4569, Z => n3551);
   U2722 : MUX2_X1 port map( A => n4477, B => n4604, S => n4569, Z => n3550);
   U2723 : OAI21_X1 port map( B1 => n4605, B2 => n4609, A => n4607, ZN => n4608
                           );
   U2724 : MUX2_X1 port map( A => n6098, B => n4572, S => n4571, Z => n3549);
   U2725 : MUX2_X1 port map( A => n6094, B => n4574, S => n4571, Z => n3548);
   U2726 : MUX2_X1 port map( A => n6090, B => n4575, S => n4571, Z => n3547);
   U2727 : MUX2_X1 port map( A => n6086, B => n4576, S => n4571, Z => n3546);
   U2728 : MUX2_X1 port map( A => n6082, B => n4577, S => n4571, Z => n3545);
   U2729 : MUX2_X1 port map( A => n6078, B => n4578, S => n4571, Z => n3544);
   U2730 : MUX2_X1 port map( A => n6074, B => n4579, S => n4571, Z => n3543);
   U2731 : MUX2_X1 port map( A => n6070, B => n4580, S => n4571, Z => n3542);
   U2732 : MUX2_X1 port map( A => n6066, B => n4581, S => n4571, Z => n3541);
   U2733 : MUX2_X1 port map( A => n6062, B => n4582, S => n4571, Z => n3540);
   U2734 : MUX2_X1 port map( A => n6058, B => n4583, S => n4571, Z => n3539);
   U2735 : MUX2_X1 port map( A => n6054, B => n4584, S => n4571, Z => n3538);
   U2736 : MUX2_X1 port map( A => n6050, B => n4585, S => n4571, Z => n3537);
   U2737 : MUX2_X1 port map( A => n6046, B => n4586, S => n4571, Z => n3536);
   U2738 : MUX2_X1 port map( A => n6042, B => n4587, S => n4571, Z => n3535);
   U2739 : MUX2_X1 port map( A => n6038, B => n4588, S => n4571, Z => n3534);
   U2740 : MUX2_X1 port map( A => n6034, B => n4589, S => n4571, Z => n3533);
   U2741 : MUX2_X1 port map( A => n6030, B => n4590, S => n4571, Z => n3532);
   U2742 : MUX2_X1 port map( A => n6026, B => n4591, S => n4571, Z => n3531);
   U2743 : MUX2_X1 port map( A => n6022, B => n4592, S => n4571, Z => n3530);
   U2744 : MUX2_X1 port map( A => n6018, B => n4593, S => n4571, Z => n3529);
   U2745 : MUX2_X1 port map( A => n6014, B => n4594, S => n4571, Z => n3528);
   U2746 : MUX2_X1 port map( A => n6010, B => n4595, S => n4571, Z => n3527);
   U2747 : MUX2_X1 port map( A => n6006, B => n4596, S => n4571, Z => n3526);
   U2748 : MUX2_X1 port map( A => n6002, B => n4597, S => n4571, Z => n3525);
   U2749 : MUX2_X1 port map( A => n5998, B => n4598, S => n4571, Z => n3524);
   U2750 : MUX2_X1 port map( A => n5994, B => n4599, S => n4571, Z => n3523);
   U2751 : MUX2_X1 port map( A => n5990, B => n4600, S => n4571, Z => n3522);
   U2752 : MUX2_X1 port map( A => n5986, B => n4601, S => n4571, Z => n3521);
   U2753 : MUX2_X1 port map( A => n5982, B => n4602, S => n4571, Z => n3520);
   U2754 : MUX2_X1 port map( A => n5978, B => n4603, S => n4571, Z => n3519);
   U2755 : MUX2_X1 port map( A => n5974, B => n4604, S => n4571, Z => n3518);
   U2756 : OAI21_X1 port map( B1 => n4605, B2 => n4611, A => n4607, ZN => n4610
                           );
   U2757 : MUX2_X1 port map( A => n6097, B => n4572, S => n4565, Z => n3517);
   U2758 : MUX2_X1 port map( A => n6093, B => n4574, S => n4565, Z => n3516);
   U2759 : MUX2_X1 port map( A => n6089, B => n4575, S => n4565, Z => n3515);
   U2760 : MUX2_X1 port map( A => n6085, B => n4576, S => n4565, Z => n3514);
   U2761 : MUX2_X1 port map( A => n6081, B => n4577, S => n4565, Z => n3513);
   U2762 : MUX2_X1 port map( A => n6077, B => n4578, S => n4565, Z => n3512);
   U2763 : MUX2_X1 port map( A => n6073, B => n4579, S => n4565, Z => n3511);
   U2764 : MUX2_X1 port map( A => n6069, B => n4580, S => n4565, Z => n3510);
   U2765 : MUX2_X1 port map( A => n6065, B => n4581, S => n4565, Z => n3509);
   U2766 : MUX2_X1 port map( A => n6061, B => n4582, S => n4565, Z => n3508);
   U2767 : MUX2_X1 port map( A => n6057, B => n4583, S => n4565, Z => n3507);
   U2768 : MUX2_X1 port map( A => n6053, B => n4584, S => n4565, Z => n3506);
   U2769 : MUX2_X1 port map( A => n6049, B => n4585, S => n4565, Z => n3505);
   U2770 : MUX2_X1 port map( A => n6045, B => n4586, S => n4565, Z => n3504);
   U2771 : MUX2_X1 port map( A => n6041, B => n4587, S => n4565, Z => n3503);
   U2772 : MUX2_X1 port map( A => n6037, B => n4588, S => n4565, Z => n3502);
   U2773 : MUX2_X1 port map( A => n6033, B => n4589, S => n4565, Z => n3501);
   U2774 : MUX2_X1 port map( A => n6029, B => n4590, S => n4565, Z => n3500);
   U2775 : MUX2_X1 port map( A => n6025, B => n4591, S => n4565, Z => n3499);
   U2776 : MUX2_X1 port map( A => n6021, B => n4592, S => n4565, Z => n3498);
   U2777 : MUX2_X1 port map( A => n6017, B => n4593, S => n4565, Z => n3497);
   U2778 : MUX2_X1 port map( A => n6013, B => n4594, S => n4565, Z => n3496);
   U2779 : MUX2_X1 port map( A => n6009, B => n4595, S => n4565, Z => n3495);
   U2780 : MUX2_X1 port map( A => n6005, B => n4596, S => n4565, Z => n3494);
   U2781 : MUX2_X1 port map( A => n6001, B => n4597, S => n4565, Z => n3493);
   U2782 : MUX2_X1 port map( A => n5997, B => n4598, S => n4565, Z => n3492);
   U2783 : MUX2_X1 port map( A => n5993, B => n4599, S => n4565, Z => n3491);
   U2784 : MUX2_X1 port map( A => n5989, B => n4600, S => n4565, Z => n3490);
   U2785 : MUX2_X1 port map( A => n5985, B => n4601, S => n4565, Z => n3489);
   U2786 : MUX2_X1 port map( A => n5981, B => n4602, S => n4565, Z => n3488);
   U2787 : MUX2_X1 port map( A => n5977, B => n4603, S => n4565, Z => n3487);
   U2788 : MUX2_X1 port map( A => n5973, B => n4604, S => n4565, Z => n3486);
   U2789 : OAI21_X1 port map( B1 => n4605, B2 => n4613, A => n4607, ZN => n4612
                           );
   U2790 : MUX2_X1 port map( A => n4414, B => n4572, S => n4567, Z => n3485);
   U2791 : MUX2_X1 port map( A => n4415, B => n4574, S => n4567, Z => n3484);
   U2792 : MUX2_X1 port map( A => n4416, B => n4575, S => n4567, Z => n3483);
   U2793 : MUX2_X1 port map( A => n4417, B => n4576, S => n4567, Z => n3482);
   U2794 : MUX2_X1 port map( A => n4418, B => n4577, S => n4567, Z => n3481);
   U2795 : MUX2_X1 port map( A => n4419, B => n4578, S => n4567, Z => n3480);
   U2796 : MUX2_X1 port map( A => n4420, B => n4579, S => n4567, Z => n3479);
   U2797 : MUX2_X1 port map( A => n4421, B => n4580, S => n4567, Z => n3478);
   U2798 : MUX2_X1 port map( A => n4422, B => n4581, S => n4567, Z => n3477);
   U2799 : MUX2_X1 port map( A => n4423, B => n4582, S => n4567, Z => n3476);
   U2800 : MUX2_X1 port map( A => n4424, B => n4583, S => n4567, Z => n3475);
   U2801 : MUX2_X1 port map( A => n4425, B => n4584, S => n4567, Z => n3474);
   U2802 : MUX2_X1 port map( A => n4426, B => n4585, S => n4567, Z => n3473);
   U2803 : MUX2_X1 port map( A => n4427, B => n4586, S => n4567, Z => n3472);
   U2804 : MUX2_X1 port map( A => n4428, B => n4587, S => n4567, Z => n3471);
   U2805 : MUX2_X1 port map( A => n4429, B => n4588, S => n4567, Z => n3470);
   U2806 : MUX2_X1 port map( A => n4430, B => n4589, S => n4567, Z => n3469);
   U2807 : MUX2_X1 port map( A => n4431, B => n4590, S => n4567, Z => n3468);
   U2808 : MUX2_X1 port map( A => n4432, B => n4591, S => n4567, Z => n3467);
   U2809 : MUX2_X1 port map( A => n4433, B => n4592, S => n4567, Z => n3466);
   U2810 : MUX2_X1 port map( A => n4434, B => n4593, S => n4567, Z => n3465);
   U2811 : MUX2_X1 port map( A => n4435, B => n4594, S => n4567, Z => n3464);
   U2812 : MUX2_X1 port map( A => n4436, B => n4595, S => n4567, Z => n3463);
   U2813 : MUX2_X1 port map( A => n4437, B => n4596, S => n4567, Z => n3462);
   U2814 : MUX2_X1 port map( A => n4438, B => n4597, S => n4567, Z => n3461);
   U2815 : MUX2_X1 port map( A => n4439, B => n4598, S => n4567, Z => n3460);
   U2816 : MUX2_X1 port map( A => n4440, B => n4599, S => n4567, Z => n3459);
   U2817 : MUX2_X1 port map( A => n4441, B => n4600, S => n4567, Z => n3458);
   U2818 : MUX2_X1 port map( A => n4442, B => n4601, S => n4567, Z => n3457);
   U2819 : MUX2_X1 port map( A => n4443, B => n4602, S => n4567, Z => n3456);
   U2820 : MUX2_X1 port map( A => n4444, B => n4603, S => n4567, Z => n3455);
   U2821 : MUX2_X1 port map( A => n4445, B => n4604, S => n4567, Z => n3454);
   U2822 : OAI21_X1 port map( B1 => n4605, B2 => n4615, A => n4607, ZN => n4614
                           );
   U2823 : MUX2_X1 port map( A => n4478, B => n4572, S => n4561, Z => n3453);
   U2824 : MUX2_X1 port map( A => n4479, B => n4574, S => n4561, Z => n3452);
   U2825 : MUX2_X1 port map( A => n4480, B => n4575, S => n4561, Z => n3451);
   U2826 : MUX2_X1 port map( A => n4481, B => n4576, S => n4561, Z => n3450);
   U2827 : MUX2_X1 port map( A => n4482, B => n4577, S => n4561, Z => n3449);
   U2828 : MUX2_X1 port map( A => n4483, B => n4578, S => n4561, Z => n3448);
   U2829 : MUX2_X1 port map( A => n4484, B => n4579, S => n4561, Z => n3447);
   U2830 : MUX2_X1 port map( A => n4485, B => n4580, S => n4561, Z => n3446);
   U2831 : MUX2_X1 port map( A => n4486, B => n4581, S => n4561, Z => n3445);
   U2832 : MUX2_X1 port map( A => n4487, B => n4582, S => n4561, Z => n3444);
   U2833 : MUX2_X1 port map( A => n4488, B => n4583, S => n4561, Z => n3443);
   U2834 : MUX2_X1 port map( A => n4489, B => n4584, S => n4561, Z => n3442);
   U2835 : MUX2_X1 port map( A => n4490, B => n4585, S => n4561, Z => n3441);
   U2836 : MUX2_X1 port map( A => n4491, B => n4586, S => n4561, Z => n3440);
   U2837 : MUX2_X1 port map( A => n4492, B => n4587, S => n4561, Z => n3439);
   U2838 : MUX2_X1 port map( A => n4493, B => n4588, S => n4561, Z => n3438);
   U2839 : MUX2_X1 port map( A => n4494, B => n4589, S => n4561, Z => n3437);
   U2840 : MUX2_X1 port map( A => n4495, B => n4590, S => n4561, Z => n3436);
   U2841 : MUX2_X1 port map( A => n4496, B => n4591, S => n4561, Z => n3435);
   U2842 : MUX2_X1 port map( A => n4497, B => n4592, S => n4561, Z => n3434);
   U2843 : MUX2_X1 port map( A => n4498, B => n4593, S => n4561, Z => n3433);
   U2844 : MUX2_X1 port map( A => n4499, B => n4594, S => n4561, Z => n3432);
   U2845 : MUX2_X1 port map( A => n4500, B => n4595, S => n4561, Z => n3431);
   U2846 : MUX2_X1 port map( A => n4501, B => n4596, S => n4561, Z => n3430);
   U2847 : MUX2_X1 port map( A => n4502, B => n4597, S => n4561, Z => n3429);
   U2848 : MUX2_X1 port map( A => n4503, B => n4598, S => n4561, Z => n3428);
   U2849 : MUX2_X1 port map( A => n4504, B => n4599, S => n4561, Z => n3427);
   U2850 : MUX2_X1 port map( A => n4505, B => n4600, S => n4561, Z => n3426);
   U2851 : MUX2_X1 port map( A => n4506, B => n4601, S => n4561, Z => n3425);
   U2852 : MUX2_X1 port map( A => n4507, B => n4602, S => n4561, Z => n3424);
   U2853 : MUX2_X1 port map( A => n4508, B => n4603, S => n4561, Z => n3423);
   U2854 : MUX2_X1 port map( A => n4509, B => n4604, S => n4561, Z => n3422);
   U2855 : OAI21_X1 port map( B1 => n4605, B2 => n4617, A => n4607, ZN => n4616
                           );
   U2856 : MUX2_X1 port map( A => n6096, B => n4572, S => n4563, Z => n3421);
   U2857 : MUX2_X1 port map( A => n6092, B => n4574, S => n4563, Z => n3420);
   U2858 : MUX2_X1 port map( A => n6088, B => n4575, S => n4563, Z => n3419);
   U2859 : MUX2_X1 port map( A => n6084, B => n4576, S => n4563, Z => n3418);
   U2860 : MUX2_X1 port map( A => n6080, B => n4577, S => n4563, Z => n3417);
   U2861 : MUX2_X1 port map( A => n6076, B => n4578, S => n4563, Z => n3416);
   U2862 : MUX2_X1 port map( A => n6072, B => n4579, S => n4563, Z => n3415);
   U2863 : MUX2_X1 port map( A => n6068, B => n4580, S => n4563, Z => n3414);
   U2864 : MUX2_X1 port map( A => n6064, B => n4581, S => n4563, Z => n3413);
   U2865 : MUX2_X1 port map( A => n6060, B => n4582, S => n4563, Z => n3412);
   U2866 : MUX2_X1 port map( A => n6056, B => n4583, S => n4563, Z => n3411);
   U2867 : MUX2_X1 port map( A => n6052, B => n4584, S => n4563, Z => n3410);
   U2868 : MUX2_X1 port map( A => n6048, B => n4585, S => n4563, Z => n3409);
   U2869 : MUX2_X1 port map( A => n6044, B => n4586, S => n4563, Z => n3408);
   U2870 : MUX2_X1 port map( A => n6040, B => n4587, S => n4563, Z => n3407);
   U2871 : MUX2_X1 port map( A => n6036, B => n4588, S => n4563, Z => n3406);
   U2872 : MUX2_X1 port map( A => n6032, B => n4589, S => n4563, Z => n3405);
   U2873 : MUX2_X1 port map( A => n6028, B => n4590, S => n4563, Z => n3404);
   U2874 : MUX2_X1 port map( A => n6024, B => n4591, S => n4563, Z => n3403);
   U2875 : MUX2_X1 port map( A => n6020, B => n4592, S => n4563, Z => n3402);
   U2876 : MUX2_X1 port map( A => n6016, B => n4593, S => n4563, Z => n3401);
   U2877 : MUX2_X1 port map( A => n6012, B => n4594, S => n4563, Z => n3400);
   U2878 : MUX2_X1 port map( A => n6008, B => n4595, S => n4563, Z => n3399);
   U2879 : MUX2_X1 port map( A => n6004, B => n4596, S => n4563, Z => n3398);
   U2880 : MUX2_X1 port map( A => n6000, B => n4597, S => n4563, Z => n3397);
   U2881 : MUX2_X1 port map( A => n5996, B => n4598, S => n4563, Z => n3396);
   U2882 : MUX2_X1 port map( A => n5992, B => n4599, S => n4563, Z => n3395);
   U2883 : MUX2_X1 port map( A => n5988, B => n4600, S => n4563, Z => n3394);
   U2884 : MUX2_X1 port map( A => n5984, B => n4601, S => n4563, Z => n3393);
   U2885 : MUX2_X1 port map( A => n5980, B => n4602, S => n4563, Z => n3392);
   U2886 : MUX2_X1 port map( A => n5976, B => n4603, S => n4563, Z => n3391);
   U2887 : MUX2_X1 port map( A => n5972, B => n4604, S => n4563, Z => n3390);
   U2888 : OAI21_X1 port map( B1 => n4605, B2 => n4619, A => n4607, ZN => n4618
                           );
   U2889 : MUX2_X1 port map( A => n6095, B => n4572, S => n4557, Z => n3389);
   U2890 : MUX2_X1 port map( A => n6091, B => n4574, S => n4557, Z => n3388);
   U2891 : MUX2_X1 port map( A => n6087, B => n4575, S => n4557, Z => n3387);
   U2892 : MUX2_X1 port map( A => n6083, B => n4576, S => n4557, Z => n3386);
   U2893 : MUX2_X1 port map( A => n6079, B => n4577, S => n4557, Z => n3385);
   U2894 : MUX2_X1 port map( A => n6075, B => n4578, S => n4557, Z => n3384);
   U2895 : MUX2_X1 port map( A => n6071, B => n4579, S => n4557, Z => n3383);
   U2896 : MUX2_X1 port map( A => n6067, B => n4580, S => n4557, Z => n3382);
   U2897 : MUX2_X1 port map( A => n6063, B => n4581, S => n4557, Z => n3381);
   U2898 : MUX2_X1 port map( A => n6059, B => n4582, S => n4557, Z => n3380);
   U2899 : MUX2_X1 port map( A => n6055, B => n4583, S => n4557, Z => n3379);
   U2900 : MUX2_X1 port map( A => n6051, B => n4584, S => n4557, Z => n3378);
   U2901 : MUX2_X1 port map( A => n6047, B => n4585, S => n4557, Z => n3377);
   U2902 : MUX2_X1 port map( A => n6043, B => n4586, S => n4557, Z => n3376);
   U2903 : MUX2_X1 port map( A => n6039, B => n4587, S => n4557, Z => n3375);
   U2904 : MUX2_X1 port map( A => n6035, B => n4588, S => n4557, Z => n3374);
   U2905 : MUX2_X1 port map( A => n6031, B => n4589, S => n4557, Z => n3373);
   U2906 : MUX2_X1 port map( A => n6027, B => n4590, S => n4557, Z => n3372);
   U2907 : MUX2_X1 port map( A => n6023, B => n4591, S => n4557, Z => n3371);
   U2908 : MUX2_X1 port map( A => n6019, B => n4592, S => n4557, Z => n3370);
   U2909 : MUX2_X1 port map( A => n6015, B => n4593, S => n4557, Z => n3369);
   U2910 : MUX2_X1 port map( A => n6011, B => n4594, S => n4557, Z => n3368);
   U2911 : MUX2_X1 port map( A => n6007, B => n4595, S => n4557, Z => n3367);
   U2912 : MUX2_X1 port map( A => n6003, B => n4596, S => n4557, Z => n3366);
   U2913 : MUX2_X1 port map( A => n5999, B => n4597, S => n4557, Z => n3365);
   U2914 : MUX2_X1 port map( A => n5995, B => n4598, S => n4557, Z => n3364);
   U2915 : MUX2_X1 port map( A => n5991, B => n4599, S => n4557, Z => n3363);
   U2916 : MUX2_X1 port map( A => n5987, B => n4600, S => n4557, Z => n3362);
   U2917 : MUX2_X1 port map( A => n5983, B => n4601, S => n4557, Z => n3361);
   U2918 : MUX2_X1 port map( A => n5979, B => n4602, S => n4557, Z => n3360);
   U2919 : MUX2_X1 port map( A => n5975, B => n4603, S => n4557, Z => n3359);
   U2920 : MUX2_X1 port map( A => n5971, B => n4604, S => n4557, Z => n3358);
   U2921 : OAI21_X1 port map( B1 => n4605, B2 => n4621, A => n4607, ZN => n4620
                           );
   U2922 : NAND3_X1 port map( A1 => n4622, A2 => n4623, A3 => n4624, ZN => 
                           n4605);
   U2923 : MUX2_X1 port map( A => n3934, B => n4572, S => n4559, Z => n3357);
   U2924 : MUX2_X1 port map( A => n3935, B => n4574, S => n4559, Z => n3356);
   U2925 : MUX2_X1 port map( A => n3936, B => n4575, S => n4559, Z => n3355);
   U2926 : MUX2_X1 port map( A => n3937, B => n4576, S => n4559, Z => n3354);
   U2927 : MUX2_X1 port map( A => n3938, B => n4577, S => n4559, Z => n3353);
   U2928 : MUX2_X1 port map( A => n3939, B => n4578, S => n4559, Z => n3352);
   U2929 : MUX2_X1 port map( A => n3940, B => n4579, S => n4559, Z => n3351);
   U2930 : MUX2_X1 port map( A => n3941, B => n4580, S => n4559, Z => n3350);
   U2931 : MUX2_X1 port map( A => n3942, B => n4581, S => n4559, Z => n3349);
   U2932 : MUX2_X1 port map( A => n3943, B => n4582, S => n4559, Z => n3348);
   U2933 : MUX2_X1 port map( A => n3944, B => n4583, S => n4559, Z => n3347);
   U2934 : MUX2_X1 port map( A => n3945, B => n4584, S => n4559, Z => n3346);
   U2935 : MUX2_X1 port map( A => n3946, B => n4585, S => n4559, Z => n3345);
   U2936 : MUX2_X1 port map( A => n3947, B => n4586, S => n4559, Z => n3344);
   U2937 : MUX2_X1 port map( A => n3948, B => n4587, S => n4559, Z => n3343);
   U2938 : MUX2_X1 port map( A => n3949, B => n4588, S => n4559, Z => n3342);
   U2939 : MUX2_X1 port map( A => n3950, B => n4589, S => n4559, Z => n3341);
   U2940 : MUX2_X1 port map( A => n3951, B => n4590, S => n4559, Z => n3340);
   U2941 : MUX2_X1 port map( A => n3952, B => n4591, S => n4559, Z => n3339);
   U2942 : MUX2_X1 port map( A => n3953, B => n4592, S => n4559, Z => n3338);
   U2943 : MUX2_X1 port map( A => n3954, B => n4593, S => n4559, Z => n3337);
   U2944 : MUX2_X1 port map( A => n3955, B => n4594, S => n4559, Z => n3336);
   U2945 : MUX2_X1 port map( A => n3956, B => n4595, S => n4559, Z => n3335);
   U2946 : MUX2_X1 port map( A => n3957, B => n4596, S => n4559, Z => n3334);
   U2947 : MUX2_X1 port map( A => n3958, B => n4597, S => n4559, Z => n3333);
   U2948 : MUX2_X1 port map( A => n3959, B => n4598, S => n4559, Z => n3332);
   U2949 : MUX2_X1 port map( A => n3960, B => n4599, S => n4559, Z => n3331);
   U2950 : MUX2_X1 port map( A => n3961, B => n4600, S => n4559, Z => n3330);
   U2951 : MUX2_X1 port map( A => n3962, B => n4601, S => n4559, Z => n3329);
   U2952 : MUX2_X1 port map( A => n3963, B => n4602, S => n4559, Z => n3328);
   U2953 : MUX2_X1 port map( A => n3964, B => n4603, S => n4559, Z => n3327);
   U2954 : MUX2_X1 port map( A => n3965, B => n4604, S => n4559, Z => n3326);
   U2955 : OAI21_X1 port map( B1 => n4606, B2 => n4626, A => n4607, ZN => n4625
                           );
   U2956 : MUX2_X1 port map( A => n4318, B => n4572, S => n4553, Z => n3325);
   U2957 : MUX2_X1 port map( A => n4319, B => n4574, S => n4553, Z => n3324);
   U2958 : MUX2_X1 port map( A => n4320, B => n4575, S => n4553, Z => n3323);
   U2959 : MUX2_X1 port map( A => n4321, B => n4576, S => n4553, Z => n3322);
   U2960 : MUX2_X1 port map( A => n4322, B => n4577, S => n4553, Z => n3321);
   U2961 : MUX2_X1 port map( A => n4323, B => n4578, S => n4553, Z => n3320);
   U2962 : MUX2_X1 port map( A => n4324, B => n4579, S => n4553, Z => n3319);
   U2963 : MUX2_X1 port map( A => n4325, B => n4580, S => n4553, Z => n3318);
   U2964 : MUX2_X1 port map( A => n4326, B => n4581, S => n4553, Z => n3317);
   U2965 : MUX2_X1 port map( A => n4327, B => n4582, S => n4553, Z => n3316);
   U2966 : MUX2_X1 port map( A => n4328, B => n4583, S => n4553, Z => n3315);
   U2967 : MUX2_X1 port map( A => n4329, B => n4584, S => n4553, Z => n3314);
   U2968 : MUX2_X1 port map( A => n4330, B => n4585, S => n4553, Z => n3313);
   U2969 : MUX2_X1 port map( A => n4331, B => n4586, S => n4553, Z => n3312);
   U2970 : MUX2_X1 port map( A => n4332, B => n4587, S => n4553, Z => n3311);
   U2971 : MUX2_X1 port map( A => n4333, B => n4588, S => n4553, Z => n3310);
   U2972 : MUX2_X1 port map( A => n4334, B => n4589, S => n4553, Z => n3309);
   U2973 : MUX2_X1 port map( A => n4335, B => n4590, S => n4553, Z => n3308);
   U2974 : MUX2_X1 port map( A => n4336, B => n4591, S => n4553, Z => n3307);
   U2975 : MUX2_X1 port map( A => n4337, B => n4592, S => n4553, Z => n3306);
   U2976 : MUX2_X1 port map( A => n4338, B => n4593, S => n4553, Z => n3305);
   U2977 : MUX2_X1 port map( A => n4339, B => n4594, S => n4553, Z => n3304);
   U2978 : MUX2_X1 port map( A => n4340, B => n4595, S => n4553, Z => n3303);
   U2979 : MUX2_X1 port map( A => n4341, B => n4596, S => n4553, Z => n3302);
   U2980 : MUX2_X1 port map( A => n4342, B => n4597, S => n4553, Z => n3301);
   U2981 : MUX2_X1 port map( A => n4343, B => n4598, S => n4553, Z => n3300);
   U2982 : MUX2_X1 port map( A => n4344, B => n4599, S => n4553, Z => n3299);
   U2983 : MUX2_X1 port map( A => n4345, B => n4600, S => n4553, Z => n3298);
   U2984 : MUX2_X1 port map( A => n4346, B => n4601, S => n4553, Z => n3297);
   U2985 : MUX2_X1 port map( A => n4347, B => n4602, S => n4553, Z => n3296);
   U2986 : MUX2_X1 port map( A => n4348, B => n4603, S => n4553, Z => n3295);
   U2987 : MUX2_X1 port map( A => n4349, B => n4604, S => n4553, Z => n3294);
   U2988 : OAI21_X1 port map( B1 => n4609, B2 => n4626, A => n4607, ZN => n4627
                           );
   U2989 : MUX2_X1 port map( A => n3966, B => n4572, S => n4555, Z => n3293);
   U2990 : MUX2_X1 port map( A => n3967, B => n4574, S => n4555, Z => n3292);
   U2991 : MUX2_X1 port map( A => n3968, B => n4575, S => n4555, Z => n3291);
   U2992 : MUX2_X1 port map( A => n3969, B => n4576, S => n4555, Z => n3290);
   U2993 : MUX2_X1 port map( A => n3970, B => n4577, S => n4555, Z => n3289);
   U2994 : MUX2_X1 port map( A => n3971, B => n4578, S => n4555, Z => n3288);
   U2995 : MUX2_X1 port map( A => n3972, B => n4579, S => n4555, Z => n3287);
   U2996 : MUX2_X1 port map( A => n3973, B => n4580, S => n4555, Z => n3286);
   U2997 : MUX2_X1 port map( A => n3974, B => n4581, S => n4555, Z => n3285);
   U2998 : MUX2_X1 port map( A => n3975, B => n4582, S => n4555, Z => n3284);
   U2999 : MUX2_X1 port map( A => n3976, B => n4583, S => n4555, Z => n3283);
   U3000 : MUX2_X1 port map( A => n3977, B => n4584, S => n4555, Z => n3282);
   U3001 : MUX2_X1 port map( A => n3978, B => n4585, S => n4555, Z => n3281);
   U3002 : MUX2_X1 port map( A => n3979, B => n4586, S => n4555, Z => n3280);
   U3003 : MUX2_X1 port map( A => n3980, B => n4587, S => n4555, Z => n3279);
   U3004 : MUX2_X1 port map( A => n3981, B => n4588, S => n4555, Z => n3278);
   U3005 : MUX2_X1 port map( A => n3982, B => n4589, S => n4555, Z => n3277);
   U3006 : MUX2_X1 port map( A => n3983, B => n4590, S => n4555, Z => n3276);
   U3007 : MUX2_X1 port map( A => n3984, B => n4591, S => n4555, Z => n3275);
   U3008 : MUX2_X1 port map( A => n3985, B => n4592, S => n4555, Z => n3274);
   U3009 : MUX2_X1 port map( A => n3986, B => n4593, S => n4555, Z => n3273);
   U3010 : MUX2_X1 port map( A => n3987, B => n4594, S => n4555, Z => n3272);
   U3011 : MUX2_X1 port map( A => n3988, B => n4595, S => n4555, Z => n3271);
   U3012 : MUX2_X1 port map( A => n3989, B => n4596, S => n4555, Z => n3270);
   U3013 : MUX2_X1 port map( A => n3990, B => n4597, S => n4555, Z => n3269);
   U3014 : MUX2_X1 port map( A => n3991, B => n4598, S => n4555, Z => n3268);
   U3015 : MUX2_X1 port map( A => n3992, B => n4599, S => n4555, Z => n3267);
   U3016 : MUX2_X1 port map( A => n3993, B => n4600, S => n4555, Z => n3266);
   U3017 : MUX2_X1 port map( A => n3994, B => n4601, S => n4555, Z => n3265);
   U3018 : MUX2_X1 port map( A => n3995, B => n4602, S => n4555, Z => n3264);
   U3019 : MUX2_X1 port map( A => n3996, B => n4603, S => n4555, Z => n3263);
   U3020 : MUX2_X1 port map( A => n3997, B => n4604, S => n4555, Z => n3262);
   U3021 : OAI21_X1 port map( B1 => n4611, B2 => n4626, A => n4607, ZN => n4628
                           );
   U3022 : MUX2_X1 port map( A => n4350, B => n4572, S => n4549, Z => n3261);
   U3023 : MUX2_X1 port map( A => n4351, B => n4574, S => n4549, Z => n3260);
   U3024 : MUX2_X1 port map( A => n4352, B => n4575, S => n4549, Z => n3259);
   U3025 : MUX2_X1 port map( A => n4353, B => n4576, S => n4549, Z => n3258);
   U3026 : MUX2_X1 port map( A => n4354, B => n4577, S => n4549, Z => n3257);
   U3027 : MUX2_X1 port map( A => n4355, B => n4578, S => n4549, Z => n3256);
   U3028 : MUX2_X1 port map( A => n4356, B => n4579, S => n4549, Z => n3255);
   U3029 : MUX2_X1 port map( A => n4357, B => n4580, S => n4549, Z => n3254);
   U3030 : MUX2_X1 port map( A => n4358, B => n4581, S => n4549, Z => n3253);
   U3031 : MUX2_X1 port map( A => n4359, B => n4582, S => n4549, Z => n3252);
   U3032 : MUX2_X1 port map( A => n4360, B => n4583, S => n4549, Z => n3251);
   U3033 : MUX2_X1 port map( A => n4361, B => n4584, S => n4549, Z => n3250);
   U3034 : MUX2_X1 port map( A => n4362, B => n4585, S => n4549, Z => n3249);
   U3035 : MUX2_X1 port map( A => n4363, B => n4586, S => n4549, Z => n3248);
   U3036 : MUX2_X1 port map( A => n4364, B => n4587, S => n4549, Z => n3247);
   U3037 : MUX2_X1 port map( A => n4365, B => n4588, S => n4549, Z => n3246);
   U3038 : MUX2_X1 port map( A => n4366, B => n4589, S => n4549, Z => n3245);
   U3039 : MUX2_X1 port map( A => n4367, B => n4590, S => n4549, Z => n3244);
   U3040 : MUX2_X1 port map( A => n4368, B => n4591, S => n4549, Z => n3243);
   U3041 : MUX2_X1 port map( A => n4369, B => n4592, S => n4549, Z => n3242);
   U3042 : MUX2_X1 port map( A => n4370, B => n4593, S => n4549, Z => n3241);
   U3043 : MUX2_X1 port map( A => n4371, B => n4594, S => n4549, Z => n3240);
   U3044 : MUX2_X1 port map( A => n4372, B => n4595, S => n4549, Z => n3239);
   U3045 : MUX2_X1 port map( A => n4373, B => n4596, S => n4549, Z => n3238);
   U3046 : MUX2_X1 port map( A => n4374, B => n4597, S => n4549, Z => n3237);
   U3047 : MUX2_X1 port map( A => n4375, B => n4598, S => n4549, Z => n3236);
   U3048 : MUX2_X1 port map( A => n4376, B => n4599, S => n4549, Z => n3235);
   U3049 : MUX2_X1 port map( A => n4377, B => n4600, S => n4549, Z => n3234);
   U3050 : MUX2_X1 port map( A => n4378, B => n4601, S => n4549, Z => n3233);
   U3051 : MUX2_X1 port map( A => n4379, B => n4602, S => n4549, Z => n3232);
   U3052 : MUX2_X1 port map( A => n4380, B => n4603, S => n4549, Z => n3231);
   U3053 : MUX2_X1 port map( A => n4381, B => n4604, S => n4549, Z => n3230);
   U3054 : OAI21_X1 port map( B1 => n4613, B2 => n4626, A => n4607, ZN => n4629
                           );
   U3055 : MUX2_X1 port map( A => n3614, B => n4572, S => n4551, Z => n3229);
   U3056 : MUX2_X1 port map( A => n3619, B => n4574, S => n4551, Z => n3228);
   U3057 : MUX2_X1 port map( A => n3624, B => n4575, S => n4551, Z => n3227);
   U3058 : MUX2_X1 port map( A => n3629, B => n4576, S => n4551, Z => n3226);
   U3059 : MUX2_X1 port map( A => n3634, B => n4577, S => n4551, Z => n3225);
   U3060 : MUX2_X1 port map( A => n3639, B => n4578, S => n4551, Z => n3224);
   U3061 : MUX2_X1 port map( A => n3644, B => n4579, S => n4551, Z => n3223);
   U3062 : MUX2_X1 port map( A => n3649, B => n4580, S => n4551, Z => n3222);
   U3063 : MUX2_X1 port map( A => n3654, B => n4581, S => n4551, Z => n3221);
   U3064 : MUX2_X1 port map( A => n3659, B => n4582, S => n4551, Z => n3220);
   U3065 : MUX2_X1 port map( A => n3664, B => n4583, S => n4551, Z => n3219);
   U3066 : MUX2_X1 port map( A => n3669, B => n4584, S => n4551, Z => n3218);
   U3067 : MUX2_X1 port map( A => n3674, B => n4585, S => n4551, Z => n3217);
   U3068 : MUX2_X1 port map( A => n3679, B => n4586, S => n4551, Z => n3216);
   U3069 : MUX2_X1 port map( A => n3684, B => n4587, S => n4551, Z => n3215);
   U3070 : MUX2_X1 port map( A => n3689, B => n4588, S => n4551, Z => n3214);
   U3071 : MUX2_X1 port map( A => n3694, B => n4589, S => n4551, Z => n3213);
   U3072 : MUX2_X1 port map( A => n3699, B => n4590, S => n4551, Z => n3212);
   U3073 : MUX2_X1 port map( A => n3704, B => n4591, S => n4551, Z => n3211);
   U3074 : MUX2_X1 port map( A => n3709, B => n4592, S => n4551, Z => n3210);
   U3075 : MUX2_X1 port map( A => n3714, B => n4593, S => n4551, Z => n3209);
   U3076 : MUX2_X1 port map( A => n3719, B => n4594, S => n4551, Z => n3208);
   U3077 : MUX2_X1 port map( A => n3724, B => n4595, S => n4551, Z => n3207);
   U3078 : MUX2_X1 port map( A => n3729, B => n4596, S => n4551, Z => n3206);
   U3079 : MUX2_X1 port map( A => n3734, B => n4597, S => n4551, Z => n3205);
   U3080 : MUX2_X1 port map( A => n3739, B => n4598, S => n4551, Z => n3204);
   U3081 : MUX2_X1 port map( A => n3744, B => n4599, S => n4551, Z => n3203);
   U3082 : MUX2_X1 port map( A => n3749, B => n4600, S => n4551, Z => n3202);
   U3083 : MUX2_X1 port map( A => n3754, B => n4601, S => n4551, Z => n3201);
   U3084 : MUX2_X1 port map( A => n3759, B => n4602, S => n4551, Z => n3200);
   U3085 : MUX2_X1 port map( A => n3764, B => n4603, S => n4551, Z => n3199);
   U3086 : MUX2_X1 port map( A => n3769, B => n4604, S => n4551, Z => n3198);
   U3087 : OAI21_X1 port map( B1 => n4615, B2 => n4626, A => n4607, ZN => n4630
                           );
   U3088 : MUX2_X1 port map( A => n3998, B => n4572, S => n4545, Z => n3197);
   U3089 : MUX2_X1 port map( A => n4003, B => n4574, S => n4545, Z => n3196);
   U3090 : MUX2_X1 port map( A => n4008, B => n4575, S => n4545, Z => n3195);
   U3091 : MUX2_X1 port map( A => n4013, B => n4576, S => n4545, Z => n3194);
   U3092 : MUX2_X1 port map( A => n4018, B => n4577, S => n4545, Z => n3193);
   U3093 : MUX2_X1 port map( A => n4023, B => n4578, S => n4545, Z => n3192);
   U3094 : MUX2_X1 port map( A => n4028, B => n4579, S => n4545, Z => n3191);
   U3095 : MUX2_X1 port map( A => n4033, B => n4580, S => n4545, Z => n3190);
   U3096 : MUX2_X1 port map( A => n4038, B => n4581, S => n4545, Z => n3189);
   U3097 : MUX2_X1 port map( A => n4043, B => n4582, S => n4545, Z => n3188);
   U3098 : MUX2_X1 port map( A => n4048, B => n4583, S => n4545, Z => n3187);
   U3099 : MUX2_X1 port map( A => n4053, B => n4584, S => n4545, Z => n3186);
   U3100 : MUX2_X1 port map( A => n4058, B => n4585, S => n4545, Z => n3185);
   U3101 : MUX2_X1 port map( A => n4063, B => n4586, S => n4545, Z => n3184);
   U3102 : MUX2_X1 port map( A => n4068, B => n4587, S => n4545, Z => n3183);
   U3103 : MUX2_X1 port map( A => n4073, B => n4588, S => n4545, Z => n3182);
   U3104 : MUX2_X1 port map( A => n4078, B => n4589, S => n4545, Z => n3181);
   U3105 : MUX2_X1 port map( A => n4083, B => n4590, S => n4545, Z => n3180);
   U3106 : MUX2_X1 port map( A => n4088, B => n4591, S => n4545, Z => n3179);
   U3107 : MUX2_X1 port map( A => n4093, B => n4592, S => n4545, Z => n3178);
   U3108 : MUX2_X1 port map( A => n4098, B => n4593, S => n4545, Z => n3177);
   U3109 : MUX2_X1 port map( A => n4103, B => n4594, S => n4545, Z => n3176);
   U3110 : MUX2_X1 port map( A => n4108, B => n4595, S => n4545, Z => n3175);
   U3111 : MUX2_X1 port map( A => n4113, B => n4596, S => n4545, Z => n3174);
   U3112 : MUX2_X1 port map( A => n4118, B => n4597, S => n4545, Z => n3173);
   U3113 : MUX2_X1 port map( A => n4123, B => n4598, S => n4545, Z => n3172);
   U3114 : MUX2_X1 port map( A => n4128, B => n4599, S => n4545, Z => n3171);
   U3115 : MUX2_X1 port map( A => n4133, B => n4600, S => n4545, Z => n3170);
   U3116 : MUX2_X1 port map( A => n4138, B => n4601, S => n4545, Z => n3169);
   U3117 : MUX2_X1 port map( A => n4143, B => n4602, S => n4545, Z => n3168);
   U3118 : MUX2_X1 port map( A => n4148, B => n4603, S => n4545, Z => n3167);
   U3119 : MUX2_X1 port map( A => n4153, B => n4604, S => n4545, Z => n3166);
   U3120 : OAI21_X1 port map( B1 => n4617, B2 => n4626, A => n4607, ZN => n4631
                           );
   U3121 : MUX2_X1 port map( A => n6418, B => n4572, S => n4547, Z => n3165);
   U3122 : MUX2_X1 port map( A => n6417, B => n4574, S => n4547, Z => n3164);
   U3123 : MUX2_X1 port map( A => n6416, B => n4575, S => n4547, Z => n3163);
   U3124 : MUX2_X1 port map( A => n6415, B => n4576, S => n4547, Z => n3162);
   U3125 : MUX2_X1 port map( A => n6414, B => n4577, S => n4547, Z => n3161);
   U3126 : MUX2_X1 port map( A => n6413, B => n4578, S => n4547, Z => n3160);
   U3127 : MUX2_X1 port map( A => n6412, B => n4579, S => n4547, Z => n3159);
   U3128 : MUX2_X1 port map( A => n6411, B => n4580, S => n4547, Z => n3158);
   U3129 : MUX2_X1 port map( A => n6410, B => n4581, S => n4547, Z => n3157);
   U3130 : MUX2_X1 port map( A => n6409, B => n4582, S => n4547, Z => n3156);
   U3131 : MUX2_X1 port map( A => n6408, B => n4583, S => n4547, Z => n3155);
   U3132 : MUX2_X1 port map( A => n6407, B => n4584, S => n4547, Z => n3154);
   U3133 : MUX2_X1 port map( A => n6406, B => n4585, S => n4547, Z => n3153);
   U3134 : MUX2_X1 port map( A => n6405, B => n4586, S => n4547, Z => n3152);
   U3135 : MUX2_X1 port map( A => n6404, B => n4587, S => n4547, Z => n3151);
   U3136 : MUX2_X1 port map( A => n6403, B => n4588, S => n4547, Z => n3150);
   U3137 : MUX2_X1 port map( A => n6402, B => n4589, S => n4547, Z => n3149);
   U3138 : MUX2_X1 port map( A => n6401, B => n4590, S => n4547, Z => n3148);
   U3139 : MUX2_X1 port map( A => n6400, B => n4591, S => n4547, Z => n3147);
   U3140 : MUX2_X1 port map( A => n6399, B => n4592, S => n4547, Z => n3146);
   U3141 : MUX2_X1 port map( A => n6398, B => n4593, S => n4547, Z => n3145);
   U3142 : MUX2_X1 port map( A => n6397, B => n4594, S => n4547, Z => n3144);
   U3143 : MUX2_X1 port map( A => n6396, B => n4595, S => n4547, Z => n3143);
   U3144 : MUX2_X1 port map( A => n6395, B => n4596, S => n4547, Z => n3142);
   U3145 : MUX2_X1 port map( A => n6394, B => n4597, S => n4547, Z => n3141);
   U3146 : MUX2_X1 port map( A => n6393, B => n4598, S => n4547, Z => n3140);
   U3147 : MUX2_X1 port map( A => n6392, B => n4599, S => n4547, Z => n3139);
   U3148 : MUX2_X1 port map( A => n6391, B => n4600, S => n4547, Z => n3138);
   U3149 : MUX2_X1 port map( A => n6390, B => n4601, S => n4547, Z => n3137);
   U3150 : MUX2_X1 port map( A => n6389, B => n4602, S => n4547, Z => n3136);
   U3151 : MUX2_X1 port map( A => n6388, B => n4603, S => n4547, Z => n3135);
   U3152 : MUX2_X1 port map( A => n6387, B => n4604, S => n4547, Z => n3134);
   U3153 : OAI21_X1 port map( B1 => n4619, B2 => n4626, A => n4607, ZN => n4632
                           );
   U3154 : MUX2_X1 port map( A => n6386, B => n4572, S => n4541, Z => n3133);
   U3155 : MUX2_X1 port map( A => n6385, B => n4574, S => n4541, Z => n3132);
   U3156 : MUX2_X1 port map( A => n6384, B => n4575, S => n4541, Z => n3131);
   U3157 : MUX2_X1 port map( A => n6383, B => n4576, S => n4541, Z => n3130);
   U3158 : MUX2_X1 port map( A => n6382, B => n4577, S => n4541, Z => n3129);
   U3159 : MUX2_X1 port map( A => n6381, B => n4578, S => n4541, Z => n3128);
   U3160 : MUX2_X1 port map( A => n6380, B => n4579, S => n4541, Z => n3127);
   U3161 : MUX2_X1 port map( A => n6379, B => n4580, S => n4541, Z => n3126);
   U3162 : MUX2_X1 port map( A => n6378, B => n4581, S => n4541, Z => n3125);
   U3163 : MUX2_X1 port map( A => n6377, B => n4582, S => n4541, Z => n3124);
   U3164 : MUX2_X1 port map( A => n6376, B => n4583, S => n4541, Z => n3123);
   U3165 : MUX2_X1 port map( A => n6375, B => n4584, S => n4541, Z => n3122);
   U3166 : MUX2_X1 port map( A => n6374, B => n4585, S => n4541, Z => n3121);
   U3167 : MUX2_X1 port map( A => n6373, B => n4586, S => n4541, Z => n3120);
   U3168 : MUX2_X1 port map( A => n6372, B => n4587, S => n4541, Z => n3119);
   U3169 : MUX2_X1 port map( A => n6371, B => n4588, S => n4541, Z => n3118);
   U3170 : MUX2_X1 port map( A => n6370, B => n4589, S => n4541, Z => n3117);
   U3171 : MUX2_X1 port map( A => n6369, B => n4590, S => n4541, Z => n3116);
   U3172 : MUX2_X1 port map( A => n6368, B => n4591, S => n4541, Z => n3115);
   U3173 : MUX2_X1 port map( A => n6367, B => n4592, S => n4541, Z => n3114);
   U3174 : MUX2_X1 port map( A => n6366, B => n4593, S => n4541, Z => n3113);
   U3175 : MUX2_X1 port map( A => n6365, B => n4594, S => n4541, Z => n3112);
   U3176 : MUX2_X1 port map( A => n6364, B => n4595, S => n4541, Z => n3111);
   U3177 : MUX2_X1 port map( A => n6363, B => n4596, S => n4541, Z => n3110);
   U3178 : MUX2_X1 port map( A => n6362, B => n4597, S => n4541, Z => n3109);
   U3179 : MUX2_X1 port map( A => n6361, B => n4598, S => n4541, Z => n3108);
   U3180 : MUX2_X1 port map( A => n6360, B => n4599, S => n4541, Z => n3107);
   U3181 : MUX2_X1 port map( A => n6359, B => n4600, S => n4541, Z => n3106);
   U3182 : MUX2_X1 port map( A => n6358, B => n4601, S => n4541, Z => n3105);
   U3183 : MUX2_X1 port map( A => n6357, B => n4602, S => n4541, Z => n3104);
   U3184 : MUX2_X1 port map( A => n6356, B => n4603, S => n4541, Z => n3103);
   U3185 : MUX2_X1 port map( A => n6355, B => n4604, S => n4541, Z => n3102);
   U3186 : OAI21_X1 port map( B1 => n4621, B2 => n4626, A => n4607, ZN => n4633
                           );
   U3187 : NAND3_X1 port map( A1 => n4624, A2 => n4623, A3 => ADD_WR(3), ZN => 
                           n4626);
   U3188 : INV_X1 port map( A => ADD_WR(4), ZN => n4623);
   U3189 : MUX2_X1 port map( A => n3615, B => n4572, S => n4543, Z => n3101);
   U3190 : MUX2_X1 port map( A => n3620, B => n4574, S => n4543, Z => n3100);
   U3191 : MUX2_X1 port map( A => n3625, B => n4575, S => n4543, Z => n3099);
   U3192 : MUX2_X1 port map( A => n3630, B => n4576, S => n4543, Z => n3098);
   U3193 : MUX2_X1 port map( A => n3635, B => n4577, S => n4543, Z => n3097);
   U3194 : MUX2_X1 port map( A => n3640, B => n4578, S => n4543, Z => n3096);
   U3195 : MUX2_X1 port map( A => n3645, B => n4579, S => n4543, Z => n3095);
   U3196 : MUX2_X1 port map( A => n3650, B => n4580, S => n4543, Z => n3094);
   U3197 : MUX2_X1 port map( A => n3655, B => n4581, S => n4543, Z => n3093);
   U3198 : MUX2_X1 port map( A => n3660, B => n4582, S => n4543, Z => n3092);
   U3199 : MUX2_X1 port map( A => n3665, B => n4583, S => n4543, Z => n3091);
   U3200 : MUX2_X1 port map( A => n3670, B => n4584, S => n4543, Z => n3090);
   U3201 : MUX2_X1 port map( A => n3675, B => n4585, S => n4543, Z => n3089);
   U3202 : MUX2_X1 port map( A => n3680, B => n4586, S => n4543, Z => n3088);
   U3203 : MUX2_X1 port map( A => n3685, B => n4587, S => n4543, Z => n3087);
   U3204 : MUX2_X1 port map( A => n3690, B => n4588, S => n4543, Z => n3086);
   U3205 : MUX2_X1 port map( A => n3695, B => n4589, S => n4543, Z => n3085);
   U3206 : MUX2_X1 port map( A => n3700, B => n4590, S => n4543, Z => n3084);
   U3207 : MUX2_X1 port map( A => n3705, B => n4591, S => n4543, Z => n3083);
   U3208 : MUX2_X1 port map( A => n3710, B => n4592, S => n4543, Z => n3082);
   U3209 : MUX2_X1 port map( A => n3715, B => n4593, S => n4543, Z => n3081);
   U3210 : MUX2_X1 port map( A => n3720, B => n4594, S => n4543, Z => n3080);
   U3211 : MUX2_X1 port map( A => n3725, B => n4595, S => n4543, Z => n3079);
   U3212 : MUX2_X1 port map( A => n3730, B => n4596, S => n4543, Z => n3078);
   U3213 : MUX2_X1 port map( A => n3735, B => n4597, S => n4543, Z => n3077);
   U3214 : MUX2_X1 port map( A => n3740, B => n4598, S => n4543, Z => n3076);
   U3215 : MUX2_X1 port map( A => n3745, B => n4599, S => n4543, Z => n3075);
   U3216 : MUX2_X1 port map( A => n3750, B => n4600, S => n4543, Z => n3074);
   U3217 : MUX2_X1 port map( A => n3755, B => n4601, S => n4543, Z => n3073);
   U3218 : MUX2_X1 port map( A => n3760, B => n4602, S => n4543, Z => n3072);
   U3219 : MUX2_X1 port map( A => n3765, B => n4603, S => n4543, Z => n3071);
   U3220 : MUX2_X1 port map( A => n3770, B => n4604, S => n4543, Z => n3070);
   U3221 : OAI21_X1 port map( B1 => n4606, B2 => n4635, A => n4607, ZN => n4634
                           );
   U3222 : MUX2_X1 port map( A => n3999, B => n4572, S => n4537, Z => n3069);
   U3223 : MUX2_X1 port map( A => n4004, B => n4574, S => n4537, Z => n3068);
   U3224 : MUX2_X1 port map( A => n4009, B => n4575, S => n4537, Z => n3067);
   U3225 : MUX2_X1 port map( A => n4014, B => n4576, S => n4537, Z => n3066);
   U3226 : MUX2_X1 port map( A => n4019, B => n4577, S => n4537, Z => n3065);
   U3227 : MUX2_X1 port map( A => n4024, B => n4578, S => n4537, Z => n3064);
   U3228 : MUX2_X1 port map( A => n4029, B => n4579, S => n4537, Z => n3063);
   U3229 : MUX2_X1 port map( A => n4034, B => n4580, S => n4537, Z => n3062);
   U3230 : MUX2_X1 port map( A => n4039, B => n4581, S => n4537, Z => n3061);
   U3231 : MUX2_X1 port map( A => n4044, B => n4582, S => n4537, Z => n3060);
   U3232 : MUX2_X1 port map( A => n4049, B => n4583, S => n4537, Z => n3059);
   U3233 : MUX2_X1 port map( A => n4054, B => n4584, S => n4537, Z => n3058);
   U3234 : MUX2_X1 port map( A => n4059, B => n4585, S => n4537, Z => n3057);
   U3235 : MUX2_X1 port map( A => n4064, B => n4586, S => n4537, Z => n3056);
   U3236 : MUX2_X1 port map( A => n4069, B => n4587, S => n4537, Z => n3055);
   U3237 : MUX2_X1 port map( A => n4074, B => n4588, S => n4537, Z => n3054);
   U3238 : MUX2_X1 port map( A => n4079, B => n4589, S => n4537, Z => n3053);
   U3239 : MUX2_X1 port map( A => n4084, B => n4590, S => n4537, Z => n3052);
   U3240 : MUX2_X1 port map( A => n4089, B => n4591, S => n4537, Z => n3051);
   U3241 : MUX2_X1 port map( A => n4094, B => n4592, S => n4537, Z => n3050);
   U3242 : MUX2_X1 port map( A => n4099, B => n4593, S => n4537, Z => n3049);
   U3243 : MUX2_X1 port map( A => n4104, B => n4594, S => n4537, Z => n3048);
   U3244 : MUX2_X1 port map( A => n4109, B => n4595, S => n4537, Z => n3047);
   U3245 : MUX2_X1 port map( A => n4114, B => n4596, S => n4537, Z => n3046);
   U3246 : MUX2_X1 port map( A => n4119, B => n4597, S => n4537, Z => n3045);
   U3247 : MUX2_X1 port map( A => n4124, B => n4598, S => n4537, Z => n3044);
   U3248 : MUX2_X1 port map( A => n4129, B => n4599, S => n4537, Z => n3043);
   U3249 : MUX2_X1 port map( A => n4134, B => n4600, S => n4537, Z => n3042);
   U3250 : MUX2_X1 port map( A => n4139, B => n4601, S => n4537, Z => n3041);
   U3251 : MUX2_X1 port map( A => n4144, B => n4602, S => n4537, Z => n3040);
   U3252 : MUX2_X1 port map( A => n4149, B => n4603, S => n4537, Z => n3039);
   U3253 : MUX2_X1 port map( A => n4154, B => n4604, S => n4537, Z => n3038);
   U3254 : OAI21_X1 port map( B1 => n4609, B2 => n4635, A => n4607, ZN => n4636
                           );
   U3255 : MUX2_X1 port map( A => n6354, B => n4572, S => n4539, Z => n3037);
   U3256 : MUX2_X1 port map( A => n6353, B => n4574, S => n4539, Z => n3036);
   U3257 : MUX2_X1 port map( A => n6352, B => n4575, S => n4539, Z => n3035);
   U3258 : MUX2_X1 port map( A => n6351, B => n4576, S => n4539, Z => n3034);
   U3259 : MUX2_X1 port map( A => n6350, B => n4577, S => n4539, Z => n3033);
   U3260 : MUX2_X1 port map( A => n6349, B => n4578, S => n4539, Z => n3032);
   U3261 : MUX2_X1 port map( A => n6348, B => n4579, S => n4539, Z => n3031);
   U3262 : MUX2_X1 port map( A => n6347, B => n4580, S => n4539, Z => n3030);
   U3263 : MUX2_X1 port map( A => n6346, B => n4581, S => n4539, Z => n3029);
   U3264 : MUX2_X1 port map( A => n6345, B => n4582, S => n4539, Z => n3028);
   U3265 : MUX2_X1 port map( A => n6344, B => n4583, S => n4539, Z => n3027);
   U3266 : MUX2_X1 port map( A => n6343, B => n4584, S => n4539, Z => n3026);
   U3267 : MUX2_X1 port map( A => n6342, B => n4585, S => n4539, Z => n3025);
   U3268 : MUX2_X1 port map( A => n6341, B => n4586, S => n4539, Z => n3024);
   U3269 : MUX2_X1 port map( A => n6340, B => n4587, S => n4539, Z => n3023);
   U3270 : MUX2_X1 port map( A => n6339, B => n4588, S => n4539, Z => n3022);
   U3271 : MUX2_X1 port map( A => n6338, B => n4589, S => n4539, Z => n3021);
   U3272 : MUX2_X1 port map( A => n6337, B => n4590, S => n4539, Z => n3020);
   U3273 : MUX2_X1 port map( A => n6336, B => n4591, S => n4539, Z => n3019);
   U3274 : MUX2_X1 port map( A => n6335, B => n4592, S => n4539, Z => n3018);
   U3275 : MUX2_X1 port map( A => n6334, B => n4593, S => n4539, Z => n3017);
   U3276 : MUX2_X1 port map( A => n6333, B => n4594, S => n4539, Z => n3016);
   U3277 : MUX2_X1 port map( A => n6332, B => n4595, S => n4539, Z => n3015);
   U3278 : MUX2_X1 port map( A => n6331, B => n4596, S => n4539, Z => n3014);
   U3279 : MUX2_X1 port map( A => n6330, B => n4597, S => n4539, Z => n3013);
   U3280 : MUX2_X1 port map( A => n6329, B => n4598, S => n4539, Z => n3012);
   U3281 : MUX2_X1 port map( A => n6328, B => n4599, S => n4539, Z => n3011);
   U3282 : MUX2_X1 port map( A => n6327, B => n4600, S => n4539, Z => n3010);
   U3283 : MUX2_X1 port map( A => n6326, B => n4601, S => n4539, Z => n3009);
   U3284 : MUX2_X1 port map( A => n6325, B => n4602, S => n4539, Z => n3008);
   U3285 : MUX2_X1 port map( A => n6324, B => n4603, S => n4539, Z => n3007);
   U3286 : MUX2_X1 port map( A => n6323, B => n4604, S => n4539, Z => n3006);
   U3287 : OAI21_X1 port map( B1 => n4611, B2 => n4635, A => n4607, ZN => n4637
                           );
   U3288 : MUX2_X1 port map( A => n6322, B => n4572, S => n4533, Z => n3005);
   U3289 : MUX2_X1 port map( A => n6321, B => n4574, S => n4533, Z => n3004);
   U3290 : MUX2_X1 port map( A => n6320, B => n4575, S => n4533, Z => n3003);
   U3291 : MUX2_X1 port map( A => n6319, B => n4576, S => n4533, Z => n3002);
   U3292 : MUX2_X1 port map( A => n6318, B => n4577, S => n4533, Z => n3001);
   U3293 : MUX2_X1 port map( A => n6317, B => n4578, S => n4533, Z => n3000);
   U3294 : MUX2_X1 port map( A => n6316, B => n4579, S => n4533, Z => n2999);
   U3295 : MUX2_X1 port map( A => n6315, B => n4580, S => n4533, Z => n2998);
   U3296 : MUX2_X1 port map( A => n6314, B => n4581, S => n4533, Z => n2997);
   U3297 : MUX2_X1 port map( A => n6313, B => n4582, S => n4533, Z => n2996);
   U3298 : MUX2_X1 port map( A => n6312, B => n4583, S => n4533, Z => n2995);
   U3299 : MUX2_X1 port map( A => n6311, B => n4584, S => n4533, Z => n2994);
   U3300 : MUX2_X1 port map( A => n6310, B => n4585, S => n4533, Z => n2993);
   U3301 : MUX2_X1 port map( A => n6309, B => n4586, S => n4533, Z => n2992);
   U3302 : MUX2_X1 port map( A => n6308, B => n4587, S => n4533, Z => n2991);
   U3303 : MUX2_X1 port map( A => n6307, B => n4588, S => n4533, Z => n2990);
   U3304 : MUX2_X1 port map( A => n6306, B => n4589, S => n4533, Z => n2989);
   U3305 : MUX2_X1 port map( A => n6305, B => n4590, S => n4533, Z => n2988);
   U3306 : MUX2_X1 port map( A => n6304, B => n4591, S => n4533, Z => n2987);
   U3307 : MUX2_X1 port map( A => n6303, B => n4592, S => n4533, Z => n2986);
   U3308 : MUX2_X1 port map( A => n6302, B => n4593, S => n4533, Z => n2985);
   U3309 : MUX2_X1 port map( A => n6301, B => n4594, S => n4533, Z => n2984);
   U3310 : MUX2_X1 port map( A => n6300, B => n4595, S => n4533, Z => n2983);
   U3311 : MUX2_X1 port map( A => n6299, B => n4596, S => n4533, Z => n2982);
   U3312 : MUX2_X1 port map( A => n6298, B => n4597, S => n4533, Z => n2981);
   U3313 : MUX2_X1 port map( A => n6297, B => n4598, S => n4533, Z => n2980);
   U3314 : MUX2_X1 port map( A => n6296, B => n4599, S => n4533, Z => n2979);
   U3315 : MUX2_X1 port map( A => n6295, B => n4600, S => n4533, Z => n2978);
   U3316 : MUX2_X1 port map( A => n6294, B => n4601, S => n4533, Z => n2977);
   U3317 : MUX2_X1 port map( A => n6293, B => n4602, S => n4533, Z => n2976);
   U3318 : MUX2_X1 port map( A => n6292, B => n4603, S => n4533, Z => n2975);
   U3319 : MUX2_X1 port map( A => n6291, B => n4604, S => n4533, Z => n2974);
   U3320 : OAI21_X1 port map( B1 => n4613, B2 => n4635, A => n4607, ZN => n4638
                           );
   U3321 : MUX2_X1 port map( A => n3616, B => n4572, S => n4535, Z => n2973);
   U3322 : MUX2_X1 port map( A => n3621, B => n4574, S => n4535, Z => n2972);
   U3323 : MUX2_X1 port map( A => n3626, B => n4575, S => n4535, Z => n2971);
   U3324 : MUX2_X1 port map( A => n3631, B => n4576, S => n4535, Z => n2970);
   U3325 : MUX2_X1 port map( A => n3636, B => n4577, S => n4535, Z => n2969);
   U3326 : MUX2_X1 port map( A => n3641, B => n4578, S => n4535, Z => n2968);
   U3327 : MUX2_X1 port map( A => n3646, B => n4579, S => n4535, Z => n2967);
   U3328 : MUX2_X1 port map( A => n3651, B => n4580, S => n4535, Z => n2966);
   U3329 : MUX2_X1 port map( A => n3656, B => n4581, S => n4535, Z => n2965);
   U3330 : MUX2_X1 port map( A => n3661, B => n4582, S => n4535, Z => n2964);
   U3331 : MUX2_X1 port map( A => n3666, B => n4583, S => n4535, Z => n2963);
   U3332 : MUX2_X1 port map( A => n3671, B => n4584, S => n4535, Z => n2962);
   U3333 : MUX2_X1 port map( A => n3676, B => n4585, S => n4535, Z => n2961);
   U3334 : MUX2_X1 port map( A => n3681, B => n4586, S => n4535, Z => n2960);
   U3335 : MUX2_X1 port map( A => n3686, B => n4587, S => n4535, Z => n2959);
   U3336 : MUX2_X1 port map( A => n3691, B => n4588, S => n4535, Z => n2958);
   U3337 : MUX2_X1 port map( A => n3696, B => n4589, S => n4535, Z => n2957);
   U3338 : MUX2_X1 port map( A => n3701, B => n4590, S => n4535, Z => n2956);
   U3339 : MUX2_X1 port map( A => n3706, B => n4591, S => n4535, Z => n2955);
   U3340 : MUX2_X1 port map( A => n3711, B => n4592, S => n4535, Z => n2954);
   U3341 : MUX2_X1 port map( A => n3716, B => n4593, S => n4535, Z => n2953);
   U3342 : MUX2_X1 port map( A => n3721, B => n4594, S => n4535, Z => n2952);
   U3343 : MUX2_X1 port map( A => n3726, B => n4595, S => n4535, Z => n2951);
   U3344 : MUX2_X1 port map( A => n3731, B => n4596, S => n4535, Z => n2950);
   U3345 : MUX2_X1 port map( A => n3736, B => n4597, S => n4535, Z => n2949);
   U3346 : MUX2_X1 port map( A => n3741, B => n4598, S => n4535, Z => n2948);
   U3347 : MUX2_X1 port map( A => n3746, B => n4599, S => n4535, Z => n2947);
   U3348 : MUX2_X1 port map( A => n3751, B => n4600, S => n4535, Z => n2946);
   U3349 : MUX2_X1 port map( A => n3756, B => n4601, S => n4535, Z => n2945);
   U3350 : MUX2_X1 port map( A => n3761, B => n4602, S => n4535, Z => n2944);
   U3351 : MUX2_X1 port map( A => n3766, B => n4603, S => n4535, Z => n2943);
   U3352 : MUX2_X1 port map( A => n3771, B => n4604, S => n4535, Z => n2942);
   U3353 : OAI21_X1 port map( B1 => n4615, B2 => n4635, A => n4607, ZN => n4639
                           );
   U3354 : MUX2_X1 port map( A => n4000, B => n4572, S => n4529, Z => n2941);
   U3355 : MUX2_X1 port map( A => n4005, B => n4574, S => n4529, Z => n2940);
   U3356 : MUX2_X1 port map( A => n4010, B => n4575, S => n4529, Z => n2939);
   U3357 : MUX2_X1 port map( A => n4015, B => n4576, S => n4529, Z => n2938);
   U3358 : MUX2_X1 port map( A => n4020, B => n4577, S => n4529, Z => n2937);
   U3359 : MUX2_X1 port map( A => n4025, B => n4578, S => n4529, Z => n2936);
   U3360 : MUX2_X1 port map( A => n4030, B => n4579, S => n4529, Z => n2935);
   U3361 : MUX2_X1 port map( A => n4035, B => n4580, S => n4529, Z => n2934);
   U3362 : MUX2_X1 port map( A => n4040, B => n4581, S => n4529, Z => n2933);
   U3363 : MUX2_X1 port map( A => n4045, B => n4582, S => n4529, Z => n2932);
   U3364 : MUX2_X1 port map( A => n4050, B => n4583, S => n4529, Z => n2931);
   U3365 : MUX2_X1 port map( A => n4055, B => n4584, S => n4529, Z => n2930);
   U3366 : MUX2_X1 port map( A => n4060, B => n4585, S => n4529, Z => n2929);
   U3367 : MUX2_X1 port map( A => n4065, B => n4586, S => n4529, Z => n2928);
   U3368 : MUX2_X1 port map( A => n4070, B => n4587, S => n4529, Z => n2927);
   U3369 : MUX2_X1 port map( A => n4075, B => n4588, S => n4529, Z => n2926);
   U3370 : MUX2_X1 port map( A => n4080, B => n4589, S => n4529, Z => n2925);
   U3371 : MUX2_X1 port map( A => n4085, B => n4590, S => n4529, Z => n2924);
   U3372 : MUX2_X1 port map( A => n4090, B => n4591, S => n4529, Z => n2923);
   U3373 : MUX2_X1 port map( A => n4095, B => n4592, S => n4529, Z => n2922);
   U3374 : MUX2_X1 port map( A => n4100, B => n4593, S => n4529, Z => n2921);
   U3375 : MUX2_X1 port map( A => n4105, B => n4594, S => n4529, Z => n2920);
   U3376 : MUX2_X1 port map( A => n4110, B => n4595, S => n4529, Z => n2919);
   U3377 : MUX2_X1 port map( A => n4115, B => n4596, S => n4529, Z => n2918);
   U3378 : MUX2_X1 port map( A => n4120, B => n4597, S => n4529, Z => n2917);
   U3379 : MUX2_X1 port map( A => n4125, B => n4598, S => n4529, Z => n2916);
   U3380 : MUX2_X1 port map( A => n4130, B => n4599, S => n4529, Z => n2915);
   U3381 : MUX2_X1 port map( A => n4135, B => n4600, S => n4529, Z => n2914);
   U3382 : MUX2_X1 port map( A => n4140, B => n4601, S => n4529, Z => n2913);
   U3383 : MUX2_X1 port map( A => n4145, B => n4602, S => n4529, Z => n2912);
   U3384 : MUX2_X1 port map( A => n4150, B => n4603, S => n4529, Z => n2911);
   U3385 : MUX2_X1 port map( A => n4155, B => n4604, S => n4529, Z => n2910);
   U3386 : OAI21_X1 port map( B1 => n4617, B2 => n4635, A => n4607, ZN => n4640
                           );
   U3387 : MUX2_X1 port map( A => n6290, B => n4572, S => n4531, Z => n2909);
   U3388 : MUX2_X1 port map( A => n6289, B => n4574, S => n4531, Z => n2908);
   U3389 : MUX2_X1 port map( A => n6288, B => n4575, S => n4531, Z => n2907);
   U3390 : MUX2_X1 port map( A => n6287, B => n4576, S => n4531, Z => n2906);
   U3391 : MUX2_X1 port map( A => n6286, B => n4577, S => n4531, Z => n2905);
   U3392 : MUX2_X1 port map( A => n6285, B => n4578, S => n4531, Z => n2904);
   U3393 : MUX2_X1 port map( A => n6284, B => n4579, S => n4531, Z => n2903);
   U3394 : MUX2_X1 port map( A => n6283, B => n4580, S => n4531, Z => n2902);
   U3395 : MUX2_X1 port map( A => n6282, B => n4581, S => n4531, Z => n2901);
   U3396 : MUX2_X1 port map( A => n6281, B => n4582, S => n4531, Z => n2900);
   U3397 : MUX2_X1 port map( A => n6280, B => n4583, S => n4531, Z => n2899);
   U3398 : MUX2_X1 port map( A => n6279, B => n4584, S => n4531, Z => n2898);
   U3399 : MUX2_X1 port map( A => n6278, B => n4585, S => n4531, Z => n2897);
   U3400 : MUX2_X1 port map( A => n6277, B => n4586, S => n4531, Z => n2896);
   U3401 : MUX2_X1 port map( A => n6276, B => n4587, S => n4531, Z => n2895);
   U3402 : MUX2_X1 port map( A => n6275, B => n4588, S => n4531, Z => n2894);
   U3403 : MUX2_X1 port map( A => n6274, B => n4589, S => n4531, Z => n2893);
   U3404 : MUX2_X1 port map( A => n6273, B => n4590, S => n4531, Z => n2892);
   U3405 : MUX2_X1 port map( A => n6272, B => n4591, S => n4531, Z => n2891);
   U3406 : MUX2_X1 port map( A => n6271, B => n4592, S => n4531, Z => n2890);
   U3407 : MUX2_X1 port map( A => n6270, B => n4593, S => n4531, Z => n2889);
   U3408 : MUX2_X1 port map( A => n6269, B => n4594, S => n4531, Z => n2888);
   U3409 : MUX2_X1 port map( A => n6268, B => n4595, S => n4531, Z => n2887);
   U3410 : MUX2_X1 port map( A => n6267, B => n4596, S => n4531, Z => n2886);
   U3411 : MUX2_X1 port map( A => n6266, B => n4597, S => n4531, Z => n2885);
   U3412 : MUX2_X1 port map( A => n6265, B => n4598, S => n4531, Z => n2884);
   U3413 : MUX2_X1 port map( A => n6264, B => n4599, S => n4531, Z => n2883);
   U3414 : MUX2_X1 port map( A => n6263, B => n4600, S => n4531, Z => n2882);
   U3415 : MUX2_X1 port map( A => n6262, B => n4601, S => n4531, Z => n2881);
   U3416 : MUX2_X1 port map( A => n6261, B => n4602, S => n4531, Z => n2880);
   U3417 : MUX2_X1 port map( A => n6260, B => n4603, S => n4531, Z => n2879);
   U3418 : MUX2_X1 port map( A => n6259, B => n4604, S => n4531, Z => n2878);
   U3419 : OAI21_X1 port map( B1 => n4619, B2 => n4635, A => n4607, ZN => n4641
                           );
   U3420 : MUX2_X1 port map( A => n6258, B => n4572, S => n4511, Z => n2877);
   U3421 : MUX2_X1 port map( A => n6257, B => n4574, S => n4511, Z => n2876);
   U3422 : MUX2_X1 port map( A => n6256, B => n4575, S => n4511, Z => n2875);
   U3423 : MUX2_X1 port map( A => n6255, B => n4576, S => n4511, Z => n2874);
   U3424 : MUX2_X1 port map( A => n6254, B => n4577, S => n4511, Z => n2873);
   U3425 : MUX2_X1 port map( A => n6253, B => n4578, S => n4511, Z => n2872);
   U3426 : MUX2_X1 port map( A => n6252, B => n4579, S => n4511, Z => n2871);
   U3427 : MUX2_X1 port map( A => n6251, B => n4580, S => n4511, Z => n2870);
   U3428 : MUX2_X1 port map( A => n6250, B => n4581, S => n4511, Z => n2869);
   U3429 : MUX2_X1 port map( A => n6249, B => n4582, S => n4511, Z => n2868);
   U3430 : MUX2_X1 port map( A => n6248, B => n4583, S => n4511, Z => n2867);
   U3431 : MUX2_X1 port map( A => n6247, B => n4584, S => n4511, Z => n2866);
   U3432 : MUX2_X1 port map( A => n6246, B => n4585, S => n4511, Z => n2865);
   U3433 : MUX2_X1 port map( A => n6245, B => n4586, S => n4511, Z => n2864);
   U3434 : MUX2_X1 port map( A => n6244, B => n4587, S => n4511, Z => n2863);
   U3435 : MUX2_X1 port map( A => n6243, B => n4588, S => n4511, Z => n2862);
   U3436 : MUX2_X1 port map( A => n6242, B => n4589, S => n4511, Z => n2861);
   U3437 : MUX2_X1 port map( A => n6241, B => n4590, S => n4511, Z => n2860);
   U3438 : MUX2_X1 port map( A => n6240, B => n4591, S => n4511, Z => n2859);
   U3439 : MUX2_X1 port map( A => n6239, B => n4592, S => n4511, Z => n2858);
   U3440 : MUX2_X1 port map( A => n6238, B => n4593, S => n4511, Z => n2857);
   U3441 : MUX2_X1 port map( A => n6237, B => n4594, S => n4511, Z => n2856);
   U3442 : MUX2_X1 port map( A => n6236, B => n4595, S => n4511, Z => n2855);
   U3443 : MUX2_X1 port map( A => n6235, B => n4596, S => n4511, Z => n2854);
   U3444 : MUX2_X1 port map( A => n6234, B => n4597, S => n4511, Z => n2853);
   U3445 : MUX2_X1 port map( A => n6233, B => n4598, S => n4511, Z => n2852);
   U3446 : MUX2_X1 port map( A => n6232, B => n4599, S => n4511, Z => n2851);
   U3447 : MUX2_X1 port map( A => n6231, B => n4600, S => n4511, Z => n2850);
   U3448 : MUX2_X1 port map( A => n6230, B => n4601, S => n4511, Z => n2849);
   U3449 : MUX2_X1 port map( A => n6229, B => n4602, S => n4511, Z => n2848);
   U3450 : MUX2_X1 port map( A => n6228, B => n4603, S => n4511, Z => n2847);
   U3451 : MUX2_X1 port map( A => n6227, B => n4604, S => n4511, Z => n2846);
   U3452 : OAI21_X1 port map( B1 => n4621, B2 => n4635, A => n4607, ZN => n4642
                           );
   U3453 : NAND3_X1 port map( A1 => n4624, A2 => n4622, A3 => ADD_WR(4), ZN => 
                           n4635);
   U3454 : INV_X1 port map( A => ADD_WR(3), ZN => n4622);
   U3455 : MUX2_X1 port map( A => n6226, B => n4572, S => n4513, Z => n2845);
   U3456 : MUX2_X1 port map( A => n6225, B => n4574, S => n4513, Z => n2844);
   U3457 : MUX2_X1 port map( A => n6224, B => n4575, S => n4513, Z => n2843);
   U3458 : MUX2_X1 port map( A => n6223, B => n4576, S => n4513, Z => n2842);
   U3459 : MUX2_X1 port map( A => n6222, B => n4577, S => n4513, Z => n2841);
   U3460 : MUX2_X1 port map( A => n6221, B => n4578, S => n4513, Z => n2840);
   U3461 : MUX2_X1 port map( A => n6220, B => n4579, S => n4513, Z => n2839);
   U3462 : MUX2_X1 port map( A => n6219, B => n4580, S => n4513, Z => n2838);
   U3463 : MUX2_X1 port map( A => n6218, B => n4581, S => n4513, Z => n2837);
   U3464 : MUX2_X1 port map( A => n6217, B => n4582, S => n4513, Z => n2836);
   U3465 : MUX2_X1 port map( A => n6216, B => n4583, S => n4513, Z => n2835);
   U3466 : MUX2_X1 port map( A => n6215, B => n4584, S => n4513, Z => n2834);
   U3467 : MUX2_X1 port map( A => n6214, B => n4585, S => n4513, Z => n2833);
   U3468 : MUX2_X1 port map( A => n6213, B => n4586, S => n4513, Z => n2832);
   U3469 : MUX2_X1 port map( A => n6212, B => n4587, S => n4513, Z => n2831);
   U3470 : MUX2_X1 port map( A => n6211, B => n4588, S => n4513, Z => n2830);
   U3471 : MUX2_X1 port map( A => n6210, B => n4589, S => n4513, Z => n2829);
   U3472 : MUX2_X1 port map( A => n6209, B => n4590, S => n4513, Z => n2828);
   U3473 : MUX2_X1 port map( A => n6208, B => n4591, S => n4513, Z => n2827);
   U3474 : MUX2_X1 port map( A => n6207, B => n4592, S => n4513, Z => n2826);
   U3475 : MUX2_X1 port map( A => n6206, B => n4593, S => n4513, Z => n2825);
   U3476 : MUX2_X1 port map( A => n6205, B => n4594, S => n4513, Z => n2824);
   U3477 : MUX2_X1 port map( A => n6204, B => n4595, S => n4513, Z => n2823);
   U3478 : MUX2_X1 port map( A => n6203, B => n4596, S => n4513, Z => n2822);
   U3479 : MUX2_X1 port map( A => n6202, B => n4597, S => n4513, Z => n2821);
   U3480 : MUX2_X1 port map( A => n6201, B => n4598, S => n4513, Z => n2820);
   U3481 : MUX2_X1 port map( A => n6200, B => n4599, S => n4513, Z => n2819);
   U3482 : MUX2_X1 port map( A => n6199, B => n4600, S => n4513, Z => n2818);
   U3483 : MUX2_X1 port map( A => n6198, B => n4601, S => n4513, Z => n2817);
   U3484 : MUX2_X1 port map( A => n6197, B => n4602, S => n4513, Z => n2816);
   U3485 : MUX2_X1 port map( A => n6196, B => n4603, S => n4513, Z => n2815);
   U3486 : MUX2_X1 port map( A => n6195, B => n4604, S => n4513, Z => n2814);
   U3487 : OAI21_X1 port map( B1 => n4606, B2 => n4644, A => n4607, ZN => n4643
                           );
   U3488 : NAND3_X1 port map( A1 => n4645, A2 => n4646, A3 => n4647, ZN => 
                           n4606);
   U3489 : MUX2_X1 port map( A => n6194, B => n4572, S => n4515, Z => n2813);
   U3490 : MUX2_X1 port map( A => n6193, B => n4574, S => n4515, Z => n2812);
   U3491 : MUX2_X1 port map( A => n6192, B => n4575, S => n4515, Z => n2811);
   U3492 : MUX2_X1 port map( A => n6191, B => n4576, S => n4515, Z => n2810);
   U3493 : MUX2_X1 port map( A => n6190, B => n4577, S => n4515, Z => n2809);
   U3494 : MUX2_X1 port map( A => n6189, B => n4578, S => n4515, Z => n2808);
   U3495 : MUX2_X1 port map( A => n6188, B => n4579, S => n4515, Z => n2807);
   U3496 : MUX2_X1 port map( A => n6187, B => n4580, S => n4515, Z => n2806);
   U3497 : MUX2_X1 port map( A => n6186, B => n4581, S => n4515, Z => n2805);
   U3498 : MUX2_X1 port map( A => n6185, B => n4582, S => n4515, Z => n2804);
   U3499 : MUX2_X1 port map( A => n6184, B => n4583, S => n4515, Z => n2803);
   U3500 : MUX2_X1 port map( A => n6183, B => n4584, S => n4515, Z => n2802);
   U3501 : MUX2_X1 port map( A => n6182, B => n4585, S => n4515, Z => n2801);
   U3502 : MUX2_X1 port map( A => n6181, B => n4586, S => n4515, Z => n2800);
   U3503 : MUX2_X1 port map( A => n6180, B => n4587, S => n4515, Z => n2799);
   U3504 : MUX2_X1 port map( A => n6179, B => n4588, S => n4515, Z => n2798);
   U3505 : MUX2_X1 port map( A => n6178, B => n4589, S => n4515, Z => n2797);
   U3506 : MUX2_X1 port map( A => n6177, B => n4590, S => n4515, Z => n2796);
   U3507 : MUX2_X1 port map( A => n6176, B => n4591, S => n4515, Z => n2795);
   U3508 : MUX2_X1 port map( A => n6175, B => n4592, S => n4515, Z => n2794);
   U3509 : MUX2_X1 port map( A => n6174, B => n4593, S => n4515, Z => n2793);
   U3510 : MUX2_X1 port map( A => n6173, B => n4594, S => n4515, Z => n2792);
   U3511 : MUX2_X1 port map( A => n6172, B => n4595, S => n4515, Z => n2791);
   U3512 : MUX2_X1 port map( A => n6171, B => n4596, S => n4515, Z => n2790);
   U3513 : MUX2_X1 port map( A => n6170, B => n4597, S => n4515, Z => n2789);
   U3514 : MUX2_X1 port map( A => n6169, B => n4598, S => n4515, Z => n2788);
   U3515 : MUX2_X1 port map( A => n6168, B => n4599, S => n4515, Z => n2787);
   U3516 : MUX2_X1 port map( A => n6167, B => n4600, S => n4515, Z => n2786);
   U3517 : MUX2_X1 port map( A => n6166, B => n4601, S => n4515, Z => n2785);
   U3518 : MUX2_X1 port map( A => n6165, B => n4602, S => n4515, Z => n2784);
   U3519 : MUX2_X1 port map( A => n6164, B => n4603, S => n4515, Z => n2783);
   U3520 : MUX2_X1 port map( A => n6163, B => n4604, S => n4515, Z => n2782);
   U3521 : OAI21_X1 port map( B1 => n4609, B2 => n4644, A => n4607, ZN => n4648
                           );
   U3522 : NAND3_X1 port map( A1 => n4645, A2 => n4646, A3 => ADD_WR(0), ZN => 
                           n4609);
   U3523 : MUX2_X1 port map( A => n3617, B => n4572, S => n4517, Z => n2781);
   U3524 : MUX2_X1 port map( A => n3622, B => n4574, S => n4517, Z => n2780);
   U3525 : MUX2_X1 port map( A => n3627, B => n4575, S => n4517, Z => n2779);
   U3526 : MUX2_X1 port map( A => n3632, B => n4576, S => n4517, Z => n2778);
   U3527 : MUX2_X1 port map( A => n3637, B => n4577, S => n4517, Z => n2777);
   U3528 : MUX2_X1 port map( A => n3642, B => n4578, S => n4517, Z => n2776);
   U3529 : MUX2_X1 port map( A => n3647, B => n4579, S => n4517, Z => n2775);
   U3530 : MUX2_X1 port map( A => n3652, B => n4580, S => n4517, Z => n2774);
   U3531 : MUX2_X1 port map( A => n3657, B => n4581, S => n4517, Z => n2773);
   U3532 : MUX2_X1 port map( A => n3662, B => n4582, S => n4517, Z => n2772);
   U3533 : MUX2_X1 port map( A => n3667, B => n4583, S => n4517, Z => n2771);
   U3534 : MUX2_X1 port map( A => n3672, B => n4584, S => n4517, Z => n2770);
   U3535 : MUX2_X1 port map( A => n3677, B => n4585, S => n4517, Z => n2769);
   U3536 : MUX2_X1 port map( A => n3682, B => n4586, S => n4517, Z => n2768);
   U3537 : MUX2_X1 port map( A => n3687, B => n4587, S => n4517, Z => n2767);
   U3538 : MUX2_X1 port map( A => n3692, B => n4588, S => n4517, Z => n2766);
   U3539 : MUX2_X1 port map( A => n3697, B => n4589, S => n4517, Z => n2765);
   U3540 : MUX2_X1 port map( A => n3702, B => n4590, S => n4517, Z => n2764);
   U3541 : MUX2_X1 port map( A => n3707, B => n4591, S => n4517, Z => n2763);
   U3542 : MUX2_X1 port map( A => n3712, B => n4592, S => n4517, Z => n2762);
   U3543 : MUX2_X1 port map( A => n3717, B => n4593, S => n4517, Z => n2761);
   U3544 : MUX2_X1 port map( A => n3722, B => n4594, S => n4517, Z => n2760);
   U3545 : MUX2_X1 port map( A => n3727, B => n4595, S => n4517, Z => n2759);
   U3546 : MUX2_X1 port map( A => n3732, B => n4596, S => n4517, Z => n2758);
   U3547 : MUX2_X1 port map( A => n3737, B => n4597, S => n4517, Z => n2757);
   U3548 : MUX2_X1 port map( A => n3742, B => n4598, S => n4517, Z => n2756);
   U3549 : MUX2_X1 port map( A => n3747, B => n4599, S => n4517, Z => n2755);
   U3550 : MUX2_X1 port map( A => n3752, B => n4600, S => n4517, Z => n2754);
   U3551 : MUX2_X1 port map( A => n3757, B => n4601, S => n4517, Z => n2753);
   U3552 : MUX2_X1 port map( A => n3762, B => n4602, S => n4517, Z => n2752);
   U3553 : MUX2_X1 port map( A => n3767, B => n4603, S => n4517, Z => n2751);
   U3554 : MUX2_X1 port map( A => n3772, B => n4604, S => n4517, Z => n2750);
   U3555 : OAI21_X1 port map( B1 => n4611, B2 => n4644, A => n4607, ZN => n4649
                           );
   U3556 : NAND3_X1 port map( A1 => n4647, A2 => n4646, A3 => ADD_WR(1), ZN => 
                           n4611);
   U3557 : MUX2_X1 port map( A => n4001, B => n4572, S => n4519, Z => n2749);
   U3558 : MUX2_X1 port map( A => n4006, B => n4574, S => n4519, Z => n2748);
   U3559 : MUX2_X1 port map( A => n4011, B => n4575, S => n4519, Z => n2747);
   U3560 : MUX2_X1 port map( A => n4016, B => n4576, S => n4519, Z => n2746);
   U3561 : MUX2_X1 port map( A => n4021, B => n4577, S => n4519, Z => n2745);
   U3562 : MUX2_X1 port map( A => n4026, B => n4578, S => n4519, Z => n2744);
   U3563 : MUX2_X1 port map( A => n4031, B => n4579, S => n4519, Z => n2743);
   U3564 : MUX2_X1 port map( A => n4036, B => n4580, S => n4519, Z => n2742);
   U3565 : MUX2_X1 port map( A => n4041, B => n4581, S => n4519, Z => n2741);
   U3566 : MUX2_X1 port map( A => n4046, B => n4582, S => n4519, Z => n2740);
   U3567 : MUX2_X1 port map( A => n4051, B => n4583, S => n4519, Z => n2739);
   U3568 : MUX2_X1 port map( A => n4056, B => n4584, S => n4519, Z => n2738);
   U3569 : MUX2_X1 port map( A => n4061, B => n4585, S => n4519, Z => n2737);
   U3570 : MUX2_X1 port map( A => n4066, B => n4586, S => n4519, Z => n2736);
   U3571 : MUX2_X1 port map( A => n4071, B => n4587, S => n4519, Z => n2735);
   U3572 : MUX2_X1 port map( A => n4076, B => n4588, S => n4519, Z => n2734);
   U3573 : MUX2_X1 port map( A => n4081, B => n4589, S => n4519, Z => n2733);
   U3574 : MUX2_X1 port map( A => n4086, B => n4590, S => n4519, Z => n2732);
   U3575 : MUX2_X1 port map( A => n4091, B => n4591, S => n4519, Z => n2731);
   U3576 : MUX2_X1 port map( A => n4096, B => n4592, S => n4519, Z => n2730);
   U3577 : MUX2_X1 port map( A => n4101, B => n4593, S => n4519, Z => n2729);
   U3578 : MUX2_X1 port map( A => n4106, B => n4594, S => n4519, Z => n2728);
   U3579 : MUX2_X1 port map( A => n4111, B => n4595, S => n4519, Z => n2727);
   U3580 : MUX2_X1 port map( A => n4116, B => n4596, S => n4519, Z => n2726);
   U3581 : MUX2_X1 port map( A => n4121, B => n4597, S => n4519, Z => n2725);
   U3582 : MUX2_X1 port map( A => n4126, B => n4598, S => n4519, Z => n2724);
   U3583 : MUX2_X1 port map( A => n4131, B => n4599, S => n4519, Z => n2723);
   U3584 : MUX2_X1 port map( A => n4136, B => n4600, S => n4519, Z => n2722);
   U3585 : MUX2_X1 port map( A => n4141, B => n4601, S => n4519, Z => n2721);
   U3586 : MUX2_X1 port map( A => n4146, B => n4602, S => n4519, Z => n2720);
   U3587 : MUX2_X1 port map( A => n4151, B => n4603, S => n4519, Z => n2719);
   U3588 : MUX2_X1 port map( A => n4156, B => n4604, S => n4519, Z => n2718);
   U3589 : OAI21_X1 port map( B1 => n4613, B2 => n4644, A => n4607, ZN => n4650
                           );
   U3590 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n4646, A3 => ADD_WR(1), ZN
                           => n4613);
   U3591 : INV_X1 port map( A => ADD_WR(2), ZN => n4646);
   U3592 : MUX2_X1 port map( A => n6162, B => n4572, S => n4521, Z => n2717);
   U3593 : MUX2_X1 port map( A => n6161, B => n4574, S => n4521, Z => n2716);
   U3594 : MUX2_X1 port map( A => n6160, B => n4575, S => n4521, Z => n2715);
   U3595 : MUX2_X1 port map( A => n6159, B => n4576, S => n4521, Z => n2714);
   U3596 : MUX2_X1 port map( A => n6158, B => n4577, S => n4521, Z => n2713);
   U3597 : MUX2_X1 port map( A => n6157, B => n4578, S => n4521, Z => n2712);
   U3598 : MUX2_X1 port map( A => n6156, B => n4579, S => n4521, Z => n2711);
   U3599 : MUX2_X1 port map( A => n6155, B => n4580, S => n4521, Z => n2710);
   U3600 : MUX2_X1 port map( A => n6154, B => n4581, S => n4521, Z => n2709);
   U3601 : MUX2_X1 port map( A => n6153, B => n4582, S => n4521, Z => n2708);
   U3602 : MUX2_X1 port map( A => n6152, B => n4583, S => n4521, Z => n2707);
   U3603 : MUX2_X1 port map( A => n6151, B => n4584, S => n4521, Z => n2706);
   U3604 : MUX2_X1 port map( A => n6150, B => n4585, S => n4521, Z => n2705);
   U3605 : MUX2_X1 port map( A => n6149, B => n4586, S => n4521, Z => n2704);
   U3606 : MUX2_X1 port map( A => n6148, B => n4587, S => n4521, Z => n2703);
   U3607 : MUX2_X1 port map( A => n6147, B => n4588, S => n4521, Z => n2702);
   U3608 : MUX2_X1 port map( A => n6146, B => n4589, S => n4521, Z => n2701);
   U3609 : MUX2_X1 port map( A => n6145, B => n4590, S => n4521, Z => n2700);
   U3610 : MUX2_X1 port map( A => n6144, B => n4591, S => n4521, Z => n2699);
   U3611 : MUX2_X1 port map( A => n6143, B => n4592, S => n4521, Z => n2698);
   U3612 : MUX2_X1 port map( A => n6142, B => n4593, S => n4521, Z => n2697);
   U3613 : MUX2_X1 port map( A => n6141, B => n4594, S => n4521, Z => n2696);
   U3614 : MUX2_X1 port map( A => n6140, B => n4595, S => n4521, Z => n2695);
   U3615 : MUX2_X1 port map( A => n6139, B => n4596, S => n4521, Z => n2694);
   U3616 : MUX2_X1 port map( A => n6138, B => n4597, S => n4521, Z => n2693);
   U3617 : MUX2_X1 port map( A => n6137, B => n4598, S => n4521, Z => n2692);
   U3618 : MUX2_X1 port map( A => n6136, B => n4599, S => n4521, Z => n2691);
   U3619 : MUX2_X1 port map( A => n6135, B => n4600, S => n4521, Z => n2690);
   U3620 : MUX2_X1 port map( A => n6134, B => n4601, S => n4521, Z => n2689);
   U3621 : MUX2_X1 port map( A => n6133, B => n4602, S => n4521, Z => n2688);
   U3622 : MUX2_X1 port map( A => n6132, B => n4603, S => n4521, Z => n2687);
   U3623 : MUX2_X1 port map( A => n6131, B => n4604, S => n4521, Z => n2686);
   U3624 : OAI21_X1 port map( B1 => n4615, B2 => n4644, A => n4607, ZN => n4651
                           );
   U3625 : NAND3_X1 port map( A1 => n4647, A2 => n4645, A3 => ADD_WR(2), ZN => 
                           n4615);
   U3626 : MUX2_X1 port map( A => n6130, B => n4572, S => n4523, Z => n2685);
   U3627 : MUX2_X1 port map( A => n6129, B => n4574, S => n4523, Z => n2684);
   U3628 : MUX2_X1 port map( A => n6128, B => n4575, S => n4523, Z => n2683);
   U3629 : MUX2_X1 port map( A => n6127, B => n4576, S => n4523, Z => n2682);
   U3630 : MUX2_X1 port map( A => n6126, B => n4577, S => n4523, Z => n2681);
   U3631 : MUX2_X1 port map( A => n6125, B => n4578, S => n4523, Z => n2680);
   U3632 : MUX2_X1 port map( A => n6124, B => n4579, S => n4523, Z => n2679);
   U3633 : MUX2_X1 port map( A => n6123, B => n4580, S => n4523, Z => n2678);
   U3634 : MUX2_X1 port map( A => n6122, B => n4581, S => n4523, Z => n2677);
   U3635 : MUX2_X1 port map( A => n6121, B => n4582, S => n4523, Z => n2676);
   U3636 : MUX2_X1 port map( A => n6120, B => n4583, S => n4523, Z => n2675);
   U3637 : MUX2_X1 port map( A => n6119, B => n4584, S => n4523, Z => n2674);
   U3638 : MUX2_X1 port map( A => n6118, B => n4585, S => n4523, Z => n2673);
   U3639 : MUX2_X1 port map( A => n6117, B => n4586, S => n4523, Z => n2672);
   U3640 : MUX2_X1 port map( A => n6116, B => n4587, S => n4523, Z => n2671);
   U3641 : MUX2_X1 port map( A => n6115, B => n4588, S => n4523, Z => n2670);
   U3642 : MUX2_X1 port map( A => n6114, B => n4589, S => n4523, Z => n2669);
   U3643 : MUX2_X1 port map( A => n6113, B => n4590, S => n4523, Z => n2668);
   U3644 : MUX2_X1 port map( A => n6112, B => n4591, S => n4523, Z => n2667);
   U3645 : MUX2_X1 port map( A => n6111, B => n4592, S => n4523, Z => n2666);
   U3646 : MUX2_X1 port map( A => n6110, B => n4593, S => n4523, Z => n2665);
   U3647 : MUX2_X1 port map( A => n6109, B => n4594, S => n4523, Z => n2664);
   U3648 : MUX2_X1 port map( A => n6108, B => n4595, S => n4523, Z => n2663);
   U3649 : MUX2_X1 port map( A => n6107, B => n4596, S => n4523, Z => n2662);
   U3650 : MUX2_X1 port map( A => n6106, B => n4597, S => n4523, Z => n2661);
   U3651 : MUX2_X1 port map( A => n6105, B => n4598, S => n4523, Z => n2660);
   U3652 : MUX2_X1 port map( A => n6104, B => n4599, S => n4523, Z => n2659);
   U3653 : MUX2_X1 port map( A => n6103, B => n4600, S => n4523, Z => n2658);
   U3654 : MUX2_X1 port map( A => n6102, B => n4601, S => n4523, Z => n2657);
   U3655 : MUX2_X1 port map( A => n6101, B => n4602, S => n4523, Z => n2656);
   U3656 : MUX2_X1 port map( A => n6100, B => n4603, S => n4523, Z => n2655);
   U3657 : MUX2_X1 port map( A => n6099, B => n4604, S => n4523, Z => n2654);
   U3658 : OAI21_X1 port map( B1 => n4617, B2 => n4644, A => n4607, ZN => n4652
                           );
   U3659 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n4645, A3 => ADD_WR(2), ZN
                           => n4617);
   U3660 : INV_X1 port map( A => ADD_WR(1), ZN => n4645);
   U3661 : MUX2_X1 port map( A => n3618, B => n4572, S => n4525, Z => n2653);
   U3662 : MUX2_X1 port map( A => n3623, B => n4574, S => n4525, Z => n2652);
   U3663 : MUX2_X1 port map( A => n3628, B => n4575, S => n4525, Z => n2651);
   U3664 : MUX2_X1 port map( A => n3633, B => n4576, S => n4525, Z => n2650);
   U3665 : MUX2_X1 port map( A => n3638, B => n4577, S => n4525, Z => n2649);
   U3666 : MUX2_X1 port map( A => n3643, B => n4578, S => n4525, Z => n2648);
   U3667 : MUX2_X1 port map( A => n3648, B => n4579, S => n4525, Z => n2647);
   U3668 : MUX2_X1 port map( A => n3653, B => n4580, S => n4525, Z => n2646);
   U3669 : MUX2_X1 port map( A => n3658, B => n4581, S => n4525, Z => n2645);
   U3670 : MUX2_X1 port map( A => n3663, B => n4582, S => n4525, Z => n2644);
   U3671 : MUX2_X1 port map( A => n3668, B => n4583, S => n4525, Z => n2643);
   U3672 : MUX2_X1 port map( A => n3673, B => n4584, S => n4525, Z => n2642);
   U3673 : MUX2_X1 port map( A => n3678, B => n4585, S => n4525, Z => n2641);
   U3674 : MUX2_X1 port map( A => n3683, B => n4586, S => n4525, Z => n2640);
   U3675 : MUX2_X1 port map( A => n3688, B => n4587, S => n4525, Z => n2639);
   U3676 : MUX2_X1 port map( A => n3693, B => n4588, S => n4525, Z => n2638);
   U3677 : MUX2_X1 port map( A => n3698, B => n4589, S => n4525, Z => n2637);
   U3678 : MUX2_X1 port map( A => n3703, B => n4590, S => n4525, Z => n2636);
   U3679 : MUX2_X1 port map( A => n3708, B => n4591, S => n4525, Z => n2635);
   U3680 : MUX2_X1 port map( A => n3713, B => n4592, S => n4525, Z => n2634);
   U3681 : MUX2_X1 port map( A => n3718, B => n4593, S => n4525, Z => n2633);
   U3682 : MUX2_X1 port map( A => n3723, B => n4594, S => n4525, Z => n2632);
   U3683 : MUX2_X1 port map( A => n3728, B => n4595, S => n4525, Z => n2631);
   U3684 : MUX2_X1 port map( A => n3733, B => n4596, S => n4525, Z => n2630);
   U3685 : MUX2_X1 port map( A => n3738, B => n4597, S => n4525, Z => n2629);
   U3686 : MUX2_X1 port map( A => n3743, B => n4598, S => n4525, Z => n2628);
   U3687 : MUX2_X1 port map( A => n3748, B => n4599, S => n4525, Z => n2627);
   U3688 : MUX2_X1 port map( A => n3753, B => n4600, S => n4525, Z => n2626);
   U3689 : MUX2_X1 port map( A => n3758, B => n4601, S => n4525, Z => n2625);
   U3690 : MUX2_X1 port map( A => n3763, B => n4602, S => n4525, Z => n2624);
   U3691 : MUX2_X1 port map( A => n3768, B => n4603, S => n4525, Z => n2623);
   U3692 : MUX2_X1 port map( A => n3773, B => n4604, S => n4525, Z => n2622);
   U3693 : OAI21_X1 port map( B1 => n4619, B2 => n4644, A => n4607, ZN => n4653
                           );
   U3694 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => n4647, A3 => ADD_WR(2), ZN
                           => n4619);
   U3695 : INV_X1 port map( A => ADD_WR(0), ZN => n4647);
   U3696 : MUX2_X1 port map( A => n4002, B => n4572, S => n4527, Z => n2621);
   U3697 : AND2_X1 port map( A1 => DATAIN(31), A2 => n4607, ZN => n4572);
   U3698 : MUX2_X1 port map( A => n4007, B => n4574, S => n4527, Z => n2620);
   U3699 : AND2_X1 port map( A1 => DATAIN(30), A2 => n4607, ZN => n4574);
   U3700 : MUX2_X1 port map( A => n4012, B => n4575, S => n4527, Z => n2619);
   U3701 : AND2_X1 port map( A1 => DATAIN(29), A2 => n4607, ZN => n4575);
   U3702 : MUX2_X1 port map( A => n4017, B => n4576, S => n4527, Z => n2618);
   U3703 : AND2_X1 port map( A1 => DATAIN(28), A2 => n4607, ZN => n4576);
   U3704 : MUX2_X1 port map( A => n4022, B => n4577, S => n4527, Z => n2617);
   U3705 : AND2_X1 port map( A1 => DATAIN(27), A2 => n4607, ZN => n4577);
   U3706 : MUX2_X1 port map( A => n4027, B => n4578, S => n4527, Z => n2616);
   U3707 : AND2_X1 port map( A1 => DATAIN(26), A2 => n4607, ZN => n4578);
   U3708 : MUX2_X1 port map( A => n4032, B => n4579, S => n4527, Z => n2615);
   U3709 : AND2_X1 port map( A1 => DATAIN(25), A2 => n4607, ZN => n4579);
   U3710 : MUX2_X1 port map( A => n4037, B => n4580, S => n4527, Z => n2614);
   U3711 : AND2_X1 port map( A1 => DATAIN(24), A2 => n4607, ZN => n4580);
   U3712 : MUX2_X1 port map( A => n4042, B => n4581, S => n4527, Z => n2613);
   U3713 : AND2_X1 port map( A1 => DATAIN(23), A2 => n4607, ZN => n4581);
   U3714 : MUX2_X1 port map( A => n4047, B => n4582, S => n4527, Z => n2612);
   U3715 : AND2_X1 port map( A1 => DATAIN(22), A2 => n4607, ZN => n4582);
   U3716 : MUX2_X1 port map( A => n4052, B => n4583, S => n4527, Z => n2611);
   U3717 : AND2_X1 port map( A1 => DATAIN(21), A2 => n4607, ZN => n4583);
   U3718 : MUX2_X1 port map( A => n4057, B => n4584, S => n4527, Z => n2610);
   U3719 : AND2_X1 port map( A1 => DATAIN(20), A2 => n4607, ZN => n4584);
   U3720 : MUX2_X1 port map( A => n4062, B => n4585, S => n4527, Z => n2609);
   U3721 : AND2_X1 port map( A1 => DATAIN(19), A2 => n4607, ZN => n4585);
   U3722 : MUX2_X1 port map( A => n4067, B => n4586, S => n4527, Z => n2608);
   U3723 : AND2_X1 port map( A1 => DATAIN(18), A2 => n4607, ZN => n4586);
   U3724 : MUX2_X1 port map( A => n4072, B => n4587, S => n4527, Z => n2607);
   U3725 : AND2_X1 port map( A1 => DATAIN(17), A2 => n4607, ZN => n4587);
   U3726 : MUX2_X1 port map( A => n4077, B => n4588, S => n4527, Z => n2606);
   U3727 : AND2_X1 port map( A1 => DATAIN(16), A2 => n4607, ZN => n4588);
   U3728 : MUX2_X1 port map( A => n4082, B => n4589, S => n4527, Z => n2605);
   U3729 : AND2_X1 port map( A1 => DATAIN(15), A2 => n4607, ZN => n4589);
   U3730 : MUX2_X1 port map( A => n4087, B => n4590, S => n4527, Z => n2604);
   U3731 : AND2_X1 port map( A1 => DATAIN(14), A2 => n4607, ZN => n4590);
   U3732 : MUX2_X1 port map( A => n4092, B => n4591, S => n4527, Z => n2603);
   U3733 : AND2_X1 port map( A1 => DATAIN(13), A2 => n4607, ZN => n4591);
   U3734 : MUX2_X1 port map( A => n4097, B => n4592, S => n4527, Z => n2602);
   U3735 : AND2_X1 port map( A1 => DATAIN(12), A2 => n4607, ZN => n4592);
   U3736 : MUX2_X1 port map( A => n4102, B => n4593, S => n4527, Z => n2601);
   U3737 : AND2_X1 port map( A1 => DATAIN(11), A2 => n4607, ZN => n4593);
   U3738 : MUX2_X1 port map( A => n4107, B => n4594, S => n4527, Z => n2600);
   U3739 : AND2_X1 port map( A1 => DATAIN(10), A2 => n4607, ZN => n4594);
   U3740 : MUX2_X1 port map( A => n4112, B => n4595, S => n4527, Z => n2599);
   U3741 : AND2_X1 port map( A1 => DATAIN(9), A2 => n4607, ZN => n4595);
   U3742 : MUX2_X1 port map( A => n4117, B => n4596, S => n4527, Z => n2598);
   U3743 : AND2_X1 port map( A1 => DATAIN(8), A2 => n4607, ZN => n4596);
   U3744 : MUX2_X1 port map( A => n4122, B => n4597, S => n4527, Z => n2597);
   U3745 : AND2_X1 port map( A1 => DATAIN(7), A2 => n4607, ZN => n4597);
   U3746 : MUX2_X1 port map( A => n4127, B => n4598, S => n4527, Z => n2596);
   U3747 : AND2_X1 port map( A1 => DATAIN(6), A2 => n4607, ZN => n4598);
   U3748 : MUX2_X1 port map( A => n4132, B => n4599, S => n4527, Z => n2595);
   U3749 : AND2_X1 port map( A1 => DATAIN(5), A2 => n4607, ZN => n4599);
   U3750 : MUX2_X1 port map( A => n4137, B => n4600, S => n4527, Z => n2594);
   U3751 : AND2_X1 port map( A1 => DATAIN(4), A2 => n4607, ZN => n4600);
   U3752 : MUX2_X1 port map( A => n4142, B => n4601, S => n4527, Z => n2593);
   U3753 : AND2_X1 port map( A1 => DATAIN(3), A2 => n4607, ZN => n4601);
   U3754 : MUX2_X1 port map( A => n4147, B => n4602, S => n4527, Z => n2592);
   U3755 : AND2_X1 port map( A1 => DATAIN(2), A2 => n4607, ZN => n4602);
   U3756 : MUX2_X1 port map( A => n4152, B => n4603, S => n4527, Z => n2591);
   U3757 : AND2_X1 port map( A1 => DATAIN(1), A2 => n4607, ZN => n4603);
   U3758 : MUX2_X1 port map( A => n4157, B => n4604, S => n4527, Z => n2590);
   U3759 : OAI21_X1 port map( B1 => n4621, B2 => n4644, A => n4607, ZN => n4654
                           );
   U3760 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => n4624, A3 => ADD_WR(4), ZN
                           => n4644);
   U3761 : AND2_X1 port map( A1 => WR, A2 => ENABLE, ZN => n4624);
   U3762 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), A3 => ADD_WR(2)
                           , ZN => n4621);
   U3763 : AND2_X1 port map( A1 => DATAIN(0), A2 => n4607, ZN => n4604);
   U3764 : MUX2_X1 port map( A => OUT2_31_port, B => n4655, S => n4656, Z => 
                           n2589);
   U3765 : NAND2_X1 port map( A1 => n4657, A2 => n4658, ZN => n4655);
   U3766 : NOR4_X1 port map( A1 => n4659, A2 => n4660, A3 => n4661, A4 => n4662
                           , ZN => n4658);
   U3767 : OAI221_X1 port map( B1 => n1, B2 => n4663, C1 => n33, C2 => n4664, A
                           => n4665, ZN => n4662);
   U3768 : AOI22_X1 port map( A1 => n4666, A2 => n6097, B1 => n4667, B2 => 
                           n6098, ZN => n4665);
   U3769 : OAI221_X1 port map( B1 => n129, B2 => n4668, C1 => n161, C2 => n4669
                           , A => n4670, ZN => n4661);
   U3770 : AOI22_X1 port map( A1 => n4671, A2 => n6095, B1 => n4672, B2 => 
                           n6096, ZN => n4670);
   U3771 : OAI221_X1 port map( B1 => n353, B2 => n4673, C1 => n321, C2 => n4674
                           , A => n4675, ZN => n4660);
   U3772 : AOI22_X1 port map( A1 => n4676, A2 => n3934, B1 => n4677, B2 => 
                           n4318, ZN => n4675);
   U3773 : OAI221_X1 port map( B1 => n3774, B2 => n4678, C1 => n4158, C2 => 
                           n4679, A => n4680, ZN => n4659);
   U3774 : AOI22_X1 port map( A1 => n4681, A2 => n3614, B1 => n4682, B2 => 
                           n3998, ZN => n4680);
   U3775 : NOR4_X1 port map( A1 => n4683, A2 => n4684, A3 => n4685, A4 => n4686
                           , ZN => n4657);
   U3776 : OAI221_X1 port map( B1 => n3775, B2 => n4687, C1 => n4159, C2 => 
                           n4688, A => n4689, ZN => n4686);
   U3777 : AOI22_X1 port map( A1 => n4690, A2 => n3615, B1 => n4691, B2 => 
                           n3999, ZN => n4689);
   U3778 : OAI221_X1 port map( B1 => n3776, B2 => n4692, C1 => n4160, C2 => 
                           n4693, A => n4694, ZN => n4685);
   U3779 : AOI22_X1 port map( A1 => n4695, A2 => n3616, B1 => n4696, B2 => 
                           n4000, ZN => n4694);
   U3780 : OAI221_X1 port map( B1 => n3777, B2 => n4697, C1 => n4161, C2 => 
                           n4698, A => n4699, ZN => n4684);
   U3781 : AOI22_X1 port map( A1 => n4700, A2 => n3617, B1 => n4701, B2 => 
                           n4001, ZN => n4699);
   U3782 : OAI221_X1 port map( B1 => n3778, B2 => n4702, C1 => n4162, C2 => 
                           n4703, A => n4704, ZN => n4683);
   U3783 : AOI22_X1 port map( A1 => n4705, A2 => n3618, B1 => n4706, B2 => 
                           n4002, ZN => n4704);
   U3784 : MUX2_X1 port map( A => OUT2_30_port, B => n4707, S => n4656, Z => 
                           n2588);
   U3785 : NAND2_X1 port map( A1 => n4708, A2 => n4709, ZN => n4707);
   U3786 : NOR4_X1 port map( A1 => n4710, A2 => n4711, A3 => n4712, A4 => n4713
                           , ZN => n4709);
   U3787 : OAI221_X1 port map( B1 => n2, B2 => n4663, C1 => n34, C2 => n4664, A
                           => n4714, ZN => n4713);
   U3788 : AOI22_X1 port map( A1 => n4666, A2 => n6093, B1 => n4667, B2 => 
                           n6094, ZN => n4714);
   U3789 : OAI221_X1 port map( B1 => n130, B2 => n4668, C1 => n162, C2 => n4669
                           , A => n4715, ZN => n4712);
   U3790 : AOI22_X1 port map( A1 => n4671, A2 => n6091, B1 => n4672, B2 => 
                           n6092, ZN => n4715);
   U3791 : OAI221_X1 port map( B1 => n354, B2 => n4673, C1 => n322, C2 => n4674
                           , A => n4716, ZN => n4711);
   U3792 : AOI22_X1 port map( A1 => n4676, A2 => n3935, B1 => n4677, B2 => 
                           n4319, ZN => n4716);
   U3793 : OAI221_X1 port map( B1 => n3779, B2 => n4678, C1 => n4163, C2 => 
                           n4679, A => n4717, ZN => n4710);
   U3794 : AOI22_X1 port map( A1 => n4681, A2 => n3619, B1 => n4682, B2 => 
                           n4003, ZN => n4717);
   U3795 : NOR4_X1 port map( A1 => n4718, A2 => n4719, A3 => n4720, A4 => n4721
                           , ZN => n4708);
   U3796 : OAI221_X1 port map( B1 => n3780, B2 => n4687, C1 => n4164, C2 => 
                           n4688, A => n4722, ZN => n4721);
   U3797 : AOI22_X1 port map( A1 => n4690, A2 => n3620, B1 => n4691, B2 => 
                           n4004, ZN => n4722);
   U3798 : OAI221_X1 port map( B1 => n3781, B2 => n4692, C1 => n4165, C2 => 
                           n4693, A => n4723, ZN => n4720);
   U3799 : AOI22_X1 port map( A1 => n4695, A2 => n3621, B1 => n4696, B2 => 
                           n4005, ZN => n4723);
   U3800 : OAI221_X1 port map( B1 => n3782, B2 => n4697, C1 => n4166, C2 => 
                           n4698, A => n4724, ZN => n4719);
   U3801 : AOI22_X1 port map( A1 => n4700, A2 => n3622, B1 => n4701, B2 => 
                           n4006, ZN => n4724);
   U3802 : OAI221_X1 port map( B1 => n3783, B2 => n4702, C1 => n4167, C2 => 
                           n4703, A => n4725, ZN => n4718);
   U3803 : AOI22_X1 port map( A1 => n4705, A2 => n3623, B1 => n4706, B2 => 
                           n4007, ZN => n4725);
   U3804 : MUX2_X1 port map( A => OUT2_29_port, B => n4726, S => n4656, Z => 
                           n2587);
   U3805 : NAND2_X1 port map( A1 => n4727, A2 => n4728, ZN => n4726);
   U3806 : NOR4_X1 port map( A1 => n4729, A2 => n4730, A3 => n4731, A4 => n4732
                           , ZN => n4728);
   U3807 : OAI221_X1 port map( B1 => n3, B2 => n4663, C1 => n35, C2 => n4664, A
                           => n4733, ZN => n4732);
   U3808 : AOI22_X1 port map( A1 => n4666, A2 => n6089, B1 => n4667, B2 => 
                           n6090, ZN => n4733);
   U3809 : OAI221_X1 port map( B1 => n131, B2 => n4668, C1 => n163, C2 => n4669
                           , A => n4734, ZN => n4731);
   U3810 : AOI22_X1 port map( A1 => n4671, A2 => n6087, B1 => n4672, B2 => 
                           n6088, ZN => n4734);
   U3811 : OAI221_X1 port map( B1 => n355, B2 => n4673, C1 => n323, C2 => n4674
                           , A => n4735, ZN => n4730);
   U3812 : AOI22_X1 port map( A1 => n4676, A2 => n3936, B1 => n4677, B2 => 
                           n4320, ZN => n4735);
   U3813 : OAI221_X1 port map( B1 => n3784, B2 => n4678, C1 => n4168, C2 => 
                           n4679, A => n4736, ZN => n4729);
   U3814 : AOI22_X1 port map( A1 => n4681, A2 => n3624, B1 => n4682, B2 => 
                           n4008, ZN => n4736);
   U3815 : NOR4_X1 port map( A1 => n4737, A2 => n4738, A3 => n4739, A4 => n4740
                           , ZN => n4727);
   U3816 : OAI221_X1 port map( B1 => n3785, B2 => n4687, C1 => n4169, C2 => 
                           n4688, A => n4741, ZN => n4740);
   U3817 : AOI22_X1 port map( A1 => n4690, A2 => n3625, B1 => n4691, B2 => 
                           n4009, ZN => n4741);
   U3818 : OAI221_X1 port map( B1 => n3786, B2 => n4692, C1 => n4170, C2 => 
                           n4693, A => n4742, ZN => n4739);
   U3819 : AOI22_X1 port map( A1 => n4695, A2 => n3626, B1 => n4696, B2 => 
                           n4010, ZN => n4742);
   U3820 : OAI221_X1 port map( B1 => n3787, B2 => n4697, C1 => n4171, C2 => 
                           n4698, A => n4743, ZN => n4738);
   U3821 : AOI22_X1 port map( A1 => n4700, A2 => n3627, B1 => n4701, B2 => 
                           n4011, ZN => n4743);
   U3822 : OAI221_X1 port map( B1 => n3788, B2 => n4702, C1 => n4172, C2 => 
                           n4703, A => n4744, ZN => n4737);
   U3823 : AOI22_X1 port map( A1 => n4705, A2 => n3628, B1 => n4706, B2 => 
                           n4012, ZN => n4744);
   U3824 : MUX2_X1 port map( A => OUT2_28_port, B => n4745, S => n4656, Z => 
                           n2586);
   U3825 : NAND2_X1 port map( A1 => n4746, A2 => n4747, ZN => n4745);
   U3826 : NOR4_X1 port map( A1 => n4748, A2 => n4749, A3 => n4750, A4 => n4751
                           , ZN => n4747);
   U3827 : OAI221_X1 port map( B1 => n4, B2 => n4663, C1 => n36, C2 => n4664, A
                           => n4752, ZN => n4751);
   U3828 : AOI22_X1 port map( A1 => n4666, A2 => n6085, B1 => n4667, B2 => 
                           n6086, ZN => n4752);
   U3829 : OAI221_X1 port map( B1 => n132, B2 => n4668, C1 => n164, C2 => n4669
                           , A => n4753, ZN => n4750);
   U3830 : AOI22_X1 port map( A1 => n4671, A2 => n6083, B1 => n4672, B2 => 
                           n6084, ZN => n4753);
   U3831 : OAI221_X1 port map( B1 => n356, B2 => n4673, C1 => n324, C2 => n4674
                           , A => n4754, ZN => n4749);
   U3832 : AOI22_X1 port map( A1 => n4676, A2 => n3937, B1 => n4677, B2 => 
                           n4321, ZN => n4754);
   U3833 : OAI221_X1 port map( B1 => n3789, B2 => n4678, C1 => n4173, C2 => 
                           n4679, A => n4755, ZN => n4748);
   U3834 : AOI22_X1 port map( A1 => n4681, A2 => n3629, B1 => n4682, B2 => 
                           n4013, ZN => n4755);
   U3835 : NOR4_X1 port map( A1 => n4756, A2 => n4757, A3 => n4758, A4 => n4759
                           , ZN => n4746);
   U3836 : OAI221_X1 port map( B1 => n3790, B2 => n4687, C1 => n4174, C2 => 
                           n4688, A => n4760, ZN => n4759);
   U3837 : AOI22_X1 port map( A1 => n4690, A2 => n3630, B1 => n4691, B2 => 
                           n4014, ZN => n4760);
   U3838 : OAI221_X1 port map( B1 => n3791, B2 => n4692, C1 => n4175, C2 => 
                           n4693, A => n4761, ZN => n4758);
   U3839 : AOI22_X1 port map( A1 => n4695, A2 => n3631, B1 => n4696, B2 => 
                           n4015, ZN => n4761);
   U3840 : OAI221_X1 port map( B1 => n3792, B2 => n4697, C1 => n4176, C2 => 
                           n4698, A => n4762, ZN => n4757);
   U3841 : AOI22_X1 port map( A1 => n4700, A2 => n3632, B1 => n4701, B2 => 
                           n4016, ZN => n4762);
   U3842 : OAI221_X1 port map( B1 => n3793, B2 => n4702, C1 => n4177, C2 => 
                           n4703, A => n4763, ZN => n4756);
   U3843 : AOI22_X1 port map( A1 => n4705, A2 => n3633, B1 => n4706, B2 => 
                           n4017, ZN => n4763);
   U3844 : MUX2_X1 port map( A => OUT2_27_port, B => n4764, S => n4656, Z => 
                           n2585);
   U3845 : NAND2_X1 port map( A1 => n4765, A2 => n4766, ZN => n4764);
   U3846 : NOR4_X1 port map( A1 => n4767, A2 => n4768, A3 => n4769, A4 => n4770
                           , ZN => n4766);
   U3847 : OAI221_X1 port map( B1 => n5, B2 => n4663, C1 => n37, C2 => n4664, A
                           => n4771, ZN => n4770);
   U3848 : AOI22_X1 port map( A1 => n4666, A2 => n6081, B1 => n4667, B2 => 
                           n6082, ZN => n4771);
   U3849 : OAI221_X1 port map( B1 => n133, B2 => n4668, C1 => n165, C2 => n4669
                           , A => n4772, ZN => n4769);
   U3850 : AOI22_X1 port map( A1 => n4671, A2 => n6079, B1 => n4672, B2 => 
                           n6080, ZN => n4772);
   U3851 : OAI221_X1 port map( B1 => n357, B2 => n4673, C1 => n325, C2 => n4674
                           , A => n4773, ZN => n4768);
   U3852 : AOI22_X1 port map( A1 => n4676, A2 => n3938, B1 => n4677, B2 => 
                           n4322, ZN => n4773);
   U3853 : OAI221_X1 port map( B1 => n3794, B2 => n4678, C1 => n4178, C2 => 
                           n4679, A => n4774, ZN => n4767);
   U3854 : AOI22_X1 port map( A1 => n4681, A2 => n3634, B1 => n4682, B2 => 
                           n4018, ZN => n4774);
   U3855 : NOR4_X1 port map( A1 => n4775, A2 => n4776, A3 => n4777, A4 => n4778
                           , ZN => n4765);
   U3856 : OAI221_X1 port map( B1 => n3795, B2 => n4687, C1 => n4179, C2 => 
                           n4688, A => n4779, ZN => n4778);
   U3857 : AOI22_X1 port map( A1 => n4690, A2 => n3635, B1 => n4691, B2 => 
                           n4019, ZN => n4779);
   U3858 : OAI221_X1 port map( B1 => n3796, B2 => n4692, C1 => n4180, C2 => 
                           n4693, A => n4780, ZN => n4777);
   U3859 : AOI22_X1 port map( A1 => n4695, A2 => n3636, B1 => n4696, B2 => 
                           n4020, ZN => n4780);
   U3860 : OAI221_X1 port map( B1 => n3797, B2 => n4697, C1 => n4181, C2 => 
                           n4698, A => n4781, ZN => n4776);
   U3861 : AOI22_X1 port map( A1 => n4700, A2 => n3637, B1 => n4701, B2 => 
                           n4021, ZN => n4781);
   U3862 : OAI221_X1 port map( B1 => n3798, B2 => n4702, C1 => n4182, C2 => 
                           n4703, A => n4782, ZN => n4775);
   U3863 : AOI22_X1 port map( A1 => n4705, A2 => n3638, B1 => n4706, B2 => 
                           n4022, ZN => n4782);
   U3864 : MUX2_X1 port map( A => OUT2_26_port, B => n4783, S => n4656, Z => 
                           n2584);
   U3865 : NAND2_X1 port map( A1 => n4784, A2 => n4785, ZN => n4783);
   U3866 : NOR4_X1 port map( A1 => n4786, A2 => n4787, A3 => n4788, A4 => n4789
                           , ZN => n4785);
   U3867 : OAI221_X1 port map( B1 => n6, B2 => n4663, C1 => n38, C2 => n4664, A
                           => n4790, ZN => n4789);
   U3868 : AOI22_X1 port map( A1 => n4666, A2 => n6077, B1 => n4667, B2 => 
                           n6078, ZN => n4790);
   U3869 : OAI221_X1 port map( B1 => n134, B2 => n4668, C1 => n166, C2 => n4669
                           , A => n4791, ZN => n4788);
   U3870 : AOI22_X1 port map( A1 => n4671, A2 => n6075, B1 => n4672, B2 => 
                           n6076, ZN => n4791);
   U3871 : OAI221_X1 port map( B1 => n358, B2 => n4673, C1 => n326, C2 => n4674
                           , A => n4792, ZN => n4787);
   U3872 : AOI22_X1 port map( A1 => n4676, A2 => n3939, B1 => n4677, B2 => 
                           n4323, ZN => n4792);
   U3873 : OAI221_X1 port map( B1 => n3799, B2 => n4678, C1 => n4183, C2 => 
                           n4679, A => n4793, ZN => n4786);
   U3874 : AOI22_X1 port map( A1 => n4681, A2 => n3639, B1 => n4682, B2 => 
                           n4023, ZN => n4793);
   U3875 : NOR4_X1 port map( A1 => n4794, A2 => n4795, A3 => n4796, A4 => n4797
                           , ZN => n4784);
   U3876 : OAI221_X1 port map( B1 => n3800, B2 => n4687, C1 => n4184, C2 => 
                           n4688, A => n4798, ZN => n4797);
   U3877 : AOI22_X1 port map( A1 => n4690, A2 => n3640, B1 => n4691, B2 => 
                           n4024, ZN => n4798);
   U3878 : OAI221_X1 port map( B1 => n3801, B2 => n4692, C1 => n4185, C2 => 
                           n4693, A => n4799, ZN => n4796);
   U3879 : AOI22_X1 port map( A1 => n4695, A2 => n3641, B1 => n4696, B2 => 
                           n4025, ZN => n4799);
   U3880 : OAI221_X1 port map( B1 => n3802, B2 => n4697, C1 => n4186, C2 => 
                           n4698, A => n4800, ZN => n4795);
   U3881 : AOI22_X1 port map( A1 => n4700, A2 => n3642, B1 => n4701, B2 => 
                           n4026, ZN => n4800);
   U3882 : OAI221_X1 port map( B1 => n3803, B2 => n4702, C1 => n4187, C2 => 
                           n4703, A => n4801, ZN => n4794);
   U3883 : AOI22_X1 port map( A1 => n4705, A2 => n3643, B1 => n4706, B2 => 
                           n4027, ZN => n4801);
   U3884 : MUX2_X1 port map( A => OUT2_25_port, B => n4802, S => n4656, Z => 
                           n2583);
   U3885 : NAND2_X1 port map( A1 => n4803, A2 => n4804, ZN => n4802);
   U3886 : NOR4_X1 port map( A1 => n4805, A2 => n4806, A3 => n4807, A4 => n4808
                           , ZN => n4804);
   U3887 : OAI221_X1 port map( B1 => n7, B2 => n4663, C1 => n39, C2 => n4664, A
                           => n4809, ZN => n4808);
   U3888 : AOI22_X1 port map( A1 => n4666, A2 => n6073, B1 => n4667, B2 => 
                           n6074, ZN => n4809);
   U3889 : OAI221_X1 port map( B1 => n135, B2 => n4668, C1 => n167, C2 => n4669
                           , A => n4810, ZN => n4807);
   U3890 : AOI22_X1 port map( A1 => n4671, A2 => n6071, B1 => n4672, B2 => 
                           n6072, ZN => n4810);
   U3891 : OAI221_X1 port map( B1 => n359, B2 => n4673, C1 => n327, C2 => n4674
                           , A => n4811, ZN => n4806);
   U3892 : AOI22_X1 port map( A1 => n4676, A2 => n3940, B1 => n4677, B2 => 
                           n4324, ZN => n4811);
   U3893 : OAI221_X1 port map( B1 => n3804, B2 => n4678, C1 => n4188, C2 => 
                           n4679, A => n4812, ZN => n4805);
   U3894 : AOI22_X1 port map( A1 => n4681, A2 => n3644, B1 => n4682, B2 => 
                           n4028, ZN => n4812);
   U3895 : NOR4_X1 port map( A1 => n4813, A2 => n4814, A3 => n4815, A4 => n4816
                           , ZN => n4803);
   U3896 : OAI221_X1 port map( B1 => n3805, B2 => n4687, C1 => n4189, C2 => 
                           n4688, A => n4817, ZN => n4816);
   U3897 : AOI22_X1 port map( A1 => n4690, A2 => n3645, B1 => n4691, B2 => 
                           n4029, ZN => n4817);
   U3898 : OAI221_X1 port map( B1 => n3806, B2 => n4692, C1 => n4190, C2 => 
                           n4693, A => n4818, ZN => n4815);
   U3899 : AOI22_X1 port map( A1 => n4695, A2 => n3646, B1 => n4696, B2 => 
                           n4030, ZN => n4818);
   U3900 : OAI221_X1 port map( B1 => n3807, B2 => n4697, C1 => n4191, C2 => 
                           n4698, A => n4819, ZN => n4814);
   U3901 : AOI22_X1 port map( A1 => n4700, A2 => n3647, B1 => n4701, B2 => 
                           n4031, ZN => n4819);
   U3902 : OAI221_X1 port map( B1 => n3808, B2 => n4702, C1 => n4192, C2 => 
                           n4703, A => n4820, ZN => n4813);
   U3903 : AOI22_X1 port map( A1 => n4705, A2 => n3648, B1 => n4706, B2 => 
                           n4032, ZN => n4820);
   U3904 : MUX2_X1 port map( A => OUT2_24_port, B => n4821, S => n4656, Z => 
                           n2582);
   U3905 : NAND2_X1 port map( A1 => n4822, A2 => n4823, ZN => n4821);
   U3906 : NOR4_X1 port map( A1 => n4824, A2 => n4825, A3 => n4826, A4 => n4827
                           , ZN => n4823);
   U3907 : OAI221_X1 port map( B1 => n8, B2 => n4663, C1 => n40, C2 => n4664, A
                           => n4828, ZN => n4827);
   U3908 : AOI22_X1 port map( A1 => n4666, A2 => n6069, B1 => n4667, B2 => 
                           n6070, ZN => n4828);
   U3909 : OAI221_X1 port map( B1 => n136, B2 => n4668, C1 => n168, C2 => n4669
                           , A => n4829, ZN => n4826);
   U3910 : AOI22_X1 port map( A1 => n4671, A2 => n6067, B1 => n4672, B2 => 
                           n6068, ZN => n4829);
   U3911 : OAI221_X1 port map( B1 => n360, B2 => n4673, C1 => n328, C2 => n4674
                           , A => n4830, ZN => n4825);
   U3912 : AOI22_X1 port map( A1 => n4676, A2 => n3941, B1 => n4677, B2 => 
                           n4325, ZN => n4830);
   U3913 : OAI221_X1 port map( B1 => n3809, B2 => n4678, C1 => n4193, C2 => 
                           n4679, A => n4831, ZN => n4824);
   U3914 : AOI22_X1 port map( A1 => n4681, A2 => n3649, B1 => n4682, B2 => 
                           n4033, ZN => n4831);
   U3915 : NOR4_X1 port map( A1 => n4832, A2 => n4833, A3 => n4834, A4 => n4835
                           , ZN => n4822);
   U3916 : OAI221_X1 port map( B1 => n3810, B2 => n4687, C1 => n4194, C2 => 
                           n4688, A => n4836, ZN => n4835);
   U3917 : AOI22_X1 port map( A1 => n4690, A2 => n3650, B1 => n4691, B2 => 
                           n4034, ZN => n4836);
   U3918 : OAI221_X1 port map( B1 => n3811, B2 => n4692, C1 => n4195, C2 => 
                           n4693, A => n4837, ZN => n4834);
   U3919 : AOI22_X1 port map( A1 => n4695, A2 => n3651, B1 => n4696, B2 => 
                           n4035, ZN => n4837);
   U3920 : OAI221_X1 port map( B1 => n3812, B2 => n4697, C1 => n4196, C2 => 
                           n4698, A => n4838, ZN => n4833);
   U3921 : AOI22_X1 port map( A1 => n4700, A2 => n3652, B1 => n4701, B2 => 
                           n4036, ZN => n4838);
   U3922 : OAI221_X1 port map( B1 => n3813, B2 => n4702, C1 => n4197, C2 => 
                           n4703, A => n4839, ZN => n4832);
   U3923 : AOI22_X1 port map( A1 => n4705, A2 => n3653, B1 => n4706, B2 => 
                           n4037, ZN => n4839);
   U3924 : MUX2_X1 port map( A => OUT2_23_port, B => n4840, S => n4656, Z => 
                           n2581);
   U3925 : NAND2_X1 port map( A1 => n4841, A2 => n4842, ZN => n4840);
   U3926 : NOR4_X1 port map( A1 => n4843, A2 => n4844, A3 => n4845, A4 => n4846
                           , ZN => n4842);
   U3927 : OAI221_X1 port map( B1 => n9, B2 => n4663, C1 => n41, C2 => n4664, A
                           => n4847, ZN => n4846);
   U3928 : AOI22_X1 port map( A1 => n4666, A2 => n6065, B1 => n4667, B2 => 
                           n6066, ZN => n4847);
   U3929 : OAI221_X1 port map( B1 => n137, B2 => n4668, C1 => n169, C2 => n4669
                           , A => n4848, ZN => n4845);
   U3930 : AOI22_X1 port map( A1 => n4671, A2 => n6063, B1 => n4672, B2 => 
                           n6064, ZN => n4848);
   U3931 : OAI221_X1 port map( B1 => n361, B2 => n4673, C1 => n329, C2 => n4674
                           , A => n4849, ZN => n4844);
   U3932 : AOI22_X1 port map( A1 => n4676, A2 => n3942, B1 => n4677, B2 => 
                           n4326, ZN => n4849);
   U3933 : OAI221_X1 port map( B1 => n3814, B2 => n4678, C1 => n4198, C2 => 
                           n4679, A => n4850, ZN => n4843);
   U3934 : AOI22_X1 port map( A1 => n4681, A2 => n3654, B1 => n4682, B2 => 
                           n4038, ZN => n4850);
   U3935 : NOR4_X1 port map( A1 => n4851, A2 => n4852, A3 => n4853, A4 => n4854
                           , ZN => n4841);
   U3936 : OAI221_X1 port map( B1 => n3815, B2 => n4687, C1 => n4199, C2 => 
                           n4688, A => n4855, ZN => n4854);
   U3937 : AOI22_X1 port map( A1 => n4690, A2 => n3655, B1 => n4691, B2 => 
                           n4039, ZN => n4855);
   U3938 : OAI221_X1 port map( B1 => n3816, B2 => n4692, C1 => n4200, C2 => 
                           n4693, A => n4856, ZN => n4853);
   U3939 : AOI22_X1 port map( A1 => n4695, A2 => n3656, B1 => n4696, B2 => 
                           n4040, ZN => n4856);
   U3940 : OAI221_X1 port map( B1 => n3817, B2 => n4697, C1 => n4201, C2 => 
                           n4698, A => n4857, ZN => n4852);
   U3941 : AOI22_X1 port map( A1 => n4700, A2 => n3657, B1 => n4701, B2 => 
                           n4041, ZN => n4857);
   U3942 : OAI221_X1 port map( B1 => n3818, B2 => n4702, C1 => n4202, C2 => 
                           n4703, A => n4858, ZN => n4851);
   U3943 : AOI22_X1 port map( A1 => n4705, A2 => n3658, B1 => n4706, B2 => 
                           n4042, ZN => n4858);
   U3944 : MUX2_X1 port map( A => OUT2_22_port, B => n4859, S => n4656, Z => 
                           n2580);
   U3945 : NAND2_X1 port map( A1 => n4860, A2 => n4861, ZN => n4859);
   U3946 : NOR4_X1 port map( A1 => n4862, A2 => n4863, A3 => n4864, A4 => n4865
                           , ZN => n4861);
   U3947 : OAI221_X1 port map( B1 => n10, B2 => n4663, C1 => n42, C2 => n4664, 
                           A => n4866, ZN => n4865);
   U3948 : AOI22_X1 port map( A1 => n4666, A2 => n6061, B1 => n4667, B2 => 
                           n6062, ZN => n4866);
   U3949 : OAI221_X1 port map( B1 => n138, B2 => n4668, C1 => n170, C2 => n4669
                           , A => n4867, ZN => n4864);
   U3950 : AOI22_X1 port map( A1 => n4671, A2 => n6059, B1 => n4672, B2 => 
                           n6060, ZN => n4867);
   U3951 : OAI221_X1 port map( B1 => n362, B2 => n4673, C1 => n330, C2 => n4674
                           , A => n4868, ZN => n4863);
   U3952 : AOI22_X1 port map( A1 => n4676, A2 => n3943, B1 => n4677, B2 => 
                           n4327, ZN => n4868);
   U3953 : OAI221_X1 port map( B1 => n3819, B2 => n4678, C1 => n4203, C2 => 
                           n4679, A => n4869, ZN => n4862);
   U3954 : AOI22_X1 port map( A1 => n4681, A2 => n3659, B1 => n4682, B2 => 
                           n4043, ZN => n4869);
   U3955 : NOR4_X1 port map( A1 => n4870, A2 => n4871, A3 => n4872, A4 => n4873
                           , ZN => n4860);
   U3956 : OAI221_X1 port map( B1 => n3820, B2 => n4687, C1 => n4204, C2 => 
                           n4688, A => n4874, ZN => n4873);
   U3957 : AOI22_X1 port map( A1 => n4690, A2 => n3660, B1 => n4691, B2 => 
                           n4044, ZN => n4874);
   U3958 : OAI221_X1 port map( B1 => n3821, B2 => n4692, C1 => n4205, C2 => 
                           n4693, A => n4875, ZN => n4872);
   U3959 : AOI22_X1 port map( A1 => n4695, A2 => n3661, B1 => n4696, B2 => 
                           n4045, ZN => n4875);
   U3960 : OAI221_X1 port map( B1 => n3822, B2 => n4697, C1 => n4206, C2 => 
                           n4698, A => n4876, ZN => n4871);
   U3961 : AOI22_X1 port map( A1 => n4700, A2 => n3662, B1 => n4701, B2 => 
                           n4046, ZN => n4876);
   U3962 : OAI221_X1 port map( B1 => n3823, B2 => n4702, C1 => n4207, C2 => 
                           n4703, A => n4877, ZN => n4870);
   U3963 : AOI22_X1 port map( A1 => n4705, A2 => n3663, B1 => n4706, B2 => 
                           n4047, ZN => n4877);
   U3964 : MUX2_X1 port map( A => OUT2_21_port, B => n4878, S => n4656, Z => 
                           n2579);
   U3965 : NAND2_X1 port map( A1 => n4879, A2 => n4880, ZN => n4878);
   U3966 : NOR4_X1 port map( A1 => n4881, A2 => n4882, A3 => n4883, A4 => n4884
                           , ZN => n4880);
   U3967 : OAI221_X1 port map( B1 => n11, B2 => n4663, C1 => n43, C2 => n4664, 
                           A => n4885, ZN => n4884);
   U3968 : AOI22_X1 port map( A1 => n4666, A2 => n6057, B1 => n4667, B2 => 
                           n6058, ZN => n4885);
   U3969 : OAI221_X1 port map( B1 => n139, B2 => n4668, C1 => n171, C2 => n4669
                           , A => n4886, ZN => n4883);
   U3970 : AOI22_X1 port map( A1 => n4671, A2 => n6055, B1 => n4672, B2 => 
                           n6056, ZN => n4886);
   U3971 : OAI221_X1 port map( B1 => n363, B2 => n4673, C1 => n331, C2 => n4674
                           , A => n4887, ZN => n4882);
   U3972 : AOI22_X1 port map( A1 => n4676, A2 => n3944, B1 => n4677, B2 => 
                           n4328, ZN => n4887);
   U3973 : OAI221_X1 port map( B1 => n3824, B2 => n4678, C1 => n4208, C2 => 
                           n4679, A => n4888, ZN => n4881);
   U3974 : AOI22_X1 port map( A1 => n4681, A2 => n3664, B1 => n4682, B2 => 
                           n4048, ZN => n4888);
   U3975 : NOR4_X1 port map( A1 => n4889, A2 => n4890, A3 => n4891, A4 => n4892
                           , ZN => n4879);
   U3976 : OAI221_X1 port map( B1 => n3825, B2 => n4687, C1 => n4209, C2 => 
                           n4688, A => n4893, ZN => n4892);
   U3977 : AOI22_X1 port map( A1 => n4690, A2 => n3665, B1 => n4691, B2 => 
                           n4049, ZN => n4893);
   U3978 : OAI221_X1 port map( B1 => n3826, B2 => n4692, C1 => n4210, C2 => 
                           n4693, A => n4894, ZN => n4891);
   U3979 : AOI22_X1 port map( A1 => n4695, A2 => n3666, B1 => n4696, B2 => 
                           n4050, ZN => n4894);
   U3980 : OAI221_X1 port map( B1 => n3827, B2 => n4697, C1 => n4211, C2 => 
                           n4698, A => n4895, ZN => n4890);
   U3981 : AOI22_X1 port map( A1 => n4700, A2 => n3667, B1 => n4701, B2 => 
                           n4051, ZN => n4895);
   U3982 : OAI221_X1 port map( B1 => n3828, B2 => n4702, C1 => n4212, C2 => 
                           n4703, A => n4896, ZN => n4889);
   U3983 : AOI22_X1 port map( A1 => n4705, A2 => n3668, B1 => n4706, B2 => 
                           n4052, ZN => n4896);
   U3984 : MUX2_X1 port map( A => OUT2_20_port, B => n4897, S => n4656, Z => 
                           n2578);
   U3985 : NAND2_X1 port map( A1 => n4898, A2 => n4899, ZN => n4897);
   U3986 : NOR4_X1 port map( A1 => n4900, A2 => n4901, A3 => n4902, A4 => n4903
                           , ZN => n4899);
   U3987 : OAI221_X1 port map( B1 => n12, B2 => n4663, C1 => n44, C2 => n4664, 
                           A => n4904, ZN => n4903);
   U3988 : AOI22_X1 port map( A1 => n4666, A2 => n6053, B1 => n4667, B2 => 
                           n6054, ZN => n4904);
   U3989 : OAI221_X1 port map( B1 => n140, B2 => n4668, C1 => n172, C2 => n4669
                           , A => n4905, ZN => n4902);
   U3990 : AOI22_X1 port map( A1 => n4671, A2 => n6051, B1 => n4672, B2 => 
                           n6052, ZN => n4905);
   U3991 : OAI221_X1 port map( B1 => n364, B2 => n4673, C1 => n332, C2 => n4674
                           , A => n4906, ZN => n4901);
   U3992 : AOI22_X1 port map( A1 => n4676, A2 => n3945, B1 => n4677, B2 => 
                           n4329, ZN => n4906);
   U3993 : OAI221_X1 port map( B1 => n3829, B2 => n4678, C1 => n4213, C2 => 
                           n4679, A => n4907, ZN => n4900);
   U3994 : AOI22_X1 port map( A1 => n4681, A2 => n3669, B1 => n4682, B2 => 
                           n4053, ZN => n4907);
   U3995 : NOR4_X1 port map( A1 => n4908, A2 => n4909, A3 => n4910, A4 => n4911
                           , ZN => n4898);
   U3996 : OAI221_X1 port map( B1 => n3830, B2 => n4687, C1 => n4214, C2 => 
                           n4688, A => n4912, ZN => n4911);
   U3997 : AOI22_X1 port map( A1 => n4690, A2 => n3670, B1 => n4691, B2 => 
                           n4054, ZN => n4912);
   U3998 : OAI221_X1 port map( B1 => n3831, B2 => n4692, C1 => n4215, C2 => 
                           n4693, A => n4913, ZN => n4910);
   U3999 : AOI22_X1 port map( A1 => n4695, A2 => n3671, B1 => n4696, B2 => 
                           n4055, ZN => n4913);
   U4000 : OAI221_X1 port map( B1 => n3832, B2 => n4697, C1 => n4216, C2 => 
                           n4698, A => n4914, ZN => n4909);
   U4001 : AOI22_X1 port map( A1 => n4700, A2 => n3672, B1 => n4701, B2 => 
                           n4056, ZN => n4914);
   U4002 : OAI221_X1 port map( B1 => n3833, B2 => n4702, C1 => n4217, C2 => 
                           n4703, A => n4915, ZN => n4908);
   U4003 : AOI22_X1 port map( A1 => n4705, A2 => n3673, B1 => n4706, B2 => 
                           n4057, ZN => n4915);
   U4004 : MUX2_X1 port map( A => OUT2_19_port, B => n4916, S => n4656, Z => 
                           n2577);
   U4005 : NAND2_X1 port map( A1 => n4917, A2 => n4918, ZN => n4916);
   U4006 : NOR4_X1 port map( A1 => n4919, A2 => n4920, A3 => n4921, A4 => n4922
                           , ZN => n4918);
   U4007 : OAI221_X1 port map( B1 => n13, B2 => n4663, C1 => n45, C2 => n4664, 
                           A => n4923, ZN => n4922);
   U4008 : AOI22_X1 port map( A1 => n4666, A2 => n6049, B1 => n4667, B2 => 
                           n6050, ZN => n4923);
   U4009 : OAI221_X1 port map( B1 => n141, B2 => n4668, C1 => n173, C2 => n4669
                           , A => n4924, ZN => n4921);
   U4010 : AOI22_X1 port map( A1 => n4671, A2 => n6047, B1 => n4672, B2 => 
                           n6048, ZN => n4924);
   U4011 : OAI221_X1 port map( B1 => n365, B2 => n4673, C1 => n333, C2 => n4674
                           , A => n4925, ZN => n4920);
   U4012 : AOI22_X1 port map( A1 => n4676, A2 => n3946, B1 => n4677, B2 => 
                           n4330, ZN => n4925);
   U4013 : OAI221_X1 port map( B1 => n3834, B2 => n4678, C1 => n4218, C2 => 
                           n4679, A => n4926, ZN => n4919);
   U4014 : AOI22_X1 port map( A1 => n4681, A2 => n3674, B1 => n4682, B2 => 
                           n4058, ZN => n4926);
   U4015 : NOR4_X1 port map( A1 => n4927, A2 => n4928, A3 => n4929, A4 => n4930
                           , ZN => n4917);
   U4016 : OAI221_X1 port map( B1 => n3835, B2 => n4687, C1 => n4219, C2 => 
                           n4688, A => n4931, ZN => n4930);
   U4017 : AOI22_X1 port map( A1 => n4690, A2 => n3675, B1 => n4691, B2 => 
                           n4059, ZN => n4931);
   U4018 : OAI221_X1 port map( B1 => n3836, B2 => n4692, C1 => n4220, C2 => 
                           n4693, A => n4932, ZN => n4929);
   U4019 : AOI22_X1 port map( A1 => n4695, A2 => n3676, B1 => n4696, B2 => 
                           n4060, ZN => n4932);
   U4020 : OAI221_X1 port map( B1 => n3837, B2 => n4697, C1 => n4221, C2 => 
                           n4698, A => n4933, ZN => n4928);
   U4021 : AOI22_X1 port map( A1 => n4700, A2 => n3677, B1 => n4701, B2 => 
                           n4061, ZN => n4933);
   U4022 : OAI221_X1 port map( B1 => n3838, B2 => n4702, C1 => n4222, C2 => 
                           n4703, A => n4934, ZN => n4927);
   U4023 : AOI22_X1 port map( A1 => n4705, A2 => n3678, B1 => n4706, B2 => 
                           n4062, ZN => n4934);
   U4024 : MUX2_X1 port map( A => OUT2_18_port, B => n4935, S => n4656, Z => 
                           n2576);
   U4025 : NAND2_X1 port map( A1 => n4936, A2 => n4937, ZN => n4935);
   U4026 : NOR4_X1 port map( A1 => n4938, A2 => n4939, A3 => n4940, A4 => n4941
                           , ZN => n4937);
   U4027 : OAI221_X1 port map( B1 => n14, B2 => n4663, C1 => n46, C2 => n4664, 
                           A => n4942, ZN => n4941);
   U4028 : AOI22_X1 port map( A1 => n4666, A2 => n6045, B1 => n4667, B2 => 
                           n6046, ZN => n4942);
   U4029 : OAI221_X1 port map( B1 => n142, B2 => n4668, C1 => n174, C2 => n4669
                           , A => n4943, ZN => n4940);
   U4030 : AOI22_X1 port map( A1 => n4671, A2 => n6043, B1 => n4672, B2 => 
                           n6044, ZN => n4943);
   U4031 : OAI221_X1 port map( B1 => n366, B2 => n4673, C1 => n334, C2 => n4674
                           , A => n4944, ZN => n4939);
   U4032 : AOI22_X1 port map( A1 => n4676, A2 => n3947, B1 => n4677, B2 => 
                           n4331, ZN => n4944);
   U4033 : OAI221_X1 port map( B1 => n3839, B2 => n4678, C1 => n4223, C2 => 
                           n4679, A => n4945, ZN => n4938);
   U4034 : AOI22_X1 port map( A1 => n4681, A2 => n3679, B1 => n4682, B2 => 
                           n4063, ZN => n4945);
   U4035 : NOR4_X1 port map( A1 => n4946, A2 => n4947, A3 => n4948, A4 => n4949
                           , ZN => n4936);
   U4036 : OAI221_X1 port map( B1 => n3840, B2 => n4687, C1 => n4224, C2 => 
                           n4688, A => n4950, ZN => n4949);
   U4037 : AOI22_X1 port map( A1 => n4690, A2 => n3680, B1 => n4691, B2 => 
                           n4064, ZN => n4950);
   U4038 : OAI221_X1 port map( B1 => n3841, B2 => n4692, C1 => n4225, C2 => 
                           n4693, A => n4951, ZN => n4948);
   U4039 : AOI22_X1 port map( A1 => n4695, A2 => n3681, B1 => n4696, B2 => 
                           n4065, ZN => n4951);
   U4040 : OAI221_X1 port map( B1 => n3842, B2 => n4697, C1 => n4226, C2 => 
                           n4698, A => n4952, ZN => n4947);
   U4041 : AOI22_X1 port map( A1 => n4700, A2 => n3682, B1 => n4701, B2 => 
                           n4066, ZN => n4952);
   U4042 : OAI221_X1 port map( B1 => n3843, B2 => n4702, C1 => n4227, C2 => 
                           n4703, A => n4953, ZN => n4946);
   U4043 : AOI22_X1 port map( A1 => n4705, A2 => n3683, B1 => n4706, B2 => 
                           n4067, ZN => n4953);
   U4044 : MUX2_X1 port map( A => OUT2_17_port, B => n4954, S => n4656, Z => 
                           n2575);
   U4045 : NAND2_X1 port map( A1 => n4955, A2 => n4956, ZN => n4954);
   U4046 : NOR4_X1 port map( A1 => n4957, A2 => n4958, A3 => n4959, A4 => n4960
                           , ZN => n4956);
   U4047 : OAI221_X1 port map( B1 => n15, B2 => n4663, C1 => n47, C2 => n4664, 
                           A => n4961, ZN => n4960);
   U4048 : AOI22_X1 port map( A1 => n4666, A2 => n6041, B1 => n4667, B2 => 
                           n6042, ZN => n4961);
   U4049 : OAI221_X1 port map( B1 => n143, B2 => n4668, C1 => n175, C2 => n4669
                           , A => n4962, ZN => n4959);
   U4050 : AOI22_X1 port map( A1 => n4671, A2 => n6039, B1 => n4672, B2 => 
                           n6040, ZN => n4962);
   U4051 : OAI221_X1 port map( B1 => n367, B2 => n4673, C1 => n335, C2 => n4674
                           , A => n4963, ZN => n4958);
   U4052 : AOI22_X1 port map( A1 => n4676, A2 => n3948, B1 => n4677, B2 => 
                           n4332, ZN => n4963);
   U4053 : OAI221_X1 port map( B1 => n3844, B2 => n4678, C1 => n4228, C2 => 
                           n4679, A => n4964, ZN => n4957);
   U4054 : AOI22_X1 port map( A1 => n4681, A2 => n3684, B1 => n4682, B2 => 
                           n4068, ZN => n4964);
   U4055 : NOR4_X1 port map( A1 => n4965, A2 => n4966, A3 => n4967, A4 => n4968
                           , ZN => n4955);
   U4056 : OAI221_X1 port map( B1 => n3845, B2 => n4687, C1 => n4229, C2 => 
                           n4688, A => n4969, ZN => n4968);
   U4057 : AOI22_X1 port map( A1 => n4690, A2 => n3685, B1 => n4691, B2 => 
                           n4069, ZN => n4969);
   U4058 : OAI221_X1 port map( B1 => n3846, B2 => n4692, C1 => n4230, C2 => 
                           n4693, A => n4970, ZN => n4967);
   U4059 : AOI22_X1 port map( A1 => n4695, A2 => n3686, B1 => n4696, B2 => 
                           n4070, ZN => n4970);
   U4060 : OAI221_X1 port map( B1 => n3847, B2 => n4697, C1 => n4231, C2 => 
                           n4698, A => n4971, ZN => n4966);
   U4061 : AOI22_X1 port map( A1 => n4700, A2 => n3687, B1 => n4701, B2 => 
                           n4071, ZN => n4971);
   U4062 : OAI221_X1 port map( B1 => n3848, B2 => n4702, C1 => n4232, C2 => 
                           n4703, A => n4972, ZN => n4965);
   U4063 : AOI22_X1 port map( A1 => n4705, A2 => n3688, B1 => n4706, B2 => 
                           n4072, ZN => n4972);
   U4064 : MUX2_X1 port map( A => OUT2_16_port, B => n4973, S => n4656, Z => 
                           n2574);
   U4065 : NAND2_X1 port map( A1 => n4974, A2 => n4975, ZN => n4973);
   U4066 : NOR4_X1 port map( A1 => n4976, A2 => n4977, A3 => n4978, A4 => n4979
                           , ZN => n4975);
   U4067 : OAI221_X1 port map( B1 => n16, B2 => n4663, C1 => n48, C2 => n4664, 
                           A => n4980, ZN => n4979);
   U4068 : AOI22_X1 port map( A1 => n4666, A2 => n6037, B1 => n4667, B2 => 
                           n6038, ZN => n4980);
   U4069 : OAI221_X1 port map( B1 => n144, B2 => n4668, C1 => n176, C2 => n4669
                           , A => n4981, ZN => n4978);
   U4070 : AOI22_X1 port map( A1 => n4671, A2 => n6035, B1 => n4672, B2 => 
                           n6036, ZN => n4981);
   U4071 : OAI221_X1 port map( B1 => n368, B2 => n4673, C1 => n336, C2 => n4674
                           , A => n4982, ZN => n4977);
   U4072 : AOI22_X1 port map( A1 => n4676, A2 => n3949, B1 => n4677, B2 => 
                           n4333, ZN => n4982);
   U4073 : OAI221_X1 port map( B1 => n3849, B2 => n4678, C1 => n4233, C2 => 
                           n4679, A => n4983, ZN => n4976);
   U4074 : AOI22_X1 port map( A1 => n4681, A2 => n3689, B1 => n4682, B2 => 
                           n4073, ZN => n4983);
   U4075 : NOR4_X1 port map( A1 => n4984, A2 => n4985, A3 => n4986, A4 => n4987
                           , ZN => n4974);
   U4076 : OAI221_X1 port map( B1 => n3850, B2 => n4687, C1 => n4234, C2 => 
                           n4688, A => n4988, ZN => n4987);
   U4077 : AOI22_X1 port map( A1 => n4690, A2 => n3690, B1 => n4691, B2 => 
                           n4074, ZN => n4988);
   U4078 : OAI221_X1 port map( B1 => n3851, B2 => n4692, C1 => n4235, C2 => 
                           n4693, A => n4989, ZN => n4986);
   U4079 : AOI22_X1 port map( A1 => n4695, A2 => n3691, B1 => n4696, B2 => 
                           n4075, ZN => n4989);
   U4080 : OAI221_X1 port map( B1 => n3852, B2 => n4697, C1 => n4236, C2 => 
                           n4698, A => n4990, ZN => n4985);
   U4081 : AOI22_X1 port map( A1 => n4700, A2 => n3692, B1 => n4701, B2 => 
                           n4076, ZN => n4990);
   U4082 : OAI221_X1 port map( B1 => n3853, B2 => n4702, C1 => n4237, C2 => 
                           n4703, A => n4991, ZN => n4984);
   U4083 : AOI22_X1 port map( A1 => n4705, A2 => n3693, B1 => n4706, B2 => 
                           n4077, ZN => n4991);
   U4084 : MUX2_X1 port map( A => OUT2_15_port, B => n4992, S => n4656, Z => 
                           n2573);
   U4085 : NAND2_X1 port map( A1 => n4993, A2 => n4994, ZN => n4992);
   U4086 : NOR4_X1 port map( A1 => n4995, A2 => n4996, A3 => n4997, A4 => n4998
                           , ZN => n4994);
   U4087 : OAI221_X1 port map( B1 => n17, B2 => n4663, C1 => n49, C2 => n4664, 
                           A => n4999, ZN => n4998);
   U4088 : AOI22_X1 port map( A1 => n4666, A2 => n6033, B1 => n4667, B2 => 
                           n6034, ZN => n4999);
   U4089 : OAI221_X1 port map( B1 => n145, B2 => n4668, C1 => n177, C2 => n4669
                           , A => n5000, ZN => n4997);
   U4090 : AOI22_X1 port map( A1 => n4671, A2 => n6031, B1 => n4672, B2 => 
                           n6032, ZN => n5000);
   U4091 : OAI221_X1 port map( B1 => n369, B2 => n4673, C1 => n337, C2 => n4674
                           , A => n5001, ZN => n4996);
   U4092 : AOI22_X1 port map( A1 => n4676, A2 => n3950, B1 => n4677, B2 => 
                           n4334, ZN => n5001);
   U4093 : OAI221_X1 port map( B1 => n3854, B2 => n4678, C1 => n4238, C2 => 
                           n4679, A => n5002, ZN => n4995);
   U4094 : AOI22_X1 port map( A1 => n4681, A2 => n3694, B1 => n4682, B2 => 
                           n4078, ZN => n5002);
   U4095 : NOR4_X1 port map( A1 => n5003, A2 => n5004, A3 => n5005, A4 => n5006
                           , ZN => n4993);
   U4096 : OAI221_X1 port map( B1 => n3855, B2 => n4687, C1 => n4239, C2 => 
                           n4688, A => n5007, ZN => n5006);
   U4097 : AOI22_X1 port map( A1 => n4690, A2 => n3695, B1 => n4691, B2 => 
                           n4079, ZN => n5007);
   U4098 : OAI221_X1 port map( B1 => n3856, B2 => n4692, C1 => n4240, C2 => 
                           n4693, A => n5008, ZN => n5005);
   U4099 : AOI22_X1 port map( A1 => n4695, A2 => n3696, B1 => n4696, B2 => 
                           n4080, ZN => n5008);
   U4100 : OAI221_X1 port map( B1 => n3857, B2 => n4697, C1 => n4241, C2 => 
                           n4698, A => n5009, ZN => n5004);
   U4101 : AOI22_X1 port map( A1 => n4700, A2 => n3697, B1 => n4701, B2 => 
                           n4081, ZN => n5009);
   U4102 : OAI221_X1 port map( B1 => n3858, B2 => n4702, C1 => n4242, C2 => 
                           n4703, A => n5010, ZN => n5003);
   U4103 : AOI22_X1 port map( A1 => n4705, A2 => n3698, B1 => n4706, B2 => 
                           n4082, ZN => n5010);
   U4104 : MUX2_X1 port map( A => OUT2_14_port, B => n5011, S => n4656, Z => 
                           n2572);
   U4105 : NAND2_X1 port map( A1 => n5012, A2 => n5013, ZN => n5011);
   U4106 : NOR4_X1 port map( A1 => n5014, A2 => n5015, A3 => n5016, A4 => n5017
                           , ZN => n5013);
   U4107 : OAI221_X1 port map( B1 => n18, B2 => n4663, C1 => n50, C2 => n4664, 
                           A => n5018, ZN => n5017);
   U4108 : AOI22_X1 port map( A1 => n4666, A2 => n6029, B1 => n4667, B2 => 
                           n6030, ZN => n5018);
   U4109 : OAI221_X1 port map( B1 => n146, B2 => n4668, C1 => n178, C2 => n4669
                           , A => n5019, ZN => n5016);
   U4110 : AOI22_X1 port map( A1 => n4671, A2 => n6027, B1 => n4672, B2 => 
                           n6028, ZN => n5019);
   U4111 : OAI221_X1 port map( B1 => n370, B2 => n4673, C1 => n338, C2 => n4674
                           , A => n5020, ZN => n5015);
   U4112 : AOI22_X1 port map( A1 => n4676, A2 => n3951, B1 => n4677, B2 => 
                           n4335, ZN => n5020);
   U4113 : OAI221_X1 port map( B1 => n3859, B2 => n4678, C1 => n4243, C2 => 
                           n4679, A => n5021, ZN => n5014);
   U4114 : AOI22_X1 port map( A1 => n4681, A2 => n3699, B1 => n4682, B2 => 
                           n4083, ZN => n5021);
   U4115 : NOR4_X1 port map( A1 => n5022, A2 => n5023, A3 => n5024, A4 => n5025
                           , ZN => n5012);
   U4116 : OAI221_X1 port map( B1 => n3860, B2 => n4687, C1 => n4244, C2 => 
                           n4688, A => n5026, ZN => n5025);
   U4117 : AOI22_X1 port map( A1 => n4690, A2 => n3700, B1 => n4691, B2 => 
                           n4084, ZN => n5026);
   U4118 : OAI221_X1 port map( B1 => n3861, B2 => n4692, C1 => n4245, C2 => 
                           n4693, A => n5027, ZN => n5024);
   U4119 : AOI22_X1 port map( A1 => n4695, A2 => n3701, B1 => n4696, B2 => 
                           n4085, ZN => n5027);
   U4120 : OAI221_X1 port map( B1 => n3862, B2 => n4697, C1 => n4246, C2 => 
                           n4698, A => n5028, ZN => n5023);
   U4121 : AOI22_X1 port map( A1 => n4700, A2 => n3702, B1 => n4701, B2 => 
                           n4086, ZN => n5028);
   U4122 : OAI221_X1 port map( B1 => n3863, B2 => n4702, C1 => n4247, C2 => 
                           n4703, A => n5029, ZN => n5022);
   U4123 : AOI22_X1 port map( A1 => n4705, A2 => n3703, B1 => n4706, B2 => 
                           n4087, ZN => n5029);
   U4124 : MUX2_X1 port map( A => OUT2_13_port, B => n5030, S => n4656, Z => 
                           n2571);
   U4125 : NAND2_X1 port map( A1 => n5031, A2 => n5032, ZN => n5030);
   U4126 : NOR4_X1 port map( A1 => n5033, A2 => n5034, A3 => n5035, A4 => n5036
                           , ZN => n5032);
   U4127 : OAI221_X1 port map( B1 => n19, B2 => n4663, C1 => n51, C2 => n4664, 
                           A => n5037, ZN => n5036);
   U4128 : AOI22_X1 port map( A1 => n4666, A2 => n6025, B1 => n4667, B2 => 
                           n6026, ZN => n5037);
   U4129 : OAI221_X1 port map( B1 => n147, B2 => n4668, C1 => n179, C2 => n4669
                           , A => n5038, ZN => n5035);
   U4130 : AOI22_X1 port map( A1 => n4671, A2 => n6023, B1 => n4672, B2 => 
                           n6024, ZN => n5038);
   U4131 : OAI221_X1 port map( B1 => n371, B2 => n4673, C1 => n339, C2 => n4674
                           , A => n5039, ZN => n5034);
   U4132 : AOI22_X1 port map( A1 => n4676, A2 => n3952, B1 => n4677, B2 => 
                           n4336, ZN => n5039);
   U4133 : OAI221_X1 port map( B1 => n3864, B2 => n4678, C1 => n4248, C2 => 
                           n4679, A => n5040, ZN => n5033);
   U4134 : AOI22_X1 port map( A1 => n4681, A2 => n3704, B1 => n4682, B2 => 
                           n4088, ZN => n5040);
   U4135 : NOR4_X1 port map( A1 => n5041, A2 => n5042, A3 => n5043, A4 => n5044
                           , ZN => n5031);
   U4136 : OAI221_X1 port map( B1 => n3865, B2 => n4687, C1 => n4249, C2 => 
                           n4688, A => n5045, ZN => n5044);
   U4137 : AOI22_X1 port map( A1 => n4690, A2 => n3705, B1 => n4691, B2 => 
                           n4089, ZN => n5045);
   U4138 : OAI221_X1 port map( B1 => n3866, B2 => n4692, C1 => n4250, C2 => 
                           n4693, A => n5046, ZN => n5043);
   U4139 : AOI22_X1 port map( A1 => n4695, A2 => n3706, B1 => n4696, B2 => 
                           n4090, ZN => n5046);
   U4140 : OAI221_X1 port map( B1 => n3867, B2 => n4697, C1 => n4251, C2 => 
                           n4698, A => n5047, ZN => n5042);
   U4141 : AOI22_X1 port map( A1 => n4700, A2 => n3707, B1 => n4701, B2 => 
                           n4091, ZN => n5047);
   U4142 : OAI221_X1 port map( B1 => n3868, B2 => n4702, C1 => n4252, C2 => 
                           n4703, A => n5048, ZN => n5041);
   U4143 : AOI22_X1 port map( A1 => n4705, A2 => n3708, B1 => n4706, B2 => 
                           n4092, ZN => n5048);
   U4144 : MUX2_X1 port map( A => OUT2_12_port, B => n5049, S => n4656, Z => 
                           n2570);
   U4145 : NAND2_X1 port map( A1 => n5050, A2 => n5051, ZN => n5049);
   U4146 : NOR4_X1 port map( A1 => n5052, A2 => n5053, A3 => n5054, A4 => n5055
                           , ZN => n5051);
   U4147 : OAI221_X1 port map( B1 => n20, B2 => n4663, C1 => n52, C2 => n4664, 
                           A => n5056, ZN => n5055);
   U4148 : AOI22_X1 port map( A1 => n4666, A2 => n6021, B1 => n4667, B2 => 
                           n6022, ZN => n5056);
   U4149 : OAI221_X1 port map( B1 => n148, B2 => n4668, C1 => n180, C2 => n4669
                           , A => n5057, ZN => n5054);
   U4150 : AOI22_X1 port map( A1 => n4671, A2 => n6019, B1 => n4672, B2 => 
                           n6020, ZN => n5057);
   U4151 : OAI221_X1 port map( B1 => n372, B2 => n4673, C1 => n340, C2 => n4674
                           , A => n5058, ZN => n5053);
   U4152 : AOI22_X1 port map( A1 => n4676, A2 => n3953, B1 => n4677, B2 => 
                           n4337, ZN => n5058);
   U4153 : OAI221_X1 port map( B1 => n3869, B2 => n4678, C1 => n4253, C2 => 
                           n4679, A => n5059, ZN => n5052);
   U4154 : AOI22_X1 port map( A1 => n4681, A2 => n3709, B1 => n4682, B2 => 
                           n4093, ZN => n5059);
   U4155 : NOR4_X1 port map( A1 => n5060, A2 => n5061, A3 => n5062, A4 => n5063
                           , ZN => n5050);
   U4156 : OAI221_X1 port map( B1 => n3870, B2 => n4687, C1 => n4254, C2 => 
                           n4688, A => n5064, ZN => n5063);
   U4157 : AOI22_X1 port map( A1 => n4690, A2 => n3710, B1 => n4691, B2 => 
                           n4094, ZN => n5064);
   U4158 : OAI221_X1 port map( B1 => n3871, B2 => n4692, C1 => n4255, C2 => 
                           n4693, A => n5065, ZN => n5062);
   U4159 : AOI22_X1 port map( A1 => n4695, A2 => n3711, B1 => n4696, B2 => 
                           n4095, ZN => n5065);
   U4160 : OAI221_X1 port map( B1 => n3872, B2 => n4697, C1 => n4256, C2 => 
                           n4698, A => n5066, ZN => n5061);
   U4161 : AOI22_X1 port map( A1 => n4700, A2 => n3712, B1 => n4701, B2 => 
                           n4096, ZN => n5066);
   U4162 : OAI221_X1 port map( B1 => n3873, B2 => n4702, C1 => n4257, C2 => 
                           n4703, A => n5067, ZN => n5060);
   U4163 : AOI22_X1 port map( A1 => n4705, A2 => n3713, B1 => n4706, B2 => 
                           n4097, ZN => n5067);
   U4164 : MUX2_X1 port map( A => OUT2_11_port, B => n5068, S => n4656, Z => 
                           n2569);
   U4165 : NAND2_X1 port map( A1 => n5069, A2 => n5070, ZN => n5068);
   U4166 : NOR4_X1 port map( A1 => n5071, A2 => n5072, A3 => n5073, A4 => n5074
                           , ZN => n5070);
   U4167 : OAI221_X1 port map( B1 => n21, B2 => n4663, C1 => n53, C2 => n4664, 
                           A => n5075, ZN => n5074);
   U4168 : AOI22_X1 port map( A1 => n4666, A2 => n6017, B1 => n4667, B2 => 
                           n6018, ZN => n5075);
   U4169 : OAI221_X1 port map( B1 => n149, B2 => n4668, C1 => n181, C2 => n4669
                           , A => n5076, ZN => n5073);
   U4170 : AOI22_X1 port map( A1 => n4671, A2 => n6015, B1 => n4672, B2 => 
                           n6016, ZN => n5076);
   U4171 : OAI221_X1 port map( B1 => n373, B2 => n4673, C1 => n341, C2 => n4674
                           , A => n5077, ZN => n5072);
   U4172 : AOI22_X1 port map( A1 => n4676, A2 => n3954, B1 => n4677, B2 => 
                           n4338, ZN => n5077);
   U4173 : OAI221_X1 port map( B1 => n3874, B2 => n4678, C1 => n4258, C2 => 
                           n4679, A => n5078, ZN => n5071);
   U4174 : AOI22_X1 port map( A1 => n4681, A2 => n3714, B1 => n4682, B2 => 
                           n4098, ZN => n5078);
   U4175 : NOR4_X1 port map( A1 => n5079, A2 => n5080, A3 => n5081, A4 => n5082
                           , ZN => n5069);
   U4176 : OAI221_X1 port map( B1 => n3875, B2 => n4687, C1 => n4259, C2 => 
                           n4688, A => n5083, ZN => n5082);
   U4177 : AOI22_X1 port map( A1 => n4690, A2 => n3715, B1 => n4691, B2 => 
                           n4099, ZN => n5083);
   U4178 : OAI221_X1 port map( B1 => n3876, B2 => n4692, C1 => n4260, C2 => 
                           n4693, A => n5084, ZN => n5081);
   U4179 : AOI22_X1 port map( A1 => n4695, A2 => n3716, B1 => n4696, B2 => 
                           n4100, ZN => n5084);
   U4180 : OAI221_X1 port map( B1 => n3877, B2 => n4697, C1 => n4261, C2 => 
                           n4698, A => n5085, ZN => n5080);
   U4181 : AOI22_X1 port map( A1 => n4700, A2 => n3717, B1 => n4701, B2 => 
                           n4101, ZN => n5085);
   U4182 : OAI221_X1 port map( B1 => n3878, B2 => n4702, C1 => n4262, C2 => 
                           n4703, A => n5086, ZN => n5079);
   U4183 : AOI22_X1 port map( A1 => n4705, A2 => n3718, B1 => n4706, B2 => 
                           n4102, ZN => n5086);
   U4184 : MUX2_X1 port map( A => OUT2_10_port, B => n5087, S => n4656, Z => 
                           n2568);
   U4185 : NAND2_X1 port map( A1 => n5088, A2 => n5089, ZN => n5087);
   U4186 : NOR4_X1 port map( A1 => n5090, A2 => n5091, A3 => n5092, A4 => n5093
                           , ZN => n5089);
   U4187 : OAI221_X1 port map( B1 => n22, B2 => n4663, C1 => n54, C2 => n4664, 
                           A => n5094, ZN => n5093);
   U4188 : AOI22_X1 port map( A1 => n4666, A2 => n6013, B1 => n4667, B2 => 
                           n6014, ZN => n5094);
   U4189 : OAI221_X1 port map( B1 => n150, B2 => n4668, C1 => n182, C2 => n4669
                           , A => n5095, ZN => n5092);
   U4190 : AOI22_X1 port map( A1 => n4671, A2 => n6011, B1 => n4672, B2 => 
                           n6012, ZN => n5095);
   U4191 : OAI221_X1 port map( B1 => n374, B2 => n4673, C1 => n342, C2 => n4674
                           , A => n5096, ZN => n5091);
   U4192 : AOI22_X1 port map( A1 => n4676, A2 => n3955, B1 => n4677, B2 => 
                           n4339, ZN => n5096);
   U4193 : OAI221_X1 port map( B1 => n3879, B2 => n4678, C1 => n4263, C2 => 
                           n4679, A => n5097, ZN => n5090);
   U4194 : AOI22_X1 port map( A1 => n4681, A2 => n3719, B1 => n4682, B2 => 
                           n4103, ZN => n5097);
   U4195 : NOR4_X1 port map( A1 => n5098, A2 => n5099, A3 => n5100, A4 => n5101
                           , ZN => n5088);
   U4196 : OAI221_X1 port map( B1 => n3880, B2 => n4687, C1 => n4264, C2 => 
                           n4688, A => n5102, ZN => n5101);
   U4197 : AOI22_X1 port map( A1 => n4690, A2 => n3720, B1 => n4691, B2 => 
                           n4104, ZN => n5102);
   U4198 : OAI221_X1 port map( B1 => n3881, B2 => n4692, C1 => n4265, C2 => 
                           n4693, A => n5103, ZN => n5100);
   U4199 : AOI22_X1 port map( A1 => n4695, A2 => n3721, B1 => n4696, B2 => 
                           n4105, ZN => n5103);
   U4200 : OAI221_X1 port map( B1 => n3882, B2 => n4697, C1 => n4266, C2 => 
                           n4698, A => n5104, ZN => n5099);
   U4201 : AOI22_X1 port map( A1 => n4700, A2 => n3722, B1 => n4701, B2 => 
                           n4106, ZN => n5104);
   U4202 : OAI221_X1 port map( B1 => n3883, B2 => n4702, C1 => n4267, C2 => 
                           n4703, A => n5105, ZN => n5098);
   U4203 : AOI22_X1 port map( A1 => n4705, A2 => n3723, B1 => n4706, B2 => 
                           n4107, ZN => n5105);
   U4204 : MUX2_X1 port map( A => OUT2_9_port, B => n5106, S => n4656, Z => 
                           n2567);
   U4205 : NAND2_X1 port map( A1 => n5107, A2 => n5108, ZN => n5106);
   U4206 : NOR4_X1 port map( A1 => n5109, A2 => n5110, A3 => n5111, A4 => n5112
                           , ZN => n5108);
   U4207 : OAI221_X1 port map( B1 => n23, B2 => n4663, C1 => n55, C2 => n4664, 
                           A => n5113, ZN => n5112);
   U4208 : AOI22_X1 port map( A1 => n4666, A2 => n6009, B1 => n4667, B2 => 
                           n6010, ZN => n5113);
   U4209 : OAI221_X1 port map( B1 => n151, B2 => n4668, C1 => n183, C2 => n4669
                           , A => n5114, ZN => n5111);
   U4210 : AOI22_X1 port map( A1 => n4671, A2 => n6007, B1 => n4672, B2 => 
                           n6008, ZN => n5114);
   U4211 : OAI221_X1 port map( B1 => n375, B2 => n4673, C1 => n343, C2 => n4674
                           , A => n5115, ZN => n5110);
   U4212 : AOI22_X1 port map( A1 => n4676, A2 => n3956, B1 => n4677, B2 => 
                           n4340, ZN => n5115);
   U4213 : OAI221_X1 port map( B1 => n3884, B2 => n4678, C1 => n4268, C2 => 
                           n4679, A => n5116, ZN => n5109);
   U4214 : AOI22_X1 port map( A1 => n4681, A2 => n3724, B1 => n4682, B2 => 
                           n4108, ZN => n5116);
   U4215 : NOR4_X1 port map( A1 => n5117, A2 => n5118, A3 => n5119, A4 => n5120
                           , ZN => n5107);
   U4216 : OAI221_X1 port map( B1 => n3885, B2 => n4687, C1 => n4269, C2 => 
                           n4688, A => n5121, ZN => n5120);
   U4217 : AOI22_X1 port map( A1 => n4690, A2 => n3725, B1 => n4691, B2 => 
                           n4109, ZN => n5121);
   U4218 : OAI221_X1 port map( B1 => n3886, B2 => n4692, C1 => n4270, C2 => 
                           n4693, A => n5122, ZN => n5119);
   U4219 : AOI22_X1 port map( A1 => n4695, A2 => n3726, B1 => n4696, B2 => 
                           n4110, ZN => n5122);
   U4220 : OAI221_X1 port map( B1 => n3887, B2 => n4697, C1 => n4271, C2 => 
                           n4698, A => n5123, ZN => n5118);
   U4221 : AOI22_X1 port map( A1 => n4700, A2 => n3727, B1 => n4701, B2 => 
                           n4111, ZN => n5123);
   U4222 : OAI221_X1 port map( B1 => n3888, B2 => n4702, C1 => n4272, C2 => 
                           n4703, A => n5124, ZN => n5117);
   U4223 : AOI22_X1 port map( A1 => n4705, A2 => n3728, B1 => n4706, B2 => 
                           n4112, ZN => n5124);
   U4224 : MUX2_X1 port map( A => OUT2_8_port, B => n5125, S => n4656, Z => 
                           n2566);
   U4225 : NAND2_X1 port map( A1 => n5126, A2 => n5127, ZN => n5125);
   U4226 : NOR4_X1 port map( A1 => n5128, A2 => n5129, A3 => n5130, A4 => n5131
                           , ZN => n5127);
   U4227 : OAI221_X1 port map( B1 => n24, B2 => n4663, C1 => n56, C2 => n4664, 
                           A => n5132, ZN => n5131);
   U4228 : AOI22_X1 port map( A1 => n4666, A2 => n6005, B1 => n4667, B2 => 
                           n6006, ZN => n5132);
   U4229 : OAI221_X1 port map( B1 => n152, B2 => n4668, C1 => n184, C2 => n4669
                           , A => n5133, ZN => n5130);
   U4230 : AOI22_X1 port map( A1 => n4671, A2 => n6003, B1 => n4672, B2 => 
                           n6004, ZN => n5133);
   U4231 : OAI221_X1 port map( B1 => n376, B2 => n4673, C1 => n344, C2 => n4674
                           , A => n5134, ZN => n5129);
   U4232 : AOI22_X1 port map( A1 => n4676, A2 => n3957, B1 => n4677, B2 => 
                           n4341, ZN => n5134);
   U4233 : OAI221_X1 port map( B1 => n3889, B2 => n4678, C1 => n4273, C2 => 
                           n4679, A => n5135, ZN => n5128);
   U4234 : AOI22_X1 port map( A1 => n4681, A2 => n3729, B1 => n4682, B2 => 
                           n4113, ZN => n5135);
   U4235 : NOR4_X1 port map( A1 => n5136, A2 => n5137, A3 => n5138, A4 => n5139
                           , ZN => n5126);
   U4236 : OAI221_X1 port map( B1 => n3890, B2 => n4687, C1 => n4274, C2 => 
                           n4688, A => n5140, ZN => n5139);
   U4237 : AOI22_X1 port map( A1 => n4690, A2 => n3730, B1 => n4691, B2 => 
                           n4114, ZN => n5140);
   U4238 : OAI221_X1 port map( B1 => n3891, B2 => n4692, C1 => n4275, C2 => 
                           n4693, A => n5141, ZN => n5138);
   U4239 : AOI22_X1 port map( A1 => n4695, A2 => n3731, B1 => n4696, B2 => 
                           n4115, ZN => n5141);
   U4240 : OAI221_X1 port map( B1 => n3892, B2 => n4697, C1 => n4276, C2 => 
                           n4698, A => n5142, ZN => n5137);
   U4241 : AOI22_X1 port map( A1 => n4700, A2 => n3732, B1 => n4701, B2 => 
                           n4116, ZN => n5142);
   U4242 : OAI221_X1 port map( B1 => n3893, B2 => n4702, C1 => n4277, C2 => 
                           n4703, A => n5143, ZN => n5136);
   U4243 : AOI22_X1 port map( A1 => n4705, A2 => n3733, B1 => n4706, B2 => 
                           n4117, ZN => n5143);
   U4244 : MUX2_X1 port map( A => OUT2_7_port, B => n5144, S => n4656, Z => 
                           n2565);
   U4245 : NAND2_X1 port map( A1 => n5145, A2 => n5146, ZN => n5144);
   U4246 : NOR4_X1 port map( A1 => n5147, A2 => n5148, A3 => n5149, A4 => n5150
                           , ZN => n5146);
   U4247 : OAI221_X1 port map( B1 => n25, B2 => n4663, C1 => n57, C2 => n4664, 
                           A => n5151, ZN => n5150);
   U4248 : AOI22_X1 port map( A1 => n4666, A2 => n6001, B1 => n4667, B2 => 
                           n6002, ZN => n5151);
   U4249 : OAI221_X1 port map( B1 => n153, B2 => n4668, C1 => n185, C2 => n4669
                           , A => n5152, ZN => n5149);
   U4250 : AOI22_X1 port map( A1 => n4671, A2 => n5999, B1 => n4672, B2 => 
                           n6000, ZN => n5152);
   U4251 : OAI221_X1 port map( B1 => n377, B2 => n4673, C1 => n345, C2 => n4674
                           , A => n5153, ZN => n5148);
   U4252 : AOI22_X1 port map( A1 => n4676, A2 => n3958, B1 => n4677, B2 => 
                           n4342, ZN => n5153);
   U4253 : OAI221_X1 port map( B1 => n3894, B2 => n4678, C1 => n4278, C2 => 
                           n4679, A => n5154, ZN => n5147);
   U4254 : AOI22_X1 port map( A1 => n4681, A2 => n3734, B1 => n4682, B2 => 
                           n4118, ZN => n5154);
   U4255 : NOR4_X1 port map( A1 => n5155, A2 => n5156, A3 => n5157, A4 => n5158
                           , ZN => n5145);
   U4256 : OAI221_X1 port map( B1 => n3895, B2 => n4687, C1 => n4279, C2 => 
                           n4688, A => n5159, ZN => n5158);
   U4257 : AOI22_X1 port map( A1 => n4690, A2 => n3735, B1 => n4691, B2 => 
                           n4119, ZN => n5159);
   U4258 : OAI221_X1 port map( B1 => n3896, B2 => n4692, C1 => n4280, C2 => 
                           n4693, A => n5160, ZN => n5157);
   U4259 : AOI22_X1 port map( A1 => n4695, A2 => n3736, B1 => n4696, B2 => 
                           n4120, ZN => n5160);
   U4260 : OAI221_X1 port map( B1 => n3897, B2 => n4697, C1 => n4281, C2 => 
                           n4698, A => n5161, ZN => n5156);
   U4261 : AOI22_X1 port map( A1 => n4700, A2 => n3737, B1 => n4701, B2 => 
                           n4121, ZN => n5161);
   U4262 : OAI221_X1 port map( B1 => n3898, B2 => n4702, C1 => n4282, C2 => 
                           n4703, A => n5162, ZN => n5155);
   U4263 : AOI22_X1 port map( A1 => n4705, A2 => n3738, B1 => n4706, B2 => 
                           n4122, ZN => n5162);
   U4264 : MUX2_X1 port map( A => OUT2_6_port, B => n5163, S => n4656, Z => 
                           n2564);
   U4265 : NAND2_X1 port map( A1 => n5164, A2 => n5165, ZN => n5163);
   U4266 : NOR4_X1 port map( A1 => n5166, A2 => n5167, A3 => n5168, A4 => n5169
                           , ZN => n5165);
   U4267 : OAI221_X1 port map( B1 => n26, B2 => n4663, C1 => n58, C2 => n4664, 
                           A => n5170, ZN => n5169);
   U4268 : AOI22_X1 port map( A1 => n4666, A2 => n5997, B1 => n4667, B2 => 
                           n5998, ZN => n5170);
   U4269 : OAI221_X1 port map( B1 => n154, B2 => n4668, C1 => n186, C2 => n4669
                           , A => n5171, ZN => n5168);
   U4270 : AOI22_X1 port map( A1 => n4671, A2 => n5995, B1 => n4672, B2 => 
                           n5996, ZN => n5171);
   U4271 : OAI221_X1 port map( B1 => n378, B2 => n4673, C1 => n346, C2 => n4674
                           , A => n5172, ZN => n5167);
   U4272 : AOI22_X1 port map( A1 => n4676, A2 => n3959, B1 => n4677, B2 => 
                           n4343, ZN => n5172);
   U4273 : OAI221_X1 port map( B1 => n3899, B2 => n4678, C1 => n4283, C2 => 
                           n4679, A => n5173, ZN => n5166);
   U4274 : AOI22_X1 port map( A1 => n4681, A2 => n3739, B1 => n4682, B2 => 
                           n4123, ZN => n5173);
   U4275 : NOR4_X1 port map( A1 => n5174, A2 => n5175, A3 => n5176, A4 => n5177
                           , ZN => n5164);
   U4276 : OAI221_X1 port map( B1 => n3900, B2 => n4687, C1 => n4284, C2 => 
                           n4688, A => n5178, ZN => n5177);
   U4277 : AOI22_X1 port map( A1 => n4690, A2 => n3740, B1 => n4691, B2 => 
                           n4124, ZN => n5178);
   U4278 : OAI221_X1 port map( B1 => n3901, B2 => n4692, C1 => n4285, C2 => 
                           n4693, A => n5179, ZN => n5176);
   U4279 : AOI22_X1 port map( A1 => n4695, A2 => n3741, B1 => n4696, B2 => 
                           n4125, ZN => n5179);
   U4280 : OAI221_X1 port map( B1 => n3902, B2 => n4697, C1 => n4286, C2 => 
                           n4698, A => n5180, ZN => n5175);
   U4281 : AOI22_X1 port map( A1 => n4700, A2 => n3742, B1 => n4701, B2 => 
                           n4126, ZN => n5180);
   U4282 : OAI221_X1 port map( B1 => n3903, B2 => n4702, C1 => n4287, C2 => 
                           n4703, A => n5181, ZN => n5174);
   U4283 : AOI22_X1 port map( A1 => n4705, A2 => n3743, B1 => n4706, B2 => 
                           n4127, ZN => n5181);
   U4284 : MUX2_X1 port map( A => OUT2_5_port, B => n5182, S => n4656, Z => 
                           n2563);
   U4285 : NAND2_X1 port map( A1 => n5183, A2 => n5184, ZN => n5182);
   U4286 : NOR4_X1 port map( A1 => n5185, A2 => n5186, A3 => n5187, A4 => n5188
                           , ZN => n5184);
   U4287 : OAI221_X1 port map( B1 => n27, B2 => n4663, C1 => n59, C2 => n4664, 
                           A => n5189, ZN => n5188);
   U4288 : AOI22_X1 port map( A1 => n4666, A2 => n5993, B1 => n4667, B2 => 
                           n5994, ZN => n5189);
   U4289 : OAI221_X1 port map( B1 => n155, B2 => n4668, C1 => n187, C2 => n4669
                           , A => n5190, ZN => n5187);
   U4290 : AOI22_X1 port map( A1 => n4671, A2 => n5991, B1 => n4672, B2 => 
                           n5992, ZN => n5190);
   U4291 : OAI221_X1 port map( B1 => n379, B2 => n4673, C1 => n347, C2 => n4674
                           , A => n5191, ZN => n5186);
   U4292 : AOI22_X1 port map( A1 => n4676, A2 => n3960, B1 => n4677, B2 => 
                           n4344, ZN => n5191);
   U4293 : OAI221_X1 port map( B1 => n3904, B2 => n4678, C1 => n4288, C2 => 
                           n4679, A => n5192, ZN => n5185);
   U4294 : AOI22_X1 port map( A1 => n4681, A2 => n3744, B1 => n4682, B2 => 
                           n4128, ZN => n5192);
   U4295 : NOR4_X1 port map( A1 => n5193, A2 => n5194, A3 => n5195, A4 => n5196
                           , ZN => n5183);
   U4296 : OAI221_X1 port map( B1 => n3905, B2 => n4687, C1 => n4289, C2 => 
                           n4688, A => n5197, ZN => n5196);
   U4297 : AOI22_X1 port map( A1 => n4690, A2 => n3745, B1 => n4691, B2 => 
                           n4129, ZN => n5197);
   U4298 : OAI221_X1 port map( B1 => n3906, B2 => n4692, C1 => n4290, C2 => 
                           n4693, A => n5198, ZN => n5195);
   U4299 : AOI22_X1 port map( A1 => n4695, A2 => n3746, B1 => n4696, B2 => 
                           n4130, ZN => n5198);
   U4300 : OAI221_X1 port map( B1 => n3907, B2 => n4697, C1 => n4291, C2 => 
                           n4698, A => n5199, ZN => n5194);
   U4301 : AOI22_X1 port map( A1 => n4700, A2 => n3747, B1 => n4701, B2 => 
                           n4131, ZN => n5199);
   U4302 : OAI221_X1 port map( B1 => n3908, B2 => n4702, C1 => n4292, C2 => 
                           n4703, A => n5200, ZN => n5193);
   U4303 : AOI22_X1 port map( A1 => n4705, A2 => n3748, B1 => n4706, B2 => 
                           n4132, ZN => n5200);
   U4304 : MUX2_X1 port map( A => OUT2_4_port, B => n5201, S => n4656, Z => 
                           n2562);
   U4305 : NAND2_X1 port map( A1 => n5202, A2 => n5203, ZN => n5201);
   U4306 : NOR4_X1 port map( A1 => n5204, A2 => n5205, A3 => n5206, A4 => n5207
                           , ZN => n5203);
   U4307 : OAI221_X1 port map( B1 => n28, B2 => n4663, C1 => n60, C2 => n4664, 
                           A => n5208, ZN => n5207);
   U4308 : AOI22_X1 port map( A1 => n4666, A2 => n5989, B1 => n4667, B2 => 
                           n5990, ZN => n5208);
   U4309 : OAI221_X1 port map( B1 => n156, B2 => n4668, C1 => n188, C2 => n4669
                           , A => n5209, ZN => n5206);
   U4310 : AOI22_X1 port map( A1 => n4671, A2 => n5987, B1 => n4672, B2 => 
                           n5988, ZN => n5209);
   U4311 : OAI221_X1 port map( B1 => n380, B2 => n4673, C1 => n348, C2 => n4674
                           , A => n5210, ZN => n5205);
   U4312 : AOI22_X1 port map( A1 => n4676, A2 => n3961, B1 => n4677, B2 => 
                           n4345, ZN => n5210);
   U4313 : OAI221_X1 port map( B1 => n3909, B2 => n4678, C1 => n4293, C2 => 
                           n4679, A => n5211, ZN => n5204);
   U4314 : AOI22_X1 port map( A1 => n4681, A2 => n3749, B1 => n4682, B2 => 
                           n4133, ZN => n5211);
   U4315 : NOR4_X1 port map( A1 => n5212, A2 => n5213, A3 => n5214, A4 => n5215
                           , ZN => n5202);
   U4316 : OAI221_X1 port map( B1 => n3910, B2 => n4687, C1 => n4294, C2 => 
                           n4688, A => n5216, ZN => n5215);
   U4317 : AOI22_X1 port map( A1 => n4690, A2 => n3750, B1 => n4691, B2 => 
                           n4134, ZN => n5216);
   U4318 : OAI221_X1 port map( B1 => n3911, B2 => n4692, C1 => n4295, C2 => 
                           n4693, A => n5217, ZN => n5214);
   U4319 : AOI22_X1 port map( A1 => n4695, A2 => n3751, B1 => n4696, B2 => 
                           n4135, ZN => n5217);
   U4320 : OAI221_X1 port map( B1 => n3912, B2 => n4697, C1 => n4296, C2 => 
                           n4698, A => n5218, ZN => n5213);
   U4321 : AOI22_X1 port map( A1 => n4700, A2 => n3752, B1 => n4701, B2 => 
                           n4136, ZN => n5218);
   U4322 : OAI221_X1 port map( B1 => n3913, B2 => n4702, C1 => n4297, C2 => 
                           n4703, A => n5219, ZN => n5212);
   U4323 : AOI22_X1 port map( A1 => n4705, A2 => n3753, B1 => n4706, B2 => 
                           n4137, ZN => n5219);
   U4324 : MUX2_X1 port map( A => OUT2_3_port, B => n5220, S => n4656, Z => 
                           n2561);
   U4325 : NAND2_X1 port map( A1 => n5221, A2 => n5222, ZN => n5220);
   U4326 : NOR4_X1 port map( A1 => n5223, A2 => n5224, A3 => n5225, A4 => n5226
                           , ZN => n5222);
   U4327 : OAI221_X1 port map( B1 => n29, B2 => n4663, C1 => n61, C2 => n4664, 
                           A => n5227, ZN => n5226);
   U4328 : AOI22_X1 port map( A1 => n4666, A2 => n5985, B1 => n4667, B2 => 
                           n5986, ZN => n5227);
   U4329 : OAI221_X1 port map( B1 => n157, B2 => n4668, C1 => n189, C2 => n4669
                           , A => n5228, ZN => n5225);
   U4330 : AOI22_X1 port map( A1 => n4671, A2 => n5983, B1 => n4672, B2 => 
                           n5984, ZN => n5228);
   U4331 : OAI221_X1 port map( B1 => n381, B2 => n4673, C1 => n349, C2 => n4674
                           , A => n5229, ZN => n5224);
   U4332 : AOI22_X1 port map( A1 => n4676, A2 => n3962, B1 => n4677, B2 => 
                           n4346, ZN => n5229);
   U4333 : OAI221_X1 port map( B1 => n3914, B2 => n4678, C1 => n4298, C2 => 
                           n4679, A => n5230, ZN => n5223);
   U4334 : AOI22_X1 port map( A1 => n4681, A2 => n3754, B1 => n4682, B2 => 
                           n4138, ZN => n5230);
   U4335 : NOR4_X1 port map( A1 => n5231, A2 => n5232, A3 => n5233, A4 => n5234
                           , ZN => n5221);
   U4336 : OAI221_X1 port map( B1 => n3915, B2 => n4687, C1 => n4299, C2 => 
                           n4688, A => n5235, ZN => n5234);
   U4337 : AOI22_X1 port map( A1 => n4690, A2 => n3755, B1 => n4691, B2 => 
                           n4139, ZN => n5235);
   U4338 : OAI221_X1 port map( B1 => n3916, B2 => n4692, C1 => n4300, C2 => 
                           n4693, A => n5236, ZN => n5233);
   U4339 : AOI22_X1 port map( A1 => n4695, A2 => n3756, B1 => n4696, B2 => 
                           n4140, ZN => n5236);
   U4340 : OAI221_X1 port map( B1 => n3917, B2 => n4697, C1 => n4301, C2 => 
                           n4698, A => n5237, ZN => n5232);
   U4341 : AOI22_X1 port map( A1 => n4700, A2 => n3757, B1 => n4701, B2 => 
                           n4141, ZN => n5237);
   U4342 : OAI221_X1 port map( B1 => n3918, B2 => n4702, C1 => n4302, C2 => 
                           n4703, A => n5238, ZN => n5231);
   U4343 : AOI22_X1 port map( A1 => n4705, A2 => n3758, B1 => n4706, B2 => 
                           n4142, ZN => n5238);
   U4344 : MUX2_X1 port map( A => OUT2_2_port, B => n5239, S => n4656, Z => 
                           n2560);
   U4345 : NAND2_X1 port map( A1 => n5240, A2 => n5241, ZN => n5239);
   U4346 : NOR4_X1 port map( A1 => n5242, A2 => n5243, A3 => n5244, A4 => n5245
                           , ZN => n5241);
   U4347 : OAI221_X1 port map( B1 => n30, B2 => n4663, C1 => n62, C2 => n4664, 
                           A => n5246, ZN => n5245);
   U4348 : AOI22_X1 port map( A1 => n4666, A2 => n5981, B1 => n4667, B2 => 
                           n5982, ZN => n5246);
   U4349 : OAI221_X1 port map( B1 => n158, B2 => n4668, C1 => n190, C2 => n4669
                           , A => n5247, ZN => n5244);
   U4350 : AOI22_X1 port map( A1 => n4671, A2 => n5979, B1 => n4672, B2 => 
                           n5980, ZN => n5247);
   U4351 : OAI221_X1 port map( B1 => n382, B2 => n4673, C1 => n350, C2 => n4674
                           , A => n5248, ZN => n5243);
   U4352 : AOI22_X1 port map( A1 => n4676, A2 => n3963, B1 => n4677, B2 => 
                           n4347, ZN => n5248);
   U4353 : OAI221_X1 port map( B1 => n3919, B2 => n4678, C1 => n4303, C2 => 
                           n4679, A => n5249, ZN => n5242);
   U4354 : AOI22_X1 port map( A1 => n4681, A2 => n3759, B1 => n4682, B2 => 
                           n4143, ZN => n5249);
   U4355 : NOR4_X1 port map( A1 => n5250, A2 => n5251, A3 => n5252, A4 => n5253
                           , ZN => n5240);
   U4356 : OAI221_X1 port map( B1 => n3920, B2 => n4687, C1 => n4304, C2 => 
                           n4688, A => n5254, ZN => n5253);
   U4357 : AOI22_X1 port map( A1 => n4690, A2 => n3760, B1 => n4691, B2 => 
                           n4144, ZN => n5254);
   U4358 : OAI221_X1 port map( B1 => n3921, B2 => n4692, C1 => n4305, C2 => 
                           n4693, A => n5255, ZN => n5252);
   U4359 : AOI22_X1 port map( A1 => n4695, A2 => n3761, B1 => n4696, B2 => 
                           n4145, ZN => n5255);
   U4360 : OAI221_X1 port map( B1 => n3922, B2 => n4697, C1 => n4306, C2 => 
                           n4698, A => n5256, ZN => n5251);
   U4361 : AOI22_X1 port map( A1 => n4700, A2 => n3762, B1 => n4701, B2 => 
                           n4146, ZN => n5256);
   U4362 : OAI221_X1 port map( B1 => n3923, B2 => n4702, C1 => n4307, C2 => 
                           n4703, A => n5257, ZN => n5250);
   U4363 : AOI22_X1 port map( A1 => n4705, A2 => n3763, B1 => n4706, B2 => 
                           n4147, ZN => n5257);
   U4364 : MUX2_X1 port map( A => OUT2_1_port, B => n5258, S => n4656, Z => 
                           n2559);
   U4365 : NAND2_X1 port map( A1 => n5259, A2 => n5260, ZN => n5258);
   U4366 : NOR4_X1 port map( A1 => n5261, A2 => n5262, A3 => n5263, A4 => n5264
                           , ZN => n5260);
   U4367 : OAI221_X1 port map( B1 => n31, B2 => n4663, C1 => n63, C2 => n4664, 
                           A => n5265, ZN => n5264);
   U4368 : AOI22_X1 port map( A1 => n4666, A2 => n5977, B1 => n4667, B2 => 
                           n5978, ZN => n5265);
   U4369 : OAI221_X1 port map( B1 => n159, B2 => n4668, C1 => n191, C2 => n4669
                           , A => n5266, ZN => n5263);
   U4370 : AOI22_X1 port map( A1 => n4671, A2 => n5975, B1 => n4672, B2 => 
                           n5976, ZN => n5266);
   U4371 : OAI221_X1 port map( B1 => n383, B2 => n4673, C1 => n351, C2 => n4674
                           , A => n5267, ZN => n5262);
   U4372 : AOI22_X1 port map( A1 => n4676, A2 => n3964, B1 => n4677, B2 => 
                           n4348, ZN => n5267);
   U4373 : OAI221_X1 port map( B1 => n3924, B2 => n4678, C1 => n4308, C2 => 
                           n4679, A => n5268, ZN => n5261);
   U4374 : AOI22_X1 port map( A1 => n4681, A2 => n3764, B1 => n4682, B2 => 
                           n4148, ZN => n5268);
   U4375 : NOR4_X1 port map( A1 => n5269, A2 => n5270, A3 => n5271, A4 => n5272
                           , ZN => n5259);
   U4376 : OAI221_X1 port map( B1 => n3925, B2 => n4687, C1 => n4309, C2 => 
                           n4688, A => n5273, ZN => n5272);
   U4377 : AOI22_X1 port map( A1 => n4690, A2 => n3765, B1 => n4691, B2 => 
                           n4149, ZN => n5273);
   U4378 : OAI221_X1 port map( B1 => n3926, B2 => n4692, C1 => n4310, C2 => 
                           n4693, A => n5274, ZN => n5271);
   U4379 : AOI22_X1 port map( A1 => n4695, A2 => n3766, B1 => n4696, B2 => 
                           n4150, ZN => n5274);
   U4380 : OAI221_X1 port map( B1 => n3927, B2 => n4697, C1 => n4311, C2 => 
                           n4698, A => n5275, ZN => n5270);
   U4381 : AOI22_X1 port map( A1 => n4700, A2 => n3767, B1 => n4701, B2 => 
                           n4151, ZN => n5275);
   U4382 : OAI221_X1 port map( B1 => n3928, B2 => n4702, C1 => n4312, C2 => 
                           n4703, A => n5276, ZN => n5269);
   U4383 : AOI22_X1 port map( A1 => n4705, A2 => n3768, B1 => n4706, B2 => 
                           n4152, ZN => n5276);
   U4384 : MUX2_X1 port map( A => OUT2_0_port, B => n5277, S => n4656, Z => 
                           n2558);
   U4385 : NAND2_X1 port map( A1 => n5278, A2 => n5279, ZN => n5277);
   U4386 : NOR4_X1 port map( A1 => n5280, A2 => n5281, A3 => n5282, A4 => n5283
                           , ZN => n5279);
   U4387 : OAI221_X1 port map( B1 => n32, B2 => n4663, C1 => n64, C2 => n4664, 
                           A => n5284, ZN => n5283);
   U4388 : AOI22_X1 port map( A1 => n4666, A2 => n5973, B1 => n4667, B2 => 
                           n5974, ZN => n5284);
   U4389 : OAI221_X1 port map( B1 => n160, B2 => n4668, C1 => n192, C2 => n4669
                           , A => n5289, ZN => n5282);
   U4390 : AOI22_X1 port map( A1 => n4671, A2 => n5971, B1 => n4672, B2 => 
                           n5972, ZN => n5289);
   U4391 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => n5292, 
                           ZN => n5287);
   U4392 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => 
                           ADD_RD2(0), ZN => n5285);
   U4393 : OAI221_X1 port map( B1 => n384, B2 => n4673, C1 => n352, C2 => n4674
                           , A => n5293, ZN => n5281);
   U4394 : AOI22_X1 port map( A1 => n4676, A2 => n3965, B1 => n4677, B2 => 
                           n4349, ZN => n5293);
   U4395 : OAI221_X1 port map( B1 => n3929, B2 => n4678, C1 => n4313, C2 => 
                           n4679, A => n5296, ZN => n5280);
   U4396 : AOI22_X1 port map( A1 => n4681, A2 => n3769, B1 => n4682, B2 => 
                           n4153, ZN => n5296);
   U4397 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(4), A3 => n5297, 
                           ZN => n5295);
   U4398 : NOR3_X1 port map( A1 => n5292, A2 => ADD_RD2(4), A3 => n5297, ZN => 
                           n5294);
   U4399 : NOR4_X1 port map( A1 => n5298, A2 => n5299, A3 => n5300, A4 => n5301
                           , ZN => n5278);
   U4400 : OAI221_X1 port map( B1 => n3930, B2 => n4687, C1 => n4314, C2 => 
                           n4688, A => n5302, ZN => n5301);
   U4401 : AOI22_X1 port map( A1 => n4690, A2 => n3770, B1 => n4691, B2 => 
                           n4154, ZN => n5302);
   U4402 : OAI221_X1 port map( B1 => n3931, B2 => n4692, C1 => n4315, C2 => 
                           n4693, A => n5305, ZN => n5300);
   U4403 : AOI22_X1 port map( A1 => n4695, A2 => n3771, B1 => n4696, B2 => 
                           n4155, ZN => n5305);
   U4404 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(3), A3 => n5306, 
                           ZN => n5304);
   U4405 : NOR3_X1 port map( A1 => n5292, A2 => ADD_RD2(3), A3 => n5306, ZN => 
                           n5303);
   U4406 : OAI221_X1 port map( B1 => n3932, B2 => n4697, C1 => n4316, C2 => 
                           n4698, A => n5307, ZN => n5299);
   U4407 : AOI22_X1 port map( A1 => n4700, A2 => n3772, B1 => n4701, B2 => 
                           n4156, ZN => n5307);
   U4408 : NOR2_X1 port map( A1 => n5310, A2 => ADD_RD2(2), ZN => n5286);
   U4409 : NOR2_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), ZN => n5288);
   U4410 : OAI221_X1 port map( B1 => n3933, B2 => n4702, C1 => n4317, C2 => 
                           n4703, A => n5311, ZN => n5298);
   U4411 : AOI22_X1 port map( A1 => n4705, A2 => n3773, B1 => n4706, B2 => 
                           n4157, ZN => n5311);
   U4412 : NOR2_X1 port map( A1 => n5312, A2 => n5310, ZN => n5290);
   U4413 : INV_X1 port map( A => ADD_RD2(1), ZN => n5310);
   U4414 : NOR3_X1 port map( A1 => n5297, A2 => ADD_RD2(0), A3 => n5306, ZN => 
                           n5309);
   U4415 : NOR2_X1 port map( A1 => n5312, A2 => ADD_RD2(1), ZN => n5291);
   U4416 : INV_X1 port map( A => ADD_RD2(2), ZN => n5312);
   U4417 : NOR3_X1 port map( A1 => n5297, A2 => n5292, A3 => n5306, ZN => n5308
                           );
   U4418 : INV_X1 port map( A => ADD_RD2(4), ZN => n5306);
   U4419 : INV_X1 port map( A => ADD_RD2(0), ZN => n5292);
   U4420 : INV_X1 port map( A => ADD_RD2(3), ZN => n5297);
   U4421 : MUX2_X1 port map( A => OUT1_31_port, B => n5313, S => n5314, Z => 
                           n2557);
   U4422 : NAND2_X1 port map( A1 => n5315, A2 => n5316, ZN => n5313);
   U4423 : NOR4_X1 port map( A1 => n5317, A2 => n5318, A3 => n5319, A4 => n5320
                           , ZN => n5316);
   U4424 : OAI221_X1 port map( B1 => n1, B2 => n5321, C1 => n33, C2 => n5322, A
                           => n5323, ZN => n5320);
   U4425 : AOI22_X1 port map( A1 => n5324, A2 => n6097, B1 => n5325, B2 => 
                           n6098, ZN => n5323);
   U4426 : OAI221_X1 port map( B1 => n129, B2 => n5326, C1 => n161, C2 => n5327
                           , A => n5328, ZN => n5319);
   U4427 : AOI22_X1 port map( A1 => n5329, A2 => n6095, B1 => n5330, B2 => 
                           n6096, ZN => n5328);
   U4428 : OAI221_X1 port map( B1 => n289, B2 => n5331, C1 => n257, C2 => n5332
                           , A => n5333, ZN => n5318);
   U4429 : AOI22_X1 port map( A1 => n5334, A2 => n3966, B1 => n5335, B2 => 
                           n4350, ZN => n5333);
   U4430 : OAI221_X1 port map( B1 => n3774, B2 => n5336, C1 => n4158, C2 => 
                           n5337, A => n5338, ZN => n5317);
   U4431 : AOI22_X1 port map( A1 => n5339, A2 => n3614, B1 => n5340, B2 => 
                           n3998, ZN => n5338);
   U4432 : NOR4_X1 port map( A1 => n5341, A2 => n5342, A3 => n5343, A4 => n5344
                           , ZN => n5315);
   U4433 : OAI221_X1 port map( B1 => n3775, B2 => n5345, C1 => n4159, C2 => 
                           n5346, A => n5347, ZN => n5344);
   U4434 : AOI22_X1 port map( A1 => n5348, A2 => n3615, B1 => n5349, B2 => 
                           n3999, ZN => n5347);
   U4435 : OAI221_X1 port map( B1 => n3776, B2 => n5350, C1 => n4160, C2 => 
                           n5351, A => n5352, ZN => n5343);
   U4436 : AOI22_X1 port map( A1 => n5353, A2 => n3616, B1 => n5354, B2 => 
                           n4000, ZN => n5352);
   U4437 : OAI221_X1 port map( B1 => n3777, B2 => n5355, C1 => n4161, C2 => 
                           n5356, A => n5357, ZN => n5342);
   U4438 : AOI22_X1 port map( A1 => n5358, A2 => n3617, B1 => n5359, B2 => 
                           n4001, ZN => n5357);
   U4439 : OAI221_X1 port map( B1 => n3778, B2 => n5360, C1 => n4162, C2 => 
                           n5361, A => n5362, ZN => n5341);
   U4440 : AOI22_X1 port map( A1 => n5363, A2 => n3618, B1 => n5364, B2 => 
                           n4002, ZN => n5362);
   U4441 : MUX2_X1 port map( A => OUT1_30_port, B => n5365, S => n5314, Z => 
                           n2556);
   U4442 : NAND2_X1 port map( A1 => n5366, A2 => n5367, ZN => n5365);
   U4443 : NOR4_X1 port map( A1 => n5368, A2 => n5369, A3 => n5370, A4 => n5371
                           , ZN => n5367);
   U4444 : OAI221_X1 port map( B1 => n2, B2 => n5321, C1 => n34, C2 => n5322, A
                           => n5372, ZN => n5371);
   U4445 : AOI22_X1 port map( A1 => n5324, A2 => n6093, B1 => n5325, B2 => 
                           n6094, ZN => n5372);
   U4446 : OAI221_X1 port map( B1 => n130, B2 => n5326, C1 => n162, C2 => n5327
                           , A => n5373, ZN => n5370);
   U4447 : AOI22_X1 port map( A1 => n5329, A2 => n6091, B1 => n5330, B2 => 
                           n6092, ZN => n5373);
   U4448 : OAI221_X1 port map( B1 => n290, B2 => n5331, C1 => n258, C2 => n5332
                           , A => n5374, ZN => n5369);
   U4449 : AOI22_X1 port map( A1 => n5334, A2 => n3967, B1 => n5335, B2 => 
                           n4351, ZN => n5374);
   U4450 : OAI221_X1 port map( B1 => n3779, B2 => n5336, C1 => n4163, C2 => 
                           n5337, A => n5375, ZN => n5368);
   U4451 : AOI22_X1 port map( A1 => n5339, A2 => n3619, B1 => n5340, B2 => 
                           n4003, ZN => n5375);
   U4452 : NOR4_X1 port map( A1 => n5376, A2 => n5377, A3 => n5378, A4 => n5379
                           , ZN => n5366);
   U4453 : OAI221_X1 port map( B1 => n3780, B2 => n5345, C1 => n4164, C2 => 
                           n5346, A => n5380, ZN => n5379);
   U4454 : AOI22_X1 port map( A1 => n5348, A2 => n3620, B1 => n5349, B2 => 
                           n4004, ZN => n5380);
   U4455 : OAI221_X1 port map( B1 => n3781, B2 => n5350, C1 => n4165, C2 => 
                           n5351, A => n5381, ZN => n5378);
   U4456 : AOI22_X1 port map( A1 => n5353, A2 => n3621, B1 => n5354, B2 => 
                           n4005, ZN => n5381);
   U4457 : OAI221_X1 port map( B1 => n3782, B2 => n5355, C1 => n4166, C2 => 
                           n5356, A => n5382, ZN => n5377);
   U4458 : AOI22_X1 port map( A1 => n5358, A2 => n3622, B1 => n5359, B2 => 
                           n4006, ZN => n5382);
   U4459 : OAI221_X1 port map( B1 => n3783, B2 => n5360, C1 => n4167, C2 => 
                           n5361, A => n5383, ZN => n5376);
   U4460 : AOI22_X1 port map( A1 => n5363, A2 => n3623, B1 => n5364, B2 => 
                           n4007, ZN => n5383);
   U4461 : MUX2_X1 port map( A => OUT1_29_port, B => n5384, S => n5314, Z => 
                           n2555);
   U4462 : NAND2_X1 port map( A1 => n5385, A2 => n5386, ZN => n5384);
   U4463 : NOR4_X1 port map( A1 => n5387, A2 => n5388, A3 => n5389, A4 => n5390
                           , ZN => n5386);
   U4464 : OAI221_X1 port map( B1 => n3, B2 => n5321, C1 => n35, C2 => n5322, A
                           => n5391, ZN => n5390);
   U4465 : AOI22_X1 port map( A1 => n5324, A2 => n6089, B1 => n5325, B2 => 
                           n6090, ZN => n5391);
   U4466 : OAI221_X1 port map( B1 => n131, B2 => n5326, C1 => n163, C2 => n5327
                           , A => n5392, ZN => n5389);
   U4467 : AOI22_X1 port map( A1 => n5329, A2 => n6087, B1 => n5330, B2 => 
                           n6088, ZN => n5392);
   U4468 : OAI221_X1 port map( B1 => n291, B2 => n5331, C1 => n259, C2 => n5332
                           , A => n5393, ZN => n5388);
   U4469 : AOI22_X1 port map( A1 => n5334, A2 => n3968, B1 => n5335, B2 => 
                           n4352, ZN => n5393);
   U4470 : OAI221_X1 port map( B1 => n3784, B2 => n5336, C1 => n4168, C2 => 
                           n5337, A => n5394, ZN => n5387);
   U4471 : AOI22_X1 port map( A1 => n5339, A2 => n3624, B1 => n5340, B2 => 
                           n4008, ZN => n5394);
   U4472 : NOR4_X1 port map( A1 => n5395, A2 => n5396, A3 => n5397, A4 => n5398
                           , ZN => n5385);
   U4473 : OAI221_X1 port map( B1 => n3785, B2 => n5345, C1 => n4169, C2 => 
                           n5346, A => n5399, ZN => n5398);
   U4474 : AOI22_X1 port map( A1 => n5348, A2 => n3625, B1 => n5349, B2 => 
                           n4009, ZN => n5399);
   U4475 : OAI221_X1 port map( B1 => n3786, B2 => n5350, C1 => n4170, C2 => 
                           n5351, A => n5400, ZN => n5397);
   U4476 : AOI22_X1 port map( A1 => n5353, A2 => n3626, B1 => n5354, B2 => 
                           n4010, ZN => n5400);
   U4477 : OAI221_X1 port map( B1 => n3787, B2 => n5355, C1 => n4171, C2 => 
                           n5356, A => n5401, ZN => n5396);
   U4478 : AOI22_X1 port map( A1 => n5358, A2 => n3627, B1 => n5359, B2 => 
                           n4011, ZN => n5401);
   U4479 : OAI221_X1 port map( B1 => n3788, B2 => n5360, C1 => n4172, C2 => 
                           n5361, A => n5402, ZN => n5395);
   U4480 : AOI22_X1 port map( A1 => n5363, A2 => n3628, B1 => n5364, B2 => 
                           n4012, ZN => n5402);
   U4481 : MUX2_X1 port map( A => OUT1_28_port, B => n5403, S => n5314, Z => 
                           n2554);
   U4482 : NAND2_X1 port map( A1 => n5404, A2 => n5405, ZN => n5403);
   U4483 : NOR4_X1 port map( A1 => n5406, A2 => n5407, A3 => n5408, A4 => n5409
                           , ZN => n5405);
   U4484 : OAI221_X1 port map( B1 => n4, B2 => n5321, C1 => n36, C2 => n5322, A
                           => n5410, ZN => n5409);
   U4485 : AOI22_X1 port map( A1 => n5324, A2 => n6085, B1 => n5325, B2 => 
                           n6086, ZN => n5410);
   U4486 : OAI221_X1 port map( B1 => n132, B2 => n5326, C1 => n164, C2 => n5327
                           , A => n5411, ZN => n5408);
   U4487 : AOI22_X1 port map( A1 => n5329, A2 => n6083, B1 => n5330, B2 => 
                           n6084, ZN => n5411);
   U4488 : OAI221_X1 port map( B1 => n292, B2 => n5331, C1 => n260, C2 => n5332
                           , A => n5412, ZN => n5407);
   U4489 : AOI22_X1 port map( A1 => n5334, A2 => n3969, B1 => n5335, B2 => 
                           n4353, ZN => n5412);
   U4490 : OAI221_X1 port map( B1 => n3789, B2 => n5336, C1 => n4173, C2 => 
                           n5337, A => n5413, ZN => n5406);
   U4491 : AOI22_X1 port map( A1 => n5339, A2 => n3629, B1 => n5340, B2 => 
                           n4013, ZN => n5413);
   U4492 : NOR4_X1 port map( A1 => n5414, A2 => n5415, A3 => n5416, A4 => n5417
                           , ZN => n5404);
   U4493 : OAI221_X1 port map( B1 => n3790, B2 => n5345, C1 => n4174, C2 => 
                           n5346, A => n5418, ZN => n5417);
   U4494 : AOI22_X1 port map( A1 => n5348, A2 => n3630, B1 => n5349, B2 => 
                           n4014, ZN => n5418);
   U4495 : OAI221_X1 port map( B1 => n3791, B2 => n5350, C1 => n4175, C2 => 
                           n5351, A => n5419, ZN => n5416);
   U4496 : AOI22_X1 port map( A1 => n5353, A2 => n3631, B1 => n5354, B2 => 
                           n4015, ZN => n5419);
   U4497 : OAI221_X1 port map( B1 => n3792, B2 => n5355, C1 => n4176, C2 => 
                           n5356, A => n5420, ZN => n5415);
   U4498 : AOI22_X1 port map( A1 => n5358, A2 => n3632, B1 => n5359, B2 => 
                           n4016, ZN => n5420);
   U4499 : OAI221_X1 port map( B1 => n3793, B2 => n5360, C1 => n4177, C2 => 
                           n5361, A => n5421, ZN => n5414);
   U4500 : AOI22_X1 port map( A1 => n5363, A2 => n3633, B1 => n5364, B2 => 
                           n4017, ZN => n5421);
   U4501 : MUX2_X1 port map( A => OUT1_27_port, B => n5422, S => n5314, Z => 
                           n2553);
   U4502 : NAND2_X1 port map( A1 => n5423, A2 => n5424, ZN => n5422);
   U4503 : NOR4_X1 port map( A1 => n5425, A2 => n5426, A3 => n5427, A4 => n5428
                           , ZN => n5424);
   U4504 : OAI221_X1 port map( B1 => n5, B2 => n5321, C1 => n37, C2 => n5322, A
                           => n5429, ZN => n5428);
   U4505 : AOI22_X1 port map( A1 => n5324, A2 => n6081, B1 => n5325, B2 => 
                           n6082, ZN => n5429);
   U4506 : OAI221_X1 port map( B1 => n133, B2 => n5326, C1 => n165, C2 => n5327
                           , A => n5430, ZN => n5427);
   U4507 : AOI22_X1 port map( A1 => n5329, A2 => n6079, B1 => n5330, B2 => 
                           n6080, ZN => n5430);
   U4508 : OAI221_X1 port map( B1 => n293, B2 => n5331, C1 => n261, C2 => n5332
                           , A => n5431, ZN => n5426);
   U4509 : AOI22_X1 port map( A1 => n5334, A2 => n3970, B1 => n5335, B2 => 
                           n4354, ZN => n5431);
   U4510 : OAI221_X1 port map( B1 => n3794, B2 => n5336, C1 => n4178, C2 => 
                           n5337, A => n5432, ZN => n5425);
   U4511 : AOI22_X1 port map( A1 => n5339, A2 => n3634, B1 => n5340, B2 => 
                           n4018, ZN => n5432);
   U4512 : NOR4_X1 port map( A1 => n5433, A2 => n5434, A3 => n5435, A4 => n5436
                           , ZN => n5423);
   U4513 : OAI221_X1 port map( B1 => n3795, B2 => n5345, C1 => n4179, C2 => 
                           n5346, A => n5437, ZN => n5436);
   U4514 : AOI22_X1 port map( A1 => n5348, A2 => n3635, B1 => n5349, B2 => 
                           n4019, ZN => n5437);
   U4515 : OAI221_X1 port map( B1 => n3796, B2 => n5350, C1 => n4180, C2 => 
                           n5351, A => n5438, ZN => n5435);
   U4516 : AOI22_X1 port map( A1 => n5353, A2 => n3636, B1 => n5354, B2 => 
                           n4020, ZN => n5438);
   U4517 : OAI221_X1 port map( B1 => n3797, B2 => n5355, C1 => n4181, C2 => 
                           n5356, A => n5439, ZN => n5434);
   U4518 : AOI22_X1 port map( A1 => n5358, A2 => n3637, B1 => n5359, B2 => 
                           n4021, ZN => n5439);
   U4519 : OAI221_X1 port map( B1 => n3798, B2 => n5360, C1 => n4182, C2 => 
                           n5361, A => n5440, ZN => n5433);
   U4520 : AOI22_X1 port map( A1 => n5363, A2 => n3638, B1 => n5364, B2 => 
                           n4022, ZN => n5440);
   U4521 : MUX2_X1 port map( A => OUT1_26_port, B => n5441, S => n5314, Z => 
                           n2552);
   U4522 : NAND2_X1 port map( A1 => n5442, A2 => n5443, ZN => n5441);
   U4523 : NOR4_X1 port map( A1 => n5444, A2 => n5445, A3 => n5446, A4 => n5447
                           , ZN => n5443);
   U4524 : OAI221_X1 port map( B1 => n6, B2 => n5321, C1 => n38, C2 => n5322, A
                           => n5448, ZN => n5447);
   U4525 : AOI22_X1 port map( A1 => n5324, A2 => n6077, B1 => n5325, B2 => 
                           n6078, ZN => n5448);
   U4526 : OAI221_X1 port map( B1 => n134, B2 => n5326, C1 => n166, C2 => n5327
                           , A => n5449, ZN => n5446);
   U4527 : AOI22_X1 port map( A1 => n5329, A2 => n6075, B1 => n5330, B2 => 
                           n6076, ZN => n5449);
   U4528 : OAI221_X1 port map( B1 => n294, B2 => n5331, C1 => n262, C2 => n5332
                           , A => n5450, ZN => n5445);
   U4529 : AOI22_X1 port map( A1 => n5334, A2 => n3971, B1 => n5335, B2 => 
                           n4355, ZN => n5450);
   U4530 : OAI221_X1 port map( B1 => n3799, B2 => n5336, C1 => n4183, C2 => 
                           n5337, A => n5451, ZN => n5444);
   U4531 : AOI22_X1 port map( A1 => n5339, A2 => n3639, B1 => n5340, B2 => 
                           n4023, ZN => n5451);
   U4532 : NOR4_X1 port map( A1 => n5452, A2 => n5453, A3 => n5454, A4 => n5455
                           , ZN => n5442);
   U4533 : OAI221_X1 port map( B1 => n3800, B2 => n5345, C1 => n4184, C2 => 
                           n5346, A => n5456, ZN => n5455);
   U4534 : AOI22_X1 port map( A1 => n5348, A2 => n3640, B1 => n5349, B2 => 
                           n4024, ZN => n5456);
   U4535 : OAI221_X1 port map( B1 => n3801, B2 => n5350, C1 => n4185, C2 => 
                           n5351, A => n5457, ZN => n5454);
   U4536 : AOI22_X1 port map( A1 => n5353, A2 => n3641, B1 => n5354, B2 => 
                           n4025, ZN => n5457);
   U4537 : OAI221_X1 port map( B1 => n3802, B2 => n5355, C1 => n4186, C2 => 
                           n5356, A => n5458, ZN => n5453);
   U4538 : AOI22_X1 port map( A1 => n5358, A2 => n3642, B1 => n5359, B2 => 
                           n4026, ZN => n5458);
   U4539 : OAI221_X1 port map( B1 => n3803, B2 => n5360, C1 => n4187, C2 => 
                           n5361, A => n5459, ZN => n5452);
   U4540 : AOI22_X1 port map( A1 => n5363, A2 => n3643, B1 => n5364, B2 => 
                           n4027, ZN => n5459);
   U4541 : MUX2_X1 port map( A => OUT1_25_port, B => n5460, S => n5314, Z => 
                           n2551);
   U4542 : NAND2_X1 port map( A1 => n5461, A2 => n5462, ZN => n5460);
   U4543 : NOR4_X1 port map( A1 => n5463, A2 => n5464, A3 => n5465, A4 => n5466
                           , ZN => n5462);
   U4544 : OAI221_X1 port map( B1 => n7, B2 => n5321, C1 => n39, C2 => n5322, A
                           => n5467, ZN => n5466);
   U4545 : AOI22_X1 port map( A1 => n5324, A2 => n6073, B1 => n5325, B2 => 
                           n6074, ZN => n5467);
   U4546 : OAI221_X1 port map( B1 => n135, B2 => n5326, C1 => n167, C2 => n5327
                           , A => n5468, ZN => n5465);
   U4547 : AOI22_X1 port map( A1 => n5329, A2 => n6071, B1 => n5330, B2 => 
                           n6072, ZN => n5468);
   U4548 : OAI221_X1 port map( B1 => n295, B2 => n5331, C1 => n263, C2 => n5332
                           , A => n5469, ZN => n5464);
   U4549 : AOI22_X1 port map( A1 => n5334, A2 => n3972, B1 => n5335, B2 => 
                           n4356, ZN => n5469);
   U4550 : OAI221_X1 port map( B1 => n3804, B2 => n5336, C1 => n4188, C2 => 
                           n5337, A => n5470, ZN => n5463);
   U4551 : AOI22_X1 port map( A1 => n5339, A2 => n3644, B1 => n5340, B2 => 
                           n4028, ZN => n5470);
   U4552 : NOR4_X1 port map( A1 => n5471, A2 => n5472, A3 => n5473, A4 => n5474
                           , ZN => n5461);
   U4553 : OAI221_X1 port map( B1 => n3805, B2 => n5345, C1 => n4189, C2 => 
                           n5346, A => n5475, ZN => n5474);
   U4554 : AOI22_X1 port map( A1 => n5348, A2 => n3645, B1 => n5349, B2 => 
                           n4029, ZN => n5475);
   U4555 : OAI221_X1 port map( B1 => n3806, B2 => n5350, C1 => n4190, C2 => 
                           n5351, A => n5476, ZN => n5473);
   U4556 : AOI22_X1 port map( A1 => n5353, A2 => n3646, B1 => n5354, B2 => 
                           n4030, ZN => n5476);
   U4557 : OAI221_X1 port map( B1 => n3807, B2 => n5355, C1 => n4191, C2 => 
                           n5356, A => n5477, ZN => n5472);
   U4558 : AOI22_X1 port map( A1 => n5358, A2 => n3647, B1 => n5359, B2 => 
                           n4031, ZN => n5477);
   U4559 : OAI221_X1 port map( B1 => n3808, B2 => n5360, C1 => n4192, C2 => 
                           n5361, A => n5478, ZN => n5471);
   U4560 : AOI22_X1 port map( A1 => n5363, A2 => n3648, B1 => n5364, B2 => 
                           n4032, ZN => n5478);
   U4561 : MUX2_X1 port map( A => OUT1_24_port, B => n5479, S => n5314, Z => 
                           n2550);
   U4562 : NAND2_X1 port map( A1 => n5480, A2 => n5481, ZN => n5479);
   U4563 : NOR4_X1 port map( A1 => n5482, A2 => n5483, A3 => n5484, A4 => n5485
                           , ZN => n5481);
   U4564 : OAI221_X1 port map( B1 => n8, B2 => n5321, C1 => n40, C2 => n5322, A
                           => n5486, ZN => n5485);
   U4565 : AOI22_X1 port map( A1 => n5324, A2 => n6069, B1 => n5325, B2 => 
                           n6070, ZN => n5486);
   U4566 : OAI221_X1 port map( B1 => n136, B2 => n5326, C1 => n168, C2 => n5327
                           , A => n5487, ZN => n5484);
   U4567 : AOI22_X1 port map( A1 => n5329, A2 => n6067, B1 => n5330, B2 => 
                           n6068, ZN => n5487);
   U4568 : OAI221_X1 port map( B1 => n296, B2 => n5331, C1 => n264, C2 => n5332
                           , A => n5488, ZN => n5483);
   U4569 : AOI22_X1 port map( A1 => n5334, A2 => n3973, B1 => n5335, B2 => 
                           n4357, ZN => n5488);
   U4570 : OAI221_X1 port map( B1 => n3809, B2 => n5336, C1 => n4193, C2 => 
                           n5337, A => n5489, ZN => n5482);
   U4571 : AOI22_X1 port map( A1 => n5339, A2 => n3649, B1 => n5340, B2 => 
                           n4033, ZN => n5489);
   U4572 : NOR4_X1 port map( A1 => n5490, A2 => n5491, A3 => n5492, A4 => n5493
                           , ZN => n5480);
   U4573 : OAI221_X1 port map( B1 => n3810, B2 => n5345, C1 => n4194, C2 => 
                           n5346, A => n5494, ZN => n5493);
   U4574 : AOI22_X1 port map( A1 => n5348, A2 => n3650, B1 => n5349, B2 => 
                           n4034, ZN => n5494);
   U4575 : OAI221_X1 port map( B1 => n3811, B2 => n5350, C1 => n4195, C2 => 
                           n5351, A => n5495, ZN => n5492);
   U4576 : AOI22_X1 port map( A1 => n5353, A2 => n3651, B1 => n5354, B2 => 
                           n4035, ZN => n5495);
   U4577 : OAI221_X1 port map( B1 => n3812, B2 => n5355, C1 => n4196, C2 => 
                           n5356, A => n5496, ZN => n5491);
   U4578 : AOI22_X1 port map( A1 => n5358, A2 => n3652, B1 => n5359, B2 => 
                           n4036, ZN => n5496);
   U4579 : OAI221_X1 port map( B1 => n3813, B2 => n5360, C1 => n4197, C2 => 
                           n5361, A => n5497, ZN => n5490);
   U4580 : AOI22_X1 port map( A1 => n5363, A2 => n3653, B1 => n5364, B2 => 
                           n4037, ZN => n5497);
   U4581 : MUX2_X1 port map( A => OUT1_23_port, B => n5498, S => n5314, Z => 
                           n2549);
   U4582 : NAND2_X1 port map( A1 => n5499, A2 => n5500, ZN => n5498);
   U4583 : NOR4_X1 port map( A1 => n5501, A2 => n5502, A3 => n5503, A4 => n5504
                           , ZN => n5500);
   U4584 : OAI221_X1 port map( B1 => n9, B2 => n5321, C1 => n41, C2 => n5322, A
                           => n5505, ZN => n5504);
   U4585 : AOI22_X1 port map( A1 => n5324, A2 => n6065, B1 => n5325, B2 => 
                           n6066, ZN => n5505);
   U4586 : OAI221_X1 port map( B1 => n137, B2 => n5326, C1 => n169, C2 => n5327
                           , A => n5506, ZN => n5503);
   U4587 : AOI22_X1 port map( A1 => n5329, A2 => n6063, B1 => n5330, B2 => 
                           n6064, ZN => n5506);
   U4588 : OAI221_X1 port map( B1 => n297, B2 => n5331, C1 => n265, C2 => n5332
                           , A => n5507, ZN => n5502);
   U4589 : AOI22_X1 port map( A1 => n5334, A2 => n3974, B1 => n5335, B2 => 
                           n4358, ZN => n5507);
   U4590 : OAI221_X1 port map( B1 => n3814, B2 => n5336, C1 => n4198, C2 => 
                           n5337, A => n5508, ZN => n5501);
   U4591 : AOI22_X1 port map( A1 => n5339, A2 => n3654, B1 => n5340, B2 => 
                           n4038, ZN => n5508);
   U4592 : NOR4_X1 port map( A1 => n5509, A2 => n5510, A3 => n5511, A4 => n5512
                           , ZN => n5499);
   U4593 : OAI221_X1 port map( B1 => n3815, B2 => n5345, C1 => n4199, C2 => 
                           n5346, A => n5513, ZN => n5512);
   U4594 : AOI22_X1 port map( A1 => n5348, A2 => n3655, B1 => n5349, B2 => 
                           n4039, ZN => n5513);
   U4595 : OAI221_X1 port map( B1 => n3816, B2 => n5350, C1 => n4200, C2 => 
                           n5351, A => n5514, ZN => n5511);
   U4596 : AOI22_X1 port map( A1 => n5353, A2 => n3656, B1 => n5354, B2 => 
                           n4040, ZN => n5514);
   U4597 : OAI221_X1 port map( B1 => n3817, B2 => n5355, C1 => n4201, C2 => 
                           n5356, A => n5515, ZN => n5510);
   U4598 : AOI22_X1 port map( A1 => n5358, A2 => n3657, B1 => n5359, B2 => 
                           n4041, ZN => n5515);
   U4599 : OAI221_X1 port map( B1 => n3818, B2 => n5360, C1 => n4202, C2 => 
                           n5361, A => n5516, ZN => n5509);
   U4600 : AOI22_X1 port map( A1 => n5363, A2 => n3658, B1 => n5364, B2 => 
                           n4042, ZN => n5516);
   U4601 : MUX2_X1 port map( A => OUT1_22_port, B => n5517, S => n5314, Z => 
                           n2548);
   U4602 : NAND2_X1 port map( A1 => n5518, A2 => n5519, ZN => n5517);
   U4603 : NOR4_X1 port map( A1 => n5520, A2 => n5521, A3 => n5522, A4 => n5523
                           , ZN => n5519);
   U4604 : OAI221_X1 port map( B1 => n10, B2 => n5321, C1 => n42, C2 => n5322, 
                           A => n5524, ZN => n5523);
   U4605 : AOI22_X1 port map( A1 => n5324, A2 => n6061, B1 => n5325, B2 => 
                           n6062, ZN => n5524);
   U4606 : OAI221_X1 port map( B1 => n138, B2 => n5326, C1 => n170, C2 => n5327
                           , A => n5525, ZN => n5522);
   U4607 : AOI22_X1 port map( A1 => n5329, A2 => n6059, B1 => n5330, B2 => 
                           n6060, ZN => n5525);
   U4608 : OAI221_X1 port map( B1 => n298, B2 => n5331, C1 => n266, C2 => n5332
                           , A => n5526, ZN => n5521);
   U4609 : AOI22_X1 port map( A1 => n5334, A2 => n3975, B1 => n5335, B2 => 
                           n4359, ZN => n5526);
   U4610 : OAI221_X1 port map( B1 => n3819, B2 => n5336, C1 => n4203, C2 => 
                           n5337, A => n5527, ZN => n5520);
   U4611 : AOI22_X1 port map( A1 => n5339, A2 => n3659, B1 => n5340, B2 => 
                           n4043, ZN => n5527);
   U4612 : NOR4_X1 port map( A1 => n5528, A2 => n5529, A3 => n5530, A4 => n5531
                           , ZN => n5518);
   U4613 : OAI221_X1 port map( B1 => n3820, B2 => n5345, C1 => n4204, C2 => 
                           n5346, A => n5532, ZN => n5531);
   U4614 : AOI22_X1 port map( A1 => n5348, A2 => n3660, B1 => n5349, B2 => 
                           n4044, ZN => n5532);
   U4615 : OAI221_X1 port map( B1 => n3821, B2 => n5350, C1 => n4205, C2 => 
                           n5351, A => n5533, ZN => n5530);
   U4616 : AOI22_X1 port map( A1 => n5353, A2 => n3661, B1 => n5354, B2 => 
                           n4045, ZN => n5533);
   U4617 : OAI221_X1 port map( B1 => n3822, B2 => n5355, C1 => n4206, C2 => 
                           n5356, A => n5534, ZN => n5529);
   U4618 : AOI22_X1 port map( A1 => n5358, A2 => n3662, B1 => n5359, B2 => 
                           n4046, ZN => n5534);
   U4619 : OAI221_X1 port map( B1 => n3823, B2 => n5360, C1 => n4207, C2 => 
                           n5361, A => n5535, ZN => n5528);
   U4620 : AOI22_X1 port map( A1 => n5363, A2 => n3663, B1 => n5364, B2 => 
                           n4047, ZN => n5535);
   U4621 : MUX2_X1 port map( A => OUT1_21_port, B => n5536, S => n5314, Z => 
                           n2547);
   U4622 : NAND2_X1 port map( A1 => n5537, A2 => n5538, ZN => n5536);
   U4623 : NOR4_X1 port map( A1 => n5539, A2 => n5540, A3 => n5541, A4 => n5542
                           , ZN => n5538);
   U4624 : OAI221_X1 port map( B1 => n11, B2 => n5321, C1 => n43, C2 => n5322, 
                           A => n5543, ZN => n5542);
   U4625 : AOI22_X1 port map( A1 => n5324, A2 => n6057, B1 => n5325, B2 => 
                           n6058, ZN => n5543);
   U4626 : OAI221_X1 port map( B1 => n139, B2 => n5326, C1 => n171, C2 => n5327
                           , A => n5544, ZN => n5541);
   U4627 : AOI22_X1 port map( A1 => n5329, A2 => n6055, B1 => n5330, B2 => 
                           n6056, ZN => n5544);
   U4628 : OAI221_X1 port map( B1 => n299, B2 => n5331, C1 => n267, C2 => n5332
                           , A => n5545, ZN => n5540);
   U4629 : AOI22_X1 port map( A1 => n5334, A2 => n3976, B1 => n5335, B2 => 
                           n4360, ZN => n5545);
   U4630 : OAI221_X1 port map( B1 => n3824, B2 => n5336, C1 => n4208, C2 => 
                           n5337, A => n5546, ZN => n5539);
   U4631 : AOI22_X1 port map( A1 => n5339, A2 => n3664, B1 => n5340, B2 => 
                           n4048, ZN => n5546);
   U4632 : NOR4_X1 port map( A1 => n5547, A2 => n5548, A3 => n5549, A4 => n5550
                           , ZN => n5537);
   U4633 : OAI221_X1 port map( B1 => n3825, B2 => n5345, C1 => n4209, C2 => 
                           n5346, A => n5551, ZN => n5550);
   U4634 : AOI22_X1 port map( A1 => n5348, A2 => n3665, B1 => n5349, B2 => 
                           n4049, ZN => n5551);
   U4635 : OAI221_X1 port map( B1 => n3826, B2 => n5350, C1 => n4210, C2 => 
                           n5351, A => n5552, ZN => n5549);
   U4636 : AOI22_X1 port map( A1 => n5353, A2 => n3666, B1 => n5354, B2 => 
                           n4050, ZN => n5552);
   U4637 : OAI221_X1 port map( B1 => n3827, B2 => n5355, C1 => n4211, C2 => 
                           n5356, A => n5553, ZN => n5548);
   U4638 : AOI22_X1 port map( A1 => n5358, A2 => n3667, B1 => n5359, B2 => 
                           n4051, ZN => n5553);
   U4639 : OAI221_X1 port map( B1 => n3828, B2 => n5360, C1 => n4212, C2 => 
                           n5361, A => n5554, ZN => n5547);
   U4640 : AOI22_X1 port map( A1 => n5363, A2 => n3668, B1 => n5364, B2 => 
                           n4052, ZN => n5554);
   U4641 : MUX2_X1 port map( A => OUT1_20_port, B => n5555, S => n5314, Z => 
                           n2546);
   U4642 : NAND2_X1 port map( A1 => n5556, A2 => n5557, ZN => n5555);
   U4643 : NOR4_X1 port map( A1 => n5558, A2 => n5559, A3 => n5560, A4 => n5561
                           , ZN => n5557);
   U4644 : OAI221_X1 port map( B1 => n12, B2 => n5321, C1 => n44, C2 => n5322, 
                           A => n5562, ZN => n5561);
   U4645 : AOI22_X1 port map( A1 => n5324, A2 => n6053, B1 => n5325, B2 => 
                           n6054, ZN => n5562);
   U4646 : OAI221_X1 port map( B1 => n140, B2 => n5326, C1 => n172, C2 => n5327
                           , A => n5563, ZN => n5560);
   U4647 : AOI22_X1 port map( A1 => n5329, A2 => n6051, B1 => n5330, B2 => 
                           n6052, ZN => n5563);
   U4648 : OAI221_X1 port map( B1 => n300, B2 => n5331, C1 => n268, C2 => n5332
                           , A => n5564, ZN => n5559);
   U4649 : AOI22_X1 port map( A1 => n5334, A2 => n3977, B1 => n5335, B2 => 
                           n4361, ZN => n5564);
   U4650 : OAI221_X1 port map( B1 => n3829, B2 => n5336, C1 => n4213, C2 => 
                           n5337, A => n5565, ZN => n5558);
   U4651 : AOI22_X1 port map( A1 => n5339, A2 => n3669, B1 => n5340, B2 => 
                           n4053, ZN => n5565);
   U4652 : NOR4_X1 port map( A1 => n5566, A2 => n5567, A3 => n5568, A4 => n5569
                           , ZN => n5556);
   U4653 : OAI221_X1 port map( B1 => n3830, B2 => n5345, C1 => n4214, C2 => 
                           n5346, A => n5570, ZN => n5569);
   U4654 : AOI22_X1 port map( A1 => n5348, A2 => n3670, B1 => n5349, B2 => 
                           n4054, ZN => n5570);
   U4655 : OAI221_X1 port map( B1 => n3831, B2 => n5350, C1 => n4215, C2 => 
                           n5351, A => n5571, ZN => n5568);
   U4656 : AOI22_X1 port map( A1 => n5353, A2 => n3671, B1 => n5354, B2 => 
                           n4055, ZN => n5571);
   U4657 : OAI221_X1 port map( B1 => n3832, B2 => n5355, C1 => n4216, C2 => 
                           n5356, A => n5572, ZN => n5567);
   U4658 : AOI22_X1 port map( A1 => n5358, A2 => n3672, B1 => n5359, B2 => 
                           n4056, ZN => n5572);
   U4659 : OAI221_X1 port map( B1 => n3833, B2 => n5360, C1 => n4217, C2 => 
                           n5361, A => n5573, ZN => n5566);
   U4660 : AOI22_X1 port map( A1 => n5363, A2 => n3673, B1 => n5364, B2 => 
                           n4057, ZN => n5573);
   U4661 : MUX2_X1 port map( A => OUT1_19_port, B => n5574, S => n5314, Z => 
                           n2545);
   U4662 : NAND2_X1 port map( A1 => n5575, A2 => n5576, ZN => n5574);
   U4663 : NOR4_X1 port map( A1 => n5577, A2 => n5578, A3 => n5579, A4 => n5580
                           , ZN => n5576);
   U4664 : OAI221_X1 port map( B1 => n13, B2 => n5321, C1 => n45, C2 => n5322, 
                           A => n5581, ZN => n5580);
   U4665 : AOI22_X1 port map( A1 => n5324, A2 => n6049, B1 => n5325, B2 => 
                           n6050, ZN => n5581);
   U4666 : OAI221_X1 port map( B1 => n141, B2 => n5326, C1 => n173, C2 => n5327
                           , A => n5582, ZN => n5579);
   U4667 : AOI22_X1 port map( A1 => n5329, A2 => n6047, B1 => n5330, B2 => 
                           n6048, ZN => n5582);
   U4668 : OAI221_X1 port map( B1 => n301, B2 => n5331, C1 => n269, C2 => n5332
                           , A => n5583, ZN => n5578);
   U4669 : AOI22_X1 port map( A1 => n5334, A2 => n3978, B1 => n5335, B2 => 
                           n4362, ZN => n5583);
   U4670 : OAI221_X1 port map( B1 => n3834, B2 => n5336, C1 => n4218, C2 => 
                           n5337, A => n5584, ZN => n5577);
   U4671 : AOI22_X1 port map( A1 => n5339, A2 => n3674, B1 => n5340, B2 => 
                           n4058, ZN => n5584);
   U4672 : NOR4_X1 port map( A1 => n5585, A2 => n5586, A3 => n5587, A4 => n5588
                           , ZN => n5575);
   U4673 : OAI221_X1 port map( B1 => n3835, B2 => n5345, C1 => n4219, C2 => 
                           n5346, A => n5589, ZN => n5588);
   U4674 : AOI22_X1 port map( A1 => n5348, A2 => n3675, B1 => n5349, B2 => 
                           n4059, ZN => n5589);
   U4675 : OAI221_X1 port map( B1 => n3836, B2 => n5350, C1 => n4220, C2 => 
                           n5351, A => n5590, ZN => n5587);
   U4676 : AOI22_X1 port map( A1 => n5353, A2 => n3676, B1 => n5354, B2 => 
                           n4060, ZN => n5590);
   U4677 : OAI221_X1 port map( B1 => n3837, B2 => n5355, C1 => n4221, C2 => 
                           n5356, A => n5591, ZN => n5586);
   U4678 : AOI22_X1 port map( A1 => n5358, A2 => n3677, B1 => n5359, B2 => 
                           n4061, ZN => n5591);
   U4679 : OAI221_X1 port map( B1 => n3838, B2 => n5360, C1 => n4222, C2 => 
                           n5361, A => n5592, ZN => n5585);
   U4680 : AOI22_X1 port map( A1 => n5363, A2 => n3678, B1 => n5364, B2 => 
                           n4062, ZN => n5592);
   U4681 : MUX2_X1 port map( A => OUT1_18_port, B => n5593, S => n5314, Z => 
                           n2544);
   U4682 : NAND2_X1 port map( A1 => n5594, A2 => n5595, ZN => n5593);
   U4683 : NOR4_X1 port map( A1 => n5596, A2 => n5597, A3 => n5598, A4 => n5599
                           , ZN => n5595);
   U4684 : OAI221_X1 port map( B1 => n14, B2 => n5321, C1 => n46, C2 => n5322, 
                           A => n5600, ZN => n5599);
   U4685 : AOI22_X1 port map( A1 => n5324, A2 => n6045, B1 => n5325, B2 => 
                           n6046, ZN => n5600);
   U4686 : OAI221_X1 port map( B1 => n142, B2 => n5326, C1 => n174, C2 => n5327
                           , A => n5601, ZN => n5598);
   U4687 : AOI22_X1 port map( A1 => n5329, A2 => n6043, B1 => n5330, B2 => 
                           n6044, ZN => n5601);
   U4688 : OAI221_X1 port map( B1 => n302, B2 => n5331, C1 => n270, C2 => n5332
                           , A => n5602, ZN => n5597);
   U4689 : AOI22_X1 port map( A1 => n5334, A2 => n3979, B1 => n5335, B2 => 
                           n4363, ZN => n5602);
   U4690 : OAI221_X1 port map( B1 => n3839, B2 => n5336, C1 => n4223, C2 => 
                           n5337, A => n5603, ZN => n5596);
   U4691 : AOI22_X1 port map( A1 => n5339, A2 => n3679, B1 => n5340, B2 => 
                           n4063, ZN => n5603);
   U4692 : NOR4_X1 port map( A1 => n5604, A2 => n5605, A3 => n5606, A4 => n5607
                           , ZN => n5594);
   U4693 : OAI221_X1 port map( B1 => n3840, B2 => n5345, C1 => n4224, C2 => 
                           n5346, A => n5608, ZN => n5607);
   U4694 : AOI22_X1 port map( A1 => n5348, A2 => n3680, B1 => n5349, B2 => 
                           n4064, ZN => n5608);
   U4695 : OAI221_X1 port map( B1 => n3841, B2 => n5350, C1 => n4225, C2 => 
                           n5351, A => n5609, ZN => n5606);
   U4696 : AOI22_X1 port map( A1 => n5353, A2 => n3681, B1 => n5354, B2 => 
                           n4065, ZN => n5609);
   U4697 : OAI221_X1 port map( B1 => n3842, B2 => n5355, C1 => n4226, C2 => 
                           n5356, A => n5610, ZN => n5605);
   U4698 : AOI22_X1 port map( A1 => n5358, A2 => n3682, B1 => n5359, B2 => 
                           n4066, ZN => n5610);
   U4699 : OAI221_X1 port map( B1 => n3843, B2 => n5360, C1 => n4227, C2 => 
                           n5361, A => n5611, ZN => n5604);
   U4700 : AOI22_X1 port map( A1 => n5363, A2 => n3683, B1 => n5364, B2 => 
                           n4067, ZN => n5611);
   U4701 : MUX2_X1 port map( A => OUT1_17_port, B => n5612, S => n5314, Z => 
                           n2543);
   U4702 : NAND2_X1 port map( A1 => n5613, A2 => n5614, ZN => n5612);
   U4703 : NOR4_X1 port map( A1 => n5615, A2 => n5616, A3 => n5617, A4 => n5618
                           , ZN => n5614);
   U4704 : OAI221_X1 port map( B1 => n15, B2 => n5321, C1 => n47, C2 => n5322, 
                           A => n5619, ZN => n5618);
   U4705 : AOI22_X1 port map( A1 => n5324, A2 => n6041, B1 => n5325, B2 => 
                           n6042, ZN => n5619);
   U4706 : OAI221_X1 port map( B1 => n143, B2 => n5326, C1 => n175, C2 => n5327
                           , A => n5620, ZN => n5617);
   U4707 : AOI22_X1 port map( A1 => n5329, A2 => n6039, B1 => n5330, B2 => 
                           n6040, ZN => n5620);
   U4708 : OAI221_X1 port map( B1 => n303, B2 => n5331, C1 => n271, C2 => n5332
                           , A => n5621, ZN => n5616);
   U4709 : AOI22_X1 port map( A1 => n5334, A2 => n3980, B1 => n5335, B2 => 
                           n4364, ZN => n5621);
   U4710 : OAI221_X1 port map( B1 => n3844, B2 => n5336, C1 => n4228, C2 => 
                           n5337, A => n5622, ZN => n5615);
   U4711 : AOI22_X1 port map( A1 => n5339, A2 => n3684, B1 => n5340, B2 => 
                           n4068, ZN => n5622);
   U4712 : NOR4_X1 port map( A1 => n5623, A2 => n5624, A3 => n5625, A4 => n5626
                           , ZN => n5613);
   U4713 : OAI221_X1 port map( B1 => n3845, B2 => n5345, C1 => n4229, C2 => 
                           n5346, A => n5627, ZN => n5626);
   U4714 : AOI22_X1 port map( A1 => n5348, A2 => n3685, B1 => n5349, B2 => 
                           n4069, ZN => n5627);
   U4715 : OAI221_X1 port map( B1 => n3846, B2 => n5350, C1 => n4230, C2 => 
                           n5351, A => n5628, ZN => n5625);
   U4716 : AOI22_X1 port map( A1 => n5353, A2 => n3686, B1 => n5354, B2 => 
                           n4070, ZN => n5628);
   U4717 : OAI221_X1 port map( B1 => n3847, B2 => n5355, C1 => n4231, C2 => 
                           n5356, A => n5629, ZN => n5624);
   U4718 : AOI22_X1 port map( A1 => n5358, A2 => n3687, B1 => n5359, B2 => 
                           n4071, ZN => n5629);
   U4719 : OAI221_X1 port map( B1 => n3848, B2 => n5360, C1 => n4232, C2 => 
                           n5361, A => n5630, ZN => n5623);
   U4720 : AOI22_X1 port map( A1 => n5363, A2 => n3688, B1 => n5364, B2 => 
                           n4072, ZN => n5630);
   U4721 : MUX2_X1 port map( A => OUT1_16_port, B => n5631, S => n5314, Z => 
                           n2542);
   U4722 : NAND2_X1 port map( A1 => n5632, A2 => n5633, ZN => n5631);
   U4723 : NOR4_X1 port map( A1 => n5634, A2 => n5635, A3 => n5636, A4 => n5637
                           , ZN => n5633);
   U4724 : OAI221_X1 port map( B1 => n16, B2 => n5321, C1 => n48, C2 => n5322, 
                           A => n5638, ZN => n5637);
   U4725 : AOI22_X1 port map( A1 => n5324, A2 => n6037, B1 => n5325, B2 => 
                           n6038, ZN => n5638);
   U4726 : OAI221_X1 port map( B1 => n144, B2 => n5326, C1 => n176, C2 => n5327
                           , A => n5639, ZN => n5636);
   U4727 : AOI22_X1 port map( A1 => n5329, A2 => n6035, B1 => n5330, B2 => 
                           n6036, ZN => n5639);
   U4728 : OAI221_X1 port map( B1 => n304, B2 => n5331, C1 => n272, C2 => n5332
                           , A => n5640, ZN => n5635);
   U4729 : AOI22_X1 port map( A1 => n5334, A2 => n3981, B1 => n5335, B2 => 
                           n4365, ZN => n5640);
   U4730 : OAI221_X1 port map( B1 => n3849, B2 => n5336, C1 => n4233, C2 => 
                           n5337, A => n5641, ZN => n5634);
   U4731 : AOI22_X1 port map( A1 => n5339, A2 => n3689, B1 => n5340, B2 => 
                           n4073, ZN => n5641);
   U4732 : NOR4_X1 port map( A1 => n5642, A2 => n5643, A3 => n5644, A4 => n5645
                           , ZN => n5632);
   U4733 : OAI221_X1 port map( B1 => n3850, B2 => n5345, C1 => n4234, C2 => 
                           n5346, A => n5646, ZN => n5645);
   U4734 : AOI22_X1 port map( A1 => n5348, A2 => n3690, B1 => n5349, B2 => 
                           n4074, ZN => n5646);
   U4735 : OAI221_X1 port map( B1 => n3851, B2 => n5350, C1 => n4235, C2 => 
                           n5351, A => n5647, ZN => n5644);
   U4736 : AOI22_X1 port map( A1 => n5353, A2 => n3691, B1 => n5354, B2 => 
                           n4075, ZN => n5647);
   U4737 : OAI221_X1 port map( B1 => n3852, B2 => n5355, C1 => n4236, C2 => 
                           n5356, A => n5648, ZN => n5643);
   U4738 : AOI22_X1 port map( A1 => n5358, A2 => n3692, B1 => n5359, B2 => 
                           n4076, ZN => n5648);
   U4739 : OAI221_X1 port map( B1 => n3853, B2 => n5360, C1 => n4237, C2 => 
                           n5361, A => n5649, ZN => n5642);
   U4740 : AOI22_X1 port map( A1 => n5363, A2 => n3693, B1 => n5364, B2 => 
                           n4077, ZN => n5649);
   U4741 : MUX2_X1 port map( A => OUT1_15_port, B => n5650, S => n5314, Z => 
                           n2541);
   U4742 : NAND2_X1 port map( A1 => n5651, A2 => n5652, ZN => n5650);
   U4743 : NOR4_X1 port map( A1 => n5653, A2 => n5654, A3 => n5655, A4 => n5656
                           , ZN => n5652);
   U4744 : OAI221_X1 port map( B1 => n17, B2 => n5321, C1 => n49, C2 => n5322, 
                           A => n5657, ZN => n5656);
   U4745 : AOI22_X1 port map( A1 => n5324, A2 => n6033, B1 => n5325, B2 => 
                           n6034, ZN => n5657);
   U4746 : OAI221_X1 port map( B1 => n145, B2 => n5326, C1 => n177, C2 => n5327
                           , A => n5658, ZN => n5655);
   U4747 : AOI22_X1 port map( A1 => n5329, A2 => n6031, B1 => n5330, B2 => 
                           n6032, ZN => n5658);
   U4748 : OAI221_X1 port map( B1 => n305, B2 => n5331, C1 => n273, C2 => n5332
                           , A => n5659, ZN => n5654);
   U4749 : AOI22_X1 port map( A1 => n5334, A2 => n3982, B1 => n5335, B2 => 
                           n4366, ZN => n5659);
   U4750 : OAI221_X1 port map( B1 => n3854, B2 => n5336, C1 => n4238, C2 => 
                           n5337, A => n5660, ZN => n5653);
   U4751 : AOI22_X1 port map( A1 => n5339, A2 => n3694, B1 => n5340, B2 => 
                           n4078, ZN => n5660);
   U4752 : NOR4_X1 port map( A1 => n5661, A2 => n5662, A3 => n5663, A4 => n5664
                           , ZN => n5651);
   U4753 : OAI221_X1 port map( B1 => n3855, B2 => n5345, C1 => n4239, C2 => 
                           n5346, A => n5665, ZN => n5664);
   U4754 : AOI22_X1 port map( A1 => n5348, A2 => n3695, B1 => n5349, B2 => 
                           n4079, ZN => n5665);
   U4755 : OAI221_X1 port map( B1 => n3856, B2 => n5350, C1 => n4240, C2 => 
                           n5351, A => n5666, ZN => n5663);
   U4756 : AOI22_X1 port map( A1 => n5353, A2 => n3696, B1 => n5354, B2 => 
                           n4080, ZN => n5666);
   U4757 : OAI221_X1 port map( B1 => n3857, B2 => n5355, C1 => n4241, C2 => 
                           n5356, A => n5667, ZN => n5662);
   U4758 : AOI22_X1 port map( A1 => n5358, A2 => n3697, B1 => n5359, B2 => 
                           n4081, ZN => n5667);
   U4759 : OAI221_X1 port map( B1 => n3858, B2 => n5360, C1 => n4242, C2 => 
                           n5361, A => n5668, ZN => n5661);
   U4760 : AOI22_X1 port map( A1 => n5363, A2 => n3698, B1 => n5364, B2 => 
                           n4082, ZN => n5668);
   U4761 : MUX2_X1 port map( A => OUT1_14_port, B => n5669, S => n5314, Z => 
                           n2540);
   U4762 : NAND2_X1 port map( A1 => n5670, A2 => n5671, ZN => n5669);
   U4763 : NOR4_X1 port map( A1 => n5672, A2 => n5673, A3 => n5674, A4 => n5675
                           , ZN => n5671);
   U4764 : OAI221_X1 port map( B1 => n18, B2 => n5321, C1 => n50, C2 => n5322, 
                           A => n5676, ZN => n5675);
   U4765 : AOI22_X1 port map( A1 => n5324, A2 => n6029, B1 => n5325, B2 => 
                           n6030, ZN => n5676);
   U4766 : OAI221_X1 port map( B1 => n146, B2 => n5326, C1 => n178, C2 => n5327
                           , A => n5677, ZN => n5674);
   U4767 : AOI22_X1 port map( A1 => n5329, A2 => n6027, B1 => n5330, B2 => 
                           n6028, ZN => n5677);
   U4768 : OAI221_X1 port map( B1 => n306, B2 => n5331, C1 => n274, C2 => n5332
                           , A => n5678, ZN => n5673);
   U4769 : AOI22_X1 port map( A1 => n5334, A2 => n3983, B1 => n5335, B2 => 
                           n4367, ZN => n5678);
   U4770 : OAI221_X1 port map( B1 => n3859, B2 => n5336, C1 => n4243, C2 => 
                           n5337, A => n5679, ZN => n5672);
   U4771 : AOI22_X1 port map( A1 => n5339, A2 => n3699, B1 => n5340, B2 => 
                           n4083, ZN => n5679);
   U4772 : NOR4_X1 port map( A1 => n5680, A2 => n5681, A3 => n5682, A4 => n5683
                           , ZN => n5670);
   U4773 : OAI221_X1 port map( B1 => n3860, B2 => n5345, C1 => n4244, C2 => 
                           n5346, A => n5684, ZN => n5683);
   U4774 : AOI22_X1 port map( A1 => n5348, A2 => n3700, B1 => n5349, B2 => 
                           n4084, ZN => n5684);
   U4775 : OAI221_X1 port map( B1 => n3861, B2 => n5350, C1 => n4245, C2 => 
                           n5351, A => n5685, ZN => n5682);
   U4776 : AOI22_X1 port map( A1 => n5353, A2 => n3701, B1 => n5354, B2 => 
                           n4085, ZN => n5685);
   U4777 : OAI221_X1 port map( B1 => n3862, B2 => n5355, C1 => n4246, C2 => 
                           n5356, A => n5686, ZN => n5681);
   U4778 : AOI22_X1 port map( A1 => n5358, A2 => n3702, B1 => n5359, B2 => 
                           n4086, ZN => n5686);
   U4779 : OAI221_X1 port map( B1 => n3863, B2 => n5360, C1 => n4247, C2 => 
                           n5361, A => n5687, ZN => n5680);
   U4780 : AOI22_X1 port map( A1 => n5363, A2 => n3703, B1 => n5364, B2 => 
                           n4087, ZN => n5687);
   U4781 : MUX2_X1 port map( A => OUT1_13_port, B => n5688, S => n5314, Z => 
                           n2539);
   U4782 : NAND2_X1 port map( A1 => n5689, A2 => n5690, ZN => n5688);
   U4783 : NOR4_X1 port map( A1 => n5691, A2 => n5692, A3 => n5693, A4 => n5694
                           , ZN => n5690);
   U4784 : OAI221_X1 port map( B1 => n19, B2 => n5321, C1 => n51, C2 => n5322, 
                           A => n5695, ZN => n5694);
   U4785 : AOI22_X1 port map( A1 => n5324, A2 => n6025, B1 => n5325, B2 => 
                           n6026, ZN => n5695);
   U4786 : OAI221_X1 port map( B1 => n147, B2 => n5326, C1 => n179, C2 => n5327
                           , A => n5696, ZN => n5693);
   U4787 : AOI22_X1 port map( A1 => n5329, A2 => n6023, B1 => n5330, B2 => 
                           n6024, ZN => n5696);
   U4788 : OAI221_X1 port map( B1 => n307, B2 => n5331, C1 => n275, C2 => n5332
                           , A => n5697, ZN => n5692);
   U4789 : AOI22_X1 port map( A1 => n5334, A2 => n3984, B1 => n5335, B2 => 
                           n4368, ZN => n5697);
   U4790 : OAI221_X1 port map( B1 => n3864, B2 => n5336, C1 => n4248, C2 => 
                           n5337, A => n5698, ZN => n5691);
   U4791 : AOI22_X1 port map( A1 => n5339, A2 => n3704, B1 => n5340, B2 => 
                           n4088, ZN => n5698);
   U4792 : NOR4_X1 port map( A1 => n5699, A2 => n5700, A3 => n5701, A4 => n5702
                           , ZN => n5689);
   U4793 : OAI221_X1 port map( B1 => n3865, B2 => n5345, C1 => n4249, C2 => 
                           n5346, A => n5703, ZN => n5702);
   U4794 : AOI22_X1 port map( A1 => n5348, A2 => n3705, B1 => n5349, B2 => 
                           n4089, ZN => n5703);
   U4795 : OAI221_X1 port map( B1 => n3866, B2 => n5350, C1 => n4250, C2 => 
                           n5351, A => n5704, ZN => n5701);
   U4796 : AOI22_X1 port map( A1 => n5353, A2 => n3706, B1 => n5354, B2 => 
                           n4090, ZN => n5704);
   U4797 : OAI221_X1 port map( B1 => n3867, B2 => n5355, C1 => n4251, C2 => 
                           n5356, A => n5705, ZN => n5700);
   U4798 : AOI22_X1 port map( A1 => n5358, A2 => n3707, B1 => n5359, B2 => 
                           n4091, ZN => n5705);
   U4799 : OAI221_X1 port map( B1 => n3868, B2 => n5360, C1 => n4252, C2 => 
                           n5361, A => n5706, ZN => n5699);
   U4800 : AOI22_X1 port map( A1 => n5363, A2 => n3708, B1 => n5364, B2 => 
                           n4092, ZN => n5706);
   U4801 : MUX2_X1 port map( A => OUT1_12_port, B => n5707, S => n5314, Z => 
                           n2538);
   U4802 : NAND2_X1 port map( A1 => n5708, A2 => n5709, ZN => n5707);
   U4803 : NOR4_X1 port map( A1 => n5710, A2 => n5711, A3 => n5712, A4 => n5713
                           , ZN => n5709);
   U4804 : OAI221_X1 port map( B1 => n20, B2 => n5321, C1 => n52, C2 => n5322, 
                           A => n5714, ZN => n5713);
   U4805 : AOI22_X1 port map( A1 => n5324, A2 => n6021, B1 => n5325, B2 => 
                           n6022, ZN => n5714);
   U4806 : OAI221_X1 port map( B1 => n148, B2 => n5326, C1 => n180, C2 => n5327
                           , A => n5715, ZN => n5712);
   U4807 : AOI22_X1 port map( A1 => n5329, A2 => n6019, B1 => n5330, B2 => 
                           n6020, ZN => n5715);
   U4808 : OAI221_X1 port map( B1 => n308, B2 => n5331, C1 => n276, C2 => n5332
                           , A => n5716, ZN => n5711);
   U4809 : AOI22_X1 port map( A1 => n5334, A2 => n3985, B1 => n5335, B2 => 
                           n4369, ZN => n5716);
   U4810 : OAI221_X1 port map( B1 => n3869, B2 => n5336, C1 => n4253, C2 => 
                           n5337, A => n5717, ZN => n5710);
   U4811 : AOI22_X1 port map( A1 => n5339, A2 => n3709, B1 => n5340, B2 => 
                           n4093, ZN => n5717);
   U4812 : NOR4_X1 port map( A1 => n5718, A2 => n5719, A3 => n5720, A4 => n5721
                           , ZN => n5708);
   U4813 : OAI221_X1 port map( B1 => n3870, B2 => n5345, C1 => n4254, C2 => 
                           n5346, A => n5722, ZN => n5721);
   U4814 : AOI22_X1 port map( A1 => n5348, A2 => n3710, B1 => n5349, B2 => 
                           n4094, ZN => n5722);
   U4815 : OAI221_X1 port map( B1 => n3871, B2 => n5350, C1 => n4255, C2 => 
                           n5351, A => n5723, ZN => n5720);
   U4816 : AOI22_X1 port map( A1 => n5353, A2 => n3711, B1 => n5354, B2 => 
                           n4095, ZN => n5723);
   U4817 : OAI221_X1 port map( B1 => n3872, B2 => n5355, C1 => n4256, C2 => 
                           n5356, A => n5724, ZN => n5719);
   U4818 : AOI22_X1 port map( A1 => n5358, A2 => n3712, B1 => n5359, B2 => 
                           n4096, ZN => n5724);
   U4819 : OAI221_X1 port map( B1 => n3873, B2 => n5360, C1 => n4257, C2 => 
                           n5361, A => n5725, ZN => n5718);
   U4820 : AOI22_X1 port map( A1 => n5363, A2 => n3713, B1 => n5364, B2 => 
                           n4097, ZN => n5725);
   U4821 : MUX2_X1 port map( A => OUT1_11_port, B => n5726, S => n5314, Z => 
                           n2537);
   U4822 : NAND2_X1 port map( A1 => n5727, A2 => n5728, ZN => n5726);
   U4823 : NOR4_X1 port map( A1 => n5729, A2 => n5730, A3 => n5731, A4 => n5732
                           , ZN => n5728);
   U4824 : OAI221_X1 port map( B1 => n21, B2 => n5321, C1 => n53, C2 => n5322, 
                           A => n5733, ZN => n5732);
   U4825 : AOI22_X1 port map( A1 => n5324, A2 => n6017, B1 => n5325, B2 => 
                           n6018, ZN => n5733);
   U4826 : OAI221_X1 port map( B1 => n149, B2 => n5326, C1 => n181, C2 => n5327
                           , A => n5734, ZN => n5731);
   U4827 : AOI22_X1 port map( A1 => n5329, A2 => n6015, B1 => n5330, B2 => 
                           n6016, ZN => n5734);
   U4828 : OAI221_X1 port map( B1 => n309, B2 => n5331, C1 => n277, C2 => n5332
                           , A => n5735, ZN => n5730);
   U4829 : AOI22_X1 port map( A1 => n5334, A2 => n3986, B1 => n5335, B2 => 
                           n4370, ZN => n5735);
   U4830 : OAI221_X1 port map( B1 => n3874, B2 => n5336, C1 => n4258, C2 => 
                           n5337, A => n5736, ZN => n5729);
   U4831 : AOI22_X1 port map( A1 => n5339, A2 => n3714, B1 => n5340, B2 => 
                           n4098, ZN => n5736);
   U4832 : NOR4_X1 port map( A1 => n5737, A2 => n5738, A3 => n5739, A4 => n5740
                           , ZN => n5727);
   U4833 : OAI221_X1 port map( B1 => n3875, B2 => n5345, C1 => n4259, C2 => 
                           n5346, A => n5741, ZN => n5740);
   U4834 : AOI22_X1 port map( A1 => n5348, A2 => n3715, B1 => n5349, B2 => 
                           n4099, ZN => n5741);
   U4835 : OAI221_X1 port map( B1 => n3876, B2 => n5350, C1 => n4260, C2 => 
                           n5351, A => n5742, ZN => n5739);
   U4836 : AOI22_X1 port map( A1 => n5353, A2 => n3716, B1 => n5354, B2 => 
                           n4100, ZN => n5742);
   U4837 : OAI221_X1 port map( B1 => n3877, B2 => n5355, C1 => n4261, C2 => 
                           n5356, A => n5743, ZN => n5738);
   U4838 : AOI22_X1 port map( A1 => n5358, A2 => n3717, B1 => n5359, B2 => 
                           n4101, ZN => n5743);
   U4839 : OAI221_X1 port map( B1 => n3878, B2 => n5360, C1 => n4262, C2 => 
                           n5361, A => n5744, ZN => n5737);
   U4840 : AOI22_X1 port map( A1 => n5363, A2 => n3718, B1 => n5364, B2 => 
                           n4102, ZN => n5744);
   U4841 : MUX2_X1 port map( A => OUT1_10_port, B => n5745, S => n5314, Z => 
                           n2536);
   U4842 : NAND2_X1 port map( A1 => n5746, A2 => n5747, ZN => n5745);
   U4843 : NOR4_X1 port map( A1 => n5748, A2 => n5749, A3 => n5750, A4 => n5751
                           , ZN => n5747);
   U4844 : OAI221_X1 port map( B1 => n22, B2 => n5321, C1 => n54, C2 => n5322, 
                           A => n5752, ZN => n5751);
   U4845 : AOI22_X1 port map( A1 => n5324, A2 => n6013, B1 => n5325, B2 => 
                           n6014, ZN => n5752);
   U4846 : OAI221_X1 port map( B1 => n150, B2 => n5326, C1 => n182, C2 => n5327
                           , A => n5753, ZN => n5750);
   U4847 : AOI22_X1 port map( A1 => n5329, A2 => n6011, B1 => n5330, B2 => 
                           n6012, ZN => n5753);
   U4848 : OAI221_X1 port map( B1 => n310, B2 => n5331, C1 => n278, C2 => n5332
                           , A => n5754, ZN => n5749);
   U4849 : AOI22_X1 port map( A1 => n5334, A2 => n3987, B1 => n5335, B2 => 
                           n4371, ZN => n5754);
   U4850 : OAI221_X1 port map( B1 => n3879, B2 => n5336, C1 => n4263, C2 => 
                           n5337, A => n5755, ZN => n5748);
   U4851 : AOI22_X1 port map( A1 => n5339, A2 => n3719, B1 => n5340, B2 => 
                           n4103, ZN => n5755);
   U4852 : NOR4_X1 port map( A1 => n5756, A2 => n5757, A3 => n5758, A4 => n5759
                           , ZN => n5746);
   U4853 : OAI221_X1 port map( B1 => n3880, B2 => n5345, C1 => n4264, C2 => 
                           n5346, A => n5760, ZN => n5759);
   U4854 : AOI22_X1 port map( A1 => n5348, A2 => n3720, B1 => n5349, B2 => 
                           n4104, ZN => n5760);
   U4855 : OAI221_X1 port map( B1 => n3881, B2 => n5350, C1 => n4265, C2 => 
                           n5351, A => n5761, ZN => n5758);
   U4856 : AOI22_X1 port map( A1 => n5353, A2 => n3721, B1 => n5354, B2 => 
                           n4105, ZN => n5761);
   U4857 : OAI221_X1 port map( B1 => n3882, B2 => n5355, C1 => n4266, C2 => 
                           n5356, A => n5762, ZN => n5757);
   U4858 : AOI22_X1 port map( A1 => n5358, A2 => n3722, B1 => n5359, B2 => 
                           n4106, ZN => n5762);
   U4859 : OAI221_X1 port map( B1 => n3883, B2 => n5360, C1 => n4267, C2 => 
                           n5361, A => n5763, ZN => n5756);
   U4860 : AOI22_X1 port map( A1 => n5363, A2 => n3723, B1 => n5364, B2 => 
                           n4107, ZN => n5763);
   U4861 : MUX2_X1 port map( A => OUT1_9_port, B => n5764, S => n5314, Z => 
                           n2535);
   U4862 : NAND2_X1 port map( A1 => n5765, A2 => n5766, ZN => n5764);
   U4863 : NOR4_X1 port map( A1 => n5767, A2 => n5768, A3 => n5769, A4 => n5770
                           , ZN => n5766);
   U4864 : OAI221_X1 port map( B1 => n23, B2 => n5321, C1 => n55, C2 => n5322, 
                           A => n5771, ZN => n5770);
   U4865 : AOI22_X1 port map( A1 => n5324, A2 => n6009, B1 => n5325, B2 => 
                           n6010, ZN => n5771);
   U4866 : OAI221_X1 port map( B1 => n151, B2 => n5326, C1 => n183, C2 => n5327
                           , A => n5772, ZN => n5769);
   U4867 : AOI22_X1 port map( A1 => n5329, A2 => n6007, B1 => n5330, B2 => 
                           n6008, ZN => n5772);
   U4868 : OAI221_X1 port map( B1 => n311, B2 => n5331, C1 => n279, C2 => n5332
                           , A => n5773, ZN => n5768);
   U4869 : AOI22_X1 port map( A1 => n5334, A2 => n3988, B1 => n5335, B2 => 
                           n4372, ZN => n5773);
   U4870 : OAI221_X1 port map( B1 => n3884, B2 => n5336, C1 => n4268, C2 => 
                           n5337, A => n5774, ZN => n5767);
   U4871 : AOI22_X1 port map( A1 => n5339, A2 => n3724, B1 => n5340, B2 => 
                           n4108, ZN => n5774);
   U4872 : NOR4_X1 port map( A1 => n5775, A2 => n5776, A3 => n5777, A4 => n5778
                           , ZN => n5765);
   U4873 : OAI221_X1 port map( B1 => n3885, B2 => n5345, C1 => n4269, C2 => 
                           n5346, A => n5779, ZN => n5778);
   U4874 : AOI22_X1 port map( A1 => n5348, A2 => n3725, B1 => n5349, B2 => 
                           n4109, ZN => n5779);
   U4875 : OAI221_X1 port map( B1 => n3886, B2 => n5350, C1 => n4270, C2 => 
                           n5351, A => n5780, ZN => n5777);
   U4876 : AOI22_X1 port map( A1 => n5353, A2 => n3726, B1 => n5354, B2 => 
                           n4110, ZN => n5780);
   U4877 : OAI221_X1 port map( B1 => n3887, B2 => n5355, C1 => n4271, C2 => 
                           n5356, A => n5781, ZN => n5776);
   U4878 : AOI22_X1 port map( A1 => n5358, A2 => n3727, B1 => n5359, B2 => 
                           n4111, ZN => n5781);
   U4879 : OAI221_X1 port map( B1 => n3888, B2 => n5360, C1 => n4272, C2 => 
                           n5361, A => n5782, ZN => n5775);
   U4880 : AOI22_X1 port map( A1 => n5363, A2 => n3728, B1 => n5364, B2 => 
                           n4112, ZN => n5782);
   U4881 : MUX2_X1 port map( A => OUT1_8_port, B => n5783, S => n5314, Z => 
                           n2534);
   U4882 : NAND2_X1 port map( A1 => n5784, A2 => n5785, ZN => n5783);
   U4883 : NOR4_X1 port map( A1 => n5786, A2 => n5787, A3 => n5788, A4 => n5789
                           , ZN => n5785);
   U4884 : OAI221_X1 port map( B1 => n24, B2 => n5321, C1 => n56, C2 => n5322, 
                           A => n5790, ZN => n5789);
   U4885 : AOI22_X1 port map( A1 => n5324, A2 => n6005, B1 => n5325, B2 => 
                           n6006, ZN => n5790);
   U4886 : OAI221_X1 port map( B1 => n152, B2 => n5326, C1 => n184, C2 => n5327
                           , A => n5791, ZN => n5788);
   U4887 : AOI22_X1 port map( A1 => n5329, A2 => n6003, B1 => n5330, B2 => 
                           n6004, ZN => n5791);
   U4888 : OAI221_X1 port map( B1 => n312, B2 => n5331, C1 => n280, C2 => n5332
                           , A => n5792, ZN => n5787);
   U4889 : AOI22_X1 port map( A1 => n5334, A2 => n3989, B1 => n5335, B2 => 
                           n4373, ZN => n5792);
   U4890 : OAI221_X1 port map( B1 => n3889, B2 => n5336, C1 => n4273, C2 => 
                           n5337, A => n5793, ZN => n5786);
   U4891 : AOI22_X1 port map( A1 => n5339, A2 => n3729, B1 => n5340, B2 => 
                           n4113, ZN => n5793);
   U4892 : NOR4_X1 port map( A1 => n5794, A2 => n5795, A3 => n5796, A4 => n5797
                           , ZN => n5784);
   U4893 : OAI221_X1 port map( B1 => n3890, B2 => n5345, C1 => n4274, C2 => 
                           n5346, A => n5798, ZN => n5797);
   U4894 : AOI22_X1 port map( A1 => n5348, A2 => n3730, B1 => n5349, B2 => 
                           n4114, ZN => n5798);
   U4895 : OAI221_X1 port map( B1 => n3891, B2 => n5350, C1 => n4275, C2 => 
                           n5351, A => n5799, ZN => n5796);
   U4896 : AOI22_X1 port map( A1 => n5353, A2 => n3731, B1 => n5354, B2 => 
                           n4115, ZN => n5799);
   U4897 : OAI221_X1 port map( B1 => n3892, B2 => n5355, C1 => n4276, C2 => 
                           n5356, A => n5800, ZN => n5795);
   U4898 : AOI22_X1 port map( A1 => n5358, A2 => n3732, B1 => n5359, B2 => 
                           n4116, ZN => n5800);
   U4899 : OAI221_X1 port map( B1 => n3893, B2 => n5360, C1 => n4277, C2 => 
                           n5361, A => n5801, ZN => n5794);
   U4900 : AOI22_X1 port map( A1 => n5363, A2 => n3733, B1 => n5364, B2 => 
                           n4117, ZN => n5801);
   U4901 : MUX2_X1 port map( A => OUT1_7_port, B => n5802, S => n5314, Z => 
                           n2533);
   U4902 : NAND2_X1 port map( A1 => n5803, A2 => n5804, ZN => n5802);
   U4903 : NOR4_X1 port map( A1 => n5805, A2 => n5806, A3 => n5807, A4 => n5808
                           , ZN => n5804);
   U4904 : OAI221_X1 port map( B1 => n25, B2 => n5321, C1 => n57, C2 => n5322, 
                           A => n5809, ZN => n5808);
   U4905 : AOI22_X1 port map( A1 => n5324, A2 => n6001, B1 => n5325, B2 => 
                           n6002, ZN => n5809);
   U4906 : OAI221_X1 port map( B1 => n153, B2 => n5326, C1 => n185, C2 => n5327
                           , A => n5810, ZN => n5807);
   U4907 : AOI22_X1 port map( A1 => n5329, A2 => n5999, B1 => n5330, B2 => 
                           n6000, ZN => n5810);
   U4908 : OAI221_X1 port map( B1 => n313, B2 => n5331, C1 => n281, C2 => n5332
                           , A => n5811, ZN => n5806);
   U4909 : AOI22_X1 port map( A1 => n5334, A2 => n3990, B1 => n5335, B2 => 
                           n4374, ZN => n5811);
   U4910 : OAI221_X1 port map( B1 => n3894, B2 => n5336, C1 => n4278, C2 => 
                           n5337, A => n5812, ZN => n5805);
   U4911 : AOI22_X1 port map( A1 => n5339, A2 => n3734, B1 => n5340, B2 => 
                           n4118, ZN => n5812);
   U4912 : NOR4_X1 port map( A1 => n5813, A2 => n5814, A3 => n5815, A4 => n5816
                           , ZN => n5803);
   U4913 : OAI221_X1 port map( B1 => n3895, B2 => n5345, C1 => n4279, C2 => 
                           n5346, A => n5817, ZN => n5816);
   U4914 : AOI22_X1 port map( A1 => n5348, A2 => n3735, B1 => n5349, B2 => 
                           n4119, ZN => n5817);
   U4915 : OAI221_X1 port map( B1 => n3896, B2 => n5350, C1 => n4280, C2 => 
                           n5351, A => n5818, ZN => n5815);
   U4916 : AOI22_X1 port map( A1 => n5353, A2 => n3736, B1 => n5354, B2 => 
                           n4120, ZN => n5818);
   U4917 : OAI221_X1 port map( B1 => n3897, B2 => n5355, C1 => n4281, C2 => 
                           n5356, A => n5819, ZN => n5814);
   U4918 : AOI22_X1 port map( A1 => n5358, A2 => n3737, B1 => n5359, B2 => 
                           n4121, ZN => n5819);
   U4919 : OAI221_X1 port map( B1 => n3898, B2 => n5360, C1 => n4282, C2 => 
                           n5361, A => n5820, ZN => n5813);
   U4920 : AOI22_X1 port map( A1 => n5363, A2 => n3738, B1 => n5364, B2 => 
                           n4122, ZN => n5820);
   U4921 : MUX2_X1 port map( A => OUT1_6_port, B => n5821, S => n5314, Z => 
                           n2532);
   U4922 : NAND2_X1 port map( A1 => n5822, A2 => n5823, ZN => n5821);
   U4923 : NOR4_X1 port map( A1 => n5824, A2 => n5825, A3 => n5826, A4 => n5827
                           , ZN => n5823);
   U4924 : OAI221_X1 port map( B1 => n26, B2 => n5321, C1 => n58, C2 => n5322, 
                           A => n5828, ZN => n5827);
   U4925 : AOI22_X1 port map( A1 => n5324, A2 => n5997, B1 => n5325, B2 => 
                           n5998, ZN => n5828);
   U4926 : OAI221_X1 port map( B1 => n154, B2 => n5326, C1 => n186, C2 => n5327
                           , A => n5829, ZN => n5826);
   U4927 : AOI22_X1 port map( A1 => n5329, A2 => n5995, B1 => n5330, B2 => 
                           n5996, ZN => n5829);
   U4928 : OAI221_X1 port map( B1 => n314, B2 => n5331, C1 => n282, C2 => n5332
                           , A => n5830, ZN => n5825);
   U4929 : AOI22_X1 port map( A1 => n5334, A2 => n3991, B1 => n5335, B2 => 
                           n4375, ZN => n5830);
   U4930 : OAI221_X1 port map( B1 => n3899, B2 => n5336, C1 => n4283, C2 => 
                           n5337, A => n5831, ZN => n5824);
   U4931 : AOI22_X1 port map( A1 => n5339, A2 => n3739, B1 => n5340, B2 => 
                           n4123, ZN => n5831);
   U4932 : NOR4_X1 port map( A1 => n5832, A2 => n5833, A3 => n5834, A4 => n5835
                           , ZN => n5822);
   U4933 : OAI221_X1 port map( B1 => n3900, B2 => n5345, C1 => n4284, C2 => 
                           n5346, A => n5836, ZN => n5835);
   U4934 : AOI22_X1 port map( A1 => n5348, A2 => n3740, B1 => n5349, B2 => 
                           n4124, ZN => n5836);
   U4935 : OAI221_X1 port map( B1 => n3901, B2 => n5350, C1 => n4285, C2 => 
                           n5351, A => n5837, ZN => n5834);
   U4936 : AOI22_X1 port map( A1 => n5353, A2 => n3741, B1 => n5354, B2 => 
                           n4125, ZN => n5837);
   U4937 : OAI221_X1 port map( B1 => n3902, B2 => n5355, C1 => n4286, C2 => 
                           n5356, A => n5838, ZN => n5833);
   U4938 : AOI22_X1 port map( A1 => n5358, A2 => n3742, B1 => n5359, B2 => 
                           n4126, ZN => n5838);
   U4939 : OAI221_X1 port map( B1 => n3903, B2 => n5360, C1 => n4287, C2 => 
                           n5361, A => n5839, ZN => n5832);
   U4940 : AOI22_X1 port map( A1 => n5363, A2 => n3743, B1 => n5364, B2 => 
                           n4127, ZN => n5839);
   U4941 : MUX2_X1 port map( A => OUT1_5_port, B => n5840, S => n5314, Z => 
                           n2531);
   U4942 : NAND2_X1 port map( A1 => n5841, A2 => n5842, ZN => n5840);
   U4943 : NOR4_X1 port map( A1 => n5843, A2 => n5844, A3 => n5845, A4 => n5846
                           , ZN => n5842);
   U4944 : OAI221_X1 port map( B1 => n27, B2 => n5321, C1 => n59, C2 => n5322, 
                           A => n5847, ZN => n5846);
   U4945 : AOI22_X1 port map( A1 => n5324, A2 => n5993, B1 => n5325, B2 => 
                           n5994, ZN => n5847);
   U4946 : OAI221_X1 port map( B1 => n155, B2 => n5326, C1 => n187, C2 => n5327
                           , A => n5848, ZN => n5845);
   U4947 : AOI22_X1 port map( A1 => n5329, A2 => n5991, B1 => n5330, B2 => 
                           n5992, ZN => n5848);
   U4948 : OAI221_X1 port map( B1 => n315, B2 => n5331, C1 => n283, C2 => n5332
                           , A => n5849, ZN => n5844);
   U4949 : AOI22_X1 port map( A1 => n5334, A2 => n3992, B1 => n5335, B2 => 
                           n4376, ZN => n5849);
   U4950 : OAI221_X1 port map( B1 => n3904, B2 => n5336, C1 => n4288, C2 => 
                           n5337, A => n5850, ZN => n5843);
   U4951 : AOI22_X1 port map( A1 => n5339, A2 => n3744, B1 => n5340, B2 => 
                           n4128, ZN => n5850);
   U4952 : NOR4_X1 port map( A1 => n5851, A2 => n5852, A3 => n5853, A4 => n5854
                           , ZN => n5841);
   U4953 : OAI221_X1 port map( B1 => n3905, B2 => n5345, C1 => n4289, C2 => 
                           n5346, A => n5855, ZN => n5854);
   U4954 : AOI22_X1 port map( A1 => n5348, A2 => n3745, B1 => n5349, B2 => 
                           n4129, ZN => n5855);
   U4955 : OAI221_X1 port map( B1 => n3906, B2 => n5350, C1 => n4290, C2 => 
                           n5351, A => n5856, ZN => n5853);
   U4956 : AOI22_X1 port map( A1 => n5353, A2 => n3746, B1 => n5354, B2 => 
                           n4130, ZN => n5856);
   U4957 : OAI221_X1 port map( B1 => n3907, B2 => n5355, C1 => n4291, C2 => 
                           n5356, A => n5857, ZN => n5852);
   U4958 : AOI22_X1 port map( A1 => n5358, A2 => n3747, B1 => n5359, B2 => 
                           n4131, ZN => n5857);
   U4959 : OAI221_X1 port map( B1 => n3908, B2 => n5360, C1 => n4292, C2 => 
                           n5361, A => n5858, ZN => n5851);
   U4960 : AOI22_X1 port map( A1 => n5363, A2 => n3748, B1 => n5364, B2 => 
                           n4132, ZN => n5858);
   U4961 : MUX2_X1 port map( A => OUT1_4_port, B => n5859, S => n5314, Z => 
                           n2530);
   U4962 : NAND2_X1 port map( A1 => n5860, A2 => n5861, ZN => n5859);
   U4963 : NOR4_X1 port map( A1 => n5862, A2 => n5863, A3 => n5864, A4 => n5865
                           , ZN => n5861);
   U4964 : OAI221_X1 port map( B1 => n28, B2 => n5321, C1 => n60, C2 => n5322, 
                           A => n5866, ZN => n5865);
   U4965 : AOI22_X1 port map( A1 => n5324, A2 => n5989, B1 => n5325, B2 => 
                           n5990, ZN => n5866);
   U4966 : OAI221_X1 port map( B1 => n156, B2 => n5326, C1 => n188, C2 => n5327
                           , A => n5867, ZN => n5864);
   U4967 : AOI22_X1 port map( A1 => n5329, A2 => n5987, B1 => n5330, B2 => 
                           n5988, ZN => n5867);
   U4968 : OAI221_X1 port map( B1 => n316, B2 => n5331, C1 => n284, C2 => n5332
                           , A => n5868, ZN => n5863);
   U4969 : AOI22_X1 port map( A1 => n5334, A2 => n3993, B1 => n5335, B2 => 
                           n4377, ZN => n5868);
   U4970 : OAI221_X1 port map( B1 => n3909, B2 => n5336, C1 => n4293, C2 => 
                           n5337, A => n5869, ZN => n5862);
   U4971 : AOI22_X1 port map( A1 => n5339, A2 => n3749, B1 => n5340, B2 => 
                           n4133, ZN => n5869);
   U4972 : NOR4_X1 port map( A1 => n5870, A2 => n5871, A3 => n5872, A4 => n5873
                           , ZN => n5860);
   U4973 : OAI221_X1 port map( B1 => n3910, B2 => n5345, C1 => n4294, C2 => 
                           n5346, A => n5874, ZN => n5873);
   U4974 : AOI22_X1 port map( A1 => n5348, A2 => n3750, B1 => n5349, B2 => 
                           n4134, ZN => n5874);
   U4975 : OAI221_X1 port map( B1 => n3911, B2 => n5350, C1 => n4295, C2 => 
                           n5351, A => n5875, ZN => n5872);
   U4976 : AOI22_X1 port map( A1 => n5353, A2 => n3751, B1 => n5354, B2 => 
                           n4135, ZN => n5875);
   U4977 : OAI221_X1 port map( B1 => n3912, B2 => n5355, C1 => n4296, C2 => 
                           n5356, A => n5876, ZN => n5871);
   U4978 : AOI22_X1 port map( A1 => n5358, A2 => n3752, B1 => n5359, B2 => 
                           n4136, ZN => n5876);
   U4979 : OAI221_X1 port map( B1 => n3913, B2 => n5360, C1 => n4297, C2 => 
                           n5361, A => n5877, ZN => n5870);
   U4980 : AOI22_X1 port map( A1 => n5363, A2 => n3753, B1 => n5364, B2 => 
                           n4137, ZN => n5877);
   U4981 : MUX2_X1 port map( A => OUT1_3_port, B => n5878, S => n5314, Z => 
                           n2529);
   U4982 : NAND2_X1 port map( A1 => n5879, A2 => n5880, ZN => n5878);
   U4983 : NOR4_X1 port map( A1 => n5881, A2 => n5882, A3 => n5883, A4 => n5884
                           , ZN => n5880);
   U4984 : OAI221_X1 port map( B1 => n29, B2 => n5321, C1 => n61, C2 => n5322, 
                           A => n5885, ZN => n5884);
   U4985 : AOI22_X1 port map( A1 => n5324, A2 => n5985, B1 => n5325, B2 => 
                           n5986, ZN => n5885);
   U4986 : OAI221_X1 port map( B1 => n157, B2 => n5326, C1 => n189, C2 => n5327
                           , A => n5886, ZN => n5883);
   U4987 : AOI22_X1 port map( A1 => n5329, A2 => n5983, B1 => n5330, B2 => 
                           n5984, ZN => n5886);
   U4988 : OAI221_X1 port map( B1 => n317, B2 => n5331, C1 => n285, C2 => n5332
                           , A => n5887, ZN => n5882);
   U4989 : AOI22_X1 port map( A1 => n5334, A2 => n3994, B1 => n5335, B2 => 
                           n4378, ZN => n5887);
   U4990 : OAI221_X1 port map( B1 => n3914, B2 => n5336, C1 => n4298, C2 => 
                           n5337, A => n5888, ZN => n5881);
   U4991 : AOI22_X1 port map( A1 => n5339, A2 => n3754, B1 => n5340, B2 => 
                           n4138, ZN => n5888);
   U4992 : NOR4_X1 port map( A1 => n5889, A2 => n5890, A3 => n5891, A4 => n5892
                           , ZN => n5879);
   U4993 : OAI221_X1 port map( B1 => n3915, B2 => n5345, C1 => n4299, C2 => 
                           n5346, A => n5893, ZN => n5892);
   U4994 : AOI22_X1 port map( A1 => n5348, A2 => n3755, B1 => n5349, B2 => 
                           n4139, ZN => n5893);
   U4995 : OAI221_X1 port map( B1 => n3916, B2 => n5350, C1 => n4300, C2 => 
                           n5351, A => n5894, ZN => n5891);
   U4996 : AOI22_X1 port map( A1 => n5353, A2 => n3756, B1 => n5354, B2 => 
                           n4140, ZN => n5894);
   U4997 : OAI221_X1 port map( B1 => n3917, B2 => n5355, C1 => n4301, C2 => 
                           n5356, A => n5895, ZN => n5890);
   U4998 : AOI22_X1 port map( A1 => n5358, A2 => n3757, B1 => n5359, B2 => 
                           n4141, ZN => n5895);
   U4999 : OAI221_X1 port map( B1 => n3918, B2 => n5360, C1 => n4302, C2 => 
                           n5361, A => n5896, ZN => n5889);
   U5000 : AOI22_X1 port map( A1 => n5363, A2 => n3758, B1 => n5364, B2 => 
                           n4142, ZN => n5896);
   U5001 : MUX2_X1 port map( A => OUT1_2_port, B => n5897, S => n5314, Z => 
                           n2528);
   U5002 : NAND2_X1 port map( A1 => n5898, A2 => n5899, ZN => n5897);
   U5003 : NOR4_X1 port map( A1 => n5900, A2 => n5901, A3 => n5902, A4 => n5903
                           , ZN => n5899);
   U5004 : OAI221_X1 port map( B1 => n30, B2 => n5321, C1 => n62, C2 => n5322, 
                           A => n5904, ZN => n5903);
   U5005 : AOI22_X1 port map( A1 => n5324, A2 => n5981, B1 => n5325, B2 => 
                           n5982, ZN => n5904);
   U5006 : OAI221_X1 port map( B1 => n158, B2 => n5326, C1 => n190, C2 => n5327
                           , A => n5905, ZN => n5902);
   U5007 : AOI22_X1 port map( A1 => n5329, A2 => n5979, B1 => n5330, B2 => 
                           n5980, ZN => n5905);
   U5008 : OAI221_X1 port map( B1 => n318, B2 => n5331, C1 => n286, C2 => n5332
                           , A => n5906, ZN => n5901);
   U5009 : AOI22_X1 port map( A1 => n5334, A2 => n3995, B1 => n5335, B2 => 
                           n4379, ZN => n5906);
   U5010 : OAI221_X1 port map( B1 => n3919, B2 => n5336, C1 => n4303, C2 => 
                           n5337, A => n5907, ZN => n5900);
   U5011 : AOI22_X1 port map( A1 => n5339, A2 => n3759, B1 => n5340, B2 => 
                           n4143, ZN => n5907);
   U5012 : NOR4_X1 port map( A1 => n5908, A2 => n5909, A3 => n5910, A4 => n5911
                           , ZN => n5898);
   U5013 : OAI221_X1 port map( B1 => n3920, B2 => n5345, C1 => n4304, C2 => 
                           n5346, A => n5912, ZN => n5911);
   U5014 : AOI22_X1 port map( A1 => n5348, A2 => n3760, B1 => n5349, B2 => 
                           n4144, ZN => n5912);
   U5015 : OAI221_X1 port map( B1 => n3921, B2 => n5350, C1 => n4305, C2 => 
                           n5351, A => n5913, ZN => n5910);
   U5016 : AOI22_X1 port map( A1 => n5353, A2 => n3761, B1 => n5354, B2 => 
                           n4145, ZN => n5913);
   U5017 : OAI221_X1 port map( B1 => n3922, B2 => n5355, C1 => n4306, C2 => 
                           n5356, A => n5914, ZN => n5909);
   U5018 : AOI22_X1 port map( A1 => n5358, A2 => n3762, B1 => n5359, B2 => 
                           n4146, ZN => n5914);
   U5019 : OAI221_X1 port map( B1 => n3923, B2 => n5360, C1 => n4307, C2 => 
                           n5361, A => n5915, ZN => n5908);
   U5020 : AOI22_X1 port map( A1 => n5363, A2 => n3763, B1 => n5364, B2 => 
                           n4147, ZN => n5915);
   U5021 : MUX2_X1 port map( A => OUT1_1_port, B => n5916, S => n5314, Z => 
                           n2527);
   U5022 : NAND2_X1 port map( A1 => n5917, A2 => n5918, ZN => n5916);
   U5023 : NOR4_X1 port map( A1 => n5919, A2 => n5920, A3 => n5921, A4 => n5922
                           , ZN => n5918);
   U5024 : OAI221_X1 port map( B1 => n31, B2 => n5321, C1 => n63, C2 => n5322, 
                           A => n5923, ZN => n5922);
   U5025 : AOI22_X1 port map( A1 => n5324, A2 => n5977, B1 => n5325, B2 => 
                           n5978, ZN => n5923);
   U5026 : OAI221_X1 port map( B1 => n159, B2 => n5326, C1 => n191, C2 => n5327
                           , A => n5924, ZN => n5921);
   U5027 : AOI22_X1 port map( A1 => n5329, A2 => n5975, B1 => n5330, B2 => 
                           n5976, ZN => n5924);
   U5028 : OAI221_X1 port map( B1 => n319, B2 => n5331, C1 => n287, C2 => n5332
                           , A => n5925, ZN => n5920);
   U5029 : AOI22_X1 port map( A1 => n5334, A2 => n3996, B1 => n5335, B2 => 
                           n4380, ZN => n5925);
   U5030 : OAI221_X1 port map( B1 => n3924, B2 => n5336, C1 => n4308, C2 => 
                           n5337, A => n5926, ZN => n5919);
   U5031 : AOI22_X1 port map( A1 => n5339, A2 => n3764, B1 => n5340, B2 => 
                           n4148, ZN => n5926);
   U5032 : NOR4_X1 port map( A1 => n5927, A2 => n5928, A3 => n5929, A4 => n5930
                           , ZN => n5917);
   U5033 : OAI221_X1 port map( B1 => n3925, B2 => n5345, C1 => n4309, C2 => 
                           n5346, A => n5931, ZN => n5930);
   U5034 : AOI22_X1 port map( A1 => n5348, A2 => n3765, B1 => n5349, B2 => 
                           n4149, ZN => n5931);
   U5035 : OAI221_X1 port map( B1 => n3926, B2 => n5350, C1 => n4310, C2 => 
                           n5351, A => n5932, ZN => n5929);
   U5036 : AOI22_X1 port map( A1 => n5353, A2 => n3766, B1 => n5354, B2 => 
                           n4150, ZN => n5932);
   U5037 : OAI221_X1 port map( B1 => n3927, B2 => n5355, C1 => n4311, C2 => 
                           n5356, A => n5933, ZN => n5928);
   U5038 : AOI22_X1 port map( A1 => n5358, A2 => n3767, B1 => n5359, B2 => 
                           n4151, ZN => n5933);
   U5039 : OAI221_X1 port map( B1 => n3928, B2 => n5360, C1 => n4312, C2 => 
                           n5361, A => n5934, ZN => n5927);
   U5040 : AOI22_X1 port map( A1 => n5363, A2 => n3768, B1 => n5364, B2 => 
                           n4152, ZN => n5934);
   U5041 : MUX2_X1 port map( A => OUT1_0_port, B => n5935, S => n5314, Z => 
                           n2526);
   U5042 : NAND2_X1 port map( A1 => n5936, A2 => n5937, ZN => n5935);
   U5043 : NOR4_X1 port map( A1 => n5938, A2 => n5939, A3 => n5940, A4 => n5941
                           , ZN => n5937);
   U5044 : OAI221_X1 port map( B1 => n32, B2 => n5321, C1 => n64, C2 => n5322, 
                           A => n5942, ZN => n5941);
   U5045 : AOI22_X1 port map( A1 => n5324, A2 => n5973, B1 => n5325, B2 => 
                           n5974, ZN => n5942);
   U5046 : OAI221_X1 port map( B1 => n160, B2 => n5326, C1 => n192, C2 => n5327
                           , A => n5947, ZN => n5940);
   U5047 : AOI22_X1 port map( A1 => n5329, A2 => n5971, B1 => n5330, B2 => 
                           n5972, ZN => n5947);
   U5048 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => n5950, 
                           ZN => n5945);
   U5049 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => 
                           ADD_RD1(0), ZN => n5943);
   U5050 : OAI221_X1 port map( B1 => n320, B2 => n5331, C1 => n288, C2 => n5332
                           , A => n5951, ZN => n5939);
   U5051 : AOI22_X1 port map( A1 => n5334, A2 => n3997, B1 => n5335, B2 => 
                           n4381, ZN => n5951);
   U5052 : OAI221_X1 port map( B1 => n3929, B2 => n5336, C1 => n4313, C2 => 
                           n5337, A => n5954, ZN => n5938);
   U5053 : AOI22_X1 port map( A1 => n5339, A2 => n3769, B1 => n5340, B2 => 
                           n4153, ZN => n5954);
   U5054 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(4), A3 => n5955, 
                           ZN => n5953);
   U5055 : NOR3_X1 port map( A1 => n5950, A2 => ADD_RD1(4), A3 => n5955, ZN => 
                           n5952);
   U5056 : NOR4_X1 port map( A1 => n5956, A2 => n5957, A3 => n5958, A4 => n5959
                           , ZN => n5936);
   U5057 : OAI221_X1 port map( B1 => n3930, B2 => n5345, C1 => n4314, C2 => 
                           n5346, A => n5960, ZN => n5959);
   U5058 : AOI22_X1 port map( A1 => n5348, A2 => n3770, B1 => n5349, B2 => 
                           n4154, ZN => n5960);
   U5059 : OAI221_X1 port map( B1 => n3931, B2 => n5350, C1 => n4315, C2 => 
                           n5351, A => n5963, ZN => n5958);
   U5060 : AOI22_X1 port map( A1 => n5353, A2 => n3771, B1 => n5354, B2 => 
                           n4155, ZN => n5963);
   U5061 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(3), A3 => n5964, 
                           ZN => n5962);
   U5062 : NOR3_X1 port map( A1 => n5950, A2 => ADD_RD1(3), A3 => n5964, ZN => 
                           n5961);
   U5063 : OAI221_X1 port map( B1 => n3932, B2 => n5355, C1 => n4316, C2 => 
                           n5356, A => n5965, ZN => n5957);
   U5064 : AOI22_X1 port map( A1 => n5358, A2 => n3772, B1 => n5359, B2 => 
                           n4156, ZN => n5965);
   U5065 : NOR2_X1 port map( A1 => n5968, A2 => ADD_RD1(2), ZN => n5944);
   U5066 : OAI221_X1 port map( B1 => n3933, B2 => n5360, C1 => n4317, C2 => 
                           n5361, A => n5969, ZN => n5956);
   U5067 : AOI22_X1 port map( A1 => n5363, A2 => n3773, B1 => n5364, B2 => 
                           n4157, ZN => n5969);
   U5068 : NOR2_X1 port map( A1 => n5970, A2 => n5968, ZN => n5948);
   U5069 : INV_X1 port map( A => ADD_RD1(1), ZN => n5968);
   U5070 : NOR3_X1 port map( A1 => n5955, A2 => ADD_RD1(0), A3 => n5964, ZN => 
                           n5967);
   U5071 : NOR2_X1 port map( A1 => n5970, A2 => ADD_RD1(1), ZN => n5949);
   U5072 : INV_X1 port map( A => ADD_RD1(2), ZN => n5970);
   U5073 : NOR3_X1 port map( A1 => n5955, A2 => n5950, A3 => n5964, ZN => n5966
                           );
   U5074 : INV_X1 port map( A => ADD_RD1(4), ZN => n5964);
   U5075 : INV_X1 port map( A => ADD_RD1(0), ZN => n5950);
   U5076 : INV_X1 port map( A => ADD_RD1(3), ZN => n5955);

end SYN_Behavioural;
