
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_WRF_DATA_W8_N_WIN3_N_REG_PER_WIN5_N_GLOBAL_REG5 is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type wrf_op is (WRF_NO_OP, WRF_OPN_CTX, WRF_CLS_CTX);
attribute ENUM_ENCODING of wrf_op : type is "00 01 10";
type wrf_state is (INACTIVE_s, READY_s, FILL_s, SPILL_s);
attribute ENUM_ENCODING of wrf_state : type is "00 01 10 11";
   
   -- Declarations for conversion functions.
   function wrf_op_to_std_logic_vector(arg : in wrf_op) return std_logic_vector
               ;
   function std_logic_vector_to_wrf_state(arg : in std_logic_vector( 1 to 2 )) 
               return wrf_state;

end CONV_PACK_WRF_DATA_W8_N_WIN3_N_REG_PER_WIN5_N_GLOBAL_REG5;

package body CONV_PACK_WRF_DATA_W8_N_WIN3_N_REG_PER_WIN5_N_GLOBAL_REG5 is
   
   -- enum type to std_logic_vector function
   function wrf_op_to_std_logic_vector(arg : in wrf_op) return std_logic_vector
   is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when WRF_NO_OP => return "00";
         when WRF_OPN_CTX => return "01";
         when WRF_CLS_CTX => return "10";
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return "00";
      end case;
   end;
   
   -- std_logic_vector to enum type function
   function std_logic_vector_to_wrf_state(arg : in std_logic_vector( 1 to 2 )) 
   return wrf_state is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when "00" => return INACTIVE_s;
         when "01" => return READY_s;
         when "10" => return FILL_s;
         when "11" => return SPILL_s;
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return INACTIVE_s;
      end case;
   end;

end CONV_PACK_WRF_DATA_W8_N_WIN3_N_REG_PER_WIN5_N_GLOBAL_REG5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_WRF_DATA_W8_N_WIN3_N_REG_PER_WIN5_N_GLOBAL_REG5.all;

entity ADDR_DEC_N_GLOBAL_REG5_N_REG_PER_WIN5_N_WIN3_0_DW01_add_0 is

   port( A, B : in std_logic_vector (5 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (5 downto 0);  CO : out std_logic);

end ADDR_DEC_N_GLOBAL_REG5_N_REG_PER_WIN5_N_WIN3_0_DW01_add_0;

architecture SYN_rpl of 
   ADDR_DEC_N_GLOBAL_REG5_N_REG_PER_WIN5_N_WIN3_0_DW01_add_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_4_port, carry_3_port, carry_2_port, n2, n5 : std_logic;

begin
   
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n2, CO => carry_2_port, S
                           => SUM(1));
   U1 : XNOR2_X1 port map( A => B(5), B => n5, ZN => SUM(5));
   U2 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n2);
   U3 : NAND2_X1 port map( A1 => B(4), A2 => carry_4_port, ZN => n5);
   U4 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U5 : XOR2_X1 port map( A => B(4), B => carry_4_port, Z => SUM(4));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_WRF_DATA_W8_N_WIN3_N_REG_PER_WIN5_N_GLOBAL_REG5.all;

entity ADDR_DEC_N_GLOBAL_REG5_N_REG_PER_WIN5_N_WIN3_2_DW01_add_0 is

   port( A, B : in std_logic_vector (5 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (5 downto 0);  CO : out std_logic);

end ADDR_DEC_N_GLOBAL_REG5_N_REG_PER_WIN5_N_WIN3_2_DW01_add_0;

architecture SYN_rpl of 
   ADDR_DEC_N_GLOBAL_REG5_N_REG_PER_WIN5_N_WIN3_2_DW01_add_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_4_port, carry_3_port, carry_2_port, n2, n5 : std_logic;

begin
   
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n2, CO => carry_2_port, S
                           => SUM(1));
   U1 : XNOR2_X1 port map( A => B(5), B => n5, ZN => SUM(5));
   U2 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n2);
   U3 : NAND2_X1 port map( A1 => B(4), A2 => carry_4_port, ZN => n5);
   U4 : XOR2_X1 port map( A => B(4), B => carry_4_port, Z => SUM(4));
   U5 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_WRF_DATA_W8_N_WIN3_N_REG_PER_WIN5_N_GLOBAL_REG5.all;

entity ADDR_DEC_N_GLOBAL_REG5_N_REG_PER_WIN5_N_WIN3_1_DW01_add_0 is

   port( A, B : in std_logic_vector (5 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (5 downto 0);  CO : out std_logic);

end ADDR_DEC_N_GLOBAL_REG5_N_REG_PER_WIN5_N_WIN3_1_DW01_add_0;

architecture SYN_rpl of 
   ADDR_DEC_N_GLOBAL_REG5_N_REG_PER_WIN5_N_WIN3_1_DW01_add_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_4_port, carry_3_port, carry_2_port, n2, n5 : std_logic;

begin
   
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => n2, CO => carry_2_port, S
                           => SUM(1));
   U1 : XNOR2_X1 port map( A => B(5), B => n5, ZN => SUM(5));
   U2 : AND2_X1 port map( A1 => B(0), A2 => A(0), ZN => n2);
   U3 : NAND2_X1 port map( A1 => B(4), A2 => carry_4_port, ZN => n5);
   U4 : XOR2_X1 port map( A => B(4), B => carry_4_port, Z => SUM(4));
   U5 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_WRF_DATA_W8_N_WIN3_N_REG_PER_WIN5_N_GLOBAL_REG5.all;

entity ADDR_DEC_N_GLOBAL_REG5_N_REG_PER_WIN5_N_WIN3_2 is

   port( VIRT_ADDR : in std_logic_vector (4 downto 0);  CWP : in 
         std_logic_vector (5 downto 0);  PHY_ADDR : out std_logic_vector (5 
         downto 0));

end ADDR_DEC_N_GLOBAL_REG5_N_REG_PER_WIN5_N_WIN3_2;

architecture SYN_Behavioural2 of ADDR_DEC_N_GLOBAL_REG5_N_REG_PER_WIN5_N_WIN3_2
   is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component ADDR_DEC_N_GLOBAL_REG5_N_REG_PER_WIN5_N_WIN3_2_DW01_add_0
      port( A, B : in std_logic_vector (5 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (5 downto 0);  CO : out std_logic);
   end component;
   
   signal N6, N7, N8, N9, N10, N31, U3_U1_Z_0, U3_U1_Z_1, U3_U1_Z_2, U3_U1_Z_3,
      U3_U2_Z_5, N16, N15, N14, sub_109_carry_3_port, sub_109_carry_4_port, 
      sub_109_carry_5_port, n1, n2, n3, n4, n5, n6_port, n7_port, n8_port, 
      n9_port, n10_port, n11, n12, n13, n14_port, n15_port, n16_port, n17, n18,
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n35, n36, n37, n38
      , n39, n40, n_1012 : std_logic;

begin
   
   n40 <= '0';
   r21 : ADDR_DEC_N_GLOBAL_REG5_N_REG_PER_WIN5_N_WIN3_2_DW01_add_0 port map( 
                           A(5) => n40, A(4) => n9_port, A(3) => U3_U1_Z_3, 
                           A(2) => U3_U1_Z_2, A(1) => U3_U1_Z_1, A(0) => 
                           U3_U1_Z_0, B(5) => U3_U2_Z_5, B(4) => n38, B(3) => 
                           n37, B(2) => n39, B(1) => n36, B(0) => n35, CI => 
                           n40, SUM(5) => N10, SUM(4) => N9, SUM(3) => N8, 
                           SUM(2) => N7, SUM(1) => N6, SUM(0) => PHY_ADDR(0), 
                           CO => n_1012);
   U3 : XOR2_X1 port map( A => n29, B => sub_109_carry_5_port, Z => n1);
   U4 : XOR2_X1 port map( A => N10, B => n8_port, Z => N31);
   U5 : XOR2_X1 port map( A => N9, B => n6_port, Z => n2);
   U6 : NAND2_X1 port map( A1 => N9, A2 => n6_port, ZN => n8_port);
   U7 : XOR2_X1 port map( A => N8, B => n5, Z => n3);
   U8 : XNOR2_X1 port map( A => n27, B => sub_109_carry_3_port, ZN => N15);
   U9 : XNOR2_X1 port map( A => n25, B => n28, ZN => N14);
   U10 : XOR2_X1 port map( A => N7, B => N6, Z => n4);
   U11 : OR2_X1 port map( A1 => n25, A2 => n28, ZN => sub_109_carry_3_port);
   U12 : OR2_X1 port map( A1 => n27, A2 => sub_109_carry_3_port, ZN => 
                           sub_109_carry_4_port);
   U13 : XNOR2_X1 port map( A => n26, B => sub_109_carry_4_port, ZN => N16);
   U14 : AND2_X1 port map( A1 => N7, A2 => N6, ZN => n5);
   U15 : AND2_X1 port map( A1 => N8, A2 => n5, ZN => n6_port);
   U17 : NAND2_X1 port map( A1 => CWP(4), A2 => n7_port, ZN => 
                           sub_109_carry_5_port);
   U18 : INV_X1 port map( A => sub_109_carry_4_port, ZN => n7_port);
   U19 : INV_X1 port map( A => CWP(3), ZN => n27);
   U20 : INV_X1 port map( A => CWP(2), ZN => n25);
   U21 : MUX2_X1 port map( A => N10, B => N31, S => n10_port, Z => PHY_ADDR(5))
                           ;
   U22 : MUX2_X1 port map( A => N9, B => n2, S => n10_port, Z => PHY_ADDR(4));
   U23 : MUX2_X1 port map( A => N8, B => n3, S => n10_port, Z => PHY_ADDR(3));
   U24 : MUX2_X1 port map( A => N7, B => n4, S => n10_port, Z => PHY_ADDR(2));
   U25 : XOR2_X1 port map( A => N6, B => n10_port, Z => PHY_ADDR(1));
   U26 : AOI211_X1 port map( C1 => n11, C2 => N15, A => n12, B => n13, ZN => 
                           n10_port);
   U27 : OR3_X1 port map( A1 => n14_port, A2 => n1, A3 => N16, ZN => n13);
   U28 : INV_X1 port map( A => n15_port, ZN => n14_port);
   U29 : OAI221_X1 port map( B1 => n11, B2 => N15, C1 => n16_port, C2 => N14, A
                           => n17, ZN => n15_port);
   U30 : INV_X1 port map( A => n18, ZN => n17);
   U31 : AOI221_X1 port map( B1 => N14, B2 => n16_port, C1 => n19, C2 => n20, A
                           => n21, ZN => n18);
   U32 : AOI21_X1 port map( B1 => CWP(0), B2 => VIRT_ADDR(0), A => n28, ZN => 
                           n21);
   U33 : NAND3_X1 port map( A1 => VIRT_ADDR(0), A2 => n28, A3 => CWP(0), ZN => 
                           n19);
   U34 : INV_X1 port map( A => CWP(1), ZN => n28);
   U35 : MUX2_X1 port map( A => VIRT_ADDR(0), B => CWP(0), S => n22, Z => n35);
   U36 : MUX2_X1 port map( A => VIRT_ADDR(1), B => CWP(1), S => n22, Z => n36);
   U37 : MUX2_X1 port map( A => VIRT_ADDR(3), B => CWP(3), S => n22, Z => n37);
   U38 : OAI21_X1 port map( B1 => n26, B2 => n12, A => n23, ZN => n38);
   U39 : INV_X1 port map( A => CWP(4), ZN => n26);
   U40 : MUX2_X1 port map( A => VIRT_ADDR(2), B => CWP(2), S => n22, Z => n39);
   U41 : NOR2_X1 port map( A1 => n29, A2 => n12, ZN => U3_U2_Z_5);
   U42 : INV_X1 port map( A => CWP(5), ZN => n29);
   n9_port <= '0';
   U44 : NAND2_X1 port map( A1 => n22, A2 => n11, ZN => U3_U1_Z_3);
   U45 : INV_X1 port map( A => VIRT_ADDR(3), ZN => n11);
   U46 : NAND2_X1 port map( A1 => n22, A2 => n16_port, ZN => U3_U1_Z_2);
   U47 : INV_X1 port map( A => VIRT_ADDR(2), ZN => n16_port);
   U48 : NAND2_X1 port map( A1 => n22, A2 => n20, ZN => U3_U1_Z_1);
   U49 : INV_X1 port map( A => VIRT_ADDR(1), ZN => n20);
   U50 : INV_X1 port map( A => n12, ZN => n22);
   U51 : OR2_X1 port map( A1 => n12, A2 => VIRT_ADDR(0), ZN => U3_U1_Z_0);
   U52 : NAND2_X1 port map( A1 => n23, A2 => n24, ZN => n12);
   U53 : NAND4_X1 port map( A1 => VIRT_ADDR(0), A2 => VIRT_ADDR(1), A3 => 
                           VIRT_ADDR(2), A4 => VIRT_ADDR(3), ZN => n24);
   U54 : INV_X1 port map( A => VIRT_ADDR(4), ZN => n23);

end SYN_Behavioural2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_WRF_DATA_W8_N_WIN3_N_REG_PER_WIN5_N_GLOBAL_REG5.all;

entity ADDR_DEC_N_GLOBAL_REG5_N_REG_PER_WIN5_N_WIN3_1 is

   port( VIRT_ADDR : in std_logic_vector (4 downto 0);  CWP : in 
         std_logic_vector (5 downto 0);  PHY_ADDR : out std_logic_vector (5 
         downto 0));

end ADDR_DEC_N_GLOBAL_REG5_N_REG_PER_WIN5_N_WIN3_1;

architecture SYN_Behavioural2 of ADDR_DEC_N_GLOBAL_REG5_N_REG_PER_WIN5_N_WIN3_1
   is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component ADDR_DEC_N_GLOBAL_REG5_N_REG_PER_WIN5_N_WIN3_1_DW01_add_0
      port( A, B : in std_logic_vector (5 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (5 downto 0);  CO : out std_logic);
   end component;
   
   signal N6, N7, N8, N9, N10, N31, U3_U1_Z_0, U3_U1_Z_1, U3_U1_Z_2, U3_U1_Z_3,
      U3_U2_Z_5, N16, N15, N14, sub_109_carry_3_port, sub_109_carry_4_port, 
      sub_109_carry_5_port, n1, n2, n3, n4, n5, n6_port, n7_port, n8_port, 
      n9_port, n10_port, n11, n12, n13, n14_port, n15_port, n16_port, n17, n18,
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n35, n36, n37, n38
      , n39, n40, n_1013 : std_logic;

begin
   
   n40 <= '0';
   r21 : ADDR_DEC_N_GLOBAL_REG5_N_REG_PER_WIN5_N_WIN3_1_DW01_add_0 port map( 
                           A(5) => n40, A(4) => n9_port, A(3) => U3_U1_Z_3, 
                           A(2) => U3_U1_Z_2, A(1) => U3_U1_Z_1, A(0) => 
                           U3_U1_Z_0, B(5) => U3_U2_Z_5, B(4) => n38, B(3) => 
                           n37, B(2) => n39, B(1) => n36, B(0) => n35, CI => 
                           n40, SUM(5) => N10, SUM(4) => N9, SUM(3) => N8, 
                           SUM(2) => N7, SUM(1) => N6, SUM(0) => PHY_ADDR(0), 
                           CO => n_1013);
   U3 : XOR2_X1 port map( A => n29, B => sub_109_carry_5_port, Z => n1);
   U4 : XOR2_X1 port map( A => N10, B => n8_port, Z => N31);
   U5 : XOR2_X1 port map( A => N9, B => n6_port, Z => n2);
   U6 : NAND2_X1 port map( A1 => N9, A2 => n6_port, ZN => n8_port);
   U7 : XOR2_X1 port map( A => N8, B => n5, Z => n3);
   U8 : XNOR2_X1 port map( A => n27, B => sub_109_carry_3_port, ZN => N15);
   U9 : XNOR2_X1 port map( A => n25, B => n28, ZN => N14);
   U10 : XOR2_X1 port map( A => N7, B => N6, Z => n4);
   U11 : OR2_X1 port map( A1 => n25, A2 => n28, ZN => sub_109_carry_3_port);
   U12 : OR2_X1 port map( A1 => n27, A2 => sub_109_carry_3_port, ZN => 
                           sub_109_carry_4_port);
   U13 : XNOR2_X1 port map( A => n26, B => sub_109_carry_4_port, ZN => N16);
   U14 : AND2_X1 port map( A1 => N7, A2 => N6, ZN => n5);
   U15 : AND2_X1 port map( A1 => N8, A2 => n5, ZN => n6_port);
   U17 : NAND2_X1 port map( A1 => CWP(4), A2 => n7_port, ZN => 
                           sub_109_carry_5_port);
   U18 : INV_X1 port map( A => sub_109_carry_4_port, ZN => n7_port);
   U19 : INV_X1 port map( A => CWP(3), ZN => n27);
   U20 : INV_X1 port map( A => CWP(2), ZN => n25);
   U21 : MUX2_X1 port map( A => N10, B => N31, S => n10_port, Z => PHY_ADDR(5))
                           ;
   U22 : MUX2_X1 port map( A => N9, B => n2, S => n10_port, Z => PHY_ADDR(4));
   U23 : MUX2_X1 port map( A => N8, B => n3, S => n10_port, Z => PHY_ADDR(3));
   U24 : MUX2_X1 port map( A => N7, B => n4, S => n10_port, Z => PHY_ADDR(2));
   U25 : XOR2_X1 port map( A => N6, B => n10_port, Z => PHY_ADDR(1));
   U26 : AOI211_X1 port map( C1 => n11, C2 => N15, A => n12, B => n13, ZN => 
                           n10_port);
   U27 : OR3_X1 port map( A1 => n14_port, A2 => n1, A3 => N16, ZN => n13);
   U28 : INV_X1 port map( A => n15_port, ZN => n14_port);
   U29 : OAI221_X1 port map( B1 => n11, B2 => N15, C1 => n16_port, C2 => N14, A
                           => n17, ZN => n15_port);
   U30 : INV_X1 port map( A => n18, ZN => n17);
   U31 : AOI221_X1 port map( B1 => N14, B2 => n16_port, C1 => n19, C2 => n20, A
                           => n21, ZN => n18);
   U32 : AOI21_X1 port map( B1 => CWP(0), B2 => VIRT_ADDR(0), A => n28, ZN => 
                           n21);
   U33 : NAND3_X1 port map( A1 => VIRT_ADDR(0), A2 => n28, A3 => CWP(0), ZN => 
                           n19);
   U34 : INV_X1 port map( A => CWP(1), ZN => n28);
   U35 : MUX2_X1 port map( A => VIRT_ADDR(0), B => CWP(0), S => n22, Z => n35);
   U36 : MUX2_X1 port map( A => VIRT_ADDR(1), B => CWP(1), S => n22, Z => n36);
   U37 : MUX2_X1 port map( A => VIRT_ADDR(3), B => CWP(3), S => n22, Z => n37);
   U38 : OAI21_X1 port map( B1 => n26, B2 => n12, A => n23, ZN => n38);
   U39 : INV_X1 port map( A => CWP(4), ZN => n26);
   U40 : MUX2_X1 port map( A => VIRT_ADDR(2), B => CWP(2), S => n22, Z => n39);
   U41 : NOR2_X1 port map( A1 => n29, A2 => n12, ZN => U3_U2_Z_5);
   U42 : INV_X1 port map( A => CWP(5), ZN => n29);
   n9_port <= '0';
   U44 : NAND2_X1 port map( A1 => n22, A2 => n11, ZN => U3_U1_Z_3);
   U45 : INV_X1 port map( A => VIRT_ADDR(3), ZN => n11);
   U46 : NAND2_X1 port map( A1 => n22, A2 => n16_port, ZN => U3_U1_Z_2);
   U47 : INV_X1 port map( A => VIRT_ADDR(2), ZN => n16_port);
   U48 : NAND2_X1 port map( A1 => n22, A2 => n20, ZN => U3_U1_Z_1);
   U49 : INV_X1 port map( A => VIRT_ADDR(1), ZN => n20);
   U50 : INV_X1 port map( A => n12, ZN => n22);
   U51 : OR2_X1 port map( A1 => n12, A2 => VIRT_ADDR(0), ZN => U3_U1_Z_0);
   U52 : NAND2_X1 port map( A1 => n23, A2 => n24, ZN => n12);
   U53 : NAND4_X1 port map( A1 => VIRT_ADDR(0), A2 => VIRT_ADDR(1), A3 => 
                           VIRT_ADDR(2), A4 => VIRT_ADDR(3), ZN => n24);
   U54 : INV_X1 port map( A => VIRT_ADDR(4), ZN => n23);

end SYN_Behavioural2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_WRF_DATA_W8_N_WIN3_N_REG_PER_WIN5_N_GLOBAL_REG5.all;

entity RF_ADDR_W6_DATA_W8 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (5 downto 0);  DATAIN : in 
         std_logic_vector (7 downto 0);  OUT1, OUT2 : out std_logic_vector (7 
         downto 0));

end RF_ADDR_W6_DATA_W8;

architecture SYN_Behavioural of RF_ADDR_W6_DATA_W8 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal OUT1_7_port, OUT1_6_port, OUT1_5_port, OUT1_4_port, OUT1_3_port, 
      OUT1_2_port, OUT1_1_port, OUT1_0_port, OUT2_7_port, OUT2_6_port, 
      OUT2_5_port, OUT2_4_port, OUT2_3_port, OUT2_2_port, OUT2_1_port, 
      OUT2_0_port, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, 
      n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, 
      n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, 
      n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, 
      n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, 
      n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, 
      n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, 
      n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, 
      n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, 
      n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, 
      n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, 
      n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, 
      n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, 
      n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, 
      n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, 
      n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, 
      n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, 
      n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, 
      n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, 
      n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, 
      n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, 
      n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, 
      n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, 
      n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, 
      n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, 
      n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, 
      n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, 
      n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, 
      n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, 
      n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, 
      n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, 
      n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, 
      n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, 
      n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, 
      n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, 
      n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, 
      n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, 
      n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, 
      n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, 
      n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, 
      n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, 
      n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, 
      n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, 
      n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, 
      n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, 
      n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, 
      n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, 
      n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, 
      n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, 
      n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, 
      n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, 
      n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, 
      n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, 
      n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, 
      n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, 
      n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, 
      n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, 
      n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, 
      n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, 
      n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, 
      n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, 
      n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, 
      n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, 
      n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, 
      n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, 
      n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, 
      n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, 
      n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, 
      n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, 
      n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, 
      n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, 
      n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, 
      n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, 
      n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, 
      n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, 
      n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, 
      n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, 
      n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, 
      n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, 
      n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, 
      n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, 
      n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, 
      n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, 
      n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, 
      n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, 
      n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, 
      n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, 
      n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, 
      n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, 
      n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, 
      n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, 
      n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, 
      n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, 
      n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, 
      n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, 
      n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, 
      n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, 
      n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, 
      n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, 
      n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, 
      n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, 
      n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, 
      n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, 
      n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, 
      n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, 
      n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, 
      n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, 
      n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, 
      n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, 
      n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, 
      n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, 
      n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, 
      n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, 
      n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, 
      n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, 
      n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, 
      n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, 
      n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, 
      n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, 
      n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, 
      n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, 
      n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, 
      n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, 
      n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, 
      n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, 
      n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, 
      n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, 
      n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, 
      n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, 
      n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, 
      n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, 
      n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, 
      n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, 
      n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, 
      n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, 
      n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, 
      n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, 
      n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, 
      n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, 
      n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, 
      n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, 
      n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, 
      n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, 
      n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, 
      n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, 
      n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, 
      n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, 
      n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, 
      n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, 
      n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, 
      n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, 
      n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, 
      n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, 
      n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, 
      n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, 
      n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, 
      n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, 
      n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, 
      n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, 
      n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, 
      n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, 
      n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, 
      n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, 
      n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, 
      n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, 
      n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, 
      n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, 
      n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, 
      n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, 
      n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, 
      n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, 
      n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, 
      n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, 
      n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, 
      n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, 
      n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, 
      n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, 
      n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, 
      n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, 
      n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, 
      n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, 
      n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, 
      n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, 
      n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, 
      n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, 
      n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, 
      n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, 
      n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, 
      n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, 
      n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, 
      n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, 
      n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, 
      n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, 
      n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, 
      n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, 
      n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, 
      n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, 
      n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, 
      n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, 
      n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, 
      n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, 
      n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, 
      n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, 
      n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, 
      n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, 
      n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, 
      n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, 
      n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, 
      n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, 
      n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, 
      n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, 
      n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, 
      n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, 
      n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, 
      n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, 
      n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, 
      n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, 
      n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n_1014, 
      n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, 
      n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, 
      n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, 
      n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, 
      n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, 
      n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, 
      n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, 
      n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, 
      n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, 
      n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, 
      n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, 
      n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, 
      n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, 
      n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, 
      n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, 
      n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, 
      n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, 
      n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, 
      n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, 
      n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, 
      n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, 
      n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, 
      n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, 
      n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, 
      n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, 
      n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, 
      n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, 
      n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, 
      n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, 
      n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, 
      n_1285 : std_logic;

begin
   OUT1 <= ( OUT1_7_port, OUT1_6_port, OUT1_5_port, OUT1_4_port, OUT1_3_port, 
      OUT1_2_port, OUT1_1_port, OUT1_0_port );
   OUT2 <= ( OUT2_7_port, OUT2_6_port, OUT2_5_port, OUT2_4_port, OUT2_3_port, 
      OUT2_2_port, OUT2_1_port, OUT2_0_port );
   
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n2002, CK => CLK, Q => n2306,
                           QN => n3831);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n2001, CK => CLK, Q => n3830,
                           QN => n2221);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n2000, CK => CLK, Q => n3829,
                           QN => n2233);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n1999, CK => CLK, Q => n3828,
                           QN => n2244);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n1998, CK => CLK, Q => n3827,
                           QN => n2255);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n1997, CK => CLK, Q => n3826,
                           QN => n2266);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n1996, CK => CLK, Q => n3825,
                           QN => n2277);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n1995, CK => CLK, Q => n3824,
                           QN => n2288);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n1994, CK => CLK, Q => n3823,
                           QN => n2291);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n1993, CK => CLK, Q => n2328,
                           QN => n3822);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n1992, CK => CLK, Q => n2329,
                           QN => n3821);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n1991, CK => CLK, Q => n2330,
                           QN => n3820);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n1990, CK => CLK, Q => n2331,
                           QN => n3819);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n1989, CK => CLK, Q => n2332,
                           QN => n3818);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n1988, CK => CLK, Q => n2333,
                           QN => n3817);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n1987, CK => CLK, Q => n2334,
                           QN => n3816);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n1986, CK => CLK, Q => n3344,
                           QN => n_1014);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n1985, CK => CLK, Q => n3376,
                           QN => n_1015);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n1984, CK => CLK, Q => n3408,
                           QN => n_1016);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n1983, CK => CLK, Q => n3440,
                           QN => n_1017);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n1982, CK => CLK, Q => n3472,
                           QN => n_1018);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n1981, CK => CLK, Q => n3504,
                           QN => n_1019);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n1980, CK => CLK, Q => n3536,
                           QN => n_1020);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n1979, CK => CLK, Q => n3568,
                           QN => n_1021);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n1978, CK => CLK, Q => n3345,
                           QN => n_1022);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n1977, CK => CLK, Q => n3377,
                           QN => n_1023);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n1976, CK => CLK, Q => n3409,
                           QN => n_1024);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n1975, CK => CLK, Q => n3441,
                           QN => n_1025);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n1974, CK => CLK, Q => n3473,
                           QN => n_1026);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n1973, CK => CLK, Q => n3505,
                           QN => n_1027);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n1972, CK => CLK, Q => n3537,
                           QN => n_1028);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n1971, CK => CLK, Q => n3569,
                           QN => n_1029);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n1970, CK => CLK, Q => n3815,
                           QN => n2184);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n1969, CK => CLK, Q => n3814,
                           QN => n2186);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n1968, CK => CLK, Q => n3813,
                           QN => n2188);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n1967, CK => CLK, Q => n3812,
                           QN => n2190);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n1966, CK => CLK, Q => n3811,
                           QN => n2192);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n1965, CK => CLK, Q => n3810,
                           QN => n2194);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n1964, CK => CLK, Q => n3809,
                           QN => n2196);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n1963, CK => CLK, Q => n3808,
                           QN => n2198);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n1962, CK => CLK, Q => n3807,
                           QN => n2290);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n1961, CK => CLK, Q => n3806,
                           QN => n2293);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n1960, CK => CLK, Q => n3805,
                           QN => n2295);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n1959, CK => CLK, Q => n3804,
                           QN => n2297);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n1958, CK => CLK, Q => n3803,
                           QN => n2299);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n1957, CK => CLK, Q => n3802,
                           QN => n2301);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n1956, CK => CLK, Q => n3801,
                           QN => n2303);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n1955, CK => CLK, Q => n3800,
                           QN => n2305);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n1954, CK => CLK, Q => n3346,
                           QN => n_1030);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n1953, CK => CLK, Q => n3378,
                           QN => n_1031);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n1952, CK => CLK, Q => n3410,
                           QN => n_1032);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n1951, CK => CLK, Q => n3442,
                           QN => n_1033);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n1950, CK => CLK, Q => n3474,
                           QN => n_1034);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n1949, CK => CLK, Q => n3506,
                           QN => n_1035);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n1948, CK => CLK, Q => n3538,
                           QN => n_1036);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n1947, CK => CLK, Q => n3570,
                           QN => n_1037);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n1946, CK => CLK, Q => n3347,
                           QN => n_1038);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n1945, CK => CLK, Q => n3379,
                           QN => n_1039);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n1944, CK => CLK, Q => n3411,
                           QN => n_1040);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n1943, CK => CLK, Q => n3443,
                           QN => n_1041);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n1942, CK => CLK, Q => n3475,
                           QN => n_1042);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n1941, CK => CLK, Q => n3507,
                           QN => n_1043);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n1940, CK => CLK, Q => n3539,
                           QN => n_1044);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n1939, CK => CLK, Q => n3571,
                           QN => n_1045);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n1938, CK => CLK, Q => n3799,
                           QN => n2183);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n1937, CK => CLK, Q => n3798,
                           QN => n2185);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n1936, CK => CLK, Q => n3797,
                           QN => n2187);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n1935, CK => CLK, Q => n3796,
                           QN => n2189);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n1934, CK => CLK, Q => n3795,
                           QN => n2191);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n1933, CK => CLK, Q => n3794,
                           QN => n2193);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n1932, CK => CLK, Q => n3793,
                           QN => n2195);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n1931, CK => CLK, Q => n3792,
                           QN => n2197);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n1930, CK => CLK, Q => n3791,
                           QN => n2289);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n1929, CK => CLK, Q => n3790,
                           QN => n2292);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n1928, CK => CLK, Q => n3789,
                           QN => n2294);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n1927, CK => CLK, Q => n3788,
                           QN => n2296);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n1926, CK => CLK, Q => n3787,
                           QN => n2298);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n1925, CK => CLK, Q => n3786,
                           QN => n2300);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n1924, CK => CLK, Q => n3785,
                           QN => n2302);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n1923, CK => CLK, Q => n3784,
                           QN => n2304);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n1922, CK => CLK, Q => n3348
                           , QN => n_1046);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n1921, CK => CLK, Q => n3380
                           , QN => n_1047);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n1920, CK => CLK, Q => n3412
                           , QN => n_1048);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n1919, CK => CLK, Q => n3444
                           , QN => n_1049);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n1918, CK => CLK, Q => n3476
                           , QN => n_1050);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n1917, CK => CLK, Q => n3508
                           , QN => n_1051);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n1916, CK => CLK, Q => n3540
                           , QN => n_1052);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n1915, CK => CLK, Q => n3572
                           , QN => n_1053);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n1914, CK => CLK, Q => n3349
                           , QN => n_1054);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n1913, CK => CLK, Q => n3381
                           , QN => n_1055);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n1912, CK => CLK, Q => n3413
                           , QN => n_1056);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n1911, CK => CLK, Q => n3445
                           , QN => n_1057);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n1910, CK => CLK, Q => n3477
                           , QN => n_1058);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n1909, CK => CLK, Q => n3509
                           , QN => n_1059);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n1908, CK => CLK, Q => n3541
                           , QN => n_1060);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n1907, CK => CLK, Q => n3573
                           , QN => n_1061);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n1906, CK => CLK, Q => n3783
                           , QN => n2209);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n1905, CK => CLK, Q => n3782
                           , QN => n2220);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n1904, CK => CLK, Q => n3781
                           , QN => n2232);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n1903, CK => CLK, Q => n2307
                           , QN => n3780);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n1902, CK => CLK, Q => n2308
                           , QN => n3779);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n1901, CK => CLK, Q => n2309
                           , QN => n3778);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n1900, CK => CLK, Q => n2310
                           , QN => n3777);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n1899, CK => CLK, Q => n2311
                           , QN => n3776);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n1898, CK => CLK, Q => n2335
                           , QN => n3775);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n1897, CK => CLK, Q => n2336
                           , QN => n3774);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n1896, CK => CLK, Q => n2337
                           , QN => n3773);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n1895, CK => CLK, Q => n2338
                           , QN => n3772);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n1894, CK => CLK, Q => n2339
                           , QN => n3771);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n1893, CK => CLK, Q => n2340
                           , QN => n3770);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n1892, CK => CLK, Q => n2341
                           , QN => n3769);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n1891, CK => CLK, Q => n2342
                           , QN => n3768);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n1890, CK => CLK, Q => n3350
                           , QN => n_1062);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n1889, CK => CLK, Q => n3382
                           , QN => n_1063);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n1888, CK => CLK, Q => n3414
                           , QN => n_1064);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n1887, CK => CLK, Q => n3446
                           , QN => n_1065);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n1886, CK => CLK, Q => n3478
                           , QN => n_1066);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n1885, CK => CLK, Q => n3510
                           , QN => n_1067);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n1884, CK => CLK, Q => n3542
                           , QN => n_1068);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n1883, CK => CLK, Q => n3574
                           , QN => n_1069);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n1882, CK => CLK, Q => n3351
                           , QN => n_1070);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n1881, CK => CLK, Q => n3383
                           , QN => n_1071);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n1880, CK => CLK, Q => n3415
                           , QN => n_1072);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n1879, CK => CLK, Q => n3447
                           , QN => n_1073);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n1878, CK => CLK, Q => n3479
                           , QN => n_1074);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n1877, CK => CLK, Q => n3511
                           , QN => n_1075);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n1876, CK => CLK, Q => n3543
                           , QN => n_1076);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n1875, CK => CLK, Q => n3575
                           , QN => n_1077);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n1874, CK => CLK, Q => n2312
                           , QN => n3767);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n1873, CK => CLK, Q => n2313
                           , QN => n3766);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n1872, CK => CLK, Q => n2314
                           , QN => n3765);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n1871, CK => CLK, Q => n2315
                           , QN => n3764);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n1870, CK => CLK, Q => n2316
                           , QN => n3763);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n1869, CK => CLK, Q => n2317
                           , QN => n3762);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n1868, CK => CLK, Q => n2318
                           , QN => n3761);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n1867, CK => CLK, Q => n2319
                           , QN => n3760);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n1866, CK => CLK, Q => n2343
                           , QN => n3759);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n1865, CK => CLK, Q => n2344
                           , QN => n3758);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n1864, CK => CLK, Q => n2345
                           , QN => n3757);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n1863, CK => CLK, Q => n2346
                           , QN => n3756);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n1862, CK => CLK, Q => n2347
                           , QN => n3755);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n1861, CK => CLK, Q => n2348
                           , QN => n3754);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n1860, CK => CLK, Q => n2349
                           , QN => n3753);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n1859, CK => CLK, Q => n2350
                           , QN => n3752);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n1858, CK => CLK, Q => n3336
                           , QN => n_1078);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n1857, CK => CLK, Q => n3368
                           , QN => n_1079);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n1856, CK => CLK, Q => n3400
                           , QN => n_1080);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n1855, CK => CLK, Q => n3432
                           , QN => n_1081);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n1854, CK => CLK, Q => n3464
                           , QN => n_1082);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n1853, CK => CLK, Q => n3496
                           , QN => n_1083);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n1852, CK => CLK, Q => n3528
                           , QN => n_1084);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n1851, CK => CLK, Q => n3560
                           , QN => n_1085);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n1850, CK => CLK, Q => n3337
                           , QN => n_1086);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n1849, CK => CLK, Q => n3369
                           , QN => n_1087);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n1848, CK => CLK, Q => n3401
                           , QN => n_1088);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n1847, CK => CLK, Q => n3433
                           , QN => n_1089);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n1846, CK => CLK, Q => n3465
                           , QN => n_1090);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n1845, CK => CLK, Q => n3497
                           , QN => n_1091);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n1844, CK => CLK, Q => n3529
                           , QN => n_1092);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n1843, CK => CLK, Q => n3561
                           , QN => n_1093);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n1842, CK => CLK, Q => n2320
                           , QN => n3751);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n1841, CK => CLK, Q => n2321
                           , QN => n3750);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n1840, CK => CLK, Q => n2322
                           , QN => n3749);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n1839, CK => CLK, Q => n2323
                           , QN => n3748);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n1838, CK => CLK, Q => n2324
                           , QN => n3747);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n1837, CK => CLK, Q => n2325
                           , QN => n3746);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n1836, CK => CLK, Q => n2326
                           , QN => n3745);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n1835, CK => CLK, Q => n2327
                           , QN => n3744);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n1834, CK => CLK, Q => n2351
                           , QN => n3743);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n1833, CK => CLK, Q => n2352
                           , QN => n3742);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n1832, CK => CLK, Q => n2353
                           , QN => n3741);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n1831, CK => CLK, Q => n2354
                           , QN => n3740);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n1830, CK => CLK, Q => n2355
                           , QN => n3739);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n1829, CK => CLK, Q => n2356
                           , QN => n3738);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n1828, CK => CLK, Q => n2357
                           , QN => n3737);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n1827, CK => CLK, Q => n2358
                           , QN => n3736);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n1826, CK => CLK, Q => n3338
                           , QN => n_1094);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n1825, CK => CLK, Q => n3370
                           , QN => n_1095);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n1824, CK => CLK, Q => n3402
                           , QN => n_1096);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n1823, CK => CLK, Q => n3434
                           , QN => n_1097);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n1822, CK => CLK, Q => n3466
                           , QN => n_1098);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n1821, CK => CLK, Q => n3498
                           , QN => n_1099);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n1820, CK => CLK, Q => n3530
                           , QN => n_1100);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n1819, CK => CLK, Q => n3562
                           , QN => n_1101);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n1818, CK => CLK, Q => n3339
                           , QN => n_1102);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n1817, CK => CLK, Q => n3371
                           , QN => n_1103);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n1816, CK => CLK, Q => n3403
                           , QN => n_1104);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n1815, CK => CLK, Q => n3435
                           , QN => n_1105);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n1814, CK => CLK, Q => n3467
                           , QN => n_1106);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n1813, CK => CLK, Q => n3499
                           , QN => n_1107);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n1812, CK => CLK, Q => n3531
                           , QN => n_1108);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n1811, CK => CLK, Q => n3563
                           , QN => n_1109);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n1810, CK => CLK, Q => n3735
                           , QN => n2208);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n1809, CK => CLK, Q => n3734
                           , QN => n2219);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n1808, CK => CLK, Q => n3733
                           , QN => n2231);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n1807, CK => CLK, Q => n3732
                           , QN => n2243);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n1806, CK => CLK, Q => n3731
                           , QN => n2254);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n1805, CK => CLK, Q => n3730
                           , QN => n2265);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n1804, CK => CLK, Q => n3729
                           , QN => n2276);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n1803, CK => CLK, Q => n3728
                           , QN => n2287);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n1802, CK => CLK, Q => n2359
                           , QN => n3727);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n1801, CK => CLK, Q => n2360
                           , QN => n3726);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n1800, CK => CLK, Q => n2361
                           , QN => n3725);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n1799, CK => CLK, Q => n2362
                           , QN => n3724);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n1798, CK => CLK, Q => n2363
                           , QN => n3723);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n1797, CK => CLK, Q => n2364
                           , QN => n3722);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n1796, CK => CLK, Q => n2365
                           , QN => n3721);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n1795, CK => CLK, Q => n2366
                           , QN => n3720);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n1794, CK => CLK, Q => n3340
                           , QN => n_1110);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n1793, CK => CLK, Q => n3372
                           , QN => n_1111);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n1792, CK => CLK, Q => n3404
                           , QN => n_1112);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n1791, CK => CLK, Q => n3436
                           , QN => n_1113);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n1790, CK => CLK, Q => n3468
                           , QN => n_1114);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n1789, CK => CLK, Q => n3500
                           , QN => n_1115);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n1788, CK => CLK, Q => n3532
                           , QN => n_1116);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n1787, CK => CLK, Q => n3564
                           , QN => n_1117);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n1786, CK => CLK, Q => n3341
                           , QN => n_1118);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n1785, CK => CLK, Q => n3373
                           , QN => n_1119);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n1784, CK => CLK, Q => n3405
                           , QN => n_1120);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n1783, CK => CLK, Q => n3437
                           , QN => n_1121);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n1782, CK => CLK, Q => n3469
                           , QN => n_1122);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n1781, CK => CLK, Q => n3501
                           , QN => n_1123);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n1780, CK => CLK, Q => n3533
                           , QN => n_1124);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n1779, CK => CLK, Q => n3565
                           , QN => n_1125);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n1778, CK => CLK, Q => n3719
                           , QN => n2207);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n1777, CK => CLK, Q => n3718
                           , QN => n2218);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n1776, CK => CLK, Q => n3717
                           , QN => n2230);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n1775, CK => CLK, Q => n3716
                           , QN => n2242);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n1774, CK => CLK, Q => n3715
                           , QN => n2253);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n1773, CK => CLK, Q => n3714
                           , QN => n2264);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n1772, CK => CLK, Q => n3713
                           , QN => n2275);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n1771, CK => CLK, Q => n3712
                           , QN => n2286);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n1770, CK => CLK, Q => n2367
                           , QN => n3711);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n1769, CK => CLK, Q => n2368
                           , QN => n3710);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n1768, CK => CLK, Q => n2369
                           , QN => n3709);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n1767, CK => CLK, Q => n2370
                           , QN => n3708);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n1766, CK => CLK, Q => n2371
                           , QN => n3707);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n1765, CK => CLK, Q => n2372
                           , QN => n3706);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n1764, CK => CLK, Q => n2373
                           , QN => n3705);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n1763, CK => CLK, Q => n2374
                           , QN => n3704);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n1762, CK => CLK, Q => n3342
                           , QN => n_1126);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n1761, CK => CLK, Q => n3374
                           , QN => n_1127);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n1760, CK => CLK, Q => n3406
                           , QN => n_1128);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n1759, CK => CLK, Q => n3438
                           , QN => n_1129);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n1758, CK => CLK, Q => n3470
                           , QN => n_1130);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n1757, CK => CLK, Q => n3502
                           , QN => n_1131);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n1756, CK => CLK, Q => n3534
                           , QN => n_1132);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n1755, CK => CLK, Q => n3566
                           , QN => n_1133);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n1754, CK => CLK, Q => n3343
                           , QN => n_1134);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n1753, CK => CLK, Q => n3375
                           , QN => n_1135);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n1752, CK => CLK, Q => n3407
                           , QN => n_1136);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n1751, CK => CLK, Q => n3439
                           , QN => n_1137);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n1750, CK => CLK, Q => n3471
                           , QN => n_1138);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n1749, CK => CLK, Q => n3503
                           , QN => n_1139);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n1748, CK => CLK, Q => n3535
                           , QN => n_1140);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n1747, CK => CLK, Q => n3567
                           , QN => n_1141);
   REGISTERS_reg_32_7_inst : DFF_X1 port map( D => n1746, CK => CLK, Q => n3703
                           , QN => n2206);
   REGISTERS_reg_32_6_inst : DFF_X1 port map( D => n1745, CK => CLK, Q => n3702
                           , QN => n2217);
   REGISTERS_reg_32_5_inst : DFF_X1 port map( D => n1744, CK => CLK, Q => n3701
                           , QN => n2229);
   REGISTERS_reg_32_4_inst : DFF_X1 port map( D => n1743, CK => CLK, Q => n3700
                           , QN => n2241);
   REGISTERS_reg_32_3_inst : DFF_X1 port map( D => n1742, CK => CLK, Q => n3699
                           , QN => n2252);
   REGISTERS_reg_32_2_inst : DFF_X1 port map( D => n1741, CK => CLK, Q => n3698
                           , QN => n2263);
   REGISTERS_reg_32_1_inst : DFF_X1 port map( D => n1740, CK => CLK, Q => n3697
                           , QN => n2274);
   REGISTERS_reg_32_0_inst : DFF_X1 port map( D => n1739, CK => CLK, Q => n3696
                           , QN => n2285);
   REGISTERS_reg_33_7_inst : DFF_X1 port map( D => n1738, CK => CLK, Q => n2375
                           , QN => n3695);
   REGISTERS_reg_33_6_inst : DFF_X1 port map( D => n1737, CK => CLK, Q => n2376
                           , QN => n3694);
   REGISTERS_reg_33_5_inst : DFF_X1 port map( D => n1736, CK => CLK, Q => n2377
                           , QN => n3693);
   REGISTERS_reg_33_4_inst : DFF_X1 port map( D => n1735, CK => CLK, Q => n2378
                           , QN => n3692);
   REGISTERS_reg_33_3_inst : DFF_X1 port map( D => n1734, CK => CLK, Q => n2379
                           , QN => n3691);
   REGISTERS_reg_33_2_inst : DFF_X1 port map( D => n1733, CK => CLK, Q => n2380
                           , QN => n3690);
   REGISTERS_reg_33_1_inst : DFF_X1 port map( D => n1732, CK => CLK, Q => n2381
                           , QN => n3689);
   REGISTERS_reg_33_0_inst : DFF_X1 port map( D => n1731, CK => CLK, Q => n2382
                           , QN => n3688);
   REGISTERS_reg_34_7_inst : DFF_X1 port map( D => n1730, CK => CLK, Q => n3328
                           , QN => n_1142);
   REGISTERS_reg_34_6_inst : DFF_X1 port map( D => n1729, CK => CLK, Q => n3360
                           , QN => n_1143);
   REGISTERS_reg_34_5_inst : DFF_X1 port map( D => n1728, CK => CLK, Q => n3392
                           , QN => n_1144);
   REGISTERS_reg_34_4_inst : DFF_X1 port map( D => n1727, CK => CLK, Q => n3424
                           , QN => n_1145);
   REGISTERS_reg_34_3_inst : DFF_X1 port map( D => n1726, CK => CLK, Q => n3456
                           , QN => n_1146);
   REGISTERS_reg_34_2_inst : DFF_X1 port map( D => n1725, CK => CLK, Q => n3488
                           , QN => n_1147);
   REGISTERS_reg_34_1_inst : DFF_X1 port map( D => n1724, CK => CLK, Q => n3520
                           , QN => n_1148);
   REGISTERS_reg_34_0_inst : DFF_X1 port map( D => n1723, CK => CLK, Q => n3552
                           , QN => n_1149);
   REGISTERS_reg_35_7_inst : DFF_X1 port map( D => n1722, CK => CLK, Q => n3329
                           , QN => n_1150);
   REGISTERS_reg_35_6_inst : DFF_X1 port map( D => n1721, CK => CLK, Q => n3361
                           , QN => n_1151);
   REGISTERS_reg_35_5_inst : DFF_X1 port map( D => n1720, CK => CLK, Q => n3393
                           , QN => n_1152);
   REGISTERS_reg_35_4_inst : DFF_X1 port map( D => n1719, CK => CLK, Q => n3425
                           , QN => n_1153);
   REGISTERS_reg_35_3_inst : DFF_X1 port map( D => n1718, CK => CLK, Q => n3457
                           , QN => n_1154);
   REGISTERS_reg_35_2_inst : DFF_X1 port map( D => n1717, CK => CLK, Q => n3489
                           , QN => n_1155);
   REGISTERS_reg_35_1_inst : DFF_X1 port map( D => n1716, CK => CLK, Q => n3521
                           , QN => n_1156);
   REGISTERS_reg_35_0_inst : DFF_X1 port map( D => n1715, CK => CLK, Q => n3553
                           , QN => n_1157);
   REGISTERS_reg_36_7_inst : DFF_X1 port map( D => n1714, CK => CLK, Q => n3687
                           , QN => n2205);
   REGISTERS_reg_36_6_inst : DFF_X1 port map( D => n1713, CK => CLK, Q => n3686
                           , QN => n2216);
   REGISTERS_reg_36_5_inst : DFF_X1 port map( D => n1712, CK => CLK, Q => n3685
                           , QN => n2228);
   REGISTERS_reg_36_4_inst : DFF_X1 port map( D => n1711, CK => CLK, Q => n3684
                           , QN => n2240);
   REGISTERS_reg_36_3_inst : DFF_X1 port map( D => n1710, CK => CLK, Q => n3683
                           , QN => n2251);
   REGISTERS_reg_36_2_inst : DFF_X1 port map( D => n1709, CK => CLK, Q => n3682
                           , QN => n2262);
   REGISTERS_reg_36_1_inst : DFF_X1 port map( D => n1708, CK => CLK, Q => n3681
                           , QN => n2273);
   REGISTERS_reg_36_0_inst : DFF_X1 port map( D => n1707, CK => CLK, Q => n3680
                           , QN => n2284);
   REGISTERS_reg_37_7_inst : DFF_X1 port map( D => n1706, CK => CLK, Q => n2383
                           , QN => n3679);
   REGISTERS_reg_37_6_inst : DFF_X1 port map( D => n1705, CK => CLK, Q => n2384
                           , QN => n3678);
   REGISTERS_reg_37_5_inst : DFF_X1 port map( D => n1704, CK => CLK, Q => n2385
                           , QN => n3677);
   REGISTERS_reg_37_4_inst : DFF_X1 port map( D => n1703, CK => CLK, Q => n2386
                           , QN => n3676);
   REGISTERS_reg_37_3_inst : DFF_X1 port map( D => n1702, CK => CLK, Q => n2387
                           , QN => n3675);
   REGISTERS_reg_37_2_inst : DFF_X1 port map( D => n1701, CK => CLK, Q => n2388
                           , QN => n3674);
   REGISTERS_reg_37_1_inst : DFF_X1 port map( D => n1700, CK => CLK, Q => n2389
                           , QN => n3673);
   REGISTERS_reg_37_0_inst : DFF_X1 port map( D => n1699, CK => CLK, Q => n2390
                           , QN => n3672);
   REGISTERS_reg_38_7_inst : DFF_X1 port map( D => n1698, CK => CLK, Q => n3330
                           , QN => n_1158);
   REGISTERS_reg_38_6_inst : DFF_X1 port map( D => n1697, CK => CLK, Q => n3362
                           , QN => n_1159);
   REGISTERS_reg_38_5_inst : DFF_X1 port map( D => n1696, CK => CLK, Q => n3394
                           , QN => n_1160);
   REGISTERS_reg_38_4_inst : DFF_X1 port map( D => n1695, CK => CLK, Q => n3426
                           , QN => n_1161);
   REGISTERS_reg_38_3_inst : DFF_X1 port map( D => n1694, CK => CLK, Q => n3458
                           , QN => n_1162);
   REGISTERS_reg_38_2_inst : DFF_X1 port map( D => n1693, CK => CLK, Q => n3490
                           , QN => n_1163);
   REGISTERS_reg_38_1_inst : DFF_X1 port map( D => n1692, CK => CLK, Q => n3522
                           , QN => n_1164);
   REGISTERS_reg_38_0_inst : DFF_X1 port map( D => n1691, CK => CLK, Q => n3554
                           , QN => n_1165);
   REGISTERS_reg_39_7_inst : DFF_X1 port map( D => n1690, CK => CLK, Q => n3331
                           , QN => n_1166);
   REGISTERS_reg_39_6_inst : DFF_X1 port map( D => n1689, CK => CLK, Q => n3363
                           , QN => n_1167);
   REGISTERS_reg_39_5_inst : DFF_X1 port map( D => n1688, CK => CLK, Q => n3395
                           , QN => n_1168);
   REGISTERS_reg_39_4_inst : DFF_X1 port map( D => n1687, CK => CLK, Q => n3427
                           , QN => n_1169);
   REGISTERS_reg_39_3_inst : DFF_X1 port map( D => n1686, CK => CLK, Q => n3459
                           , QN => n_1170);
   REGISTERS_reg_39_2_inst : DFF_X1 port map( D => n1685, CK => CLK, Q => n3491
                           , QN => n_1171);
   REGISTERS_reg_39_1_inst : DFF_X1 port map( D => n1684, CK => CLK, Q => n3523
                           , QN => n_1172);
   REGISTERS_reg_39_0_inst : DFF_X1 port map( D => n1683, CK => CLK, Q => n3555
                           , QN => n_1173);
   REGISTERS_reg_40_7_inst : DFF_X1 port map( D => n1682, CK => CLK, Q => n3671
                           , QN => n2204);
   REGISTERS_reg_40_6_inst : DFF_X1 port map( D => n1681, CK => CLK, Q => n3670
                           , QN => n2215);
   REGISTERS_reg_40_5_inst : DFF_X1 port map( D => n1680, CK => CLK, Q => n3669
                           , QN => n2227);
   REGISTERS_reg_40_4_inst : DFF_X1 port map( D => n1679, CK => CLK, Q => n3668
                           , QN => n2239);
   REGISTERS_reg_40_3_inst : DFF_X1 port map( D => n1678, CK => CLK, Q => n3667
                           , QN => n2250);
   REGISTERS_reg_40_2_inst : DFF_X1 port map( D => n1677, CK => CLK, Q => n3666
                           , QN => n2261);
   REGISTERS_reg_40_1_inst : DFF_X1 port map( D => n1676, CK => CLK, Q => n3665
                           , QN => n2272);
   REGISTERS_reg_40_0_inst : DFF_X1 port map( D => n1675, CK => CLK, Q => n3664
                           , QN => n2283);
   REGISTERS_reg_41_7_inst : DFF_X1 port map( D => n1674, CK => CLK, Q => n2391
                           , QN => n3663);
   REGISTERS_reg_41_6_inst : DFF_X1 port map( D => n1673, CK => CLK, Q => n2392
                           , QN => n3662);
   REGISTERS_reg_41_5_inst : DFF_X1 port map( D => n1672, CK => CLK, Q => n2393
                           , QN => n3661);
   REGISTERS_reg_41_4_inst : DFF_X1 port map( D => n1671, CK => CLK, Q => n2394
                           , QN => n3660);
   REGISTERS_reg_41_3_inst : DFF_X1 port map( D => n1670, CK => CLK, Q => n2395
                           , QN => n3659);
   REGISTERS_reg_41_2_inst : DFF_X1 port map( D => n1669, CK => CLK, Q => n2396
                           , QN => n3658);
   REGISTERS_reg_41_1_inst : DFF_X1 port map( D => n1668, CK => CLK, Q => n2397
                           , QN => n3657);
   REGISTERS_reg_41_0_inst : DFF_X1 port map( D => n1667, CK => CLK, Q => n2398
                           , QN => n3656);
   REGISTERS_reg_42_7_inst : DFF_X1 port map( D => n1666, CK => CLK, Q => n3332
                           , QN => n_1174);
   REGISTERS_reg_42_6_inst : DFF_X1 port map( D => n1665, CK => CLK, Q => n3364
                           , QN => n_1175);
   REGISTERS_reg_42_5_inst : DFF_X1 port map( D => n1664, CK => CLK, Q => n3396
                           , QN => n_1176);
   REGISTERS_reg_42_4_inst : DFF_X1 port map( D => n1663, CK => CLK, Q => n3428
                           , QN => n_1177);
   REGISTERS_reg_42_3_inst : DFF_X1 port map( D => n1662, CK => CLK, Q => n3460
                           , QN => n_1178);
   REGISTERS_reg_42_2_inst : DFF_X1 port map( D => n1661, CK => CLK, Q => n3492
                           , QN => n_1179);
   REGISTERS_reg_42_1_inst : DFF_X1 port map( D => n1660, CK => CLK, Q => n3524
                           , QN => n_1180);
   REGISTERS_reg_42_0_inst : DFF_X1 port map( D => n1659, CK => CLK, Q => n3556
                           , QN => n_1181);
   REGISTERS_reg_43_7_inst : DFF_X1 port map( D => n1658, CK => CLK, Q => n3333
                           , QN => n_1182);
   REGISTERS_reg_43_6_inst : DFF_X1 port map( D => n1657, CK => CLK, Q => n3365
                           , QN => n_1183);
   REGISTERS_reg_43_5_inst : DFF_X1 port map( D => n1656, CK => CLK, Q => n3397
                           , QN => n_1184);
   REGISTERS_reg_43_4_inst : DFF_X1 port map( D => n1655, CK => CLK, Q => n3429
                           , QN => n_1185);
   REGISTERS_reg_43_3_inst : DFF_X1 port map( D => n1654, CK => CLK, Q => n3461
                           , QN => n_1186);
   REGISTERS_reg_43_2_inst : DFF_X1 port map( D => n1653, CK => CLK, Q => n3493
                           , QN => n_1187);
   REGISTERS_reg_43_1_inst : DFF_X1 port map( D => n1652, CK => CLK, Q => n3525
                           , QN => n_1188);
   REGISTERS_reg_43_0_inst : DFF_X1 port map( D => n1651, CK => CLK, Q => n3557
                           , QN => n_1189);
   REGISTERS_reg_44_7_inst : DFF_X1 port map( D => n1650, CK => CLK, Q => n3655
                           , QN => n2203);
   REGISTERS_reg_44_6_inst : DFF_X1 port map( D => n1649, CK => CLK, Q => n3654
                           , QN => n2214);
   REGISTERS_reg_44_5_inst : DFF_X1 port map( D => n1648, CK => CLK, Q => n3653
                           , QN => n2226);
   REGISTERS_reg_44_4_inst : DFF_X1 port map( D => n1647, CK => CLK, Q => n3652
                           , QN => n2238);
   REGISTERS_reg_44_3_inst : DFF_X1 port map( D => n1646, CK => CLK, Q => n3651
                           , QN => n2249);
   REGISTERS_reg_44_2_inst : DFF_X1 port map( D => n1645, CK => CLK, Q => n3650
                           , QN => n2260);
   REGISTERS_reg_44_1_inst : DFF_X1 port map( D => n1644, CK => CLK, Q => n3649
                           , QN => n2271);
   REGISTERS_reg_44_0_inst : DFF_X1 port map( D => n1643, CK => CLK, Q => n3648
                           , QN => n2282);
   REGISTERS_reg_45_7_inst : DFF_X1 port map( D => n1642, CK => CLK, Q => n2399
                           , QN => n3647);
   REGISTERS_reg_45_6_inst : DFF_X1 port map( D => n1641, CK => CLK, Q => n2400
                           , QN => n3646);
   REGISTERS_reg_45_5_inst : DFF_X1 port map( D => n1640, CK => CLK, Q => n2401
                           , QN => n3645);
   REGISTERS_reg_45_4_inst : DFF_X1 port map( D => n1639, CK => CLK, Q => n2402
                           , QN => n3644);
   REGISTERS_reg_45_3_inst : DFF_X1 port map( D => n1638, CK => CLK, Q => n2403
                           , QN => n3643);
   REGISTERS_reg_45_2_inst : DFF_X1 port map( D => n1637, CK => CLK, Q => n2404
                           , QN => n3642);
   REGISTERS_reg_45_1_inst : DFF_X1 port map( D => n1636, CK => CLK, Q => n2405
                           , QN => n3641);
   REGISTERS_reg_45_0_inst : DFF_X1 port map( D => n1635, CK => CLK, Q => n2406
                           , QN => n3640);
   REGISTERS_reg_46_7_inst : DFF_X1 port map( D => n1634, CK => CLK, Q => n3334
                           , QN => n_1190);
   REGISTERS_reg_46_6_inst : DFF_X1 port map( D => n1633, CK => CLK, Q => n3366
                           , QN => n_1191);
   REGISTERS_reg_46_5_inst : DFF_X1 port map( D => n1632, CK => CLK, Q => n3398
                           , QN => n_1192);
   REGISTERS_reg_46_4_inst : DFF_X1 port map( D => n1631, CK => CLK, Q => n3430
                           , QN => n_1193);
   REGISTERS_reg_46_3_inst : DFF_X1 port map( D => n1630, CK => CLK, Q => n3462
                           , QN => n_1194);
   REGISTERS_reg_46_2_inst : DFF_X1 port map( D => n1629, CK => CLK, Q => n3494
                           , QN => n_1195);
   REGISTERS_reg_46_1_inst : DFF_X1 port map( D => n1628, CK => CLK, Q => n3526
                           , QN => n_1196);
   REGISTERS_reg_46_0_inst : DFF_X1 port map( D => n1627, CK => CLK, Q => n3558
                           , QN => n_1197);
   REGISTERS_reg_47_7_inst : DFF_X1 port map( D => n1626, CK => CLK, Q => n3335
                           , QN => n_1198);
   REGISTERS_reg_47_6_inst : DFF_X1 port map( D => n1625, CK => CLK, Q => n3367
                           , QN => n_1199);
   REGISTERS_reg_47_5_inst : DFF_X1 port map( D => n1624, CK => CLK, Q => n3399
                           , QN => n_1200);
   REGISTERS_reg_47_4_inst : DFF_X1 port map( D => n1623, CK => CLK, Q => n3431
                           , QN => n_1201);
   REGISTERS_reg_47_3_inst : DFF_X1 port map( D => n1622, CK => CLK, Q => n3463
                           , QN => n_1202);
   REGISTERS_reg_47_2_inst : DFF_X1 port map( D => n1621, CK => CLK, Q => n3495
                           , QN => n_1203);
   REGISTERS_reg_47_1_inst : DFF_X1 port map( D => n1620, CK => CLK, Q => n3527
                           , QN => n_1204);
   REGISTERS_reg_47_0_inst : DFF_X1 port map( D => n1619, CK => CLK, Q => n3559
                           , QN => n_1205);
   REGISTERS_reg_48_7_inst : DFF_X1 port map( D => n1618, CK => CLK, Q => n3639
                           , QN => n2202);
   REGISTERS_reg_48_6_inst : DFF_X1 port map( D => n1617, CK => CLK, Q => n3638
                           , QN => n2213);
   REGISTERS_reg_48_5_inst : DFF_X1 port map( D => n1616, CK => CLK, Q => n3637
                           , QN => n2225);
   REGISTERS_reg_48_4_inst : DFF_X1 port map( D => n1615, CK => CLK, Q => n3636
                           , QN => n2237);
   REGISTERS_reg_48_3_inst : DFF_X1 port map( D => n1614, CK => CLK, Q => n3635
                           , QN => n2248);
   REGISTERS_reg_48_2_inst : DFF_X1 port map( D => n1613, CK => CLK, Q => n3634
                           , QN => n2259);
   REGISTERS_reg_48_1_inst : DFF_X1 port map( D => n1612, CK => CLK, Q => n3633
                           , QN => n2270);
   REGISTERS_reg_48_0_inst : DFF_X1 port map( D => n1611, CK => CLK, Q => n3632
                           , QN => n2281);
   REGISTERS_reg_49_7_inst : DFF_X1 port map( D => n1610, CK => CLK, Q => n2407
                           , QN => n3631);
   REGISTERS_reg_49_6_inst : DFF_X1 port map( D => n1609, CK => CLK, Q => n2408
                           , QN => n3630);
   REGISTERS_reg_49_5_inst : DFF_X1 port map( D => n1608, CK => CLK, Q => n2409
                           , QN => n3629);
   REGISTERS_reg_49_4_inst : DFF_X1 port map( D => n1607, CK => CLK, Q => n2410
                           , QN => n3628);
   REGISTERS_reg_49_3_inst : DFF_X1 port map( D => n1606, CK => CLK, Q => n2411
                           , QN => n3627);
   REGISTERS_reg_49_2_inst : DFF_X1 port map( D => n1605, CK => CLK, Q => n2412
                           , QN => n3626);
   REGISTERS_reg_49_1_inst : DFF_X1 port map( D => n1604, CK => CLK, Q => n2413
                           , QN => n3625);
   REGISTERS_reg_49_0_inst : DFF_X1 port map( D => n1603, CK => CLK, Q => n2414
                           , QN => n3624);
   REGISTERS_reg_50_7_inst : DFF_X1 port map( D => n1602, CK => CLK, Q => n3320
                           , QN => n_1206);
   REGISTERS_reg_50_6_inst : DFF_X1 port map( D => n1601, CK => CLK, Q => n3352
                           , QN => n_1207);
   REGISTERS_reg_50_5_inst : DFF_X1 port map( D => n1600, CK => CLK, Q => n3384
                           , QN => n_1208);
   REGISTERS_reg_50_4_inst : DFF_X1 port map( D => n1599, CK => CLK, Q => n3416
                           , QN => n_1209);
   REGISTERS_reg_50_3_inst : DFF_X1 port map( D => n1598, CK => CLK, Q => n3448
                           , QN => n_1210);
   REGISTERS_reg_50_2_inst : DFF_X1 port map( D => n1597, CK => CLK, Q => n3480
                           , QN => n_1211);
   REGISTERS_reg_50_1_inst : DFF_X1 port map( D => n1596, CK => CLK, Q => n3512
                           , QN => n_1212);
   REGISTERS_reg_50_0_inst : DFF_X1 port map( D => n1595, CK => CLK, Q => n3544
                           , QN => n_1213);
   REGISTERS_reg_51_7_inst : DFF_X1 port map( D => n1594, CK => CLK, Q => n3321
                           , QN => n_1214);
   REGISTERS_reg_51_6_inst : DFF_X1 port map( D => n1593, CK => CLK, Q => n3353
                           , QN => n_1215);
   REGISTERS_reg_51_5_inst : DFF_X1 port map( D => n1592, CK => CLK, Q => n3385
                           , QN => n_1216);
   REGISTERS_reg_51_4_inst : DFF_X1 port map( D => n1591, CK => CLK, Q => n3417
                           , QN => n_1217);
   REGISTERS_reg_51_3_inst : DFF_X1 port map( D => n1590, CK => CLK, Q => n3449
                           , QN => n_1218);
   REGISTERS_reg_51_2_inst : DFF_X1 port map( D => n1589, CK => CLK, Q => n3481
                           , QN => n_1219);
   REGISTERS_reg_51_1_inst : DFF_X1 port map( D => n1588, CK => CLK, Q => n3513
                           , QN => n_1220);
   REGISTERS_reg_51_0_inst : DFF_X1 port map( D => n1587, CK => CLK, Q => n3545
                           , QN => n_1221);
   REGISTERS_reg_52_7_inst : DFF_X1 port map( D => n1586, CK => CLK, Q => n3623
                           , QN => n2201);
   REGISTERS_reg_52_6_inst : DFF_X1 port map( D => n1585, CK => CLK, Q => n3622
                           , QN => n2212);
   REGISTERS_reg_52_5_inst : DFF_X1 port map( D => n1584, CK => CLK, Q => n3621
                           , QN => n2224);
   REGISTERS_reg_52_4_inst : DFF_X1 port map( D => n1583, CK => CLK, Q => n3620
                           , QN => n2236);
   REGISTERS_reg_52_3_inst : DFF_X1 port map( D => n1582, CK => CLK, Q => n3619
                           , QN => n2247);
   REGISTERS_reg_52_2_inst : DFF_X1 port map( D => n1581, CK => CLK, Q => n3618
                           , QN => n2258);
   REGISTERS_reg_52_1_inst : DFF_X1 port map( D => n1580, CK => CLK, Q => n3617
                           , QN => n2269);
   REGISTERS_reg_52_0_inst : DFF_X1 port map( D => n1579, CK => CLK, Q => n3616
                           , QN => n2280);
   REGISTERS_reg_53_7_inst : DFF_X1 port map( D => n1578, CK => CLK, Q => n2415
                           , QN => n3615);
   REGISTERS_reg_53_6_inst : DFF_X1 port map( D => n1577, CK => CLK, Q => n2416
                           , QN => n3614);
   REGISTERS_reg_53_5_inst : DFF_X1 port map( D => n1576, CK => CLK, Q => n2417
                           , QN => n3613);
   REGISTERS_reg_53_4_inst : DFF_X1 port map( D => n1575, CK => CLK, Q => n2418
                           , QN => n3612);
   REGISTERS_reg_53_3_inst : DFF_X1 port map( D => n1574, CK => CLK, Q => n2419
                           , QN => n3611);
   REGISTERS_reg_53_2_inst : DFF_X1 port map( D => n1573, CK => CLK, Q => n2420
                           , QN => n3610);
   REGISTERS_reg_53_1_inst : DFF_X1 port map( D => n1572, CK => CLK, Q => n2421
                           , QN => n3609);
   REGISTERS_reg_53_0_inst : DFF_X1 port map( D => n1571, CK => CLK, Q => n2422
                           , QN => n3608);
   REGISTERS_reg_54_7_inst : DFF_X1 port map( D => n1570, CK => CLK, Q => n3322
                           , QN => n_1222);
   REGISTERS_reg_54_6_inst : DFF_X1 port map( D => n1569, CK => CLK, Q => n3354
                           , QN => n_1223);
   REGISTERS_reg_54_5_inst : DFF_X1 port map( D => n1568, CK => CLK, Q => n3386
                           , QN => n_1224);
   REGISTERS_reg_54_4_inst : DFF_X1 port map( D => n1567, CK => CLK, Q => n3418
                           , QN => n_1225);
   REGISTERS_reg_54_3_inst : DFF_X1 port map( D => n1566, CK => CLK, Q => n3450
                           , QN => n_1226);
   REGISTERS_reg_54_2_inst : DFF_X1 port map( D => n1565, CK => CLK, Q => n3482
                           , QN => n_1227);
   REGISTERS_reg_54_1_inst : DFF_X1 port map( D => n1564, CK => CLK, Q => n3514
                           , QN => n_1228);
   REGISTERS_reg_54_0_inst : DFF_X1 port map( D => n1563, CK => CLK, Q => n3546
                           , QN => n_1229);
   REGISTERS_reg_55_7_inst : DFF_X1 port map( D => n1562, CK => CLK, Q => n3323
                           , QN => n_1230);
   REGISTERS_reg_55_6_inst : DFF_X1 port map( D => n1561, CK => CLK, Q => n3355
                           , QN => n_1231);
   REGISTERS_reg_55_5_inst : DFF_X1 port map( D => n1560, CK => CLK, Q => n3387
                           , QN => n_1232);
   REGISTERS_reg_55_4_inst : DFF_X1 port map( D => n1559, CK => CLK, Q => n3419
                           , QN => n_1233);
   REGISTERS_reg_55_3_inst : DFF_X1 port map( D => n1558, CK => CLK, Q => n3451
                           , QN => n_1234);
   REGISTERS_reg_55_2_inst : DFF_X1 port map( D => n1557, CK => CLK, Q => n3483
                           , QN => n_1235);
   REGISTERS_reg_55_1_inst : DFF_X1 port map( D => n1556, CK => CLK, Q => n3515
                           , QN => n_1236);
   REGISTERS_reg_55_0_inst : DFF_X1 port map( D => n1555, CK => CLK, Q => n3547
                           , QN => n_1237);
   REGISTERS_reg_56_7_inst : DFF_X1 port map( D => n1554, CK => CLK, Q => n3607
                           , QN => n2200);
   REGISTERS_reg_56_6_inst : DFF_X1 port map( D => n1553, CK => CLK, Q => n3606
                           , QN => n2211);
   REGISTERS_reg_56_5_inst : DFF_X1 port map( D => n1552, CK => CLK, Q => n3605
                           , QN => n2223);
   REGISTERS_reg_56_4_inst : DFF_X1 port map( D => n1551, CK => CLK, Q => n3604
                           , QN => n2235);
   REGISTERS_reg_56_3_inst : DFF_X1 port map( D => n1550, CK => CLK, Q => n3603
                           , QN => n2246);
   REGISTERS_reg_56_2_inst : DFF_X1 port map( D => n1549, CK => CLK, Q => n3602
                           , QN => n2257);
   REGISTERS_reg_56_1_inst : DFF_X1 port map( D => n1548, CK => CLK, Q => n3601
                           , QN => n2268);
   REGISTERS_reg_56_0_inst : DFF_X1 port map( D => n1547, CK => CLK, Q => n3600
                           , QN => n2279);
   REGISTERS_reg_57_7_inst : DFF_X1 port map( D => n1546, CK => CLK, Q => n2423
                           , QN => n3599);
   REGISTERS_reg_57_6_inst : DFF_X1 port map( D => n1545, CK => CLK, Q => n2424
                           , QN => n3598);
   REGISTERS_reg_57_5_inst : DFF_X1 port map( D => n1544, CK => CLK, Q => n2425
                           , QN => n3597);
   REGISTERS_reg_57_4_inst : DFF_X1 port map( D => n1543, CK => CLK, Q => n2426
                           , QN => n3596);
   REGISTERS_reg_57_3_inst : DFF_X1 port map( D => n1542, CK => CLK, Q => n2427
                           , QN => n3595);
   REGISTERS_reg_57_2_inst : DFF_X1 port map( D => n1541, CK => CLK, Q => n2428
                           , QN => n3594);
   REGISTERS_reg_57_1_inst : DFF_X1 port map( D => n1540, CK => CLK, Q => n2429
                           , QN => n3593);
   REGISTERS_reg_57_0_inst : DFF_X1 port map( D => n1539, CK => CLK, Q => n2430
                           , QN => n3592);
   REGISTERS_reg_58_7_inst : DFF_X1 port map( D => n1538, CK => CLK, Q => n3324
                           , QN => n_1238);
   REGISTERS_reg_58_6_inst : DFF_X1 port map( D => n1537, CK => CLK, Q => n3356
                           , QN => n_1239);
   REGISTERS_reg_58_5_inst : DFF_X1 port map( D => n1536, CK => CLK, Q => n3388
                           , QN => n_1240);
   REGISTERS_reg_58_4_inst : DFF_X1 port map( D => n1535, CK => CLK, Q => n3420
                           , QN => n_1241);
   REGISTERS_reg_58_3_inst : DFF_X1 port map( D => n1534, CK => CLK, Q => n3452
                           , QN => n_1242);
   REGISTERS_reg_58_2_inst : DFF_X1 port map( D => n1533, CK => CLK, Q => n3484
                           , QN => n_1243);
   REGISTERS_reg_58_1_inst : DFF_X1 port map( D => n1532, CK => CLK, Q => n3516
                           , QN => n_1244);
   REGISTERS_reg_58_0_inst : DFF_X1 port map( D => n1531, CK => CLK, Q => n3548
                           , QN => n_1245);
   REGISTERS_reg_59_7_inst : DFF_X1 port map( D => n1530, CK => CLK, Q => n3325
                           , QN => n_1246);
   REGISTERS_reg_59_6_inst : DFF_X1 port map( D => n1529, CK => CLK, Q => n3357
                           , QN => n_1247);
   REGISTERS_reg_59_5_inst : DFF_X1 port map( D => n1528, CK => CLK, Q => n3389
                           , QN => n_1248);
   REGISTERS_reg_59_4_inst : DFF_X1 port map( D => n1527, CK => CLK, Q => n3421
                           , QN => n_1249);
   REGISTERS_reg_59_3_inst : DFF_X1 port map( D => n1526, CK => CLK, Q => n3453
                           , QN => n_1250);
   REGISTERS_reg_59_2_inst : DFF_X1 port map( D => n1525, CK => CLK, Q => n3485
                           , QN => n_1251);
   REGISTERS_reg_59_1_inst : DFF_X1 port map( D => n1524, CK => CLK, Q => n3517
                           , QN => n_1252);
   REGISTERS_reg_59_0_inst : DFF_X1 port map( D => n1523, CK => CLK, Q => n3549
                           , QN => n_1253);
   REGISTERS_reg_60_7_inst : DFF_X1 port map( D => n1522, CK => CLK, Q => n3591
                           , QN => n2199);
   REGISTERS_reg_60_6_inst : DFF_X1 port map( D => n1521, CK => CLK, Q => n3590
                           , QN => n2210);
   REGISTERS_reg_60_5_inst : DFF_X1 port map( D => n1520, CK => CLK, Q => n3589
                           , QN => n2222);
   REGISTERS_reg_60_4_inst : DFF_X1 port map( D => n1519, CK => CLK, Q => n3588
                           , QN => n2234);
   REGISTERS_reg_60_3_inst : DFF_X1 port map( D => n1518, CK => CLK, Q => n3587
                           , QN => n2245);
   REGISTERS_reg_60_2_inst : DFF_X1 port map( D => n1517, CK => CLK, Q => n3586
                           , QN => n2256);
   REGISTERS_reg_60_1_inst : DFF_X1 port map( D => n1516, CK => CLK, Q => n3585
                           , QN => n2267);
   REGISTERS_reg_60_0_inst : DFF_X1 port map( D => n1515, CK => CLK, Q => n3584
                           , QN => n2278);
   REGISTERS_reg_61_7_inst : DFF_X1 port map( D => n1514, CK => CLK, Q => n2431
                           , QN => n3583);
   REGISTERS_reg_61_6_inst : DFF_X1 port map( D => n1513, CK => CLK, Q => n2432
                           , QN => n3582);
   REGISTERS_reg_61_5_inst : DFF_X1 port map( D => n1512, CK => CLK, Q => n2433
                           , QN => n3581);
   REGISTERS_reg_61_4_inst : DFF_X1 port map( D => n1511, CK => CLK, Q => n2434
                           , QN => n3580);
   REGISTERS_reg_61_3_inst : DFF_X1 port map( D => n1510, CK => CLK, Q => n2435
                           , QN => n3579);
   REGISTERS_reg_61_2_inst : DFF_X1 port map( D => n1509, CK => CLK, Q => n2436
                           , QN => n3578);
   REGISTERS_reg_61_1_inst : DFF_X1 port map( D => n1508, CK => CLK, Q => n2437
                           , QN => n3577);
   REGISTERS_reg_61_0_inst : DFF_X1 port map( D => n1507, CK => CLK, Q => n2438
                           , QN => n3576);
   REGISTERS_reg_62_7_inst : DFF_X1 port map( D => n1506, CK => CLK, Q => n3326
                           , QN => n_1254);
   REGISTERS_reg_62_6_inst : DFF_X1 port map( D => n1505, CK => CLK, Q => n3358
                           , QN => n_1255);
   REGISTERS_reg_62_5_inst : DFF_X1 port map( D => n1504, CK => CLK, Q => n3390
                           , QN => n_1256);
   REGISTERS_reg_62_4_inst : DFF_X1 port map( D => n1503, CK => CLK, Q => n3422
                           , QN => n_1257);
   REGISTERS_reg_62_3_inst : DFF_X1 port map( D => n1502, CK => CLK, Q => n3454
                           , QN => n_1258);
   REGISTERS_reg_62_2_inst : DFF_X1 port map( D => n1501, CK => CLK, Q => n3486
                           , QN => n_1259);
   REGISTERS_reg_62_1_inst : DFF_X1 port map( D => n1500, CK => CLK, Q => n3518
                           , QN => n_1260);
   REGISTERS_reg_62_0_inst : DFF_X1 port map( D => n1499, CK => CLK, Q => n3550
                           , QN => n_1261);
   REGISTERS_reg_63_7_inst : DFF_X1 port map( D => n1498, CK => CLK, Q => n3327
                           , QN => n_1262);
   REGISTERS_reg_63_6_inst : DFF_X1 port map( D => n1497, CK => CLK, Q => n3359
                           , QN => n_1263);
   REGISTERS_reg_63_5_inst : DFF_X1 port map( D => n1496, CK => CLK, Q => n3391
                           , QN => n_1264);
   REGISTERS_reg_63_4_inst : DFF_X1 port map( D => n1495, CK => CLK, Q => n3423
                           , QN => n_1265);
   REGISTERS_reg_63_3_inst : DFF_X1 port map( D => n1494, CK => CLK, Q => n3455
                           , QN => n_1266);
   REGISTERS_reg_63_2_inst : DFF_X1 port map( D => n1493, CK => CLK, Q => n3487
                           , QN => n_1267);
   REGISTERS_reg_63_1_inst : DFF_X1 port map( D => n1492, CK => CLK, Q => n3519
                           , QN => n_1268);
   REGISTERS_reg_63_0_inst : DFF_X1 port map( D => n1491, CK => CLK, Q => n3551
                           , QN => n_1269);
   OUT2_reg_7_inst : DFF_X1 port map( D => n1490, CK => CLK, Q => OUT2_7_port, 
                           QN => n_1270);
   OUT2_reg_6_inst : DFF_X1 port map( D => n1489, CK => CLK, Q => OUT2_6_port, 
                           QN => n_1271);
   OUT2_reg_5_inst : DFF_X1 port map( D => n1488, CK => CLK, Q => OUT2_5_port, 
                           QN => n_1272);
   OUT2_reg_4_inst : DFF_X1 port map( D => n1487, CK => CLK, Q => OUT2_4_port, 
                           QN => n_1273);
   OUT2_reg_3_inst : DFF_X1 port map( D => n1486, CK => CLK, Q => OUT2_3_port, 
                           QN => n_1274);
   OUT2_reg_2_inst : DFF_X1 port map( D => n1485, CK => CLK, Q => OUT2_2_port, 
                           QN => n_1275);
   OUT2_reg_1_inst : DFF_X1 port map( D => n1484, CK => CLK, Q => OUT2_1_port, 
                           QN => n_1276);
   OUT2_reg_0_inst : DFF_X1 port map( D => n1483, CK => CLK, Q => OUT2_0_port, 
                           QN => n_1277);
   OUT1_reg_7_inst : DFF_X1 port map( D => n1482, CK => CLK, Q => OUT1_7_port, 
                           QN => n_1278);
   OUT1_reg_6_inst : DFF_X1 port map( D => n1481, CK => CLK, Q => OUT1_6_port, 
                           QN => n_1279);
   OUT1_reg_5_inst : DFF_X1 port map( D => n1480, CK => CLK, Q => OUT1_5_port, 
                           QN => n_1280);
   OUT1_reg_4_inst : DFF_X1 port map( D => n1479, CK => CLK, Q => OUT1_4_port, 
                           QN => n_1281);
   OUT1_reg_3_inst : DFF_X1 port map( D => n1478, CK => CLK, Q => OUT1_3_port, 
                           QN => n_1282);
   OUT1_reg_2_inst : DFF_X1 port map( D => n1477, CK => CLK, Q => OUT1_2_port, 
                           QN => n_1283);
   OUT1_reg_1_inst : DFF_X1 port map( D => n1476, CK => CLK, Q => OUT1_1_port, 
                           QN => n_1284);
   OUT1_reg_0_inst : DFF_X1 port map( D => n1475, CK => CLK, Q => OUT1_0_port, 
                           QN => n_1285);
   U3 : AND2_X2 port map( A1 => DATAIN(7), A2 => n2450, ZN => n2439);
   U4 : AND2_X2 port map( A1 => DATAIN(6), A2 => n2450, ZN => n2441);
   U5 : AND2_X2 port map( A1 => DATAIN(5), A2 => n2450, ZN => n2442);
   U6 : AND2_X2 port map( A1 => DATAIN(4), A2 => n2450, ZN => n2443);
   U7 : AND2_X2 port map( A1 => DATAIN(3), A2 => n2450, ZN => n2444);
   U8 : AND2_X2 port map( A1 => DATAIN(2), A2 => n2450, ZN => n2445);
   U9 : AND2_X2 port map( A1 => DATAIN(1), A2 => n2450, ZN => n2446);
   U10 : AND2_X2 port map( A1 => DATAIN(0), A2 => n2450, ZN => n2447);
   U11 : INV_X4 port map( A => RESET, ZN => n2450);
   U12 : NOR2_X2 port map( A1 => n2927, A2 => ADD_RD2(1), ZN => n2873);
   U13 : NOR2_X2 port map( A1 => n3319, A2 => ADD_RD1(1), ZN => n3265);
   U14 : NOR2_X2 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(1), ZN => n2874);
   U15 : NOR2_X2 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(1), ZN => n3266);
   U16 : MUX2_X1 port map( A => n2306, B => n2439, S => n2440, Z => n2002);
   U17 : MUX2_X1 port map( A => n3830, B => n2441, S => n2440, Z => n2001);
   U18 : MUX2_X1 port map( A => n3829, B => n2442, S => n2440, Z => n2000);
   U19 : MUX2_X1 port map( A => n3828, B => n2443, S => n2440, Z => n1999);
   U20 : MUX2_X1 port map( A => n3827, B => n2444, S => n2440, Z => n1998);
   U21 : MUX2_X1 port map( A => n3826, B => n2445, S => n2440, Z => n1997);
   U22 : MUX2_X1 port map( A => n3825, B => n2446, S => n2440, Z => n1996);
   U23 : MUX2_X1 port map( A => n3824, B => n2447, S => n2440, Z => n1995);
   U24 : OAI21_X1 port map( B1 => n2448, B2 => n2449, A => n2450, ZN => n2440);
   U25 : MUX2_X1 port map( A => n3823, B => n2439, S => n2451, Z => n1994);
   U26 : MUX2_X1 port map( A => n2328, B => n2441, S => n2451, Z => n1993);
   U27 : MUX2_X1 port map( A => n2329, B => n2442, S => n2451, Z => n1992);
   U28 : MUX2_X1 port map( A => n2330, B => n2443, S => n2451, Z => n1991);
   U29 : MUX2_X1 port map( A => n2331, B => n2444, S => n2451, Z => n1990);
   U30 : MUX2_X1 port map( A => n2332, B => n2445, S => n2451, Z => n1989);
   U31 : MUX2_X1 port map( A => n2333, B => n2446, S => n2451, Z => n1988);
   U32 : MUX2_X1 port map( A => n2334, B => n2447, S => n2451, Z => n1987);
   U33 : OAI21_X1 port map( B1 => n2448, B2 => n2452, A => n2450, ZN => n2451);
   U34 : MUX2_X1 port map( A => n3344, B => n2439, S => n2453, Z => n1986);
   U35 : MUX2_X1 port map( A => n3376, B => n2441, S => n2453, Z => n1985);
   U36 : MUX2_X1 port map( A => n3408, B => n2442, S => n2453, Z => n1984);
   U37 : MUX2_X1 port map( A => n3440, B => n2443, S => n2453, Z => n1983);
   U38 : MUX2_X1 port map( A => n3472, B => n2444, S => n2453, Z => n1982);
   U39 : MUX2_X1 port map( A => n3504, B => n2445, S => n2453, Z => n1981);
   U40 : MUX2_X1 port map( A => n3536, B => n2446, S => n2453, Z => n1980);
   U41 : MUX2_X1 port map( A => n3568, B => n2447, S => n2453, Z => n1979);
   U42 : OAI21_X1 port map( B1 => n2448, B2 => n2454, A => n2450, ZN => n2453);
   U43 : MUX2_X1 port map( A => n3345, B => n2439, S => n2455, Z => n1978);
   U44 : MUX2_X1 port map( A => n3377, B => n2441, S => n2455, Z => n1977);
   U45 : MUX2_X1 port map( A => n3409, B => n2442, S => n2455, Z => n1976);
   U46 : MUX2_X1 port map( A => n3441, B => n2443, S => n2455, Z => n1975);
   U47 : MUX2_X1 port map( A => n3473, B => n2444, S => n2455, Z => n1974);
   U48 : MUX2_X1 port map( A => n3505, B => n2445, S => n2455, Z => n1973);
   U49 : MUX2_X1 port map( A => n3537, B => n2446, S => n2455, Z => n1972);
   U50 : MUX2_X1 port map( A => n3569, B => n2447, S => n2455, Z => n1971);
   U51 : OAI21_X1 port map( B1 => n2448, B2 => n2456, A => n2450, ZN => n2455);
   U52 : MUX2_X1 port map( A => n3815, B => n2439, S => n2457, Z => n1970);
   U53 : MUX2_X1 port map( A => n3814, B => n2441, S => n2457, Z => n1969);
   U54 : MUX2_X1 port map( A => n3813, B => n2442, S => n2457, Z => n1968);
   U55 : MUX2_X1 port map( A => n3812, B => n2443, S => n2457, Z => n1967);
   U56 : MUX2_X1 port map( A => n3811, B => n2444, S => n2457, Z => n1966);
   U57 : MUX2_X1 port map( A => n3810, B => n2445, S => n2457, Z => n1965);
   U58 : MUX2_X1 port map( A => n3809, B => n2446, S => n2457, Z => n1964);
   U59 : MUX2_X1 port map( A => n3808, B => n2447, S => n2457, Z => n1963);
   U60 : OAI21_X1 port map( B1 => n2448, B2 => n2458, A => n2450, ZN => n2457);
   U61 : MUX2_X1 port map( A => n3807, B => n2439, S => n2459, Z => n1962);
   U62 : MUX2_X1 port map( A => n3806, B => n2441, S => n2459, Z => n1961);
   U63 : MUX2_X1 port map( A => n3805, B => n2442, S => n2459, Z => n1960);
   U64 : MUX2_X1 port map( A => n3804, B => n2443, S => n2459, Z => n1959);
   U65 : MUX2_X1 port map( A => n3803, B => n2444, S => n2459, Z => n1958);
   U66 : MUX2_X1 port map( A => n3802, B => n2445, S => n2459, Z => n1957);
   U67 : MUX2_X1 port map( A => n3801, B => n2446, S => n2459, Z => n1956);
   U68 : MUX2_X1 port map( A => n3800, B => n2447, S => n2459, Z => n1955);
   U69 : OAI21_X1 port map( B1 => n2448, B2 => n2460, A => n2450, ZN => n2459);
   U70 : MUX2_X1 port map( A => n3346, B => n2439, S => n2461, Z => n1954);
   U71 : MUX2_X1 port map( A => n3378, B => n2441, S => n2461, Z => n1953);
   U72 : MUX2_X1 port map( A => n3410, B => n2442, S => n2461, Z => n1952);
   U73 : MUX2_X1 port map( A => n3442, B => n2443, S => n2461, Z => n1951);
   U74 : MUX2_X1 port map( A => n3474, B => n2444, S => n2461, Z => n1950);
   U75 : MUX2_X1 port map( A => n3506, B => n2445, S => n2461, Z => n1949);
   U76 : MUX2_X1 port map( A => n3538, B => n2446, S => n2461, Z => n1948);
   U77 : MUX2_X1 port map( A => n3570, B => n2447, S => n2461, Z => n1947);
   U78 : OAI21_X1 port map( B1 => n2448, B2 => n2462, A => n2450, ZN => n2461);
   U79 : MUX2_X1 port map( A => n3347, B => n2439, S => n2463, Z => n1946);
   U80 : MUX2_X1 port map( A => n3379, B => n2441, S => n2463, Z => n1945);
   U81 : MUX2_X1 port map( A => n3411, B => n2442, S => n2463, Z => n1944);
   U82 : MUX2_X1 port map( A => n3443, B => n2443, S => n2463, Z => n1943);
   U83 : MUX2_X1 port map( A => n3475, B => n2444, S => n2463, Z => n1942);
   U84 : MUX2_X1 port map( A => n3507, B => n2445, S => n2463, Z => n1941);
   U85 : MUX2_X1 port map( A => n3539, B => n2446, S => n2463, Z => n1940);
   U86 : MUX2_X1 port map( A => n3571, B => n2447, S => n2463, Z => n1939);
   U87 : OAI21_X1 port map( B1 => n2448, B2 => n2464, A => n2450, ZN => n2463);
   U88 : NAND3_X1 port map( A1 => n2465, A2 => n2466, A3 => n2467, ZN => n2448)
                           ;
   U89 : MUX2_X1 port map( A => n3799, B => n2439, S => n2468, Z => n1938);
   U90 : MUX2_X1 port map( A => n3798, B => n2441, S => n2468, Z => n1937);
   U91 : MUX2_X1 port map( A => n3797, B => n2442, S => n2468, Z => n1936);
   U92 : MUX2_X1 port map( A => n3796, B => n2443, S => n2468, Z => n1935);
   U93 : MUX2_X1 port map( A => n3795, B => n2444, S => n2468, Z => n1934);
   U94 : MUX2_X1 port map( A => n3794, B => n2445, S => n2468, Z => n1933);
   U95 : MUX2_X1 port map( A => n3793, B => n2446, S => n2468, Z => n1932);
   U96 : MUX2_X1 port map( A => n3792, B => n2447, S => n2468, Z => n1931);
   U97 : OAI21_X1 port map( B1 => n2449, B2 => n2469, A => n2450, ZN => n2468);
   U98 : MUX2_X1 port map( A => n3791, B => n2439, S => n2470, Z => n1930);
   U99 : MUX2_X1 port map( A => n3790, B => n2441, S => n2470, Z => n1929);
   U100 : MUX2_X1 port map( A => n3789, B => n2442, S => n2470, Z => n1928);
   U101 : MUX2_X1 port map( A => n3788, B => n2443, S => n2470, Z => n1927);
   U102 : MUX2_X1 port map( A => n3787, B => n2444, S => n2470, Z => n1926);
   U103 : MUX2_X1 port map( A => n3786, B => n2445, S => n2470, Z => n1925);
   U104 : MUX2_X1 port map( A => n3785, B => n2446, S => n2470, Z => n1924);
   U105 : MUX2_X1 port map( A => n3784, B => n2447, S => n2470, Z => n1923);
   U106 : OAI21_X1 port map( B1 => n2452, B2 => n2469, A => n2450, ZN => n2470)
                           ;
   U107 : MUX2_X1 port map( A => n3348, B => n2439, S => n2471, Z => n1922);
   U108 : MUX2_X1 port map( A => n3380, B => n2441, S => n2471, Z => n1921);
   U109 : MUX2_X1 port map( A => n3412, B => n2442, S => n2471, Z => n1920);
   U110 : MUX2_X1 port map( A => n3444, B => n2443, S => n2471, Z => n1919);
   U111 : MUX2_X1 port map( A => n3476, B => n2444, S => n2471, Z => n1918);
   U112 : MUX2_X1 port map( A => n3508, B => n2445, S => n2471, Z => n1917);
   U113 : MUX2_X1 port map( A => n3540, B => n2446, S => n2471, Z => n1916);
   U114 : MUX2_X1 port map( A => n3572, B => n2447, S => n2471, Z => n1915);
   U115 : OAI21_X1 port map( B1 => n2454, B2 => n2469, A => n2450, ZN => n2471)
                           ;
   U116 : MUX2_X1 port map( A => n3349, B => n2439, S => n2472, Z => n1914);
   U117 : MUX2_X1 port map( A => n3381, B => n2441, S => n2472, Z => n1913);
   U118 : MUX2_X1 port map( A => n3413, B => n2442, S => n2472, Z => n1912);
   U119 : MUX2_X1 port map( A => n3445, B => n2443, S => n2472, Z => n1911);
   U120 : MUX2_X1 port map( A => n3477, B => n2444, S => n2472, Z => n1910);
   U121 : MUX2_X1 port map( A => n3509, B => n2445, S => n2472, Z => n1909);
   U122 : MUX2_X1 port map( A => n3541, B => n2446, S => n2472, Z => n1908);
   U123 : MUX2_X1 port map( A => n3573, B => n2447, S => n2472, Z => n1907);
   U124 : OAI21_X1 port map( B1 => n2456, B2 => n2469, A => n2450, ZN => n2472)
                           ;
   U125 : MUX2_X1 port map( A => n3783, B => n2439, S => n2473, Z => n1906);
   U126 : MUX2_X1 port map( A => n3782, B => n2441, S => n2473, Z => n1905);
   U127 : MUX2_X1 port map( A => n3781, B => n2442, S => n2473, Z => n1904);
   U128 : MUX2_X1 port map( A => n2307, B => n2443, S => n2473, Z => n1903);
   U129 : MUX2_X1 port map( A => n2308, B => n2444, S => n2473, Z => n1902);
   U130 : MUX2_X1 port map( A => n2309, B => n2445, S => n2473, Z => n1901);
   U131 : MUX2_X1 port map( A => n2310, B => n2446, S => n2473, Z => n1900);
   U132 : MUX2_X1 port map( A => n2311, B => n2447, S => n2473, Z => n1899);
   U133 : OAI21_X1 port map( B1 => n2458, B2 => n2469, A => n2450, ZN => n2473)
                           ;
   U134 : MUX2_X1 port map( A => n2335, B => n2439, S => n2474, Z => n1898);
   U135 : MUX2_X1 port map( A => n2336, B => n2441, S => n2474, Z => n1897);
   U136 : MUX2_X1 port map( A => n2337, B => n2442, S => n2474, Z => n1896);
   U137 : MUX2_X1 port map( A => n2338, B => n2443, S => n2474, Z => n1895);
   U138 : MUX2_X1 port map( A => n2339, B => n2444, S => n2474, Z => n1894);
   U139 : MUX2_X1 port map( A => n2340, B => n2445, S => n2474, Z => n1893);
   U140 : MUX2_X1 port map( A => n2341, B => n2446, S => n2474, Z => n1892);
   U141 : MUX2_X1 port map( A => n2342, B => n2447, S => n2474, Z => n1891);
   U142 : OAI21_X1 port map( B1 => n2460, B2 => n2469, A => n2450, ZN => n2474)
                           ;
   U143 : MUX2_X1 port map( A => n3350, B => n2439, S => n2475, Z => n1890);
   U144 : MUX2_X1 port map( A => n3382, B => n2441, S => n2475, Z => n1889);
   U145 : MUX2_X1 port map( A => n3414, B => n2442, S => n2475, Z => n1888);
   U146 : MUX2_X1 port map( A => n3446, B => n2443, S => n2475, Z => n1887);
   U147 : MUX2_X1 port map( A => n3478, B => n2444, S => n2475, Z => n1886);
   U148 : MUX2_X1 port map( A => n3510, B => n2445, S => n2475, Z => n1885);
   U149 : MUX2_X1 port map( A => n3542, B => n2446, S => n2475, Z => n1884);
   U150 : MUX2_X1 port map( A => n3574, B => n2447, S => n2475, Z => n1883);
   U151 : OAI21_X1 port map( B1 => n2462, B2 => n2469, A => n2450, ZN => n2475)
                           ;
   U152 : MUX2_X1 port map( A => n3351, B => n2439, S => n2476, Z => n1882);
   U153 : MUX2_X1 port map( A => n3383, B => n2441, S => n2476, Z => n1881);
   U154 : MUX2_X1 port map( A => n3415, B => n2442, S => n2476, Z => n1880);
   U155 : MUX2_X1 port map( A => n3447, B => n2443, S => n2476, Z => n1879);
   U156 : MUX2_X1 port map( A => n3479, B => n2444, S => n2476, Z => n1878);
   U157 : MUX2_X1 port map( A => n3511, B => n2445, S => n2476, Z => n1877);
   U158 : MUX2_X1 port map( A => n3543, B => n2446, S => n2476, Z => n1876);
   U159 : MUX2_X1 port map( A => n3575, B => n2447, S => n2476, Z => n1875);
   U160 : OAI21_X1 port map( B1 => n2464, B2 => n2469, A => n2450, ZN => n2476)
                           ;
   U161 : NAND3_X1 port map( A1 => n2467, A2 => n2466, A3 => ADD_WR(3), ZN => 
                           n2469);
   U162 : MUX2_X1 port map( A => n2312, B => n2439, S => n2477, Z => n1874);
   U163 : MUX2_X1 port map( A => n2313, B => n2441, S => n2477, Z => n1873);
   U164 : MUX2_X1 port map( A => n2314, B => n2442, S => n2477, Z => n1872);
   U165 : MUX2_X1 port map( A => n2315, B => n2443, S => n2477, Z => n1871);
   U166 : MUX2_X1 port map( A => n2316, B => n2444, S => n2477, Z => n1870);
   U167 : MUX2_X1 port map( A => n2317, B => n2445, S => n2477, Z => n1869);
   U168 : MUX2_X1 port map( A => n2318, B => n2446, S => n2477, Z => n1868);
   U169 : MUX2_X1 port map( A => n2319, B => n2447, S => n2477, Z => n1867);
   U170 : OAI21_X1 port map( B1 => n2449, B2 => n2478, A => n2450, ZN => n2477)
                           ;
   U171 : MUX2_X1 port map( A => n2343, B => n2439, S => n2479, Z => n1866);
   U172 : MUX2_X1 port map( A => n2344, B => n2441, S => n2479, Z => n1865);
   U173 : MUX2_X1 port map( A => n2345, B => n2442, S => n2479, Z => n1864);
   U174 : MUX2_X1 port map( A => n2346, B => n2443, S => n2479, Z => n1863);
   U175 : MUX2_X1 port map( A => n2347, B => n2444, S => n2479, Z => n1862);
   U176 : MUX2_X1 port map( A => n2348, B => n2445, S => n2479, Z => n1861);
   U177 : MUX2_X1 port map( A => n2349, B => n2446, S => n2479, Z => n1860);
   U178 : MUX2_X1 port map( A => n2350, B => n2447, S => n2479, Z => n1859);
   U179 : OAI21_X1 port map( B1 => n2452, B2 => n2478, A => n2450, ZN => n2479)
                           ;
   U180 : MUX2_X1 port map( A => n3336, B => n2439, S => n2480, Z => n1858);
   U181 : MUX2_X1 port map( A => n3368, B => n2441, S => n2480, Z => n1857);
   U182 : MUX2_X1 port map( A => n3400, B => n2442, S => n2480, Z => n1856);
   U183 : MUX2_X1 port map( A => n3432, B => n2443, S => n2480, Z => n1855);
   U184 : MUX2_X1 port map( A => n3464, B => n2444, S => n2480, Z => n1854);
   U185 : MUX2_X1 port map( A => n3496, B => n2445, S => n2480, Z => n1853);
   U186 : MUX2_X1 port map( A => n3528, B => n2446, S => n2480, Z => n1852);
   U187 : MUX2_X1 port map( A => n3560, B => n2447, S => n2480, Z => n1851);
   U188 : OAI21_X1 port map( B1 => n2454, B2 => n2478, A => n2450, ZN => n2480)
                           ;
   U189 : MUX2_X1 port map( A => n3337, B => n2439, S => n2481, Z => n1850);
   U190 : MUX2_X1 port map( A => n3369, B => n2441, S => n2481, Z => n1849);
   U191 : MUX2_X1 port map( A => n3401, B => n2442, S => n2481, Z => n1848);
   U192 : MUX2_X1 port map( A => n3433, B => n2443, S => n2481, Z => n1847);
   U193 : MUX2_X1 port map( A => n3465, B => n2444, S => n2481, Z => n1846);
   U194 : MUX2_X1 port map( A => n3497, B => n2445, S => n2481, Z => n1845);
   U195 : MUX2_X1 port map( A => n3529, B => n2446, S => n2481, Z => n1844);
   U196 : MUX2_X1 port map( A => n3561, B => n2447, S => n2481, Z => n1843);
   U197 : OAI21_X1 port map( B1 => n2456, B2 => n2478, A => n2450, ZN => n2481)
                           ;
   U198 : MUX2_X1 port map( A => n2320, B => n2439, S => n2482, Z => n1842);
   U199 : MUX2_X1 port map( A => n2321, B => n2441, S => n2482, Z => n1841);
   U200 : MUX2_X1 port map( A => n2322, B => n2442, S => n2482, Z => n1840);
   U201 : MUX2_X1 port map( A => n2323, B => n2443, S => n2482, Z => n1839);
   U202 : MUX2_X1 port map( A => n2324, B => n2444, S => n2482, Z => n1838);
   U203 : MUX2_X1 port map( A => n2325, B => n2445, S => n2482, Z => n1837);
   U204 : MUX2_X1 port map( A => n2326, B => n2446, S => n2482, Z => n1836);
   U205 : MUX2_X1 port map( A => n2327, B => n2447, S => n2482, Z => n1835);
   U206 : OAI21_X1 port map( B1 => n2458, B2 => n2478, A => n2450, ZN => n2482)
                           ;
   U207 : MUX2_X1 port map( A => n2351, B => n2439, S => n2483, Z => n1834);
   U208 : MUX2_X1 port map( A => n2352, B => n2441, S => n2483, Z => n1833);
   U209 : MUX2_X1 port map( A => n2353, B => n2442, S => n2483, Z => n1832);
   U210 : MUX2_X1 port map( A => n2354, B => n2443, S => n2483, Z => n1831);
   U211 : MUX2_X1 port map( A => n2355, B => n2444, S => n2483, Z => n1830);
   U212 : MUX2_X1 port map( A => n2356, B => n2445, S => n2483, Z => n1829);
   U213 : MUX2_X1 port map( A => n2357, B => n2446, S => n2483, Z => n1828);
   U214 : MUX2_X1 port map( A => n2358, B => n2447, S => n2483, Z => n1827);
   U215 : OAI21_X1 port map( B1 => n2460, B2 => n2478, A => n2450, ZN => n2483)
                           ;
   U216 : MUX2_X1 port map( A => n3338, B => n2439, S => n2484, Z => n1826);
   U217 : MUX2_X1 port map( A => n3370, B => n2441, S => n2484, Z => n1825);
   U218 : MUX2_X1 port map( A => n3402, B => n2442, S => n2484, Z => n1824);
   U219 : MUX2_X1 port map( A => n3434, B => n2443, S => n2484, Z => n1823);
   U220 : MUX2_X1 port map( A => n3466, B => n2444, S => n2484, Z => n1822);
   U221 : MUX2_X1 port map( A => n3498, B => n2445, S => n2484, Z => n1821);
   U222 : MUX2_X1 port map( A => n3530, B => n2446, S => n2484, Z => n1820);
   U223 : MUX2_X1 port map( A => n3562, B => n2447, S => n2484, Z => n1819);
   U224 : OAI21_X1 port map( B1 => n2462, B2 => n2478, A => n2450, ZN => n2484)
                           ;
   U225 : MUX2_X1 port map( A => n3339, B => n2439, S => n2485, Z => n1818);
   U226 : MUX2_X1 port map( A => n3371, B => n2441, S => n2485, Z => n1817);
   U227 : MUX2_X1 port map( A => n3403, B => n2442, S => n2485, Z => n1816);
   U228 : MUX2_X1 port map( A => n3435, B => n2443, S => n2485, Z => n1815);
   U229 : MUX2_X1 port map( A => n3467, B => n2444, S => n2485, Z => n1814);
   U230 : MUX2_X1 port map( A => n3499, B => n2445, S => n2485, Z => n1813);
   U231 : MUX2_X1 port map( A => n3531, B => n2446, S => n2485, Z => n1812);
   U232 : MUX2_X1 port map( A => n3563, B => n2447, S => n2485, Z => n1811);
   U233 : OAI21_X1 port map( B1 => n2464, B2 => n2478, A => n2450, ZN => n2485)
                           ;
   U234 : NAND3_X1 port map( A1 => n2467, A2 => n2465, A3 => ADD_WR(4), ZN => 
                           n2478);
   U235 : MUX2_X1 port map( A => n3735, B => n2439, S => n2486, Z => n1810);
   U236 : MUX2_X1 port map( A => n3734, B => n2441, S => n2486, Z => n1809);
   U237 : MUX2_X1 port map( A => n3733, B => n2442, S => n2486, Z => n1808);
   U238 : MUX2_X1 port map( A => n3732, B => n2443, S => n2486, Z => n1807);
   U239 : MUX2_X1 port map( A => n3731, B => n2444, S => n2486, Z => n1806);
   U240 : MUX2_X1 port map( A => n3730, B => n2445, S => n2486, Z => n1805);
   U241 : MUX2_X1 port map( A => n3729, B => n2446, S => n2486, Z => n1804);
   U242 : MUX2_X1 port map( A => n3728, B => n2447, S => n2486, Z => n1803);
   U243 : OAI21_X1 port map( B1 => n2449, B2 => n2487, A => n2450, ZN => n2486)
                           ;
   U244 : MUX2_X1 port map( A => n2359, B => n2439, S => n2488, Z => n1802);
   U245 : MUX2_X1 port map( A => n2360, B => n2441, S => n2488, Z => n1801);
   U246 : MUX2_X1 port map( A => n2361, B => n2442, S => n2488, Z => n1800);
   U247 : MUX2_X1 port map( A => n2362, B => n2443, S => n2488, Z => n1799);
   U248 : MUX2_X1 port map( A => n2363, B => n2444, S => n2488, Z => n1798);
   U249 : MUX2_X1 port map( A => n2364, B => n2445, S => n2488, Z => n1797);
   U250 : MUX2_X1 port map( A => n2365, B => n2446, S => n2488, Z => n1796);
   U251 : MUX2_X1 port map( A => n2366, B => n2447, S => n2488, Z => n1795);
   U252 : OAI21_X1 port map( B1 => n2452, B2 => n2487, A => n2450, ZN => n2488)
                           ;
   U253 : MUX2_X1 port map( A => n3340, B => n2439, S => n2489, Z => n1794);
   U254 : MUX2_X1 port map( A => n3372, B => n2441, S => n2489, Z => n1793);
   U255 : MUX2_X1 port map( A => n3404, B => n2442, S => n2489, Z => n1792);
   U256 : MUX2_X1 port map( A => n3436, B => n2443, S => n2489, Z => n1791);
   U257 : MUX2_X1 port map( A => n3468, B => n2444, S => n2489, Z => n1790);
   U258 : MUX2_X1 port map( A => n3500, B => n2445, S => n2489, Z => n1789);
   U259 : MUX2_X1 port map( A => n3532, B => n2446, S => n2489, Z => n1788);
   U260 : MUX2_X1 port map( A => n3564, B => n2447, S => n2489, Z => n1787);
   U261 : OAI21_X1 port map( B1 => n2454, B2 => n2487, A => n2450, ZN => n2489)
                           ;
   U262 : MUX2_X1 port map( A => n3341, B => n2439, S => n2490, Z => n1786);
   U263 : MUX2_X1 port map( A => n3373, B => n2441, S => n2490, Z => n1785);
   U264 : MUX2_X1 port map( A => n3405, B => n2442, S => n2490, Z => n1784);
   U265 : MUX2_X1 port map( A => n3437, B => n2443, S => n2490, Z => n1783);
   U266 : MUX2_X1 port map( A => n3469, B => n2444, S => n2490, Z => n1782);
   U267 : MUX2_X1 port map( A => n3501, B => n2445, S => n2490, Z => n1781);
   U268 : MUX2_X1 port map( A => n3533, B => n2446, S => n2490, Z => n1780);
   U269 : MUX2_X1 port map( A => n3565, B => n2447, S => n2490, Z => n1779);
   U270 : OAI21_X1 port map( B1 => n2456, B2 => n2487, A => n2450, ZN => n2490)
                           ;
   U271 : MUX2_X1 port map( A => n3719, B => n2439, S => n2491, Z => n1778);
   U272 : MUX2_X1 port map( A => n3718, B => n2441, S => n2491, Z => n1777);
   U273 : MUX2_X1 port map( A => n3717, B => n2442, S => n2491, Z => n1776);
   U274 : MUX2_X1 port map( A => n3716, B => n2443, S => n2491, Z => n1775);
   U275 : MUX2_X1 port map( A => n3715, B => n2444, S => n2491, Z => n1774);
   U276 : MUX2_X1 port map( A => n3714, B => n2445, S => n2491, Z => n1773);
   U277 : MUX2_X1 port map( A => n3713, B => n2446, S => n2491, Z => n1772);
   U278 : MUX2_X1 port map( A => n3712, B => n2447, S => n2491, Z => n1771);
   U279 : OAI21_X1 port map( B1 => n2458, B2 => n2487, A => n2450, ZN => n2491)
                           ;
   U280 : MUX2_X1 port map( A => n2367, B => n2439, S => n2492, Z => n1770);
   U281 : MUX2_X1 port map( A => n2368, B => n2441, S => n2492, Z => n1769);
   U282 : MUX2_X1 port map( A => n2369, B => n2442, S => n2492, Z => n1768);
   U283 : MUX2_X1 port map( A => n2370, B => n2443, S => n2492, Z => n1767);
   U284 : MUX2_X1 port map( A => n2371, B => n2444, S => n2492, Z => n1766);
   U285 : MUX2_X1 port map( A => n2372, B => n2445, S => n2492, Z => n1765);
   U286 : MUX2_X1 port map( A => n2373, B => n2446, S => n2492, Z => n1764);
   U287 : MUX2_X1 port map( A => n2374, B => n2447, S => n2492, Z => n1763);
   U288 : OAI21_X1 port map( B1 => n2460, B2 => n2487, A => n2450, ZN => n2492)
                           ;
   U289 : MUX2_X1 port map( A => n3342, B => n2439, S => n2493, Z => n1762);
   U290 : MUX2_X1 port map( A => n3374, B => n2441, S => n2493, Z => n1761);
   U291 : MUX2_X1 port map( A => n3406, B => n2442, S => n2493, Z => n1760);
   U292 : MUX2_X1 port map( A => n3438, B => n2443, S => n2493, Z => n1759);
   U293 : MUX2_X1 port map( A => n3470, B => n2444, S => n2493, Z => n1758);
   U294 : MUX2_X1 port map( A => n3502, B => n2445, S => n2493, Z => n1757);
   U295 : MUX2_X1 port map( A => n3534, B => n2446, S => n2493, Z => n1756);
   U296 : MUX2_X1 port map( A => n3566, B => n2447, S => n2493, Z => n1755);
   U297 : OAI21_X1 port map( B1 => n2462, B2 => n2487, A => n2450, ZN => n2493)
                           ;
   U298 : MUX2_X1 port map( A => n3343, B => n2439, S => n2494, Z => n1754);
   U299 : MUX2_X1 port map( A => n3375, B => n2441, S => n2494, Z => n1753);
   U300 : MUX2_X1 port map( A => n3407, B => n2442, S => n2494, Z => n1752);
   U301 : MUX2_X1 port map( A => n3439, B => n2443, S => n2494, Z => n1751);
   U302 : MUX2_X1 port map( A => n3471, B => n2444, S => n2494, Z => n1750);
   U303 : MUX2_X1 port map( A => n3503, B => n2445, S => n2494, Z => n1749);
   U304 : MUX2_X1 port map( A => n3535, B => n2446, S => n2494, Z => n1748);
   U305 : MUX2_X1 port map( A => n3567, B => n2447, S => n2494, Z => n1747);
   U306 : OAI21_X1 port map( B1 => n2464, B2 => n2487, A => n2450, ZN => n2494)
                           ;
   U307 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => n2467, A3 => ADD_WR(4), ZN 
                           => n2487);
   U308 : AND3_X1 port map( A1 => ENABLE, A2 => n2495, A3 => WR, ZN => n2467);
   U309 : INV_X1 port map( A => ADD_WR(5), ZN => n2495);
   U310 : MUX2_X1 port map( A => n3703, B => n2439, S => n2496, Z => n1746);
   U311 : MUX2_X1 port map( A => n3702, B => n2441, S => n2496, Z => n1745);
   U312 : MUX2_X1 port map( A => n3701, B => n2442, S => n2496, Z => n1744);
   U313 : MUX2_X1 port map( A => n3700, B => n2443, S => n2496, Z => n1743);
   U314 : MUX2_X1 port map( A => n3699, B => n2444, S => n2496, Z => n1742);
   U315 : MUX2_X1 port map( A => n3698, B => n2445, S => n2496, Z => n1741);
   U316 : MUX2_X1 port map( A => n3697, B => n2446, S => n2496, Z => n1740);
   U317 : MUX2_X1 port map( A => n3696, B => n2447, S => n2496, Z => n1739);
   U318 : OAI21_X1 port map( B1 => n2449, B2 => n2497, A => n2450, ZN => n2496)
                           ;
   U319 : MUX2_X1 port map( A => n2375, B => n2439, S => n2498, Z => n1738);
   U320 : MUX2_X1 port map( A => n2376, B => n2441, S => n2498, Z => n1737);
   U321 : MUX2_X1 port map( A => n2377, B => n2442, S => n2498, Z => n1736);
   U322 : MUX2_X1 port map( A => n2378, B => n2443, S => n2498, Z => n1735);
   U323 : MUX2_X1 port map( A => n2379, B => n2444, S => n2498, Z => n1734);
   U324 : MUX2_X1 port map( A => n2380, B => n2445, S => n2498, Z => n1733);
   U325 : MUX2_X1 port map( A => n2381, B => n2446, S => n2498, Z => n1732);
   U326 : MUX2_X1 port map( A => n2382, B => n2447, S => n2498, Z => n1731);
   U327 : OAI21_X1 port map( B1 => n2452, B2 => n2497, A => n2450, ZN => n2498)
                           ;
   U328 : MUX2_X1 port map( A => n3328, B => n2439, S => n2499, Z => n1730);
   U329 : MUX2_X1 port map( A => n3360, B => n2441, S => n2499, Z => n1729);
   U330 : MUX2_X1 port map( A => n3392, B => n2442, S => n2499, Z => n1728);
   U331 : MUX2_X1 port map( A => n3424, B => n2443, S => n2499, Z => n1727);
   U332 : MUX2_X1 port map( A => n3456, B => n2444, S => n2499, Z => n1726);
   U333 : MUX2_X1 port map( A => n3488, B => n2445, S => n2499, Z => n1725);
   U334 : MUX2_X1 port map( A => n3520, B => n2446, S => n2499, Z => n1724);
   U335 : MUX2_X1 port map( A => n3552, B => n2447, S => n2499, Z => n1723);
   U336 : OAI21_X1 port map( B1 => n2454, B2 => n2497, A => n2450, ZN => n2499)
                           ;
   U337 : MUX2_X1 port map( A => n3329, B => n2439, S => n2500, Z => n1722);
   U338 : MUX2_X1 port map( A => n3361, B => n2441, S => n2500, Z => n1721);
   U339 : MUX2_X1 port map( A => n3393, B => n2442, S => n2500, Z => n1720);
   U340 : MUX2_X1 port map( A => n3425, B => n2443, S => n2500, Z => n1719);
   U341 : MUX2_X1 port map( A => n3457, B => n2444, S => n2500, Z => n1718);
   U342 : MUX2_X1 port map( A => n3489, B => n2445, S => n2500, Z => n1717);
   U343 : MUX2_X1 port map( A => n3521, B => n2446, S => n2500, Z => n1716);
   U344 : MUX2_X1 port map( A => n3553, B => n2447, S => n2500, Z => n1715);
   U345 : OAI21_X1 port map( B1 => n2456, B2 => n2497, A => n2450, ZN => n2500)
                           ;
   U346 : MUX2_X1 port map( A => n3687, B => n2439, S => n2501, Z => n1714);
   U347 : MUX2_X1 port map( A => n3686, B => n2441, S => n2501, Z => n1713);
   U348 : MUX2_X1 port map( A => n3685, B => n2442, S => n2501, Z => n1712);
   U349 : MUX2_X1 port map( A => n3684, B => n2443, S => n2501, Z => n1711);
   U350 : MUX2_X1 port map( A => n3683, B => n2444, S => n2501, Z => n1710);
   U351 : MUX2_X1 port map( A => n3682, B => n2445, S => n2501, Z => n1709);
   U352 : MUX2_X1 port map( A => n3681, B => n2446, S => n2501, Z => n1708);
   U353 : MUX2_X1 port map( A => n3680, B => n2447, S => n2501, Z => n1707);
   U354 : OAI21_X1 port map( B1 => n2458, B2 => n2497, A => n2450, ZN => n2501)
                           ;
   U355 : MUX2_X1 port map( A => n2383, B => n2439, S => n2502, Z => n1706);
   U356 : MUX2_X1 port map( A => n2384, B => n2441, S => n2502, Z => n1705);
   U357 : MUX2_X1 port map( A => n2385, B => n2442, S => n2502, Z => n1704);
   U358 : MUX2_X1 port map( A => n2386, B => n2443, S => n2502, Z => n1703);
   U359 : MUX2_X1 port map( A => n2387, B => n2444, S => n2502, Z => n1702);
   U360 : MUX2_X1 port map( A => n2388, B => n2445, S => n2502, Z => n1701);
   U361 : MUX2_X1 port map( A => n2389, B => n2446, S => n2502, Z => n1700);
   U362 : MUX2_X1 port map( A => n2390, B => n2447, S => n2502, Z => n1699);
   U363 : OAI21_X1 port map( B1 => n2460, B2 => n2497, A => n2450, ZN => n2502)
                           ;
   U364 : MUX2_X1 port map( A => n3330, B => n2439, S => n2503, Z => n1698);
   U365 : MUX2_X1 port map( A => n3362, B => n2441, S => n2503, Z => n1697);
   U366 : MUX2_X1 port map( A => n3394, B => n2442, S => n2503, Z => n1696);
   U367 : MUX2_X1 port map( A => n3426, B => n2443, S => n2503, Z => n1695);
   U368 : MUX2_X1 port map( A => n3458, B => n2444, S => n2503, Z => n1694);
   U369 : MUX2_X1 port map( A => n3490, B => n2445, S => n2503, Z => n1693);
   U370 : MUX2_X1 port map( A => n3522, B => n2446, S => n2503, Z => n1692);
   U371 : MUX2_X1 port map( A => n3554, B => n2447, S => n2503, Z => n1691);
   U372 : OAI21_X1 port map( B1 => n2462, B2 => n2497, A => n2450, ZN => n2503)
                           ;
   U373 : MUX2_X1 port map( A => n3331, B => n2439, S => n2504, Z => n1690);
   U374 : MUX2_X1 port map( A => n3363, B => n2441, S => n2504, Z => n1689);
   U375 : MUX2_X1 port map( A => n3395, B => n2442, S => n2504, Z => n1688);
   U376 : MUX2_X1 port map( A => n3427, B => n2443, S => n2504, Z => n1687);
   U377 : MUX2_X1 port map( A => n3459, B => n2444, S => n2504, Z => n1686);
   U378 : MUX2_X1 port map( A => n3491, B => n2445, S => n2504, Z => n1685);
   U379 : MUX2_X1 port map( A => n3523, B => n2446, S => n2504, Z => n1684);
   U380 : MUX2_X1 port map( A => n3555, B => n2447, S => n2504, Z => n1683);
   U381 : OAI21_X1 port map( B1 => n2464, B2 => n2497, A => n2450, ZN => n2504)
                           ;
   U382 : NAND3_X1 port map( A1 => n2465, A2 => n2466, A3 => n2505, ZN => n2497
                           );
   U383 : MUX2_X1 port map( A => n3671, B => n2439, S => n2506, Z => n1682);
   U384 : MUX2_X1 port map( A => n3670, B => n2441, S => n2506, Z => n1681);
   U385 : MUX2_X1 port map( A => n3669, B => n2442, S => n2506, Z => n1680);
   U386 : MUX2_X1 port map( A => n3668, B => n2443, S => n2506, Z => n1679);
   U387 : MUX2_X1 port map( A => n3667, B => n2444, S => n2506, Z => n1678);
   U388 : MUX2_X1 port map( A => n3666, B => n2445, S => n2506, Z => n1677);
   U389 : MUX2_X1 port map( A => n3665, B => n2446, S => n2506, Z => n1676);
   U390 : MUX2_X1 port map( A => n3664, B => n2447, S => n2506, Z => n1675);
   U391 : OAI21_X1 port map( B1 => n2449, B2 => n2507, A => n2450, ZN => n2506)
                           ;
   U392 : MUX2_X1 port map( A => n2391, B => n2439, S => n2508, Z => n1674);
   U393 : MUX2_X1 port map( A => n2392, B => n2441, S => n2508, Z => n1673);
   U394 : MUX2_X1 port map( A => n2393, B => n2442, S => n2508, Z => n1672);
   U395 : MUX2_X1 port map( A => n2394, B => n2443, S => n2508, Z => n1671);
   U396 : MUX2_X1 port map( A => n2395, B => n2444, S => n2508, Z => n1670);
   U397 : MUX2_X1 port map( A => n2396, B => n2445, S => n2508, Z => n1669);
   U398 : MUX2_X1 port map( A => n2397, B => n2446, S => n2508, Z => n1668);
   U399 : MUX2_X1 port map( A => n2398, B => n2447, S => n2508, Z => n1667);
   U400 : OAI21_X1 port map( B1 => n2452, B2 => n2507, A => n2450, ZN => n2508)
                           ;
   U401 : MUX2_X1 port map( A => n3332, B => n2439, S => n2509, Z => n1666);
   U402 : MUX2_X1 port map( A => n3364, B => n2441, S => n2509, Z => n1665);
   U403 : MUX2_X1 port map( A => n3396, B => n2442, S => n2509, Z => n1664);
   U404 : MUX2_X1 port map( A => n3428, B => n2443, S => n2509, Z => n1663);
   U405 : MUX2_X1 port map( A => n3460, B => n2444, S => n2509, Z => n1662);
   U406 : MUX2_X1 port map( A => n3492, B => n2445, S => n2509, Z => n1661);
   U407 : MUX2_X1 port map( A => n3524, B => n2446, S => n2509, Z => n1660);
   U408 : MUX2_X1 port map( A => n3556, B => n2447, S => n2509, Z => n1659);
   U409 : OAI21_X1 port map( B1 => n2454, B2 => n2507, A => n2450, ZN => n2509)
                           ;
   U410 : MUX2_X1 port map( A => n3333, B => n2439, S => n2510, Z => n1658);
   U411 : MUX2_X1 port map( A => n3365, B => n2441, S => n2510, Z => n1657);
   U412 : MUX2_X1 port map( A => n3397, B => n2442, S => n2510, Z => n1656);
   U413 : MUX2_X1 port map( A => n3429, B => n2443, S => n2510, Z => n1655);
   U414 : MUX2_X1 port map( A => n3461, B => n2444, S => n2510, Z => n1654);
   U415 : MUX2_X1 port map( A => n3493, B => n2445, S => n2510, Z => n1653);
   U416 : MUX2_X1 port map( A => n3525, B => n2446, S => n2510, Z => n1652);
   U417 : MUX2_X1 port map( A => n3557, B => n2447, S => n2510, Z => n1651);
   U418 : OAI21_X1 port map( B1 => n2456, B2 => n2507, A => n2450, ZN => n2510)
                           ;
   U419 : MUX2_X1 port map( A => n3655, B => n2439, S => n2511, Z => n1650);
   U420 : MUX2_X1 port map( A => n3654, B => n2441, S => n2511, Z => n1649);
   U421 : MUX2_X1 port map( A => n3653, B => n2442, S => n2511, Z => n1648);
   U422 : MUX2_X1 port map( A => n3652, B => n2443, S => n2511, Z => n1647);
   U423 : MUX2_X1 port map( A => n3651, B => n2444, S => n2511, Z => n1646);
   U424 : MUX2_X1 port map( A => n3650, B => n2445, S => n2511, Z => n1645);
   U425 : MUX2_X1 port map( A => n3649, B => n2446, S => n2511, Z => n1644);
   U426 : MUX2_X1 port map( A => n3648, B => n2447, S => n2511, Z => n1643);
   U427 : OAI21_X1 port map( B1 => n2458, B2 => n2507, A => n2450, ZN => n2511)
                           ;
   U428 : MUX2_X1 port map( A => n2399, B => n2439, S => n2512, Z => n1642);
   U429 : MUX2_X1 port map( A => n2400, B => n2441, S => n2512, Z => n1641);
   U430 : MUX2_X1 port map( A => n2401, B => n2442, S => n2512, Z => n1640);
   U431 : MUX2_X1 port map( A => n2402, B => n2443, S => n2512, Z => n1639);
   U432 : MUX2_X1 port map( A => n2403, B => n2444, S => n2512, Z => n1638);
   U433 : MUX2_X1 port map( A => n2404, B => n2445, S => n2512, Z => n1637);
   U434 : MUX2_X1 port map( A => n2405, B => n2446, S => n2512, Z => n1636);
   U435 : MUX2_X1 port map( A => n2406, B => n2447, S => n2512, Z => n1635);
   U436 : OAI21_X1 port map( B1 => n2460, B2 => n2507, A => n2450, ZN => n2512)
                           ;
   U437 : MUX2_X1 port map( A => n3334, B => n2439, S => n2513, Z => n1634);
   U438 : MUX2_X1 port map( A => n3366, B => n2441, S => n2513, Z => n1633);
   U439 : MUX2_X1 port map( A => n3398, B => n2442, S => n2513, Z => n1632);
   U440 : MUX2_X1 port map( A => n3430, B => n2443, S => n2513, Z => n1631);
   U441 : MUX2_X1 port map( A => n3462, B => n2444, S => n2513, Z => n1630);
   U442 : MUX2_X1 port map( A => n3494, B => n2445, S => n2513, Z => n1629);
   U443 : MUX2_X1 port map( A => n3526, B => n2446, S => n2513, Z => n1628);
   U444 : MUX2_X1 port map( A => n3558, B => n2447, S => n2513, Z => n1627);
   U445 : OAI21_X1 port map( B1 => n2462, B2 => n2507, A => n2450, ZN => n2513)
                           ;
   U446 : MUX2_X1 port map( A => n3335, B => n2439, S => n2514, Z => n1626);
   U447 : MUX2_X1 port map( A => n3367, B => n2441, S => n2514, Z => n1625);
   U448 : MUX2_X1 port map( A => n3399, B => n2442, S => n2514, Z => n1624);
   U449 : MUX2_X1 port map( A => n3431, B => n2443, S => n2514, Z => n1623);
   U450 : MUX2_X1 port map( A => n3463, B => n2444, S => n2514, Z => n1622);
   U451 : MUX2_X1 port map( A => n3495, B => n2445, S => n2514, Z => n1621);
   U452 : MUX2_X1 port map( A => n3527, B => n2446, S => n2514, Z => n1620);
   U453 : MUX2_X1 port map( A => n3559, B => n2447, S => n2514, Z => n1619);
   U454 : OAI21_X1 port map( B1 => n2464, B2 => n2507, A => n2450, ZN => n2514)
                           ;
   U455 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => n2466, A3 => n2505, ZN => 
                           n2507);
   U456 : INV_X1 port map( A => ADD_WR(4), ZN => n2466);
   U457 : MUX2_X1 port map( A => n3639, B => n2439, S => n2515, Z => n1618);
   U458 : MUX2_X1 port map( A => n3638, B => n2441, S => n2515, Z => n1617);
   U459 : MUX2_X1 port map( A => n3637, B => n2442, S => n2515, Z => n1616);
   U460 : MUX2_X1 port map( A => n3636, B => n2443, S => n2515, Z => n1615);
   U461 : MUX2_X1 port map( A => n3635, B => n2444, S => n2515, Z => n1614);
   U462 : MUX2_X1 port map( A => n3634, B => n2445, S => n2515, Z => n1613);
   U463 : MUX2_X1 port map( A => n3633, B => n2446, S => n2515, Z => n1612);
   U464 : MUX2_X1 port map( A => n3632, B => n2447, S => n2515, Z => n1611);
   U465 : OAI21_X1 port map( B1 => n2449, B2 => n2516, A => n2450, ZN => n2515)
                           ;
   U466 : MUX2_X1 port map( A => n2407, B => n2439, S => n2517, Z => n1610);
   U467 : MUX2_X1 port map( A => n2408, B => n2441, S => n2517, Z => n1609);
   U468 : MUX2_X1 port map( A => n2409, B => n2442, S => n2517, Z => n1608);
   U469 : MUX2_X1 port map( A => n2410, B => n2443, S => n2517, Z => n1607);
   U470 : MUX2_X1 port map( A => n2411, B => n2444, S => n2517, Z => n1606);
   U471 : MUX2_X1 port map( A => n2412, B => n2445, S => n2517, Z => n1605);
   U472 : MUX2_X1 port map( A => n2413, B => n2446, S => n2517, Z => n1604);
   U473 : MUX2_X1 port map( A => n2414, B => n2447, S => n2517, Z => n1603);
   U474 : OAI21_X1 port map( B1 => n2452, B2 => n2516, A => n2450, ZN => n2517)
                           ;
   U475 : MUX2_X1 port map( A => n3320, B => n2439, S => n2518, Z => n1602);
   U476 : MUX2_X1 port map( A => n3352, B => n2441, S => n2518, Z => n1601);
   U477 : MUX2_X1 port map( A => n3384, B => n2442, S => n2518, Z => n1600);
   U478 : MUX2_X1 port map( A => n3416, B => n2443, S => n2518, Z => n1599);
   U479 : MUX2_X1 port map( A => n3448, B => n2444, S => n2518, Z => n1598);
   U480 : MUX2_X1 port map( A => n3480, B => n2445, S => n2518, Z => n1597);
   U481 : MUX2_X1 port map( A => n3512, B => n2446, S => n2518, Z => n1596);
   U482 : MUX2_X1 port map( A => n3544, B => n2447, S => n2518, Z => n1595);
   U483 : OAI21_X1 port map( B1 => n2454, B2 => n2516, A => n2450, ZN => n2518)
                           ;
   U484 : MUX2_X1 port map( A => n3321, B => n2439, S => n2519, Z => n1594);
   U485 : MUX2_X1 port map( A => n3353, B => n2441, S => n2519, Z => n1593);
   U486 : MUX2_X1 port map( A => n3385, B => n2442, S => n2519, Z => n1592);
   U487 : MUX2_X1 port map( A => n3417, B => n2443, S => n2519, Z => n1591);
   U488 : MUX2_X1 port map( A => n3449, B => n2444, S => n2519, Z => n1590);
   U489 : MUX2_X1 port map( A => n3481, B => n2445, S => n2519, Z => n1589);
   U490 : MUX2_X1 port map( A => n3513, B => n2446, S => n2519, Z => n1588);
   U491 : MUX2_X1 port map( A => n3545, B => n2447, S => n2519, Z => n1587);
   U492 : OAI21_X1 port map( B1 => n2456, B2 => n2516, A => n2450, ZN => n2519)
                           ;
   U493 : MUX2_X1 port map( A => n3623, B => n2439, S => n2520, Z => n1586);
   U494 : MUX2_X1 port map( A => n3622, B => n2441, S => n2520, Z => n1585);
   U495 : MUX2_X1 port map( A => n3621, B => n2442, S => n2520, Z => n1584);
   U496 : MUX2_X1 port map( A => n3620, B => n2443, S => n2520, Z => n1583);
   U497 : MUX2_X1 port map( A => n3619, B => n2444, S => n2520, Z => n1582);
   U498 : MUX2_X1 port map( A => n3618, B => n2445, S => n2520, Z => n1581);
   U499 : MUX2_X1 port map( A => n3617, B => n2446, S => n2520, Z => n1580);
   U500 : MUX2_X1 port map( A => n3616, B => n2447, S => n2520, Z => n1579);
   U501 : OAI21_X1 port map( B1 => n2458, B2 => n2516, A => n2450, ZN => n2520)
                           ;
   U502 : MUX2_X1 port map( A => n2415, B => n2439, S => n2521, Z => n1578);
   U503 : MUX2_X1 port map( A => n2416, B => n2441, S => n2521, Z => n1577);
   U504 : MUX2_X1 port map( A => n2417, B => n2442, S => n2521, Z => n1576);
   U505 : MUX2_X1 port map( A => n2418, B => n2443, S => n2521, Z => n1575);
   U506 : MUX2_X1 port map( A => n2419, B => n2444, S => n2521, Z => n1574);
   U507 : MUX2_X1 port map( A => n2420, B => n2445, S => n2521, Z => n1573);
   U508 : MUX2_X1 port map( A => n2421, B => n2446, S => n2521, Z => n1572);
   U509 : MUX2_X1 port map( A => n2422, B => n2447, S => n2521, Z => n1571);
   U510 : OAI21_X1 port map( B1 => n2460, B2 => n2516, A => n2450, ZN => n2521)
                           ;
   U511 : MUX2_X1 port map( A => n3322, B => n2439, S => n2522, Z => n1570);
   U512 : MUX2_X1 port map( A => n3354, B => n2441, S => n2522, Z => n1569);
   U513 : MUX2_X1 port map( A => n3386, B => n2442, S => n2522, Z => n1568);
   U514 : MUX2_X1 port map( A => n3418, B => n2443, S => n2522, Z => n1567);
   U515 : MUX2_X1 port map( A => n3450, B => n2444, S => n2522, Z => n1566);
   U516 : MUX2_X1 port map( A => n3482, B => n2445, S => n2522, Z => n1565);
   U517 : MUX2_X1 port map( A => n3514, B => n2446, S => n2522, Z => n1564);
   U518 : MUX2_X1 port map( A => n3546, B => n2447, S => n2522, Z => n1563);
   U519 : OAI21_X1 port map( B1 => n2462, B2 => n2516, A => n2450, ZN => n2522)
                           ;
   U520 : MUX2_X1 port map( A => n3323, B => n2439, S => n2523, Z => n1562);
   U521 : MUX2_X1 port map( A => n3355, B => n2441, S => n2523, Z => n1561);
   U522 : MUX2_X1 port map( A => n3387, B => n2442, S => n2523, Z => n1560);
   U523 : MUX2_X1 port map( A => n3419, B => n2443, S => n2523, Z => n1559);
   U524 : MUX2_X1 port map( A => n3451, B => n2444, S => n2523, Z => n1558);
   U525 : MUX2_X1 port map( A => n3483, B => n2445, S => n2523, Z => n1557);
   U526 : MUX2_X1 port map( A => n3515, B => n2446, S => n2523, Z => n1556);
   U527 : MUX2_X1 port map( A => n3547, B => n2447, S => n2523, Z => n1555);
   U528 : OAI21_X1 port map( B1 => n2464, B2 => n2516, A => n2450, ZN => n2523)
                           ;
   U529 : NAND3_X1 port map( A1 => ADD_WR(4), A2 => n2465, A3 => n2505, ZN => 
                           n2516);
   U530 : INV_X1 port map( A => ADD_WR(3), ZN => n2465);
   U531 : MUX2_X1 port map( A => n3607, B => n2439, S => n2524, Z => n1554);
   U532 : MUX2_X1 port map( A => n3606, B => n2441, S => n2524, Z => n1553);
   U533 : MUX2_X1 port map( A => n3605, B => n2442, S => n2524, Z => n1552);
   U534 : MUX2_X1 port map( A => n3604, B => n2443, S => n2524, Z => n1551);
   U535 : MUX2_X1 port map( A => n3603, B => n2444, S => n2524, Z => n1550);
   U536 : MUX2_X1 port map( A => n3602, B => n2445, S => n2524, Z => n1549);
   U537 : MUX2_X1 port map( A => n3601, B => n2446, S => n2524, Z => n1548);
   U538 : MUX2_X1 port map( A => n3600, B => n2447, S => n2524, Z => n1547);
   U539 : OAI21_X1 port map( B1 => n2449, B2 => n2525, A => n2450, ZN => n2524)
                           ;
   U540 : NAND3_X1 port map( A1 => n2526, A2 => n2527, A3 => n2528, ZN => n2449
                           );
   U541 : MUX2_X1 port map( A => n2423, B => n2439, S => n2529, Z => n1546);
   U542 : MUX2_X1 port map( A => n2424, B => n2441, S => n2529, Z => n1545);
   U543 : MUX2_X1 port map( A => n2425, B => n2442, S => n2529, Z => n1544);
   U544 : MUX2_X1 port map( A => n2426, B => n2443, S => n2529, Z => n1543);
   U545 : MUX2_X1 port map( A => n2427, B => n2444, S => n2529, Z => n1542);
   U546 : MUX2_X1 port map( A => n2428, B => n2445, S => n2529, Z => n1541);
   U547 : MUX2_X1 port map( A => n2429, B => n2446, S => n2529, Z => n1540);
   U548 : MUX2_X1 port map( A => n2430, B => n2447, S => n2529, Z => n1539);
   U549 : OAI21_X1 port map( B1 => n2452, B2 => n2525, A => n2450, ZN => n2529)
                           ;
   U550 : NAND3_X1 port map( A1 => n2526, A2 => n2527, A3 => ADD_WR(0), ZN => 
                           n2452);
   U551 : MUX2_X1 port map( A => n3324, B => n2439, S => n2530, Z => n1538);
   U552 : MUX2_X1 port map( A => n3356, B => n2441, S => n2530, Z => n1537);
   U553 : MUX2_X1 port map( A => n3388, B => n2442, S => n2530, Z => n1536);
   U554 : MUX2_X1 port map( A => n3420, B => n2443, S => n2530, Z => n1535);
   U555 : MUX2_X1 port map( A => n3452, B => n2444, S => n2530, Z => n1534);
   U556 : MUX2_X1 port map( A => n3484, B => n2445, S => n2530, Z => n1533);
   U557 : MUX2_X1 port map( A => n3516, B => n2446, S => n2530, Z => n1532);
   U558 : MUX2_X1 port map( A => n3548, B => n2447, S => n2530, Z => n1531);
   U559 : OAI21_X1 port map( B1 => n2454, B2 => n2525, A => n2450, ZN => n2530)
                           ;
   U560 : NAND3_X1 port map( A1 => n2528, A2 => n2527, A3 => ADD_WR(1), ZN => 
                           n2454);
   U561 : MUX2_X1 port map( A => n3325, B => n2439, S => n2531, Z => n1530);
   U562 : MUX2_X1 port map( A => n3357, B => n2441, S => n2531, Z => n1529);
   U563 : MUX2_X1 port map( A => n3389, B => n2442, S => n2531, Z => n1528);
   U564 : MUX2_X1 port map( A => n3421, B => n2443, S => n2531, Z => n1527);
   U565 : MUX2_X1 port map( A => n3453, B => n2444, S => n2531, Z => n1526);
   U566 : MUX2_X1 port map( A => n3485, B => n2445, S => n2531, Z => n1525);
   U567 : MUX2_X1 port map( A => n3517, B => n2446, S => n2531, Z => n1524);
   U568 : MUX2_X1 port map( A => n3549, B => n2447, S => n2531, Z => n1523);
   U569 : OAI21_X1 port map( B1 => n2456, B2 => n2525, A => n2450, ZN => n2531)
                           ;
   U570 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n2527, A3 => ADD_WR(1), ZN 
                           => n2456);
   U571 : INV_X1 port map( A => ADD_WR(2), ZN => n2527);
   U572 : MUX2_X1 port map( A => n3591, B => n2439, S => n2532, Z => n1522);
   U573 : MUX2_X1 port map( A => n3590, B => n2441, S => n2532, Z => n1521);
   U574 : MUX2_X1 port map( A => n3589, B => n2442, S => n2532, Z => n1520);
   U575 : MUX2_X1 port map( A => n3588, B => n2443, S => n2532, Z => n1519);
   U576 : MUX2_X1 port map( A => n3587, B => n2444, S => n2532, Z => n1518);
   U577 : MUX2_X1 port map( A => n3586, B => n2445, S => n2532, Z => n1517);
   U578 : MUX2_X1 port map( A => n3585, B => n2446, S => n2532, Z => n1516);
   U579 : MUX2_X1 port map( A => n3584, B => n2447, S => n2532, Z => n1515);
   U580 : OAI21_X1 port map( B1 => n2458, B2 => n2525, A => n2450, ZN => n2532)
                           ;
   U581 : NAND3_X1 port map( A1 => n2528, A2 => n2526, A3 => ADD_WR(2), ZN => 
                           n2458);
   U582 : MUX2_X1 port map( A => n2431, B => n2439, S => n2533, Z => n1514);
   U583 : MUX2_X1 port map( A => n2432, B => n2441, S => n2533, Z => n1513);
   U584 : MUX2_X1 port map( A => n2433, B => n2442, S => n2533, Z => n1512);
   U585 : MUX2_X1 port map( A => n2434, B => n2443, S => n2533, Z => n1511);
   U586 : MUX2_X1 port map( A => n2435, B => n2444, S => n2533, Z => n1510);
   U587 : MUX2_X1 port map( A => n2436, B => n2445, S => n2533, Z => n1509);
   U588 : MUX2_X1 port map( A => n2437, B => n2446, S => n2533, Z => n1508);
   U589 : MUX2_X1 port map( A => n2438, B => n2447, S => n2533, Z => n1507);
   U590 : OAI21_X1 port map( B1 => n2460, B2 => n2525, A => n2450, ZN => n2533)
                           ;
   U591 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n2526, A3 => ADD_WR(2), ZN 
                           => n2460);
   U592 : INV_X1 port map( A => ADD_WR(1), ZN => n2526);
   U593 : MUX2_X1 port map( A => n3326, B => n2439, S => n2534, Z => n1506);
   U594 : MUX2_X1 port map( A => n3358, B => n2441, S => n2534, Z => n1505);
   U595 : MUX2_X1 port map( A => n3390, B => n2442, S => n2534, Z => n1504);
   U596 : MUX2_X1 port map( A => n3422, B => n2443, S => n2534, Z => n1503);
   U597 : MUX2_X1 port map( A => n3454, B => n2444, S => n2534, Z => n1502);
   U598 : MUX2_X1 port map( A => n3486, B => n2445, S => n2534, Z => n1501);
   U599 : MUX2_X1 port map( A => n3518, B => n2446, S => n2534, Z => n1500);
   U600 : MUX2_X1 port map( A => n3550, B => n2447, S => n2534, Z => n1499);
   U601 : OAI21_X1 port map( B1 => n2462, B2 => n2525, A => n2450, ZN => n2534)
                           ;
   U602 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => n2528, A3 => ADD_WR(2), ZN 
                           => n2462);
   U603 : INV_X1 port map( A => ADD_WR(0), ZN => n2528);
   U604 : MUX2_X1 port map( A => n3327, B => n2439, S => n2535, Z => n1498);
   U605 : MUX2_X1 port map( A => n3359, B => n2441, S => n2535, Z => n1497);
   U606 : MUX2_X1 port map( A => n3391, B => n2442, S => n2535, Z => n1496);
   U607 : MUX2_X1 port map( A => n3423, B => n2443, S => n2535, Z => n1495);
   U608 : MUX2_X1 port map( A => n3455, B => n2444, S => n2535, Z => n1494);
   U609 : MUX2_X1 port map( A => n3487, B => n2445, S => n2535, Z => n1493);
   U610 : MUX2_X1 port map( A => n3519, B => n2446, S => n2535, Z => n1492);
   U611 : MUX2_X1 port map( A => n3551, B => n2447, S => n2535, Z => n1491);
   U612 : OAI21_X1 port map( B1 => n2464, B2 => n2525, A => n2450, ZN => n2535)
                           ;
   U613 : NAND3_X1 port map( A1 => ADD_WR(4), A2 => ADD_WR(3), A3 => n2505, ZN 
                           => n2525);
   U614 : AND3_X1 port map( A1 => WR, A2 => ENABLE, A3 => ADD_WR(5), ZN => 
                           n2505);
   U615 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), A3 => ADD_WR(2),
                           ZN => n2464);
   U616 : MUX2_X1 port map( A => OUT2_7_port, B => n2536, S => n2537, Z => 
                           n1490);
   U617 : NAND4_X1 port map( A1 => n2538, A2 => n2539, A3 => n2540, A4 => n2541
                           , ZN => n2536);
   U618 : NOR4_X1 port map( A1 => n2542, A2 => n2543, A3 => n2544, A4 => n2545,
                           ZN => n2541);
   U619 : OAI221_X1 port map( B1 => n2199, B2 => n2546, C1 => n3583, C2 => 
                           n2547, A => n2548, ZN => n2545);
   U620 : AOI22_X1 port map( A1 => n2549, A2 => n3326, B1 => n2550, B2 => n3327
                           , ZN => n2548);
   U621 : OAI221_X1 port map( B1 => n2200, B2 => n2551, C1 => n3599, C2 => 
                           n2552, A => n2553, ZN => n2544);
   U622 : AOI22_X1 port map( A1 => n2554, A2 => n3324, B1 => n2555, B2 => n3325
                           , ZN => n2553);
   U623 : OAI221_X1 port map( B1 => n2201, B2 => n2556, C1 => n3615, C2 => 
                           n2557, A => n2558, ZN => n2543);
   U624 : AOI22_X1 port map( A1 => n2559, A2 => n3322, B1 => n2560, B2 => n3323
                           , ZN => n2558);
   U625 : OAI221_X1 port map( B1 => n2202, B2 => n2561, C1 => n3631, C2 => 
                           n2562, A => n2563, ZN => n2542);
   U626 : AOI22_X1 port map( A1 => n2564, A2 => n3320, B1 => n2565, B2 => n3321
                           , ZN => n2563);
   U627 : NOR4_X1 port map( A1 => n2566, A2 => n2567, A3 => n2568, A4 => n2569,
                           ZN => n2540);
   U628 : OAI221_X1 port map( B1 => n2203, B2 => n2570, C1 => n3647, C2 => 
                           n2571, A => n2572, ZN => n2569);
   U629 : AOI22_X1 port map( A1 => n2573, A2 => n3334, B1 => n2574, B2 => n3335
                           , ZN => n2572);
   U630 : OAI221_X1 port map( B1 => n2204, B2 => n2575, C1 => n3663, C2 => 
                           n2576, A => n2577, ZN => n2568);
   U631 : AOI22_X1 port map( A1 => n2578, A2 => n3332, B1 => n2579, B2 => n3333
                           , ZN => n2577);
   U632 : OAI221_X1 port map( B1 => n2205, B2 => n2580, C1 => n3679, C2 => 
                           n2581, A => n2582, ZN => n2567);
   U633 : AOI22_X1 port map( A1 => n2583, A2 => n3330, B1 => n2584, B2 => n3331
                           , ZN => n2582);
   U634 : OAI221_X1 port map( B1 => n2206, B2 => n2585, C1 => n3695, C2 => 
                           n2586, A => n2587, ZN => n2566);
   U635 : AOI22_X1 port map( A1 => n2588, A2 => n3328, B1 => n2589, B2 => n3329
                           , ZN => n2587);
   U636 : NOR4_X1 port map( A1 => n2590, A2 => n2591, A3 => n2592, A4 => n2593,
                           ZN => n2539);
   U637 : OAI221_X1 port map( B1 => n2207, B2 => n2594, C1 => n3711, C2 => 
                           n2595, A => n2596, ZN => n2593);
   U638 : AOI22_X1 port map( A1 => n2597, A2 => n3342, B1 => n2598, B2 => n3343
                           , ZN => n2596);
   U639 : OAI221_X1 port map( B1 => n2208, B2 => n2599, C1 => n3727, C2 => 
                           n2600, A => n2601, ZN => n2592);
   U640 : AOI22_X1 port map( A1 => n2602, A2 => n3340, B1 => n2603, B2 => n3341
                           , ZN => n2601);
   U641 : OAI221_X1 port map( B1 => n3751, B2 => n2604, C1 => n3743, C2 => 
                           n2605, A => n2606, ZN => n2591);
   U642 : AOI22_X1 port map( A1 => n2607, A2 => n3338, B1 => n2608, B2 => n3339
                           , ZN => n2606);
   U643 : OAI221_X1 port map( B1 => n3767, B2 => n2609, C1 => n3759, C2 => 
                           n2610, A => n2611, ZN => n2590);
   U644 : AOI22_X1 port map( A1 => n2612, A2 => n3336, B1 => n2613, B2 => n3337
                           , ZN => n2611);
   U645 : NOR4_X1 port map( A1 => n2614, A2 => n2615, A3 => n2616, A4 => n2617,
                           ZN => n2538);
   U646 : OAI221_X1 port map( B1 => n2209, B2 => n2618, C1 => n3775, C2 => 
                           n2619, A => n2620, ZN => n2617);
   U647 : AOI22_X1 port map( A1 => n2621, A2 => n3350, B1 => n2622, B2 => n3351
                           , ZN => n2620);
   U648 : OAI221_X1 port map( B1 => n2183, B2 => n2623, C1 => n2289, C2 => 
                           n2624, A => n2625, ZN => n2616);
   U649 : AOI22_X1 port map( A1 => n2626, A2 => n3348, B1 => n2627, B2 => n3349
                           , ZN => n2625);
   U650 : OAI221_X1 port map( B1 => n2184, B2 => n2628, C1 => n2290, C2 => 
                           n2629, A => n2630, ZN => n2615);
   U651 : AOI22_X1 port map( A1 => n2631, A2 => n3346, B1 => n2632, B2 => n3347
                           , ZN => n2630);
   U652 : OAI221_X1 port map( B1 => n3831, B2 => n2633, C1 => n2291, C2 => 
                           n2634, A => n2635, ZN => n2614);
   U653 : AOI22_X1 port map( A1 => n2636, A2 => n3344, B1 => n2637, B2 => n3345
                           , ZN => n2635);
   U654 : MUX2_X1 port map( A => OUT2_6_port, B => n2638, S => n2537, Z => 
                           n1489);
   U655 : NAND4_X1 port map( A1 => n2639, A2 => n2640, A3 => n2641, A4 => n2642
                           , ZN => n2638);
   U656 : NOR4_X1 port map( A1 => n2643, A2 => n2644, A3 => n2645, A4 => n2646,
                           ZN => n2642);
   U657 : OAI221_X1 port map( B1 => n2210, B2 => n2546, C1 => n3582, C2 => 
                           n2547, A => n2647, ZN => n2646);
   U658 : AOI22_X1 port map( A1 => n2549, A2 => n3358, B1 => n2550, B2 => n3359
                           , ZN => n2647);
   U659 : OAI221_X1 port map( B1 => n2211, B2 => n2551, C1 => n3598, C2 => 
                           n2552, A => n2648, ZN => n2645);
   U660 : AOI22_X1 port map( A1 => n2554, A2 => n3356, B1 => n2555, B2 => n3357
                           , ZN => n2648);
   U661 : OAI221_X1 port map( B1 => n2212, B2 => n2556, C1 => n3614, C2 => 
                           n2557, A => n2649, ZN => n2644);
   U662 : AOI22_X1 port map( A1 => n2559, A2 => n3354, B1 => n2560, B2 => n3355
                           , ZN => n2649);
   U663 : OAI221_X1 port map( B1 => n2213, B2 => n2561, C1 => n3630, C2 => 
                           n2562, A => n2650, ZN => n2643);
   U664 : AOI22_X1 port map( A1 => n2564, A2 => n3352, B1 => n2565, B2 => n3353
                           , ZN => n2650);
   U665 : NOR4_X1 port map( A1 => n2651, A2 => n2652, A3 => n2653, A4 => n2654,
                           ZN => n2641);
   U666 : OAI221_X1 port map( B1 => n2214, B2 => n2570, C1 => n3646, C2 => 
                           n2571, A => n2655, ZN => n2654);
   U667 : AOI22_X1 port map( A1 => n2573, A2 => n3366, B1 => n2574, B2 => n3367
                           , ZN => n2655);
   U668 : OAI221_X1 port map( B1 => n2215, B2 => n2575, C1 => n3662, C2 => 
                           n2576, A => n2656, ZN => n2653);
   U669 : AOI22_X1 port map( A1 => n2578, A2 => n3364, B1 => n2579, B2 => n3365
                           , ZN => n2656);
   U670 : OAI221_X1 port map( B1 => n2216, B2 => n2580, C1 => n3678, C2 => 
                           n2581, A => n2657, ZN => n2652);
   U671 : AOI22_X1 port map( A1 => n2583, A2 => n3362, B1 => n2584, B2 => n3363
                           , ZN => n2657);
   U672 : OAI221_X1 port map( B1 => n2217, B2 => n2585, C1 => n3694, C2 => 
                           n2586, A => n2658, ZN => n2651);
   U673 : AOI22_X1 port map( A1 => n2588, A2 => n3360, B1 => n2589, B2 => n3361
                           , ZN => n2658);
   U674 : NOR4_X1 port map( A1 => n2659, A2 => n2660, A3 => n2661, A4 => n2662,
                           ZN => n2640);
   U675 : OAI221_X1 port map( B1 => n2218, B2 => n2594, C1 => n3710, C2 => 
                           n2595, A => n2663, ZN => n2662);
   U676 : AOI22_X1 port map( A1 => n2597, A2 => n3374, B1 => n2598, B2 => n3375
                           , ZN => n2663);
   U677 : OAI221_X1 port map( B1 => n2219, B2 => n2599, C1 => n3726, C2 => 
                           n2600, A => n2664, ZN => n2661);
   U678 : AOI22_X1 port map( A1 => n2602, A2 => n3372, B1 => n2603, B2 => n3373
                           , ZN => n2664);
   U679 : OAI221_X1 port map( B1 => n3750, B2 => n2604, C1 => n3742, C2 => 
                           n2605, A => n2665, ZN => n2660);
   U680 : AOI22_X1 port map( A1 => n2607, A2 => n3370, B1 => n2608, B2 => n3371
                           , ZN => n2665);
   U681 : OAI221_X1 port map( B1 => n3766, B2 => n2609, C1 => n3758, C2 => 
                           n2610, A => n2666, ZN => n2659);
   U682 : AOI22_X1 port map( A1 => n2612, A2 => n3368, B1 => n2613, B2 => n3369
                           , ZN => n2666);
   U683 : NOR4_X1 port map( A1 => n2667, A2 => n2668, A3 => n2669, A4 => n2670,
                           ZN => n2639);
   U684 : OAI221_X1 port map( B1 => n2220, B2 => n2618, C1 => n3774, C2 => 
                           n2619, A => n2671, ZN => n2670);
   U685 : AOI22_X1 port map( A1 => n2621, A2 => n3382, B1 => n2622, B2 => n3383
                           , ZN => n2671);
   U686 : OAI221_X1 port map( B1 => n2185, B2 => n2623, C1 => n2292, C2 => 
                           n2624, A => n2672, ZN => n2669);
   U687 : AOI22_X1 port map( A1 => n2626, A2 => n3380, B1 => n2627, B2 => n3381
                           , ZN => n2672);
   U688 : OAI221_X1 port map( B1 => n2186, B2 => n2628, C1 => n2293, C2 => 
                           n2629, A => n2673, ZN => n2668);
   U689 : AOI22_X1 port map( A1 => n2631, A2 => n3378, B1 => n2632, B2 => n3379
                           , ZN => n2673);
   U690 : OAI221_X1 port map( B1 => n2221, B2 => n2633, C1 => n3822, C2 => 
                           n2634, A => n2674, ZN => n2667);
   U691 : AOI22_X1 port map( A1 => n2636, A2 => n3376, B1 => n2637, B2 => n3377
                           , ZN => n2674);
   U692 : MUX2_X1 port map( A => OUT2_5_port, B => n2675, S => n2537, Z => 
                           n1488);
   U693 : NAND4_X1 port map( A1 => n2676, A2 => n2677, A3 => n2678, A4 => n2679
                           , ZN => n2675);
   U694 : NOR4_X1 port map( A1 => n2680, A2 => n2681, A3 => n2682, A4 => n2683,
                           ZN => n2679);
   U695 : OAI221_X1 port map( B1 => n2222, B2 => n2546, C1 => n3581, C2 => 
                           n2547, A => n2684, ZN => n2683);
   U696 : AOI22_X1 port map( A1 => n2549, A2 => n3390, B1 => n2550, B2 => n3391
                           , ZN => n2684);
   U697 : OAI221_X1 port map( B1 => n2223, B2 => n2551, C1 => n3597, C2 => 
                           n2552, A => n2685, ZN => n2682);
   U698 : AOI22_X1 port map( A1 => n2554, A2 => n3388, B1 => n2555, B2 => n3389
                           , ZN => n2685);
   U699 : OAI221_X1 port map( B1 => n2224, B2 => n2556, C1 => n3613, C2 => 
                           n2557, A => n2686, ZN => n2681);
   U700 : AOI22_X1 port map( A1 => n2559, A2 => n3386, B1 => n2560, B2 => n3387
                           , ZN => n2686);
   U701 : OAI221_X1 port map( B1 => n2225, B2 => n2561, C1 => n3629, C2 => 
                           n2562, A => n2687, ZN => n2680);
   U702 : AOI22_X1 port map( A1 => n2564, A2 => n3384, B1 => n2565, B2 => n3385
                           , ZN => n2687);
   U703 : NOR4_X1 port map( A1 => n2688, A2 => n2689, A3 => n2690, A4 => n2691,
                           ZN => n2678);
   U704 : OAI221_X1 port map( B1 => n2226, B2 => n2570, C1 => n3645, C2 => 
                           n2571, A => n2692, ZN => n2691);
   U705 : AOI22_X1 port map( A1 => n2573, A2 => n3398, B1 => n2574, B2 => n3399
                           , ZN => n2692);
   U706 : OAI221_X1 port map( B1 => n2227, B2 => n2575, C1 => n3661, C2 => 
                           n2576, A => n2693, ZN => n2690);
   U707 : AOI22_X1 port map( A1 => n2578, A2 => n3396, B1 => n2579, B2 => n3397
                           , ZN => n2693);
   U708 : OAI221_X1 port map( B1 => n2228, B2 => n2580, C1 => n3677, C2 => 
                           n2581, A => n2694, ZN => n2689);
   U709 : AOI22_X1 port map( A1 => n2583, A2 => n3394, B1 => n2584, B2 => n3395
                           , ZN => n2694);
   U710 : OAI221_X1 port map( B1 => n2229, B2 => n2585, C1 => n3693, C2 => 
                           n2586, A => n2695, ZN => n2688);
   U711 : AOI22_X1 port map( A1 => n2588, A2 => n3392, B1 => n2589, B2 => n3393
                           , ZN => n2695);
   U712 : NOR4_X1 port map( A1 => n2696, A2 => n2697, A3 => n2698, A4 => n2699,
                           ZN => n2677);
   U713 : OAI221_X1 port map( B1 => n2230, B2 => n2594, C1 => n3709, C2 => 
                           n2595, A => n2700, ZN => n2699);
   U714 : AOI22_X1 port map( A1 => n2597, A2 => n3406, B1 => n2598, B2 => n3407
                           , ZN => n2700);
   U715 : OAI221_X1 port map( B1 => n2231, B2 => n2599, C1 => n3725, C2 => 
                           n2600, A => n2701, ZN => n2698);
   U716 : AOI22_X1 port map( A1 => n2602, A2 => n3404, B1 => n2603, B2 => n3405
                           , ZN => n2701);
   U717 : OAI221_X1 port map( B1 => n3749, B2 => n2604, C1 => n3741, C2 => 
                           n2605, A => n2702, ZN => n2697);
   U718 : AOI22_X1 port map( A1 => n2607, A2 => n3402, B1 => n2608, B2 => n3403
                           , ZN => n2702);
   U719 : OAI221_X1 port map( B1 => n3765, B2 => n2609, C1 => n3757, C2 => 
                           n2610, A => n2703, ZN => n2696);
   U720 : AOI22_X1 port map( A1 => n2612, A2 => n3400, B1 => n2613, B2 => n3401
                           , ZN => n2703);
   U721 : NOR4_X1 port map( A1 => n2704, A2 => n2705, A3 => n2706, A4 => n2707,
                           ZN => n2676);
   U722 : OAI221_X1 port map( B1 => n2232, B2 => n2618, C1 => n3773, C2 => 
                           n2619, A => n2708, ZN => n2707);
   U723 : AOI22_X1 port map( A1 => n2621, A2 => n3414, B1 => n2622, B2 => n3415
                           , ZN => n2708);
   U724 : OAI221_X1 port map( B1 => n2187, B2 => n2623, C1 => n2294, C2 => 
                           n2624, A => n2709, ZN => n2706);
   U725 : AOI22_X1 port map( A1 => n2626, A2 => n3412, B1 => n2627, B2 => n3413
                           , ZN => n2709);
   U726 : OAI221_X1 port map( B1 => n2188, B2 => n2628, C1 => n2295, C2 => 
                           n2629, A => n2710, ZN => n2705);
   U727 : AOI22_X1 port map( A1 => n2631, A2 => n3410, B1 => n2632, B2 => n3411
                           , ZN => n2710);
   U728 : OAI221_X1 port map( B1 => n2233, B2 => n2633, C1 => n3821, C2 => 
                           n2634, A => n2711, ZN => n2704);
   U729 : AOI22_X1 port map( A1 => n2636, A2 => n3408, B1 => n2637, B2 => n3409
                           , ZN => n2711);
   U730 : MUX2_X1 port map( A => OUT2_4_port, B => n2712, S => n2537, Z => 
                           n1487);
   U731 : NAND4_X1 port map( A1 => n2713, A2 => n2714, A3 => n2715, A4 => n2716
                           , ZN => n2712);
   U732 : NOR4_X1 port map( A1 => n2717, A2 => n2718, A3 => n2719, A4 => n2720,
                           ZN => n2716);
   U733 : OAI221_X1 port map( B1 => n2234, B2 => n2546, C1 => n3580, C2 => 
                           n2547, A => n2721, ZN => n2720);
   U734 : AOI22_X1 port map( A1 => n2549, A2 => n3422, B1 => n2550, B2 => n3423
                           , ZN => n2721);
   U735 : OAI221_X1 port map( B1 => n2235, B2 => n2551, C1 => n3596, C2 => 
                           n2552, A => n2722, ZN => n2719);
   U736 : AOI22_X1 port map( A1 => n2554, A2 => n3420, B1 => n2555, B2 => n3421
                           , ZN => n2722);
   U737 : OAI221_X1 port map( B1 => n2236, B2 => n2556, C1 => n3612, C2 => 
                           n2557, A => n2723, ZN => n2718);
   U738 : AOI22_X1 port map( A1 => n2559, A2 => n3418, B1 => n2560, B2 => n3419
                           , ZN => n2723);
   U739 : OAI221_X1 port map( B1 => n2237, B2 => n2561, C1 => n3628, C2 => 
                           n2562, A => n2724, ZN => n2717);
   U740 : AOI22_X1 port map( A1 => n2564, A2 => n3416, B1 => n2565, B2 => n3417
                           , ZN => n2724);
   U741 : NOR4_X1 port map( A1 => n2725, A2 => n2726, A3 => n2727, A4 => n2728,
                           ZN => n2715);
   U742 : OAI221_X1 port map( B1 => n2238, B2 => n2570, C1 => n3644, C2 => 
                           n2571, A => n2729, ZN => n2728);
   U743 : AOI22_X1 port map( A1 => n2573, A2 => n3430, B1 => n2574, B2 => n3431
                           , ZN => n2729);
   U744 : OAI221_X1 port map( B1 => n2239, B2 => n2575, C1 => n3660, C2 => 
                           n2576, A => n2730, ZN => n2727);
   U745 : AOI22_X1 port map( A1 => n2578, A2 => n3428, B1 => n2579, B2 => n3429
                           , ZN => n2730);
   U746 : OAI221_X1 port map( B1 => n2240, B2 => n2580, C1 => n3676, C2 => 
                           n2581, A => n2731, ZN => n2726);
   U747 : AOI22_X1 port map( A1 => n2583, A2 => n3426, B1 => n2584, B2 => n3427
                           , ZN => n2731);
   U748 : OAI221_X1 port map( B1 => n2241, B2 => n2585, C1 => n3692, C2 => 
                           n2586, A => n2732, ZN => n2725);
   U749 : AOI22_X1 port map( A1 => n2588, A2 => n3424, B1 => n2589, B2 => n3425
                           , ZN => n2732);
   U750 : NOR4_X1 port map( A1 => n2733, A2 => n2734, A3 => n2735, A4 => n2736,
                           ZN => n2714);
   U751 : OAI221_X1 port map( B1 => n2242, B2 => n2594, C1 => n3708, C2 => 
                           n2595, A => n2737, ZN => n2736);
   U752 : AOI22_X1 port map( A1 => n2597, A2 => n3438, B1 => n2598, B2 => n3439
                           , ZN => n2737);
   U753 : OAI221_X1 port map( B1 => n2243, B2 => n2599, C1 => n3724, C2 => 
                           n2600, A => n2738, ZN => n2735);
   U754 : AOI22_X1 port map( A1 => n2602, A2 => n3436, B1 => n2603, B2 => n3437
                           , ZN => n2738);
   U755 : OAI221_X1 port map( B1 => n3748, B2 => n2604, C1 => n3740, C2 => 
                           n2605, A => n2739, ZN => n2734);
   U756 : AOI22_X1 port map( A1 => n2607, A2 => n3434, B1 => n2608, B2 => n3435
                           , ZN => n2739);
   U757 : OAI221_X1 port map( B1 => n3764, B2 => n2609, C1 => n3756, C2 => 
                           n2610, A => n2740, ZN => n2733);
   U758 : AOI22_X1 port map( A1 => n2612, A2 => n3432, B1 => n2613, B2 => n3433
                           , ZN => n2740);
   U759 : NOR4_X1 port map( A1 => n2741, A2 => n2742, A3 => n2743, A4 => n2744,
                           ZN => n2713);
   U760 : OAI221_X1 port map( B1 => n3780, B2 => n2618, C1 => n3772, C2 => 
                           n2619, A => n2745, ZN => n2744);
   U761 : AOI22_X1 port map( A1 => n2621, A2 => n3446, B1 => n2622, B2 => n3447
                           , ZN => n2745);
   U762 : OAI221_X1 port map( B1 => n2189, B2 => n2623, C1 => n2296, C2 => 
                           n2624, A => n2746, ZN => n2743);
   U763 : AOI22_X1 port map( A1 => n2626, A2 => n3444, B1 => n2627, B2 => n3445
                           , ZN => n2746);
   U764 : OAI221_X1 port map( B1 => n2190, B2 => n2628, C1 => n2297, C2 => 
                           n2629, A => n2747, ZN => n2742);
   U765 : AOI22_X1 port map( A1 => n2631, A2 => n3442, B1 => n2632, B2 => n3443
                           , ZN => n2747);
   U766 : OAI221_X1 port map( B1 => n2244, B2 => n2633, C1 => n3820, C2 => 
                           n2634, A => n2748, ZN => n2741);
   U767 : AOI22_X1 port map( A1 => n2636, A2 => n3440, B1 => n2637, B2 => n3441
                           , ZN => n2748);
   U768 : MUX2_X1 port map( A => OUT2_3_port, B => n2749, S => n2537, Z => 
                           n1486);
   U769 : NAND4_X1 port map( A1 => n2750, A2 => n2751, A3 => n2752, A4 => n2753
                           , ZN => n2749);
   U770 : NOR4_X1 port map( A1 => n2754, A2 => n2755, A3 => n2756, A4 => n2757,
                           ZN => n2753);
   U771 : OAI221_X1 port map( B1 => n2245, B2 => n2546, C1 => n3579, C2 => 
                           n2547, A => n2758, ZN => n2757);
   U772 : AOI22_X1 port map( A1 => n2549, A2 => n3454, B1 => n2550, B2 => n3455
                           , ZN => n2758);
   U773 : OAI221_X1 port map( B1 => n2246, B2 => n2551, C1 => n3595, C2 => 
                           n2552, A => n2759, ZN => n2756);
   U774 : AOI22_X1 port map( A1 => n2554, A2 => n3452, B1 => n2555, B2 => n3453
                           , ZN => n2759);
   U775 : OAI221_X1 port map( B1 => n2247, B2 => n2556, C1 => n3611, C2 => 
                           n2557, A => n2760, ZN => n2755);
   U776 : AOI22_X1 port map( A1 => n2559, A2 => n3450, B1 => n2560, B2 => n3451
                           , ZN => n2760);
   U777 : OAI221_X1 port map( B1 => n2248, B2 => n2561, C1 => n3627, C2 => 
                           n2562, A => n2761, ZN => n2754);
   U778 : AOI22_X1 port map( A1 => n2564, A2 => n3448, B1 => n2565, B2 => n3449
                           , ZN => n2761);
   U779 : NOR4_X1 port map( A1 => n2762, A2 => n2763, A3 => n2764, A4 => n2765,
                           ZN => n2752);
   U780 : OAI221_X1 port map( B1 => n2249, B2 => n2570, C1 => n3643, C2 => 
                           n2571, A => n2766, ZN => n2765);
   U781 : AOI22_X1 port map( A1 => n2573, A2 => n3462, B1 => n2574, B2 => n3463
                           , ZN => n2766);
   U782 : OAI221_X1 port map( B1 => n2250, B2 => n2575, C1 => n3659, C2 => 
                           n2576, A => n2767, ZN => n2764);
   U783 : AOI22_X1 port map( A1 => n2578, A2 => n3460, B1 => n2579, B2 => n3461
                           , ZN => n2767);
   U784 : OAI221_X1 port map( B1 => n2251, B2 => n2580, C1 => n3675, C2 => 
                           n2581, A => n2768, ZN => n2763);
   U785 : AOI22_X1 port map( A1 => n2583, A2 => n3458, B1 => n2584, B2 => n3459
                           , ZN => n2768);
   U786 : OAI221_X1 port map( B1 => n2252, B2 => n2585, C1 => n3691, C2 => 
                           n2586, A => n2769, ZN => n2762);
   U787 : AOI22_X1 port map( A1 => n2588, A2 => n3456, B1 => n2589, B2 => n3457
                           , ZN => n2769);
   U788 : NOR4_X1 port map( A1 => n2770, A2 => n2771, A3 => n2772, A4 => n2773,
                           ZN => n2751);
   U789 : OAI221_X1 port map( B1 => n2253, B2 => n2594, C1 => n3707, C2 => 
                           n2595, A => n2774, ZN => n2773);
   U790 : AOI22_X1 port map( A1 => n2597, A2 => n3470, B1 => n2598, B2 => n3471
                           , ZN => n2774);
   U791 : OAI221_X1 port map( B1 => n2254, B2 => n2599, C1 => n3723, C2 => 
                           n2600, A => n2775, ZN => n2772);
   U792 : AOI22_X1 port map( A1 => n2602, A2 => n3468, B1 => n2603, B2 => n3469
                           , ZN => n2775);
   U793 : OAI221_X1 port map( B1 => n3747, B2 => n2604, C1 => n3739, C2 => 
                           n2605, A => n2776, ZN => n2771);
   U794 : AOI22_X1 port map( A1 => n2607, A2 => n3466, B1 => n2608, B2 => n3467
                           , ZN => n2776);
   U795 : OAI221_X1 port map( B1 => n3763, B2 => n2609, C1 => n3755, C2 => 
                           n2610, A => n2777, ZN => n2770);
   U796 : AOI22_X1 port map( A1 => n2612, A2 => n3464, B1 => n2613, B2 => n3465
                           , ZN => n2777);
   U797 : NOR4_X1 port map( A1 => n2778, A2 => n2779, A3 => n2780, A4 => n2781,
                           ZN => n2750);
   U798 : OAI221_X1 port map( B1 => n3779, B2 => n2618, C1 => n3771, C2 => 
                           n2619, A => n2782, ZN => n2781);
   U799 : AOI22_X1 port map( A1 => n2621, A2 => n3478, B1 => n2622, B2 => n3479
                           , ZN => n2782);
   U800 : OAI221_X1 port map( B1 => n2191, B2 => n2623, C1 => n2298, C2 => 
                           n2624, A => n2783, ZN => n2780);
   U801 : AOI22_X1 port map( A1 => n2626, A2 => n3476, B1 => n2627, B2 => n3477
                           , ZN => n2783);
   U802 : OAI221_X1 port map( B1 => n2192, B2 => n2628, C1 => n2299, C2 => 
                           n2629, A => n2784, ZN => n2779);
   U803 : AOI22_X1 port map( A1 => n2631, A2 => n3474, B1 => n2632, B2 => n3475
                           , ZN => n2784);
   U804 : OAI221_X1 port map( B1 => n2255, B2 => n2633, C1 => n3819, C2 => 
                           n2634, A => n2785, ZN => n2778);
   U805 : AOI22_X1 port map( A1 => n2636, A2 => n3472, B1 => n2637, B2 => n3473
                           , ZN => n2785);
   U806 : MUX2_X1 port map( A => OUT2_2_port, B => n2786, S => n2537, Z => 
                           n1485);
   U807 : NAND4_X1 port map( A1 => n2787, A2 => n2788, A3 => n2789, A4 => n2790
                           , ZN => n2786);
   U808 : NOR4_X1 port map( A1 => n2791, A2 => n2792, A3 => n2793, A4 => n2794,
                           ZN => n2790);
   U809 : OAI221_X1 port map( B1 => n2256, B2 => n2546, C1 => n3578, C2 => 
                           n2547, A => n2795, ZN => n2794);
   U810 : AOI22_X1 port map( A1 => n2549, A2 => n3486, B1 => n2550, B2 => n3487
                           , ZN => n2795);
   U811 : OAI221_X1 port map( B1 => n2257, B2 => n2551, C1 => n3594, C2 => 
                           n2552, A => n2796, ZN => n2793);
   U812 : AOI22_X1 port map( A1 => n2554, A2 => n3484, B1 => n2555, B2 => n3485
                           , ZN => n2796);
   U813 : OAI221_X1 port map( B1 => n2258, B2 => n2556, C1 => n3610, C2 => 
                           n2557, A => n2797, ZN => n2792);
   U814 : AOI22_X1 port map( A1 => n2559, A2 => n3482, B1 => n2560, B2 => n3483
                           , ZN => n2797);
   U815 : OAI221_X1 port map( B1 => n2259, B2 => n2561, C1 => n3626, C2 => 
                           n2562, A => n2798, ZN => n2791);
   U816 : AOI22_X1 port map( A1 => n2564, A2 => n3480, B1 => n2565, B2 => n3481
                           , ZN => n2798);
   U817 : NOR4_X1 port map( A1 => n2799, A2 => n2800, A3 => n2801, A4 => n2802,
                           ZN => n2789);
   U818 : OAI221_X1 port map( B1 => n2260, B2 => n2570, C1 => n3642, C2 => 
                           n2571, A => n2803, ZN => n2802);
   U819 : AOI22_X1 port map( A1 => n2573, A2 => n3494, B1 => n2574, B2 => n3495
                           , ZN => n2803);
   U820 : OAI221_X1 port map( B1 => n2261, B2 => n2575, C1 => n3658, C2 => 
                           n2576, A => n2804, ZN => n2801);
   U821 : AOI22_X1 port map( A1 => n2578, A2 => n3492, B1 => n2579, B2 => n3493
                           , ZN => n2804);
   U822 : OAI221_X1 port map( B1 => n2262, B2 => n2580, C1 => n3674, C2 => 
                           n2581, A => n2805, ZN => n2800);
   U823 : AOI22_X1 port map( A1 => n2583, A2 => n3490, B1 => n2584, B2 => n3491
                           , ZN => n2805);
   U824 : OAI221_X1 port map( B1 => n2263, B2 => n2585, C1 => n3690, C2 => 
                           n2586, A => n2806, ZN => n2799);
   U825 : AOI22_X1 port map( A1 => n2588, A2 => n3488, B1 => n2589, B2 => n3489
                           , ZN => n2806);
   U826 : NOR4_X1 port map( A1 => n2807, A2 => n2808, A3 => n2809, A4 => n2810,
                           ZN => n2788);
   U827 : OAI221_X1 port map( B1 => n2264, B2 => n2594, C1 => n3706, C2 => 
                           n2595, A => n2811, ZN => n2810);
   U828 : AOI22_X1 port map( A1 => n2597, A2 => n3502, B1 => n2598, B2 => n3503
                           , ZN => n2811);
   U829 : OAI221_X1 port map( B1 => n2265, B2 => n2599, C1 => n3722, C2 => 
                           n2600, A => n2812, ZN => n2809);
   U830 : AOI22_X1 port map( A1 => n2602, A2 => n3500, B1 => n2603, B2 => n3501
                           , ZN => n2812);
   U831 : OAI221_X1 port map( B1 => n3746, B2 => n2604, C1 => n3738, C2 => 
                           n2605, A => n2813, ZN => n2808);
   U832 : AOI22_X1 port map( A1 => n2607, A2 => n3498, B1 => n2608, B2 => n3499
                           , ZN => n2813);
   U833 : OAI221_X1 port map( B1 => n3762, B2 => n2609, C1 => n3754, C2 => 
                           n2610, A => n2814, ZN => n2807);
   U834 : AOI22_X1 port map( A1 => n2612, A2 => n3496, B1 => n2613, B2 => n3497
                           , ZN => n2814);
   U835 : NOR4_X1 port map( A1 => n2815, A2 => n2816, A3 => n2817, A4 => n2818,
                           ZN => n2787);
   U836 : OAI221_X1 port map( B1 => n3778, B2 => n2618, C1 => n3770, C2 => 
                           n2619, A => n2819, ZN => n2818);
   U837 : AOI22_X1 port map( A1 => n2621, A2 => n3510, B1 => n2622, B2 => n3511
                           , ZN => n2819);
   U838 : OAI221_X1 port map( B1 => n2193, B2 => n2623, C1 => n2300, C2 => 
                           n2624, A => n2820, ZN => n2817);
   U839 : AOI22_X1 port map( A1 => n2626, A2 => n3508, B1 => n2627, B2 => n3509
                           , ZN => n2820);
   U840 : OAI221_X1 port map( B1 => n2194, B2 => n2628, C1 => n2301, C2 => 
                           n2629, A => n2821, ZN => n2816);
   U841 : AOI22_X1 port map( A1 => n2631, A2 => n3506, B1 => n2632, B2 => n3507
                           , ZN => n2821);
   U842 : OAI221_X1 port map( B1 => n2266, B2 => n2633, C1 => n3818, C2 => 
                           n2634, A => n2822, ZN => n2815);
   U843 : AOI22_X1 port map( A1 => n2636, A2 => n3504, B1 => n2637, B2 => n3505
                           , ZN => n2822);
   U844 : MUX2_X1 port map( A => OUT2_1_port, B => n2823, S => n2537, Z => 
                           n1484);
   U845 : NAND4_X1 port map( A1 => n2824, A2 => n2825, A3 => n2826, A4 => n2827
                           , ZN => n2823);
   U846 : NOR4_X1 port map( A1 => n2828, A2 => n2829, A3 => n2830, A4 => n2831,
                           ZN => n2827);
   U847 : OAI221_X1 port map( B1 => n2267, B2 => n2546, C1 => n3577, C2 => 
                           n2547, A => n2832, ZN => n2831);
   U848 : AOI22_X1 port map( A1 => n2549, A2 => n3518, B1 => n2550, B2 => n3519
                           , ZN => n2832);
   U849 : OAI221_X1 port map( B1 => n2268, B2 => n2551, C1 => n3593, C2 => 
                           n2552, A => n2833, ZN => n2830);
   U850 : AOI22_X1 port map( A1 => n2554, A2 => n3516, B1 => n2555, B2 => n3517
                           , ZN => n2833);
   U851 : OAI221_X1 port map( B1 => n2269, B2 => n2556, C1 => n3609, C2 => 
                           n2557, A => n2834, ZN => n2829);
   U852 : AOI22_X1 port map( A1 => n2559, A2 => n3514, B1 => n2560, B2 => n3515
                           , ZN => n2834);
   U853 : OAI221_X1 port map( B1 => n2270, B2 => n2561, C1 => n3625, C2 => 
                           n2562, A => n2835, ZN => n2828);
   U854 : AOI22_X1 port map( A1 => n2564, A2 => n3512, B1 => n2565, B2 => n3513
                           , ZN => n2835);
   U855 : NOR4_X1 port map( A1 => n2836, A2 => n2837, A3 => n2838, A4 => n2839,
                           ZN => n2826);
   U856 : OAI221_X1 port map( B1 => n2271, B2 => n2570, C1 => n3641, C2 => 
                           n2571, A => n2840, ZN => n2839);
   U857 : AOI22_X1 port map( A1 => n2573, A2 => n3526, B1 => n2574, B2 => n3527
                           , ZN => n2840);
   U858 : OAI221_X1 port map( B1 => n2272, B2 => n2575, C1 => n3657, C2 => 
                           n2576, A => n2841, ZN => n2838);
   U859 : AOI22_X1 port map( A1 => n2578, A2 => n3524, B1 => n2579, B2 => n3525
                           , ZN => n2841);
   U860 : OAI221_X1 port map( B1 => n2273, B2 => n2580, C1 => n3673, C2 => 
                           n2581, A => n2842, ZN => n2837);
   U861 : AOI22_X1 port map( A1 => n2583, A2 => n3522, B1 => n2584, B2 => n3523
                           , ZN => n2842);
   U862 : OAI221_X1 port map( B1 => n2274, B2 => n2585, C1 => n3689, C2 => 
                           n2586, A => n2843, ZN => n2836);
   U863 : AOI22_X1 port map( A1 => n2588, A2 => n3520, B1 => n2589, B2 => n3521
                           , ZN => n2843);
   U864 : NOR4_X1 port map( A1 => n2844, A2 => n2845, A3 => n2846, A4 => n2847,
                           ZN => n2825);
   U865 : OAI221_X1 port map( B1 => n2275, B2 => n2594, C1 => n3705, C2 => 
                           n2595, A => n2848, ZN => n2847);
   U866 : AOI22_X1 port map( A1 => n2597, A2 => n3534, B1 => n2598, B2 => n3535
                           , ZN => n2848);
   U867 : OAI221_X1 port map( B1 => n2276, B2 => n2599, C1 => n3721, C2 => 
                           n2600, A => n2849, ZN => n2846);
   U868 : AOI22_X1 port map( A1 => n2602, A2 => n3532, B1 => n2603, B2 => n3533
                           , ZN => n2849);
   U869 : OAI221_X1 port map( B1 => n3745, B2 => n2604, C1 => n3737, C2 => 
                           n2605, A => n2850, ZN => n2845);
   U870 : AOI22_X1 port map( A1 => n2607, A2 => n3530, B1 => n2608, B2 => n3531
                           , ZN => n2850);
   U871 : OAI221_X1 port map( B1 => n3761, B2 => n2609, C1 => n3753, C2 => 
                           n2610, A => n2851, ZN => n2844);
   U872 : AOI22_X1 port map( A1 => n2612, A2 => n3528, B1 => n2613, B2 => n3529
                           , ZN => n2851);
   U873 : NOR4_X1 port map( A1 => n2852, A2 => n2853, A3 => n2854, A4 => n2855,
                           ZN => n2824);
   U874 : OAI221_X1 port map( B1 => n3777, B2 => n2618, C1 => n3769, C2 => 
                           n2619, A => n2856, ZN => n2855);
   U875 : AOI22_X1 port map( A1 => n2621, A2 => n3542, B1 => n2622, B2 => n3543
                           , ZN => n2856);
   U876 : OAI221_X1 port map( B1 => n2195, B2 => n2623, C1 => n2302, C2 => 
                           n2624, A => n2857, ZN => n2854);
   U877 : AOI22_X1 port map( A1 => n2626, A2 => n3540, B1 => n2627, B2 => n3541
                           , ZN => n2857);
   U878 : OAI221_X1 port map( B1 => n2196, B2 => n2628, C1 => n2303, C2 => 
                           n2629, A => n2858, ZN => n2853);
   U879 : AOI22_X1 port map( A1 => n2631, A2 => n3538, B1 => n2632, B2 => n3539
                           , ZN => n2858);
   U880 : OAI221_X1 port map( B1 => n2277, B2 => n2633, C1 => n3817, C2 => 
                           n2634, A => n2859, ZN => n2852);
   U881 : AOI22_X1 port map( A1 => n2636, A2 => n3536, B1 => n2637, B2 => n3537
                           , ZN => n2859);
   U882 : MUX2_X1 port map( A => OUT2_0_port, B => n2860, S => n2537, Z => 
                           n1483);
   U883 : AND3_X1 port map( A1 => ENABLE, A2 => n2450, A3 => RD2, ZN => n2537);
   U884 : NAND4_X1 port map( A1 => n2861, A2 => n2862, A3 => n2863, A4 => n2864
                           , ZN => n2860);
   U885 : NOR4_X1 port map( A1 => n2865, A2 => n2866, A3 => n2867, A4 => n2868,
                           ZN => n2864);
   U886 : OAI221_X1 port map( B1 => n2278, B2 => n2546, C1 => n3576, C2 => 
                           n2547, A => n2869, ZN => n2868);
   U887 : AOI22_X1 port map( A1 => n2549, A2 => n3550, B1 => n2550, B2 => n3551
                           , ZN => n2869);
   U888 : AND2_X1 port map( A1 => n2870, A2 => n2871, ZN => n2550);
   U889 : AND2_X1 port map( A1 => n2870, A2 => n2872, ZN => n2549);
   U890 : NAND2_X1 port map( A1 => n2870, A2 => n2873, ZN => n2547);
   U891 : NAND2_X1 port map( A1 => n2870, A2 => n2874, ZN => n2546);
   U892 : AND2_X1 port map( A1 => n2875, A2 => n2876, ZN => n2870);
   U893 : OAI221_X1 port map( B1 => n2279, B2 => n2551, C1 => n3592, C2 => 
                           n2552, A => n2877, ZN => n2867);
   U894 : AOI22_X1 port map( A1 => n2554, A2 => n3548, B1 => n2555, B2 => n3549
                           , ZN => n2877);
   U895 : AND2_X1 port map( A1 => n2878, A2 => n2871, ZN => n2555);
   U896 : AND2_X1 port map( A1 => n2878, A2 => n2872, ZN => n2554);
   U897 : NAND2_X1 port map( A1 => n2878, A2 => n2873, ZN => n2552);
   U898 : NAND2_X1 port map( A1 => n2878, A2 => n2874, ZN => n2551);
   U899 : AND2_X1 port map( A1 => n2879, A2 => n2876, ZN => n2878);
   U900 : OAI221_X1 port map( B1 => n2280, B2 => n2556, C1 => n3608, C2 => 
                           n2557, A => n2880, ZN => n2866);
   U901 : AOI22_X1 port map( A1 => n2559, A2 => n3546, B1 => n2560, B2 => n3547
                           , ZN => n2880);
   U902 : AND2_X1 port map( A1 => n2881, A2 => n2871, ZN => n2560);
   U903 : AND2_X1 port map( A1 => n2881, A2 => n2872, ZN => n2559);
   U904 : NAND2_X1 port map( A1 => n2881, A2 => n2873, ZN => n2557);
   U905 : NAND2_X1 port map( A1 => n2881, A2 => n2874, ZN => n2556);
   U906 : AND2_X1 port map( A1 => n2882, A2 => n2876, ZN => n2881);
   U907 : OAI221_X1 port map( B1 => n2281, B2 => n2561, C1 => n3624, C2 => 
                           n2562, A => n2883, ZN => n2865);
   U908 : AOI22_X1 port map( A1 => n2564, A2 => n3544, B1 => n2565, B2 => n3545
                           , ZN => n2883);
   U909 : AND2_X1 port map( A1 => n2871, A2 => n2884, ZN => n2565);
   U910 : AND2_X1 port map( A1 => n2872, A2 => n2884, ZN => n2564);
   U911 : NAND2_X1 port map( A1 => n2873, A2 => n2884, ZN => n2562);
   U912 : NAND2_X1 port map( A1 => n2874, A2 => n2884, ZN => n2561);
   U913 : AND2_X1 port map( A1 => n2876, A2 => n2885, ZN => n2884);
   U914 : AND2_X1 port map( A1 => ADD_RD2(5), A2 => ADD_RD2(4), ZN => n2876);
   U915 : NOR4_X1 port map( A1 => n2886, A2 => n2887, A3 => n2888, A4 => n2889,
                           ZN => n2863);
   U916 : OAI221_X1 port map( B1 => n2282, B2 => n2570, C1 => n3640, C2 => 
                           n2571, A => n2890, ZN => n2889);
   U917 : AOI22_X1 port map( A1 => n2573, A2 => n3558, B1 => n2574, B2 => n3559
                           , ZN => n2890);
   U918 : AND2_X1 port map( A1 => n2891, A2 => n2871, ZN => n2574);
   U919 : AND2_X1 port map( A1 => n2891, A2 => n2872, ZN => n2573);
   U920 : NAND2_X1 port map( A1 => n2891, A2 => n2873, ZN => n2571);
   U921 : NAND2_X1 port map( A1 => n2891, A2 => n2874, ZN => n2570);
   U922 : AND2_X1 port map( A1 => n2892, A2 => n2875, ZN => n2891);
   U923 : OAI221_X1 port map( B1 => n2283, B2 => n2575, C1 => n3656, C2 => 
                           n2576, A => n2893, ZN => n2888);
   U924 : AOI22_X1 port map( A1 => n2578, A2 => n3556, B1 => n2579, B2 => n3557
                           , ZN => n2893);
   U925 : AND2_X1 port map( A1 => n2894, A2 => n2871, ZN => n2579);
   U926 : AND2_X1 port map( A1 => n2894, A2 => n2872, ZN => n2578);
   U927 : NAND2_X1 port map( A1 => n2894, A2 => n2873, ZN => n2576);
   U928 : NAND2_X1 port map( A1 => n2894, A2 => n2874, ZN => n2575);
   U929 : AND2_X1 port map( A1 => n2892, A2 => n2879, ZN => n2894);
   U930 : OAI221_X1 port map( B1 => n2284, B2 => n2580, C1 => n3672, C2 => 
                           n2581, A => n2895, ZN => n2887);
   U931 : AOI22_X1 port map( A1 => n2583, A2 => n3554, B1 => n2584, B2 => n3555
                           , ZN => n2895);
   U932 : AND2_X1 port map( A1 => n2896, A2 => n2871, ZN => n2584);
   U933 : AND2_X1 port map( A1 => n2896, A2 => n2872, ZN => n2583);
   U934 : NAND2_X1 port map( A1 => n2896, A2 => n2873, ZN => n2581);
   U935 : NAND2_X1 port map( A1 => n2896, A2 => n2874, ZN => n2580);
   U936 : AND2_X1 port map( A1 => n2892, A2 => n2882, ZN => n2896);
   U937 : OAI221_X1 port map( B1 => n2285, B2 => n2585, C1 => n3688, C2 => 
                           n2586, A => n2897, ZN => n2886);
   U938 : AOI22_X1 port map( A1 => n2588, A2 => n3552, B1 => n2589, B2 => n3553
                           , ZN => n2897);
   U939 : AND2_X1 port map( A1 => n2898, A2 => n2871, ZN => n2589);
   U940 : AND2_X1 port map( A1 => n2898, A2 => n2872, ZN => n2588);
   U941 : NAND2_X1 port map( A1 => n2898, A2 => n2873, ZN => n2586);
   U942 : NAND2_X1 port map( A1 => n2898, A2 => n2874, ZN => n2585);
   U943 : AND2_X1 port map( A1 => n2892, A2 => n2885, ZN => n2898);
   U944 : AND2_X1 port map( A1 => ADD_RD2(5), A2 => n2899, ZN => n2892);
   U945 : NOR4_X1 port map( A1 => n2900, A2 => n2901, A3 => n2902, A4 => n2903,
                           ZN => n2862);
   U946 : OAI221_X1 port map( B1 => n2286, B2 => n2594, C1 => n3704, C2 => 
                           n2595, A => n2904, ZN => n2903);
   U947 : AOI22_X1 port map( A1 => n2597, A2 => n3566, B1 => n2598, B2 => n3567
                           , ZN => n2904);
   U948 : AND2_X1 port map( A1 => n2905, A2 => n2871, ZN => n2598);
   U949 : AND2_X1 port map( A1 => n2905, A2 => n2872, ZN => n2597);
   U950 : NAND2_X1 port map( A1 => n2905, A2 => n2873, ZN => n2595);
   U951 : NAND2_X1 port map( A1 => n2905, A2 => n2874, ZN => n2594);
   U952 : AND2_X1 port map( A1 => n2906, A2 => n2875, ZN => n2905);
   U953 : OAI221_X1 port map( B1 => n2287, B2 => n2599, C1 => n3720, C2 => 
                           n2600, A => n2907, ZN => n2902);
   U954 : AOI22_X1 port map( A1 => n2602, A2 => n3564, B1 => n2603, B2 => n3565
                           , ZN => n2907);
   U955 : AND2_X1 port map( A1 => n2908, A2 => n2871, ZN => n2603);
   U956 : AND2_X1 port map( A1 => n2908, A2 => n2872, ZN => n2602);
   U957 : NAND2_X1 port map( A1 => n2908, A2 => n2873, ZN => n2600);
   U958 : NAND2_X1 port map( A1 => n2908, A2 => n2874, ZN => n2599);
   U959 : AND2_X1 port map( A1 => n2906, A2 => n2879, ZN => n2908);
   U960 : OAI221_X1 port map( B1 => n3744, B2 => n2604, C1 => n3736, C2 => 
                           n2605, A => n2909, ZN => n2901);
   U961 : AOI22_X1 port map( A1 => n2607, A2 => n3562, B1 => n2608, B2 => n3563
                           , ZN => n2909);
   U962 : AND2_X1 port map( A1 => n2910, A2 => n2871, ZN => n2608);
   U963 : AND2_X1 port map( A1 => n2910, A2 => n2872, ZN => n2607);
   U964 : NAND2_X1 port map( A1 => n2910, A2 => n2873, ZN => n2605);
   U965 : NAND2_X1 port map( A1 => n2910, A2 => n2874, ZN => n2604);
   U966 : AND2_X1 port map( A1 => n2906, A2 => n2882, ZN => n2910);
   U967 : OAI221_X1 port map( B1 => n3760, B2 => n2609, C1 => n3752, C2 => 
                           n2610, A => n2911, ZN => n2900);
   U968 : AOI22_X1 port map( A1 => n2612, A2 => n3560, B1 => n2613, B2 => n3561
                           , ZN => n2911);
   U969 : AND2_X1 port map( A1 => n2912, A2 => n2871, ZN => n2613);
   U970 : AND2_X1 port map( A1 => n2912, A2 => n2872, ZN => n2612);
   U971 : NAND2_X1 port map( A1 => n2912, A2 => n2873, ZN => n2610);
   U972 : NAND2_X1 port map( A1 => n2912, A2 => n2874, ZN => n2609);
   U973 : AND2_X1 port map( A1 => n2906, A2 => n2885, ZN => n2912);
   U974 : NOR2_X1 port map( A1 => n2899, A2 => ADD_RD2(5), ZN => n2906);
   U975 : INV_X1 port map( A => ADD_RD2(4), ZN => n2899);
   U976 : NOR4_X1 port map( A1 => n2913, A2 => n2914, A3 => n2915, A4 => n2916,
                           ZN => n2861);
   U977 : OAI221_X1 port map( B1 => n3776, B2 => n2618, C1 => n3768, C2 => 
                           n2619, A => n2917, ZN => n2916);
   U978 : AOI22_X1 port map( A1 => n2621, A2 => n3574, B1 => n2622, B2 => n3575
                           , ZN => n2917);
   U979 : AND2_X1 port map( A1 => n2918, A2 => n2871, ZN => n2622);
   U980 : AND2_X1 port map( A1 => n2918, A2 => n2872, ZN => n2621);
   U981 : NAND2_X1 port map( A1 => n2918, A2 => n2873, ZN => n2619);
   U982 : NAND2_X1 port map( A1 => n2918, A2 => n2874, ZN => n2618);
   U983 : AND2_X1 port map( A1 => n2919, A2 => n2875, ZN => n2918);
   U984 : AND2_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(2), ZN => n2875);
   U985 : OAI221_X1 port map( B1 => n2197, B2 => n2623, C1 => n2304, C2 => 
                           n2624, A => n2920, ZN => n2915);
   U986 : AOI22_X1 port map( A1 => n2626, A2 => n3572, B1 => n2627, B2 => n3573
                           , ZN => n2920);
   U987 : AND2_X1 port map( A1 => n2921, A2 => n2871, ZN => n2627);
   U988 : AND2_X1 port map( A1 => n2921, A2 => n2872, ZN => n2626);
   U989 : NAND2_X1 port map( A1 => n2921, A2 => n2873, ZN => n2624);
   U990 : NAND2_X1 port map( A1 => n2921, A2 => n2874, ZN => n2623);
   U991 : AND2_X1 port map( A1 => n2919, A2 => n2879, ZN => n2921);
   U992 : AND2_X1 port map( A1 => ADD_RD2(3), A2 => n2922, ZN => n2879);
   U993 : OAI221_X1 port map( B1 => n2198, B2 => n2628, C1 => n2305, C2 => 
                           n2629, A => n2923, ZN => n2914);
   U994 : AOI22_X1 port map( A1 => n2631, A2 => n3570, B1 => n2632, B2 => n3571
                           , ZN => n2923);
   U995 : AND2_X1 port map( A1 => n2924, A2 => n2871, ZN => n2632);
   U996 : AND2_X1 port map( A1 => n2924, A2 => n2872, ZN => n2631);
   U997 : NAND2_X1 port map( A1 => n2924, A2 => n2873, ZN => n2629);
   U998 : NAND2_X1 port map( A1 => n2924, A2 => n2874, ZN => n2628);
   U999 : AND2_X1 port map( A1 => n2919, A2 => n2882, ZN => n2924);
   U1000 : NOR2_X1 port map( A1 => n2922, A2 => ADD_RD2(3), ZN => n2882);
   U1001 : INV_X1 port map( A => ADD_RD2(2), ZN => n2922);
   U1002 : OAI221_X1 port map( B1 => n2288, B2 => n2633, C1 => n3816, C2 => 
                           n2634, A => n2925, ZN => n2913);
   U1003 : AOI22_X1 port map( A1 => n2636, A2 => n3568, B1 => n2637, B2 => 
                           n3569, ZN => n2925);
   U1004 : AND2_X1 port map( A1 => n2926, A2 => n2871, ZN => n2637);
   U1005 : AND2_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(1), ZN => n2871);
   U1006 : AND2_X1 port map( A1 => n2926, A2 => n2872, ZN => n2636);
   U1007 : AND2_X1 port map( A1 => ADD_RD2(1), A2 => n2927, ZN => n2872);
   U1008 : NAND2_X1 port map( A1 => n2926, A2 => n2873, ZN => n2634);
   U1009 : INV_X1 port map( A => ADD_RD2(0), ZN => n2927);
   U1010 : NAND2_X1 port map( A1 => n2926, A2 => n2874, ZN => n2633);
   U1011 : AND2_X1 port map( A1 => n2919, A2 => n2885, ZN => n2926);
   U1012 : NOR2_X1 port map( A1 => ADD_RD2(2), A2 => ADD_RD2(3), ZN => n2885);
   U1013 : NOR2_X1 port map( A1 => ADD_RD2(4), A2 => ADD_RD2(5), ZN => n2919);
   U1014 : MUX2_X1 port map( A => OUT1_7_port, B => n2928, S => n2929, Z => 
                           n1482);
   U1015 : NAND4_X1 port map( A1 => n2930, A2 => n2931, A3 => n2932, A4 => 
                           n2933, ZN => n2928);
   U1016 : NOR4_X1 port map( A1 => n2934, A2 => n2935, A3 => n2936, A4 => n2937
                           , ZN => n2933);
   U1017 : OAI221_X1 port map( B1 => n2199, B2 => n2938, C1 => n3583, C2 => 
                           n2939, A => n2940, ZN => n2937);
   U1018 : AOI22_X1 port map( A1 => n2941, A2 => n3326, B1 => n2942, B2 => 
                           n3327, ZN => n2940);
   U1019 : OAI221_X1 port map( B1 => n2200, B2 => n2943, C1 => n3599, C2 => 
                           n2944, A => n2945, ZN => n2936);
   U1020 : AOI22_X1 port map( A1 => n2946, A2 => n3324, B1 => n2947, B2 => 
                           n3325, ZN => n2945);
   U1021 : OAI221_X1 port map( B1 => n2201, B2 => n2948, C1 => n3615, C2 => 
                           n2949, A => n2950, ZN => n2935);
   U1022 : AOI22_X1 port map( A1 => n2951, A2 => n3322, B1 => n2952, B2 => 
                           n3323, ZN => n2950);
   U1023 : OAI221_X1 port map( B1 => n2202, B2 => n2953, C1 => n3631, C2 => 
                           n2954, A => n2955, ZN => n2934);
   U1024 : AOI22_X1 port map( A1 => n2956, A2 => n3320, B1 => n2957, B2 => 
                           n3321, ZN => n2955);
   U1025 : NOR4_X1 port map( A1 => n2958, A2 => n2959, A3 => n2960, A4 => n2961
                           , ZN => n2932);
   U1026 : OAI221_X1 port map( B1 => n2203, B2 => n2962, C1 => n3647, C2 => 
                           n2963, A => n2964, ZN => n2961);
   U1027 : AOI22_X1 port map( A1 => n2965, A2 => n3334, B1 => n2966, B2 => 
                           n3335, ZN => n2964);
   U1028 : OAI221_X1 port map( B1 => n2204, B2 => n2967, C1 => n3663, C2 => 
                           n2968, A => n2969, ZN => n2960);
   U1029 : AOI22_X1 port map( A1 => n2970, A2 => n3332, B1 => n2971, B2 => 
                           n3333, ZN => n2969);
   U1030 : OAI221_X1 port map( B1 => n2205, B2 => n2972, C1 => n3679, C2 => 
                           n2973, A => n2974, ZN => n2959);
   U1031 : AOI22_X1 port map( A1 => n2975, A2 => n3330, B1 => n2976, B2 => 
                           n3331, ZN => n2974);
   U1032 : OAI221_X1 port map( B1 => n2206, B2 => n2977, C1 => n3695, C2 => 
                           n2978, A => n2979, ZN => n2958);
   U1033 : AOI22_X1 port map( A1 => n2980, A2 => n3328, B1 => n2981, B2 => 
                           n3329, ZN => n2979);
   U1034 : NOR4_X1 port map( A1 => n2982, A2 => n2983, A3 => n2984, A4 => n2985
                           , ZN => n2931);
   U1035 : OAI221_X1 port map( B1 => n2207, B2 => n2986, C1 => n3711, C2 => 
                           n2987, A => n2988, ZN => n2985);
   U1036 : AOI22_X1 port map( A1 => n2989, A2 => n3342, B1 => n2990, B2 => 
                           n3343, ZN => n2988);
   U1037 : OAI221_X1 port map( B1 => n2208, B2 => n2991, C1 => n3727, C2 => 
                           n2992, A => n2993, ZN => n2984);
   U1038 : AOI22_X1 port map( A1 => n2994, A2 => n3340, B1 => n2995, B2 => 
                           n3341, ZN => n2993);
   U1039 : OAI221_X1 port map( B1 => n3751, B2 => n2996, C1 => n3743, C2 => 
                           n2997, A => n2998, ZN => n2983);
   U1040 : AOI22_X1 port map( A1 => n2999, A2 => n3338, B1 => n3000, B2 => 
                           n3339, ZN => n2998);
   U1041 : OAI221_X1 port map( B1 => n3767, B2 => n3001, C1 => n3759, C2 => 
                           n3002, A => n3003, ZN => n2982);
   U1042 : AOI22_X1 port map( A1 => n3004, A2 => n3336, B1 => n3005, B2 => 
                           n3337, ZN => n3003);
   U1043 : NOR4_X1 port map( A1 => n3006, A2 => n3007, A3 => n3008, A4 => n3009
                           , ZN => n2930);
   U1044 : OAI221_X1 port map( B1 => n2209, B2 => n3010, C1 => n3775, C2 => 
                           n3011, A => n3012, ZN => n3009);
   U1045 : AOI22_X1 port map( A1 => n3013, A2 => n3350, B1 => n3014, B2 => 
                           n3351, ZN => n3012);
   U1046 : OAI221_X1 port map( B1 => n2183, B2 => n3015, C1 => n2289, C2 => 
                           n3016, A => n3017, ZN => n3008);
   U1047 : AOI22_X1 port map( A1 => n3018, A2 => n3348, B1 => n3019, B2 => 
                           n3349, ZN => n3017);
   U1048 : OAI221_X1 port map( B1 => n2184, B2 => n3020, C1 => n2290, C2 => 
                           n3021, A => n3022, ZN => n3007);
   U1049 : AOI22_X1 port map( A1 => n3023, A2 => n3346, B1 => n3024, B2 => 
                           n3347, ZN => n3022);
   U1050 : OAI221_X1 port map( B1 => n3831, B2 => n3025, C1 => n2291, C2 => 
                           n3026, A => n3027, ZN => n3006);
   U1051 : AOI22_X1 port map( A1 => n3028, A2 => n3344, B1 => n3029, B2 => 
                           n3345, ZN => n3027);
   U1052 : MUX2_X1 port map( A => OUT1_6_port, B => n3030, S => n2929, Z => 
                           n1481);
   U1053 : NAND4_X1 port map( A1 => n3031, A2 => n3032, A3 => n3033, A4 => 
                           n3034, ZN => n3030);
   U1054 : NOR4_X1 port map( A1 => n3035, A2 => n3036, A3 => n3037, A4 => n3038
                           , ZN => n3034);
   U1055 : OAI221_X1 port map( B1 => n2210, B2 => n2938, C1 => n3582, C2 => 
                           n2939, A => n3039, ZN => n3038);
   U1056 : AOI22_X1 port map( A1 => n2941, A2 => n3358, B1 => n2942, B2 => 
                           n3359, ZN => n3039);
   U1057 : OAI221_X1 port map( B1 => n2211, B2 => n2943, C1 => n3598, C2 => 
                           n2944, A => n3040, ZN => n3037);
   U1058 : AOI22_X1 port map( A1 => n2946, A2 => n3356, B1 => n2947, B2 => 
                           n3357, ZN => n3040);
   U1059 : OAI221_X1 port map( B1 => n2212, B2 => n2948, C1 => n3614, C2 => 
                           n2949, A => n3041, ZN => n3036);
   U1060 : AOI22_X1 port map( A1 => n2951, A2 => n3354, B1 => n2952, B2 => 
                           n3355, ZN => n3041);
   U1061 : OAI221_X1 port map( B1 => n2213, B2 => n2953, C1 => n3630, C2 => 
                           n2954, A => n3042, ZN => n3035);
   U1062 : AOI22_X1 port map( A1 => n2956, A2 => n3352, B1 => n2957, B2 => 
                           n3353, ZN => n3042);
   U1063 : NOR4_X1 port map( A1 => n3043, A2 => n3044, A3 => n3045, A4 => n3046
                           , ZN => n3033);
   U1064 : OAI221_X1 port map( B1 => n2214, B2 => n2962, C1 => n3646, C2 => 
                           n2963, A => n3047, ZN => n3046);
   U1065 : AOI22_X1 port map( A1 => n2965, A2 => n3366, B1 => n2966, B2 => 
                           n3367, ZN => n3047);
   U1066 : OAI221_X1 port map( B1 => n2215, B2 => n2967, C1 => n3662, C2 => 
                           n2968, A => n3048, ZN => n3045);
   U1067 : AOI22_X1 port map( A1 => n2970, A2 => n3364, B1 => n2971, B2 => 
                           n3365, ZN => n3048);
   U1068 : OAI221_X1 port map( B1 => n2216, B2 => n2972, C1 => n3678, C2 => 
                           n2973, A => n3049, ZN => n3044);
   U1069 : AOI22_X1 port map( A1 => n2975, A2 => n3362, B1 => n2976, B2 => 
                           n3363, ZN => n3049);
   U1070 : OAI221_X1 port map( B1 => n2217, B2 => n2977, C1 => n3694, C2 => 
                           n2978, A => n3050, ZN => n3043);
   U1071 : AOI22_X1 port map( A1 => n2980, A2 => n3360, B1 => n2981, B2 => 
                           n3361, ZN => n3050);
   U1072 : NOR4_X1 port map( A1 => n3051, A2 => n3052, A3 => n3053, A4 => n3054
                           , ZN => n3032);
   U1073 : OAI221_X1 port map( B1 => n2218, B2 => n2986, C1 => n3710, C2 => 
                           n2987, A => n3055, ZN => n3054);
   U1074 : AOI22_X1 port map( A1 => n2989, A2 => n3374, B1 => n2990, B2 => 
                           n3375, ZN => n3055);
   U1075 : OAI221_X1 port map( B1 => n2219, B2 => n2991, C1 => n3726, C2 => 
                           n2992, A => n3056, ZN => n3053);
   U1076 : AOI22_X1 port map( A1 => n2994, A2 => n3372, B1 => n2995, B2 => 
                           n3373, ZN => n3056);
   U1077 : OAI221_X1 port map( B1 => n3750, B2 => n2996, C1 => n3742, C2 => 
                           n2997, A => n3057, ZN => n3052);
   U1078 : AOI22_X1 port map( A1 => n2999, A2 => n3370, B1 => n3000, B2 => 
                           n3371, ZN => n3057);
   U1079 : OAI221_X1 port map( B1 => n3766, B2 => n3001, C1 => n3758, C2 => 
                           n3002, A => n3058, ZN => n3051);
   U1080 : AOI22_X1 port map( A1 => n3004, A2 => n3368, B1 => n3005, B2 => 
                           n3369, ZN => n3058);
   U1081 : NOR4_X1 port map( A1 => n3059, A2 => n3060, A3 => n3061, A4 => n3062
                           , ZN => n3031);
   U1082 : OAI221_X1 port map( B1 => n2220, B2 => n3010, C1 => n3774, C2 => 
                           n3011, A => n3063, ZN => n3062);
   U1083 : AOI22_X1 port map( A1 => n3013, A2 => n3382, B1 => n3014, B2 => 
                           n3383, ZN => n3063);
   U1084 : OAI221_X1 port map( B1 => n2185, B2 => n3015, C1 => n2292, C2 => 
                           n3016, A => n3064, ZN => n3061);
   U1085 : AOI22_X1 port map( A1 => n3018, A2 => n3380, B1 => n3019, B2 => 
                           n3381, ZN => n3064);
   U1086 : OAI221_X1 port map( B1 => n2186, B2 => n3020, C1 => n2293, C2 => 
                           n3021, A => n3065, ZN => n3060);
   U1087 : AOI22_X1 port map( A1 => n3023, A2 => n3378, B1 => n3024, B2 => 
                           n3379, ZN => n3065);
   U1088 : OAI221_X1 port map( B1 => n2221, B2 => n3025, C1 => n3822, C2 => 
                           n3026, A => n3066, ZN => n3059);
   U1089 : AOI22_X1 port map( A1 => n3028, A2 => n3376, B1 => n3029, B2 => 
                           n3377, ZN => n3066);
   U1090 : MUX2_X1 port map( A => OUT1_5_port, B => n3067, S => n2929, Z => 
                           n1480);
   U1091 : NAND4_X1 port map( A1 => n3068, A2 => n3069, A3 => n3070, A4 => 
                           n3071, ZN => n3067);
   U1092 : NOR4_X1 port map( A1 => n3072, A2 => n3073, A3 => n3074, A4 => n3075
                           , ZN => n3071);
   U1093 : OAI221_X1 port map( B1 => n2222, B2 => n2938, C1 => n3581, C2 => 
                           n2939, A => n3076, ZN => n3075);
   U1094 : AOI22_X1 port map( A1 => n2941, A2 => n3390, B1 => n2942, B2 => 
                           n3391, ZN => n3076);
   U1095 : OAI221_X1 port map( B1 => n2223, B2 => n2943, C1 => n3597, C2 => 
                           n2944, A => n3077, ZN => n3074);
   U1096 : AOI22_X1 port map( A1 => n2946, A2 => n3388, B1 => n2947, B2 => 
                           n3389, ZN => n3077);
   U1097 : OAI221_X1 port map( B1 => n2224, B2 => n2948, C1 => n3613, C2 => 
                           n2949, A => n3078, ZN => n3073);
   U1098 : AOI22_X1 port map( A1 => n2951, A2 => n3386, B1 => n2952, B2 => 
                           n3387, ZN => n3078);
   U1099 : OAI221_X1 port map( B1 => n2225, B2 => n2953, C1 => n3629, C2 => 
                           n2954, A => n3079, ZN => n3072);
   U1100 : AOI22_X1 port map( A1 => n2956, A2 => n3384, B1 => n2957, B2 => 
                           n3385, ZN => n3079);
   U1101 : NOR4_X1 port map( A1 => n3080, A2 => n3081, A3 => n3082, A4 => n3083
                           , ZN => n3070);
   U1102 : OAI221_X1 port map( B1 => n2226, B2 => n2962, C1 => n3645, C2 => 
                           n2963, A => n3084, ZN => n3083);
   U1103 : AOI22_X1 port map( A1 => n2965, A2 => n3398, B1 => n2966, B2 => 
                           n3399, ZN => n3084);
   U1104 : OAI221_X1 port map( B1 => n2227, B2 => n2967, C1 => n3661, C2 => 
                           n2968, A => n3085, ZN => n3082);
   U1105 : AOI22_X1 port map( A1 => n2970, A2 => n3396, B1 => n2971, B2 => 
                           n3397, ZN => n3085);
   U1106 : OAI221_X1 port map( B1 => n2228, B2 => n2972, C1 => n3677, C2 => 
                           n2973, A => n3086, ZN => n3081);
   U1107 : AOI22_X1 port map( A1 => n2975, A2 => n3394, B1 => n2976, B2 => 
                           n3395, ZN => n3086);
   U1108 : OAI221_X1 port map( B1 => n2229, B2 => n2977, C1 => n3693, C2 => 
                           n2978, A => n3087, ZN => n3080);
   U1109 : AOI22_X1 port map( A1 => n2980, A2 => n3392, B1 => n2981, B2 => 
                           n3393, ZN => n3087);
   U1110 : NOR4_X1 port map( A1 => n3088, A2 => n3089, A3 => n3090, A4 => n3091
                           , ZN => n3069);
   U1111 : OAI221_X1 port map( B1 => n2230, B2 => n2986, C1 => n3709, C2 => 
                           n2987, A => n3092, ZN => n3091);
   U1112 : AOI22_X1 port map( A1 => n2989, A2 => n3406, B1 => n2990, B2 => 
                           n3407, ZN => n3092);
   U1113 : OAI221_X1 port map( B1 => n2231, B2 => n2991, C1 => n3725, C2 => 
                           n2992, A => n3093, ZN => n3090);
   U1114 : AOI22_X1 port map( A1 => n2994, A2 => n3404, B1 => n2995, B2 => 
                           n3405, ZN => n3093);
   U1115 : OAI221_X1 port map( B1 => n3749, B2 => n2996, C1 => n3741, C2 => 
                           n2997, A => n3094, ZN => n3089);
   U1116 : AOI22_X1 port map( A1 => n2999, A2 => n3402, B1 => n3000, B2 => 
                           n3403, ZN => n3094);
   U1117 : OAI221_X1 port map( B1 => n3765, B2 => n3001, C1 => n3757, C2 => 
                           n3002, A => n3095, ZN => n3088);
   U1118 : AOI22_X1 port map( A1 => n3004, A2 => n3400, B1 => n3005, B2 => 
                           n3401, ZN => n3095);
   U1119 : NOR4_X1 port map( A1 => n3096, A2 => n3097, A3 => n3098, A4 => n3099
                           , ZN => n3068);
   U1120 : OAI221_X1 port map( B1 => n2232, B2 => n3010, C1 => n3773, C2 => 
                           n3011, A => n3100, ZN => n3099);
   U1121 : AOI22_X1 port map( A1 => n3013, A2 => n3414, B1 => n3014, B2 => 
                           n3415, ZN => n3100);
   U1122 : OAI221_X1 port map( B1 => n2187, B2 => n3015, C1 => n2294, C2 => 
                           n3016, A => n3101, ZN => n3098);
   U1123 : AOI22_X1 port map( A1 => n3018, A2 => n3412, B1 => n3019, B2 => 
                           n3413, ZN => n3101);
   U1124 : OAI221_X1 port map( B1 => n2188, B2 => n3020, C1 => n2295, C2 => 
                           n3021, A => n3102, ZN => n3097);
   U1125 : AOI22_X1 port map( A1 => n3023, A2 => n3410, B1 => n3024, B2 => 
                           n3411, ZN => n3102);
   U1126 : OAI221_X1 port map( B1 => n2233, B2 => n3025, C1 => n3821, C2 => 
                           n3026, A => n3103, ZN => n3096);
   U1127 : AOI22_X1 port map( A1 => n3028, A2 => n3408, B1 => n3029, B2 => 
                           n3409, ZN => n3103);
   U1128 : MUX2_X1 port map( A => OUT1_4_port, B => n3104, S => n2929, Z => 
                           n1479);
   U1129 : NAND4_X1 port map( A1 => n3105, A2 => n3106, A3 => n3107, A4 => 
                           n3108, ZN => n3104);
   U1130 : NOR4_X1 port map( A1 => n3109, A2 => n3110, A3 => n3111, A4 => n3112
                           , ZN => n3108);
   U1131 : OAI221_X1 port map( B1 => n2234, B2 => n2938, C1 => n3580, C2 => 
                           n2939, A => n3113, ZN => n3112);
   U1132 : AOI22_X1 port map( A1 => n2941, A2 => n3422, B1 => n2942, B2 => 
                           n3423, ZN => n3113);
   U1133 : OAI221_X1 port map( B1 => n2235, B2 => n2943, C1 => n3596, C2 => 
                           n2944, A => n3114, ZN => n3111);
   U1134 : AOI22_X1 port map( A1 => n2946, A2 => n3420, B1 => n2947, B2 => 
                           n3421, ZN => n3114);
   U1135 : OAI221_X1 port map( B1 => n2236, B2 => n2948, C1 => n3612, C2 => 
                           n2949, A => n3115, ZN => n3110);
   U1136 : AOI22_X1 port map( A1 => n2951, A2 => n3418, B1 => n2952, B2 => 
                           n3419, ZN => n3115);
   U1137 : OAI221_X1 port map( B1 => n2237, B2 => n2953, C1 => n3628, C2 => 
                           n2954, A => n3116, ZN => n3109);
   U1138 : AOI22_X1 port map( A1 => n2956, A2 => n3416, B1 => n2957, B2 => 
                           n3417, ZN => n3116);
   U1139 : NOR4_X1 port map( A1 => n3117, A2 => n3118, A3 => n3119, A4 => n3120
                           , ZN => n3107);
   U1140 : OAI221_X1 port map( B1 => n2238, B2 => n2962, C1 => n3644, C2 => 
                           n2963, A => n3121, ZN => n3120);
   U1141 : AOI22_X1 port map( A1 => n2965, A2 => n3430, B1 => n2966, B2 => 
                           n3431, ZN => n3121);
   U1142 : OAI221_X1 port map( B1 => n2239, B2 => n2967, C1 => n3660, C2 => 
                           n2968, A => n3122, ZN => n3119);
   U1143 : AOI22_X1 port map( A1 => n2970, A2 => n3428, B1 => n2971, B2 => 
                           n3429, ZN => n3122);
   U1144 : OAI221_X1 port map( B1 => n2240, B2 => n2972, C1 => n3676, C2 => 
                           n2973, A => n3123, ZN => n3118);
   U1145 : AOI22_X1 port map( A1 => n2975, A2 => n3426, B1 => n2976, B2 => 
                           n3427, ZN => n3123);
   U1146 : OAI221_X1 port map( B1 => n2241, B2 => n2977, C1 => n3692, C2 => 
                           n2978, A => n3124, ZN => n3117);
   U1147 : AOI22_X1 port map( A1 => n2980, A2 => n3424, B1 => n2981, B2 => 
                           n3425, ZN => n3124);
   U1148 : NOR4_X1 port map( A1 => n3125, A2 => n3126, A3 => n3127, A4 => n3128
                           , ZN => n3106);
   U1149 : OAI221_X1 port map( B1 => n2242, B2 => n2986, C1 => n3708, C2 => 
                           n2987, A => n3129, ZN => n3128);
   U1150 : AOI22_X1 port map( A1 => n2989, A2 => n3438, B1 => n2990, B2 => 
                           n3439, ZN => n3129);
   U1151 : OAI221_X1 port map( B1 => n2243, B2 => n2991, C1 => n3724, C2 => 
                           n2992, A => n3130, ZN => n3127);
   U1152 : AOI22_X1 port map( A1 => n2994, A2 => n3436, B1 => n2995, B2 => 
                           n3437, ZN => n3130);
   U1153 : OAI221_X1 port map( B1 => n3748, B2 => n2996, C1 => n3740, C2 => 
                           n2997, A => n3131, ZN => n3126);
   U1154 : AOI22_X1 port map( A1 => n2999, A2 => n3434, B1 => n3000, B2 => 
                           n3435, ZN => n3131);
   U1155 : OAI221_X1 port map( B1 => n3764, B2 => n3001, C1 => n3756, C2 => 
                           n3002, A => n3132, ZN => n3125);
   U1156 : AOI22_X1 port map( A1 => n3004, A2 => n3432, B1 => n3005, B2 => 
                           n3433, ZN => n3132);
   U1157 : NOR4_X1 port map( A1 => n3133, A2 => n3134, A3 => n3135, A4 => n3136
                           , ZN => n3105);
   U1158 : OAI221_X1 port map( B1 => n3780, B2 => n3010, C1 => n3772, C2 => 
                           n3011, A => n3137, ZN => n3136);
   U1159 : AOI22_X1 port map( A1 => n3013, A2 => n3446, B1 => n3014, B2 => 
                           n3447, ZN => n3137);
   U1160 : OAI221_X1 port map( B1 => n2189, B2 => n3015, C1 => n2296, C2 => 
                           n3016, A => n3138, ZN => n3135);
   U1161 : AOI22_X1 port map( A1 => n3018, A2 => n3444, B1 => n3019, B2 => 
                           n3445, ZN => n3138);
   U1162 : OAI221_X1 port map( B1 => n2190, B2 => n3020, C1 => n2297, C2 => 
                           n3021, A => n3139, ZN => n3134);
   U1163 : AOI22_X1 port map( A1 => n3023, A2 => n3442, B1 => n3024, B2 => 
                           n3443, ZN => n3139);
   U1164 : OAI221_X1 port map( B1 => n2244, B2 => n3025, C1 => n3820, C2 => 
                           n3026, A => n3140, ZN => n3133);
   U1165 : AOI22_X1 port map( A1 => n3028, A2 => n3440, B1 => n3029, B2 => 
                           n3441, ZN => n3140);
   U1166 : MUX2_X1 port map( A => OUT1_3_port, B => n3141, S => n2929, Z => 
                           n1478);
   U1167 : NAND4_X1 port map( A1 => n3142, A2 => n3143, A3 => n3144, A4 => 
                           n3145, ZN => n3141);
   U1168 : NOR4_X1 port map( A1 => n3146, A2 => n3147, A3 => n3148, A4 => n3149
                           , ZN => n3145);
   U1169 : OAI221_X1 port map( B1 => n2245, B2 => n2938, C1 => n3579, C2 => 
                           n2939, A => n3150, ZN => n3149);
   U1170 : AOI22_X1 port map( A1 => n2941, A2 => n3454, B1 => n2942, B2 => 
                           n3455, ZN => n3150);
   U1171 : OAI221_X1 port map( B1 => n2246, B2 => n2943, C1 => n3595, C2 => 
                           n2944, A => n3151, ZN => n3148);
   U1172 : AOI22_X1 port map( A1 => n2946, A2 => n3452, B1 => n2947, B2 => 
                           n3453, ZN => n3151);
   U1173 : OAI221_X1 port map( B1 => n2247, B2 => n2948, C1 => n3611, C2 => 
                           n2949, A => n3152, ZN => n3147);
   U1174 : AOI22_X1 port map( A1 => n2951, A2 => n3450, B1 => n2952, B2 => 
                           n3451, ZN => n3152);
   U1175 : OAI221_X1 port map( B1 => n2248, B2 => n2953, C1 => n3627, C2 => 
                           n2954, A => n3153, ZN => n3146);
   U1176 : AOI22_X1 port map( A1 => n2956, A2 => n3448, B1 => n2957, B2 => 
                           n3449, ZN => n3153);
   U1177 : NOR4_X1 port map( A1 => n3154, A2 => n3155, A3 => n3156, A4 => n3157
                           , ZN => n3144);
   U1178 : OAI221_X1 port map( B1 => n2249, B2 => n2962, C1 => n3643, C2 => 
                           n2963, A => n3158, ZN => n3157);
   U1179 : AOI22_X1 port map( A1 => n2965, A2 => n3462, B1 => n2966, B2 => 
                           n3463, ZN => n3158);
   U1180 : OAI221_X1 port map( B1 => n2250, B2 => n2967, C1 => n3659, C2 => 
                           n2968, A => n3159, ZN => n3156);
   U1181 : AOI22_X1 port map( A1 => n2970, A2 => n3460, B1 => n2971, B2 => 
                           n3461, ZN => n3159);
   U1182 : OAI221_X1 port map( B1 => n2251, B2 => n2972, C1 => n3675, C2 => 
                           n2973, A => n3160, ZN => n3155);
   U1183 : AOI22_X1 port map( A1 => n2975, A2 => n3458, B1 => n2976, B2 => 
                           n3459, ZN => n3160);
   U1184 : OAI221_X1 port map( B1 => n2252, B2 => n2977, C1 => n3691, C2 => 
                           n2978, A => n3161, ZN => n3154);
   U1185 : AOI22_X1 port map( A1 => n2980, A2 => n3456, B1 => n2981, B2 => 
                           n3457, ZN => n3161);
   U1186 : NOR4_X1 port map( A1 => n3162, A2 => n3163, A3 => n3164, A4 => n3165
                           , ZN => n3143);
   U1187 : OAI221_X1 port map( B1 => n2253, B2 => n2986, C1 => n3707, C2 => 
                           n2987, A => n3166, ZN => n3165);
   U1188 : AOI22_X1 port map( A1 => n2989, A2 => n3470, B1 => n2990, B2 => 
                           n3471, ZN => n3166);
   U1189 : OAI221_X1 port map( B1 => n2254, B2 => n2991, C1 => n3723, C2 => 
                           n2992, A => n3167, ZN => n3164);
   U1190 : AOI22_X1 port map( A1 => n2994, A2 => n3468, B1 => n2995, B2 => 
                           n3469, ZN => n3167);
   U1191 : OAI221_X1 port map( B1 => n3747, B2 => n2996, C1 => n3739, C2 => 
                           n2997, A => n3168, ZN => n3163);
   U1192 : AOI22_X1 port map( A1 => n2999, A2 => n3466, B1 => n3000, B2 => 
                           n3467, ZN => n3168);
   U1193 : OAI221_X1 port map( B1 => n3763, B2 => n3001, C1 => n3755, C2 => 
                           n3002, A => n3169, ZN => n3162);
   U1194 : AOI22_X1 port map( A1 => n3004, A2 => n3464, B1 => n3005, B2 => 
                           n3465, ZN => n3169);
   U1195 : NOR4_X1 port map( A1 => n3170, A2 => n3171, A3 => n3172, A4 => n3173
                           , ZN => n3142);
   U1196 : OAI221_X1 port map( B1 => n3779, B2 => n3010, C1 => n3771, C2 => 
                           n3011, A => n3174, ZN => n3173);
   U1197 : AOI22_X1 port map( A1 => n3013, A2 => n3478, B1 => n3014, B2 => 
                           n3479, ZN => n3174);
   U1198 : OAI221_X1 port map( B1 => n2191, B2 => n3015, C1 => n2298, C2 => 
                           n3016, A => n3175, ZN => n3172);
   U1199 : AOI22_X1 port map( A1 => n3018, A2 => n3476, B1 => n3019, B2 => 
                           n3477, ZN => n3175);
   U1200 : OAI221_X1 port map( B1 => n2192, B2 => n3020, C1 => n2299, C2 => 
                           n3021, A => n3176, ZN => n3171);
   U1201 : AOI22_X1 port map( A1 => n3023, A2 => n3474, B1 => n3024, B2 => 
                           n3475, ZN => n3176);
   U1202 : OAI221_X1 port map( B1 => n2255, B2 => n3025, C1 => n3819, C2 => 
                           n3026, A => n3177, ZN => n3170);
   U1203 : AOI22_X1 port map( A1 => n3028, A2 => n3472, B1 => n3029, B2 => 
                           n3473, ZN => n3177);
   U1204 : MUX2_X1 port map( A => OUT1_2_port, B => n3178, S => n2929, Z => 
                           n1477);
   U1205 : NAND4_X1 port map( A1 => n3179, A2 => n3180, A3 => n3181, A4 => 
                           n3182, ZN => n3178);
   U1206 : NOR4_X1 port map( A1 => n3183, A2 => n3184, A3 => n3185, A4 => n3186
                           , ZN => n3182);
   U1207 : OAI221_X1 port map( B1 => n2256, B2 => n2938, C1 => n3578, C2 => 
                           n2939, A => n3187, ZN => n3186);
   U1208 : AOI22_X1 port map( A1 => n2941, A2 => n3486, B1 => n2942, B2 => 
                           n3487, ZN => n3187);
   U1209 : OAI221_X1 port map( B1 => n2257, B2 => n2943, C1 => n3594, C2 => 
                           n2944, A => n3188, ZN => n3185);
   U1210 : AOI22_X1 port map( A1 => n2946, A2 => n3484, B1 => n2947, B2 => 
                           n3485, ZN => n3188);
   U1211 : OAI221_X1 port map( B1 => n2258, B2 => n2948, C1 => n3610, C2 => 
                           n2949, A => n3189, ZN => n3184);
   U1212 : AOI22_X1 port map( A1 => n2951, A2 => n3482, B1 => n2952, B2 => 
                           n3483, ZN => n3189);
   U1213 : OAI221_X1 port map( B1 => n2259, B2 => n2953, C1 => n3626, C2 => 
                           n2954, A => n3190, ZN => n3183);
   U1214 : AOI22_X1 port map( A1 => n2956, A2 => n3480, B1 => n2957, B2 => 
                           n3481, ZN => n3190);
   U1215 : NOR4_X1 port map( A1 => n3191, A2 => n3192, A3 => n3193, A4 => n3194
                           , ZN => n3181);
   U1216 : OAI221_X1 port map( B1 => n2260, B2 => n2962, C1 => n3642, C2 => 
                           n2963, A => n3195, ZN => n3194);
   U1217 : AOI22_X1 port map( A1 => n2965, A2 => n3494, B1 => n2966, B2 => 
                           n3495, ZN => n3195);
   U1218 : OAI221_X1 port map( B1 => n2261, B2 => n2967, C1 => n3658, C2 => 
                           n2968, A => n3196, ZN => n3193);
   U1219 : AOI22_X1 port map( A1 => n2970, A2 => n3492, B1 => n2971, B2 => 
                           n3493, ZN => n3196);
   U1220 : OAI221_X1 port map( B1 => n2262, B2 => n2972, C1 => n3674, C2 => 
                           n2973, A => n3197, ZN => n3192);
   U1221 : AOI22_X1 port map( A1 => n2975, A2 => n3490, B1 => n2976, B2 => 
                           n3491, ZN => n3197);
   U1222 : OAI221_X1 port map( B1 => n2263, B2 => n2977, C1 => n3690, C2 => 
                           n2978, A => n3198, ZN => n3191);
   U1223 : AOI22_X1 port map( A1 => n2980, A2 => n3488, B1 => n2981, B2 => 
                           n3489, ZN => n3198);
   U1224 : NOR4_X1 port map( A1 => n3199, A2 => n3200, A3 => n3201, A4 => n3202
                           , ZN => n3180);
   U1225 : OAI221_X1 port map( B1 => n2264, B2 => n2986, C1 => n3706, C2 => 
                           n2987, A => n3203, ZN => n3202);
   U1226 : AOI22_X1 port map( A1 => n2989, A2 => n3502, B1 => n2990, B2 => 
                           n3503, ZN => n3203);
   U1227 : OAI221_X1 port map( B1 => n2265, B2 => n2991, C1 => n3722, C2 => 
                           n2992, A => n3204, ZN => n3201);
   U1228 : AOI22_X1 port map( A1 => n2994, A2 => n3500, B1 => n2995, B2 => 
                           n3501, ZN => n3204);
   U1229 : OAI221_X1 port map( B1 => n3746, B2 => n2996, C1 => n3738, C2 => 
                           n2997, A => n3205, ZN => n3200);
   U1230 : AOI22_X1 port map( A1 => n2999, A2 => n3498, B1 => n3000, B2 => 
                           n3499, ZN => n3205);
   U1231 : OAI221_X1 port map( B1 => n3762, B2 => n3001, C1 => n3754, C2 => 
                           n3002, A => n3206, ZN => n3199);
   U1232 : AOI22_X1 port map( A1 => n3004, A2 => n3496, B1 => n3005, B2 => 
                           n3497, ZN => n3206);
   U1233 : NOR4_X1 port map( A1 => n3207, A2 => n3208, A3 => n3209, A4 => n3210
                           , ZN => n3179);
   U1234 : OAI221_X1 port map( B1 => n3778, B2 => n3010, C1 => n3770, C2 => 
                           n3011, A => n3211, ZN => n3210);
   U1235 : AOI22_X1 port map( A1 => n3013, A2 => n3510, B1 => n3014, B2 => 
                           n3511, ZN => n3211);
   U1236 : OAI221_X1 port map( B1 => n2193, B2 => n3015, C1 => n2300, C2 => 
                           n3016, A => n3212, ZN => n3209);
   U1237 : AOI22_X1 port map( A1 => n3018, A2 => n3508, B1 => n3019, B2 => 
                           n3509, ZN => n3212);
   U1238 : OAI221_X1 port map( B1 => n2194, B2 => n3020, C1 => n2301, C2 => 
                           n3021, A => n3213, ZN => n3208);
   U1239 : AOI22_X1 port map( A1 => n3023, A2 => n3506, B1 => n3024, B2 => 
                           n3507, ZN => n3213);
   U1240 : OAI221_X1 port map( B1 => n2266, B2 => n3025, C1 => n3818, C2 => 
                           n3026, A => n3214, ZN => n3207);
   U1241 : AOI22_X1 port map( A1 => n3028, A2 => n3504, B1 => n3029, B2 => 
                           n3505, ZN => n3214);
   U1242 : MUX2_X1 port map( A => OUT1_1_port, B => n3215, S => n2929, Z => 
                           n1476);
   U1243 : NAND4_X1 port map( A1 => n3216, A2 => n3217, A3 => n3218, A4 => 
                           n3219, ZN => n3215);
   U1244 : NOR4_X1 port map( A1 => n3220, A2 => n3221, A3 => n3222, A4 => n3223
                           , ZN => n3219);
   U1245 : OAI221_X1 port map( B1 => n2267, B2 => n2938, C1 => n3577, C2 => 
                           n2939, A => n3224, ZN => n3223);
   U1246 : AOI22_X1 port map( A1 => n2941, A2 => n3518, B1 => n2942, B2 => 
                           n3519, ZN => n3224);
   U1247 : OAI221_X1 port map( B1 => n2268, B2 => n2943, C1 => n3593, C2 => 
                           n2944, A => n3225, ZN => n3222);
   U1248 : AOI22_X1 port map( A1 => n2946, A2 => n3516, B1 => n2947, B2 => 
                           n3517, ZN => n3225);
   U1249 : OAI221_X1 port map( B1 => n2269, B2 => n2948, C1 => n3609, C2 => 
                           n2949, A => n3226, ZN => n3221);
   U1250 : AOI22_X1 port map( A1 => n2951, A2 => n3514, B1 => n2952, B2 => 
                           n3515, ZN => n3226);
   U1251 : OAI221_X1 port map( B1 => n2270, B2 => n2953, C1 => n3625, C2 => 
                           n2954, A => n3227, ZN => n3220);
   U1252 : AOI22_X1 port map( A1 => n2956, A2 => n3512, B1 => n2957, B2 => 
                           n3513, ZN => n3227);
   U1253 : NOR4_X1 port map( A1 => n3228, A2 => n3229, A3 => n3230, A4 => n3231
                           , ZN => n3218);
   U1254 : OAI221_X1 port map( B1 => n2271, B2 => n2962, C1 => n3641, C2 => 
                           n2963, A => n3232, ZN => n3231);
   U1255 : AOI22_X1 port map( A1 => n2965, A2 => n3526, B1 => n2966, B2 => 
                           n3527, ZN => n3232);
   U1256 : OAI221_X1 port map( B1 => n2272, B2 => n2967, C1 => n3657, C2 => 
                           n2968, A => n3233, ZN => n3230);
   U1257 : AOI22_X1 port map( A1 => n2970, A2 => n3524, B1 => n2971, B2 => 
                           n3525, ZN => n3233);
   U1258 : OAI221_X1 port map( B1 => n2273, B2 => n2972, C1 => n3673, C2 => 
                           n2973, A => n3234, ZN => n3229);
   U1259 : AOI22_X1 port map( A1 => n2975, A2 => n3522, B1 => n2976, B2 => 
                           n3523, ZN => n3234);
   U1260 : OAI221_X1 port map( B1 => n2274, B2 => n2977, C1 => n3689, C2 => 
                           n2978, A => n3235, ZN => n3228);
   U1261 : AOI22_X1 port map( A1 => n2980, A2 => n3520, B1 => n2981, B2 => 
                           n3521, ZN => n3235);
   U1262 : NOR4_X1 port map( A1 => n3236, A2 => n3237, A3 => n3238, A4 => n3239
                           , ZN => n3217);
   U1263 : OAI221_X1 port map( B1 => n2275, B2 => n2986, C1 => n3705, C2 => 
                           n2987, A => n3240, ZN => n3239);
   U1264 : AOI22_X1 port map( A1 => n2989, A2 => n3534, B1 => n2990, B2 => 
                           n3535, ZN => n3240);
   U1265 : OAI221_X1 port map( B1 => n2276, B2 => n2991, C1 => n3721, C2 => 
                           n2992, A => n3241, ZN => n3238);
   U1266 : AOI22_X1 port map( A1 => n2994, A2 => n3532, B1 => n2995, B2 => 
                           n3533, ZN => n3241);
   U1267 : OAI221_X1 port map( B1 => n3745, B2 => n2996, C1 => n3737, C2 => 
                           n2997, A => n3242, ZN => n3237);
   U1268 : AOI22_X1 port map( A1 => n2999, A2 => n3530, B1 => n3000, B2 => 
                           n3531, ZN => n3242);
   U1269 : OAI221_X1 port map( B1 => n3761, B2 => n3001, C1 => n3753, C2 => 
                           n3002, A => n3243, ZN => n3236);
   U1270 : AOI22_X1 port map( A1 => n3004, A2 => n3528, B1 => n3005, B2 => 
                           n3529, ZN => n3243);
   U1271 : NOR4_X1 port map( A1 => n3244, A2 => n3245, A3 => n3246, A4 => n3247
                           , ZN => n3216);
   U1272 : OAI221_X1 port map( B1 => n3777, B2 => n3010, C1 => n3769, C2 => 
                           n3011, A => n3248, ZN => n3247);
   U1273 : AOI22_X1 port map( A1 => n3013, A2 => n3542, B1 => n3014, B2 => 
                           n3543, ZN => n3248);
   U1274 : OAI221_X1 port map( B1 => n2195, B2 => n3015, C1 => n2302, C2 => 
                           n3016, A => n3249, ZN => n3246);
   U1275 : AOI22_X1 port map( A1 => n3018, A2 => n3540, B1 => n3019, B2 => 
                           n3541, ZN => n3249);
   U1276 : OAI221_X1 port map( B1 => n2196, B2 => n3020, C1 => n2303, C2 => 
                           n3021, A => n3250, ZN => n3245);
   U1277 : AOI22_X1 port map( A1 => n3023, A2 => n3538, B1 => n3024, B2 => 
                           n3539, ZN => n3250);
   U1278 : OAI221_X1 port map( B1 => n2277, B2 => n3025, C1 => n3817, C2 => 
                           n3026, A => n3251, ZN => n3244);
   U1279 : AOI22_X1 port map( A1 => n3028, A2 => n3536, B1 => n3029, B2 => 
                           n3537, ZN => n3251);
   U1280 : MUX2_X1 port map( A => OUT1_0_port, B => n3252, S => n2929, Z => 
                           n1475);
   U1281 : AND3_X1 port map( A1 => ENABLE, A2 => n2450, A3 => RD1, ZN => n2929)
                           ;
   U1282 : NAND4_X1 port map( A1 => n3253, A2 => n3254, A3 => n3255, A4 => 
                           n3256, ZN => n3252);
   U1283 : NOR4_X1 port map( A1 => n3257, A2 => n3258, A3 => n3259, A4 => n3260
                           , ZN => n3256);
   U1284 : OAI221_X1 port map( B1 => n2278, B2 => n2938, C1 => n3576, C2 => 
                           n2939, A => n3261, ZN => n3260);
   U1285 : AOI22_X1 port map( A1 => n2941, A2 => n3550, B1 => n2942, B2 => 
                           n3551, ZN => n3261);
   U1286 : AND2_X1 port map( A1 => n3262, A2 => n3263, ZN => n2942);
   U1287 : AND2_X1 port map( A1 => n3262, A2 => n3264, ZN => n2941);
   U1288 : NAND2_X1 port map( A1 => n3262, A2 => n3265, ZN => n2939);
   U1289 : NAND2_X1 port map( A1 => n3262, A2 => n3266, ZN => n2938);
   U1290 : AND2_X1 port map( A1 => n3267, A2 => n3268, ZN => n3262);
   U1291 : OAI221_X1 port map( B1 => n2279, B2 => n2943, C1 => n3592, C2 => 
                           n2944, A => n3269, ZN => n3259);
   U1292 : AOI22_X1 port map( A1 => n2946, A2 => n3548, B1 => n2947, B2 => 
                           n3549, ZN => n3269);
   U1293 : AND2_X1 port map( A1 => n3270, A2 => n3263, ZN => n2947);
   U1294 : AND2_X1 port map( A1 => n3270, A2 => n3264, ZN => n2946);
   U1295 : NAND2_X1 port map( A1 => n3270, A2 => n3265, ZN => n2944);
   U1296 : NAND2_X1 port map( A1 => n3270, A2 => n3266, ZN => n2943);
   U1297 : AND2_X1 port map( A1 => n3271, A2 => n3268, ZN => n3270);
   U1298 : OAI221_X1 port map( B1 => n2280, B2 => n2948, C1 => n3608, C2 => 
                           n2949, A => n3272, ZN => n3258);
   U1299 : AOI22_X1 port map( A1 => n2951, A2 => n3546, B1 => n2952, B2 => 
                           n3547, ZN => n3272);
   U1300 : AND2_X1 port map( A1 => n3273, A2 => n3263, ZN => n2952);
   U1301 : AND2_X1 port map( A1 => n3273, A2 => n3264, ZN => n2951);
   U1302 : NAND2_X1 port map( A1 => n3273, A2 => n3265, ZN => n2949);
   U1303 : NAND2_X1 port map( A1 => n3273, A2 => n3266, ZN => n2948);
   U1304 : AND2_X1 port map( A1 => n3274, A2 => n3268, ZN => n3273);
   U1305 : OAI221_X1 port map( B1 => n2281, B2 => n2953, C1 => n3624, C2 => 
                           n2954, A => n3275, ZN => n3257);
   U1306 : AOI22_X1 port map( A1 => n2956, A2 => n3544, B1 => n2957, B2 => 
                           n3545, ZN => n3275);
   U1307 : AND2_X1 port map( A1 => n3263, A2 => n3276, ZN => n2957);
   U1308 : AND2_X1 port map( A1 => n3264, A2 => n3276, ZN => n2956);
   U1309 : NAND2_X1 port map( A1 => n3265, A2 => n3276, ZN => n2954);
   U1310 : NAND2_X1 port map( A1 => n3266, A2 => n3276, ZN => n2953);
   U1311 : AND2_X1 port map( A1 => n3268, A2 => n3277, ZN => n3276);
   U1312 : AND2_X1 port map( A1 => ADD_RD1(5), A2 => ADD_RD1(4), ZN => n3268);
   U1313 : NOR4_X1 port map( A1 => n3278, A2 => n3279, A3 => n3280, A4 => n3281
                           , ZN => n3255);
   U1314 : OAI221_X1 port map( B1 => n2282, B2 => n2962, C1 => n3640, C2 => 
                           n2963, A => n3282, ZN => n3281);
   U1315 : AOI22_X1 port map( A1 => n2965, A2 => n3558, B1 => n2966, B2 => 
                           n3559, ZN => n3282);
   U1316 : AND2_X1 port map( A1 => n3283, A2 => n3263, ZN => n2966);
   U1317 : AND2_X1 port map( A1 => n3283, A2 => n3264, ZN => n2965);
   U1318 : NAND2_X1 port map( A1 => n3283, A2 => n3265, ZN => n2963);
   U1319 : NAND2_X1 port map( A1 => n3283, A2 => n3266, ZN => n2962);
   U1320 : AND2_X1 port map( A1 => n3284, A2 => n3267, ZN => n3283);
   U1321 : OAI221_X1 port map( B1 => n2283, B2 => n2967, C1 => n3656, C2 => 
                           n2968, A => n3285, ZN => n3280);
   U1322 : AOI22_X1 port map( A1 => n2970, A2 => n3556, B1 => n2971, B2 => 
                           n3557, ZN => n3285);
   U1323 : AND2_X1 port map( A1 => n3286, A2 => n3263, ZN => n2971);
   U1324 : AND2_X1 port map( A1 => n3286, A2 => n3264, ZN => n2970);
   U1325 : NAND2_X1 port map( A1 => n3286, A2 => n3265, ZN => n2968);
   U1326 : NAND2_X1 port map( A1 => n3286, A2 => n3266, ZN => n2967);
   U1327 : AND2_X1 port map( A1 => n3284, A2 => n3271, ZN => n3286);
   U1328 : OAI221_X1 port map( B1 => n2284, B2 => n2972, C1 => n3672, C2 => 
                           n2973, A => n3287, ZN => n3279);
   U1329 : AOI22_X1 port map( A1 => n2975, A2 => n3554, B1 => n2976, B2 => 
                           n3555, ZN => n3287);
   U1330 : AND2_X1 port map( A1 => n3288, A2 => n3263, ZN => n2976);
   U1331 : AND2_X1 port map( A1 => n3288, A2 => n3264, ZN => n2975);
   U1332 : NAND2_X1 port map( A1 => n3288, A2 => n3265, ZN => n2973);
   U1333 : NAND2_X1 port map( A1 => n3288, A2 => n3266, ZN => n2972);
   U1334 : AND2_X1 port map( A1 => n3284, A2 => n3274, ZN => n3288);
   U1335 : OAI221_X1 port map( B1 => n2285, B2 => n2977, C1 => n3688, C2 => 
                           n2978, A => n3289, ZN => n3278);
   U1336 : AOI22_X1 port map( A1 => n2980, A2 => n3552, B1 => n2981, B2 => 
                           n3553, ZN => n3289);
   U1337 : AND2_X1 port map( A1 => n3290, A2 => n3263, ZN => n2981);
   U1338 : AND2_X1 port map( A1 => n3290, A2 => n3264, ZN => n2980);
   U1339 : NAND2_X1 port map( A1 => n3290, A2 => n3265, ZN => n2978);
   U1340 : NAND2_X1 port map( A1 => n3290, A2 => n3266, ZN => n2977);
   U1341 : AND2_X1 port map( A1 => n3284, A2 => n3277, ZN => n3290);
   U1342 : AND2_X1 port map( A1 => ADD_RD1(5), A2 => n3291, ZN => n3284);
   U1343 : NOR4_X1 port map( A1 => n3292, A2 => n3293, A3 => n3294, A4 => n3295
                           , ZN => n3254);
   U1344 : OAI221_X1 port map( B1 => n2286, B2 => n2986, C1 => n3704, C2 => 
                           n2987, A => n3296, ZN => n3295);
   U1345 : AOI22_X1 port map( A1 => n2989, A2 => n3566, B1 => n2990, B2 => 
                           n3567, ZN => n3296);
   U1346 : AND2_X1 port map( A1 => n3297, A2 => n3263, ZN => n2990);
   U1347 : AND2_X1 port map( A1 => n3297, A2 => n3264, ZN => n2989);
   U1348 : NAND2_X1 port map( A1 => n3297, A2 => n3265, ZN => n2987);
   U1349 : NAND2_X1 port map( A1 => n3297, A2 => n3266, ZN => n2986);
   U1350 : AND2_X1 port map( A1 => n3298, A2 => n3267, ZN => n3297);
   U1351 : OAI221_X1 port map( B1 => n2287, B2 => n2991, C1 => n3720, C2 => 
                           n2992, A => n3299, ZN => n3294);
   U1352 : AOI22_X1 port map( A1 => n2994, A2 => n3564, B1 => n2995, B2 => 
                           n3565, ZN => n3299);
   U1353 : AND2_X1 port map( A1 => n3300, A2 => n3263, ZN => n2995);
   U1354 : AND2_X1 port map( A1 => n3300, A2 => n3264, ZN => n2994);
   U1355 : NAND2_X1 port map( A1 => n3300, A2 => n3265, ZN => n2992);
   U1356 : NAND2_X1 port map( A1 => n3300, A2 => n3266, ZN => n2991);
   U1357 : AND2_X1 port map( A1 => n3298, A2 => n3271, ZN => n3300);
   U1358 : OAI221_X1 port map( B1 => n3744, B2 => n2996, C1 => n3736, C2 => 
                           n2997, A => n3301, ZN => n3293);
   U1359 : AOI22_X1 port map( A1 => n2999, A2 => n3562, B1 => n3000, B2 => 
                           n3563, ZN => n3301);
   U1360 : AND2_X1 port map( A1 => n3302, A2 => n3263, ZN => n3000);
   U1361 : AND2_X1 port map( A1 => n3302, A2 => n3264, ZN => n2999);
   U1362 : NAND2_X1 port map( A1 => n3302, A2 => n3265, ZN => n2997);
   U1363 : NAND2_X1 port map( A1 => n3302, A2 => n3266, ZN => n2996);
   U1364 : AND2_X1 port map( A1 => n3298, A2 => n3274, ZN => n3302);
   U1365 : OAI221_X1 port map( B1 => n3760, B2 => n3001, C1 => n3752, C2 => 
                           n3002, A => n3303, ZN => n3292);
   U1366 : AOI22_X1 port map( A1 => n3004, A2 => n3560, B1 => n3005, B2 => 
                           n3561, ZN => n3303);
   U1367 : AND2_X1 port map( A1 => n3304, A2 => n3263, ZN => n3005);
   U1368 : AND2_X1 port map( A1 => n3304, A2 => n3264, ZN => n3004);
   U1369 : NAND2_X1 port map( A1 => n3304, A2 => n3265, ZN => n3002);
   U1370 : NAND2_X1 port map( A1 => n3304, A2 => n3266, ZN => n3001);
   U1371 : AND2_X1 port map( A1 => n3298, A2 => n3277, ZN => n3304);
   U1372 : NOR2_X1 port map( A1 => n3291, A2 => ADD_RD1(5), ZN => n3298);
   U1373 : INV_X1 port map( A => ADD_RD1(4), ZN => n3291);
   U1374 : NOR4_X1 port map( A1 => n3305, A2 => n3306, A3 => n3307, A4 => n3308
                           , ZN => n3253);
   U1375 : OAI221_X1 port map( B1 => n3776, B2 => n3010, C1 => n3768, C2 => 
                           n3011, A => n3309, ZN => n3308);
   U1376 : AOI22_X1 port map( A1 => n3013, A2 => n3574, B1 => n3014, B2 => 
                           n3575, ZN => n3309);
   U1377 : AND2_X1 port map( A1 => n3310, A2 => n3263, ZN => n3014);
   U1378 : AND2_X1 port map( A1 => n3310, A2 => n3264, ZN => n3013);
   U1379 : NAND2_X1 port map( A1 => n3310, A2 => n3265, ZN => n3011);
   U1380 : NAND2_X1 port map( A1 => n3310, A2 => n3266, ZN => n3010);
   U1381 : AND2_X1 port map( A1 => n3311, A2 => n3267, ZN => n3310);
   U1382 : AND2_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(2), ZN => n3267);
   U1383 : OAI221_X1 port map( B1 => n2197, B2 => n3015, C1 => n2304, C2 => 
                           n3016, A => n3312, ZN => n3307);
   U1384 : AOI22_X1 port map( A1 => n3018, A2 => n3572, B1 => n3019, B2 => 
                           n3573, ZN => n3312);
   U1385 : AND2_X1 port map( A1 => n3313, A2 => n3263, ZN => n3019);
   U1386 : AND2_X1 port map( A1 => n3313, A2 => n3264, ZN => n3018);
   U1387 : NAND2_X1 port map( A1 => n3313, A2 => n3265, ZN => n3016);
   U1388 : NAND2_X1 port map( A1 => n3313, A2 => n3266, ZN => n3015);
   U1389 : AND2_X1 port map( A1 => n3311, A2 => n3271, ZN => n3313);
   U1390 : AND2_X1 port map( A1 => ADD_RD1(3), A2 => n3314, ZN => n3271);
   U1391 : OAI221_X1 port map( B1 => n2198, B2 => n3020, C1 => n2305, C2 => 
                           n3021, A => n3315, ZN => n3306);
   U1392 : AOI22_X1 port map( A1 => n3023, A2 => n3570, B1 => n3024, B2 => 
                           n3571, ZN => n3315);
   U1393 : AND2_X1 port map( A1 => n3316, A2 => n3263, ZN => n3024);
   U1394 : AND2_X1 port map( A1 => n3316, A2 => n3264, ZN => n3023);
   U1395 : NAND2_X1 port map( A1 => n3316, A2 => n3265, ZN => n3021);
   U1396 : NAND2_X1 port map( A1 => n3316, A2 => n3266, ZN => n3020);
   U1397 : AND2_X1 port map( A1 => n3311, A2 => n3274, ZN => n3316);
   U1398 : NOR2_X1 port map( A1 => n3314, A2 => ADD_RD1(3), ZN => n3274);
   U1399 : INV_X1 port map( A => ADD_RD1(2), ZN => n3314);
   U1400 : OAI221_X1 port map( B1 => n2288, B2 => n3025, C1 => n3816, C2 => 
                           n3026, A => n3317, ZN => n3305);
   U1401 : AOI22_X1 port map( A1 => n3028, A2 => n3568, B1 => n3029, B2 => 
                           n3569, ZN => n3317);
   U1402 : AND2_X1 port map( A1 => n3318, A2 => n3263, ZN => n3029);
   U1403 : AND2_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(1), ZN => n3263);
   U1404 : AND2_X1 port map( A1 => n3318, A2 => n3264, ZN => n3028);
   U1405 : AND2_X1 port map( A1 => ADD_RD1(1), A2 => n3319, ZN => n3264);
   U1406 : NAND2_X1 port map( A1 => n3318, A2 => n3265, ZN => n3026);
   U1407 : INV_X1 port map( A => ADD_RD1(0), ZN => n3319);
   U1408 : NAND2_X1 port map( A1 => n3318, A2 => n3266, ZN => n3025);
   U1409 : AND2_X1 port map( A1 => n3311, A2 => n3277, ZN => n3318);
   U1410 : NOR2_X1 port map( A1 => ADD_RD1(2), A2 => ADD_RD1(3), ZN => n3277);
   U1411 : NOR2_X1 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(5), ZN => n3311);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_WRF_DATA_W8_N_WIN3_N_REG_PER_WIN5_N_GLOBAL_REG5.all;

entity ADDR_DEC_N_GLOBAL_REG5_N_REG_PER_WIN5_N_WIN3_0 is

   port( VIRT_ADDR : in std_logic_vector (4 downto 0);  CWP : in 
         std_logic_vector (5 downto 0);  PHY_ADDR : out std_logic_vector (5 
         downto 0));

end ADDR_DEC_N_GLOBAL_REG5_N_REG_PER_WIN5_N_WIN3_0;

architecture SYN_Behavioural2 of ADDR_DEC_N_GLOBAL_REG5_N_REG_PER_WIN5_N_WIN3_0
   is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component ADDR_DEC_N_GLOBAL_REG5_N_REG_PER_WIN5_N_WIN3_0_DW01_add_0
      port( A, B : in std_logic_vector (5 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (5 downto 0);  CO : out std_logic);
   end component;
   
   signal N6, N7, N8, N9, N10, N31, U3_U1_Z_0, U3_U1_Z_1, U3_U1_Z_2, U3_U1_Z_3,
      U3_U2_Z_5, N16, N15, N14, n42, sub_109_carry_3_port, sub_109_carry_4_port
      , sub_109_carry_5_port, n1, n2, n3, n4, n5, n6_port, n7_port, n8_port, 
      n9_port, n10_port, n11, n12, n13, n14_port, n15_port, n16_port, n17, n18,
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n35, n36, n37, n38
      , n39, n_1286 : std_logic;

begin
   
   n42 <= '0';
   r21 : ADDR_DEC_N_GLOBAL_REG5_N_REG_PER_WIN5_N_WIN3_0_DW01_add_0 port map( 
                           A(5) => n42, A(4) => n9_port, A(3) => U3_U1_Z_3, 
                           A(2) => U3_U1_Z_2, A(1) => U3_U1_Z_1, A(0) => 
                           U3_U1_Z_0, B(5) => U3_U2_Z_5, B(4) => n38, B(3) => 
                           n37, B(2) => n39, B(1) => n36, B(0) => n35, CI => 
                           n42, SUM(5) => N10, SUM(4) => N9, SUM(3) => N8, 
                           SUM(2) => N7, SUM(1) => N6, SUM(0) => PHY_ADDR(0), 
                           CO => n_1286);
   U3 : XOR2_X1 port map( A => n29, B => sub_109_carry_5_port, Z => n1);
   U4 : XOR2_X1 port map( A => N9, B => n6_port, Z => n2);
   U5 : XOR2_X1 port map( A => N10, B => n8_port, Z => N31);
   U6 : NAND2_X1 port map( A1 => N9, A2 => n6_port, ZN => n8_port);
   U7 : XOR2_X1 port map( A => N7, B => N6, Z => n3);
   U8 : XOR2_X1 port map( A => N8, B => n5, Z => n4);
   U9 : XNOR2_X1 port map( A => n27, B => sub_109_carry_3_port, ZN => N15);
   U10 : XNOR2_X1 port map( A => n25, B => n28, ZN => N14);
   U11 : OR2_X1 port map( A1 => n25, A2 => n28, ZN => sub_109_carry_3_port);
   U12 : OR2_X1 port map( A1 => n27, A2 => sub_109_carry_3_port, ZN => 
                           sub_109_carry_4_port);
   U13 : XNOR2_X1 port map( A => n26, B => sub_109_carry_4_port, ZN => N16);
   U14 : AND2_X1 port map( A1 => N7, A2 => N6, ZN => n5);
   U15 : AND2_X1 port map( A1 => N8, A2 => n5, ZN => n6_port);
   U17 : NAND2_X1 port map( A1 => CWP(4), A2 => n7_port, ZN => 
                           sub_109_carry_5_port);
   U18 : INV_X1 port map( A => sub_109_carry_4_port, ZN => n7_port);
   U19 : INV_X1 port map( A => CWP(3), ZN => n27);
   U20 : INV_X1 port map( A => CWP(2), ZN => n25);
   U21 : MUX2_X1 port map( A => N10, B => N31, S => n10_port, Z => PHY_ADDR(5))
                           ;
   U22 : MUX2_X1 port map( A => N9, B => n2, S => n10_port, Z => PHY_ADDR(4));
   U23 : MUX2_X1 port map( A => N8, B => n4, S => n10_port, Z => PHY_ADDR(3));
   U24 : MUX2_X1 port map( A => N7, B => n3, S => n10_port, Z => PHY_ADDR(2));
   U25 : XOR2_X1 port map( A => N6, B => n10_port, Z => PHY_ADDR(1));
   U26 : AOI211_X1 port map( C1 => n11, C2 => N15, A => n12, B => n13, ZN => 
                           n10_port);
   U27 : OR3_X1 port map( A1 => n14_port, A2 => n1, A3 => N16, ZN => n13);
   U28 : INV_X1 port map( A => n15_port, ZN => n14_port);
   U29 : OAI221_X1 port map( B1 => n11, B2 => N15, C1 => n16_port, C2 => N14, A
                           => n17, ZN => n15_port);
   U30 : INV_X1 port map( A => n18, ZN => n17);
   U31 : AOI221_X1 port map( B1 => N14, B2 => n16_port, C1 => n19, C2 => n20, A
                           => n21, ZN => n18);
   U32 : AOI21_X1 port map( B1 => CWP(0), B2 => VIRT_ADDR(0), A => n28, ZN => 
                           n21);
   U33 : NAND3_X1 port map( A1 => VIRT_ADDR(0), A2 => n28, A3 => CWP(0), ZN => 
                           n19);
   U34 : INV_X1 port map( A => CWP(1), ZN => n28);
   U35 : MUX2_X1 port map( A => VIRT_ADDR(0), B => CWP(0), S => n22, Z => n35);
   U36 : MUX2_X1 port map( A => VIRT_ADDR(1), B => CWP(1), S => n22, Z => n36);
   U37 : MUX2_X1 port map( A => VIRT_ADDR(3), B => CWP(3), S => n22, Z => n37);
   U38 : OAI21_X1 port map( B1 => n26, B2 => n12, A => n23, ZN => n38);
   U39 : INV_X1 port map( A => CWP(4), ZN => n26);
   U40 : MUX2_X1 port map( A => VIRT_ADDR(2), B => CWP(2), S => n22, Z => n39);
   U41 : NOR2_X1 port map( A1 => n29, A2 => n12, ZN => U3_U2_Z_5);
   U42 : INV_X1 port map( A => CWP(5), ZN => n29);
   n9_port <= '0';
   U44 : NAND2_X1 port map( A1 => n22, A2 => n11, ZN => U3_U1_Z_3);
   U45 : INV_X1 port map( A => VIRT_ADDR(3), ZN => n11);
   U46 : NAND2_X1 port map( A1 => n22, A2 => n16_port, ZN => U3_U1_Z_2);
   U47 : INV_X1 port map( A => VIRT_ADDR(2), ZN => n16_port);
   U48 : NAND2_X1 port map( A1 => n22, A2 => n20, ZN => U3_U1_Z_1);
   U49 : INV_X1 port map( A => VIRT_ADDR(1), ZN => n20);
   U50 : INV_X1 port map( A => n12, ZN => n22);
   U51 : OR2_X1 port map( A1 => n12, A2 => VIRT_ADDR(0), ZN => U3_U1_Z_0);
   U52 : NAND2_X1 port map( A1 => n23, A2 => n24, ZN => n12);
   U53 : NAND4_X1 port map( A1 => VIRT_ADDR(0), A2 => VIRT_ADDR(1), A3 => 
                           VIRT_ADDR(2), A4 => VIRT_ADDR(3), ZN => n24);
   U54 : INV_X1 port map( A => VIRT_ADDR(4), ZN => n23);

end SYN_Behavioural2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_WRF_DATA_W8_N_WIN3_N_REG_PER_WIN5_N_GLOBAL_REG5.all;

entity WRF_CU_N_GLOBAL_REG5_N_REG_PER_WIN5_N_WIN3 is

   port( CLK, RESET, TRNSF_CPLT_ACK : in std_logic;  OP : in std_logic_vector 
         (0 to 1);  STATE : out std_logic_vector (0 to 1);  CWP, SWP : out 
         std_logic_vector (5 downto 0));

end WRF_CU_N_GLOBAL_REG5_N_REG_PER_WIN5_N_WIN3;

architecture SYN_Behavioural of WRF_CU_N_GLOBAL_REG5_N_REG_PER_WIN5_N_WIN3 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal X_Logic0_port, CWP_4_port, CWP_3_port, CWP_2_port, CWP_1_port, 
      CWP_0_port, SWP_4_port, SWP_3_port, SWP_2_port, SWP_1_port, 
      wrf_cu_cur_state_2_port, wrf_cu_cur_state_1_port, wrf_cu_cur_state_0_port
      , wrf_cu_fut_state_1_port, N66, N96, N132, N133, N134, U3_U1_Z_1, 
      U3_U1_Z_2, U3_U1_Z_3, U3_U1_Z_4, n32, n33, n34, n35, n36, n38, n39, n40, 
      n41, n92, n93, n94, n95, n96_port, n97, n98, n100, n101, n102, n103, n105
      , r34_carry_1_port, r34_carry_2_port, r34_carry_3_port, r34_carry_4_port,
      n85, n83, n84, n86, n87, n88, n89, n90, n91, n99, n104, n106, n107, n108,
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, 
      n132_port, n133_port, n134_port, n135, n136, n137, n138, n139, n140, n141
      , n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
      n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, STATE_0_port,
      n165, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293 : std_logic;

begin
   STATE <= ( N66, STATE_0_port );
   CWP <= ( X_Logic0_port, CWP_4_port, CWP_3_port, CWP_2_port, CWP_1_port, 
      CWP_0_port );
   SWP <= ( X_Logic0_port, SWP_4_port, SWP_3_port, SWP_2_port, SWP_1_port, N96 
      );
   
   X_Logic0_port <= '0';
   spill_cntr_reg_0_inst : DFFS_X1 port map( D => n105, CK => CLK, SN => n165, 
                           Q => n_1287, QN => n161);
   wrf_cu_cur_state_reg_1_inst : DFFR_X1 port map( D => wrf_cu_fut_state_1_port
                           , CK => CLK, RN => n165, Q => 
                           wrf_cu_cur_state_1_port, QN => n84);
   fill_cntr_reg_0_inst : DFFR_X1 port map( D => n93, CK => CLK, RN => n165, Q 
                           => n_1288, QN => n160);
   wrf_cu_cur_state_reg_2_inst : DFFR_X1 port map( D => n163, CK => CLK, RN => 
                           n165, Q => wrf_cu_cur_state_2_port, QN => n83);
   wrf_cu_cur_state_reg_0_inst : DFFR_X1 port map( D => n85, CK => CLK, RN => 
                           n165, Q => wrf_cu_cur_state_0_port, QN => n_1289);
   cwp_cntr_reg_1_inst : DFFR_X1 port map( D => n98, CK => CLK, RN => n165, Q 
                           => CWP_1_port, QN => n35);
   cwp_cntr_reg_3_inst : DFFR_X1 port map( D => n96_port, CK => CLK, RN => n165
                           , Q => CWP_3_port, QN => n33);
   cwp_cntr_reg_4_inst : DFFR_X1 port map( D => n95, CK => CLK, RN => n165, Q 
                           => CWP_4_port, QN => n32);
   cwp_cntr_reg_2_inst : DFFR_X1 port map( D => n97, CK => CLK, RN => n165, Q 
                           => CWP_2_port, QN => n34);
   swp_cntr_reg_4_inst : DFFR_X1 port map( D => n100, CK => CLK, RN => n165, Q 
                           => SWP_4_port, QN => n38);
   swp_cntr_reg_2_inst : DFFR_X1 port map( D => n102, CK => CLK, RN => n165, Q 
                           => SWP_2_port, QN => n40);
   swp_cntr_reg_1_inst : DFFR_X1 port map( D => n103, CK => CLK, RN => n165, Q 
                           => SWP_1_port, QN => n41);
   swp_cntr_reg_3_inst : DFFR_X1 port map( D => n101, CK => CLK, RN => n165, Q 
                           => SWP_3_port, QN => n39);
   fill_cntr_reg_1_inst : DFFS_X1 port map( D => n92, CK => CLK, SN => n165, Q 
                           => n_1290, QN => n159);
   spill_cntr_reg_1_inst : DFFR_X1 port map( D => n94, CK => CLK, RN => n165, Q
                           => n_1291, QN => n158);
   r34_U1_1 : FA_X1 port map( A => U3_U1_Z_1, B => n162, CI => r34_carry_1_port
                           , CO => r34_carry_2_port, S => n_1292);
   r34_U1_2 : FA_X1 port map( A => U3_U1_Z_2, B => r34_carry_1_port, CI => 
                           r34_carry_2_port, CO => r34_carry_3_port, S => N132)
                           ;
   r34_U1_3 : FA_X1 port map( A => U3_U1_Z_3, B => n162, CI => r34_carry_3_port
                           , CO => r34_carry_4_port, S => N133);
   r34_U1_4 : FA_X1 port map( A => U3_U1_Z_4, B => r34_carry_1_port, CI => 
                           r34_carry_4_port, CO => n_1293, S => N134);
   U3 : NAND3_X1 port map( A1 => n35, A2 => n33, A3 => n36, ZN => n151);
   U4 : NOR4_X1 port map( A1 => n149, A2 => SWP_3_port, A3 => n38, A4 => n40, 
                           ZN => n148);
   U5 : INV_X2 port map( A => SWP_1_port, ZN => n157);
   n149 <= '0';
   N96 <= '0';
   CWP_0_port <= '0';
   n36 <= '1';
   U10 : INV_X1 port map( A => n162, ZN => r34_carry_1_port);
   U11 : NOR2_X1 port map( A1 => n86, A2 => n87, ZN => n162);
   U12 : INV_X1 port map( A => RESET, ZN => n165);
   U13 : OAI22_X1 port map( A1 => U3_U1_Z_1, A2 => n88, B1 => n35, B2 => n89, 
                           ZN => n98);
   U14 : OAI221_X1 port map( B1 => n90, B2 => n91, C1 => n34, C2 => n89, A => 
                           n99, ZN => n97);
   U15 : INV_X1 port map( A => N132, ZN => n91);
   U16 : OAI22_X1 port map( A1 => n88, A2 => n104, B1 => n33, B2 => n89, ZN => 
                           n96_port);
   U17 : OAI221_X1 port map( B1 => n90, B2 => n106, C1 => n32, C2 => n89, A => 
                           n99, ZN => n95);
   U18 : NAND4_X1 port map( A1 => n107, A2 => n85, A3 => n32, A4 => n108, ZN =>
                           n99);
   U19 : AND2_X1 port map( A1 => n34, A2 => n163, ZN => n108);
   U20 : AOI21_X1 port map( B1 => n109, B2 => n110, A => n111, ZN => n89);
   U21 : INV_X1 port map( A => N134, ZN => n106);
   U22 : AOI21_X1 port map( B1 => n85, B2 => n163, A => n112, ZN => n90);
   U23 : OAI22_X1 port map( A1 => n161, A2 => n113, B1 => n158, B2 => n114, ZN 
                           => n94);
   U24 : OAI22_X1 port map( A1 => n159, A2 => n113, B1 => n160, B2 => n114, ZN 
                           => n93);
   U25 : OAI221_X1 port map( B1 => n159, B2 => n114, C1 => n160, C2 => n113, A 
                           => n115, ZN => n92);
   U26 : OAI221_X1 port map( B1 => n161, B2 => n114, C1 => n158, C2 => n113, A 
                           => n115, ZN => n105);
   U27 : NAND3_X1 port map( A1 => n116, A2 => STATE_0_port, A3 => n110, ZN => 
                           n113);
   U28 : INV_X1 port map( A => n117, ZN => n110);
   U29 : NOR3_X1 port map( A1 => n118, A2 => n119, A3 => n111, ZN => n114);
   U30 : OAI21_X1 port map( B1 => U3_U1_Z_1, B2 => n122, A => n123, ZN => n103)
                           ;
   U31 : INV_X1 port map( A => n124, ZN => n123);
   U32 : MUX2_X1 port map( A => n120, B => n121, S => n41, Z => n124);
   U33 : NAND2_X1 port map( A1 => n125, A2 => n126, ZN => n102);
   U34 : OAI21_X1 port map( B1 => n127, B2 => N132, A => n128, ZN => n126);
   U35 : MUX2_X1 port map( A => n129, B => n130, S => n40, Z => n125);
   U36 : NAND2_X1 port map( A1 => n121, A2 => SWP_1_port, ZN => n130);
   U37 : AOI21_X1 port map( B1 => n121, B2 => n41, A => n120, ZN => n129);
   U38 : OAI221_X1 port map( B1 => n39, B2 => n131, C1 => n122, C2 => n104, A 
                           => n132_port, ZN => n101);
   U39 : INV_X1 port map( A => n133_port, ZN => n132_port);
   U40 : INV_X1 port map( A => N133, ZN => n104);
   U41 : NOR2_X1 port map( A1 => n134_port, A2 => n120, ZN => n131);
   U42 : NOR3_X1 port map( A1 => n135, A2 => n41, A3 => n40, ZN => n134_port);
   U43 : NAND2_X1 port map( A1 => n136, A2 => n137, ZN => n100);
   U44 : OAI21_X1 port map( B1 => n127, B2 => N134, A => n128, ZN => n137);
   U45 : INV_X1 port map( A => n138, ZN => n128);
   U46 : MUX2_X1 port map( A => n139, B => n140, S => n38, Z => n136);
   U47 : NAND2_X1 port map( A1 => n121, A2 => n141, ZN => n140);
   U48 : NOR2_X1 port map( A1 => n133_port, A2 => n120, ZN => n139);
   U49 : NAND2_X1 port map( A1 => n117, A2 => n142, ZN => n120);
   U50 : NAND3_X1 port map( A1 => n143, A2 => n138, A3 => n111, ZN => n142);
   U51 : INV_X1 port map( A => n144, ZN => n111);
   U52 : NAND2_X1 port map( A1 => n144, A2 => n115, ZN => n117);
   U53 : OR3_X1 port map( A1 => n85, A2 => wrf_cu_fut_state_1_port, A3 => n163,
                           ZN => n115);
   U54 : NAND2_X1 port map( A1 => wrf_cu_fut_state_1_port, A2 => n85, ZN => 
                           n144);
   U55 : NAND3_X1 port map( A1 => n116, A2 => n138, A3 => n145, ZN => 
                           wrf_cu_fut_state_1_port);
   U56 : MUX2_X1 port map( A => n146, B => wrf_cu_cur_state_1_port, S => 
                           wrf_cu_cur_state_2_port, Z => n145);
   U57 : OR3_X1 port map( A1 => n147, A2 => OP(0), A3 => n84, ZN => n146);
   U58 : INV_X1 port map( A => n118, ZN => n116);
   U59 : NOR2_X1 port map( A1 => n141, A2 => n135, ZN => n133_port);
   U60 : INV_X1 port map( A => n121, ZN => n135);
   U61 : NOR2_X1 port map( A1 => n143, A2 => n148, ZN => n121);
   U62 : OAI21_X1 port map( B1 => n41, B2 => n40, A => n39, ZN => n141);
   U63 : OAI22_X1 port map( A1 => n38, A2 => n122, B1 => n32, B2 => n88, ZN => 
                           U3_U1_Z_4);
   U64 : OAI22_X1 port map( A1 => n39, A2 => n122, B1 => n33, B2 => n88, ZN => 
                           U3_U1_Z_3);
   U65 : OAI22_X1 port map( A1 => n40, A2 => n122, B1 => n34, B2 => n88, ZN => 
                           U3_U1_Z_2);
   U66 : OAI22_X1 port map( A1 => n41, A2 => n122, B1 => n35, B2 => n88, ZN => 
                           U3_U1_Z_1);
   U67 : NOR2_X1 port map( A1 => n112, A2 => n87, ZN => n88);
   U68 : AND3_X1 port map( A1 => n150, A2 => n85, A3 => n163, ZN => n87);
   U69 : INV_X1 port map( A => n109, ZN => n163);
   U70 : NAND3_X1 port map( A1 => n32, A2 => n107, A3 => n34, ZN => n150);
   U71 : INV_X1 port map( A => n151, ZN => n107);
   U72 : NOR3_X1 port map( A1 => n152, A2 => n85, A3 => n109, ZN => n112);
   U73 : NAND4_X1 port map( A1 => n153, A2 => wrf_cu_cur_state_1_port, A3 => 
                           wrf_cu_cur_state_0_port, A4 => n83, ZN => n109);
   U74 : MUX2_X1 port map( A => n147, B => n154, S => OP(0), Z => n153);
   U75 : NOR2_X1 port map( A1 => OP(1), A2 => n160, ZN => n154);
   U76 : NOR2_X1 port map( A1 => n155, A2 => n161, ZN => n147);
   U77 : NAND3_X1 port map( A1 => n156, A2 => n143, A3 => 
                           wrf_cu_cur_state_1_port, ZN => n85);
   U78 : NAND3_X1 port map( A1 => wrf_cu_cur_state_1_port, A2 => TRNSF_CPLT_ACK
                           , A3 => n118, ZN => n143);
   U79 : NOR2_X1 port map( A1 => wrf_cu_cur_state_2_port, A2 => 
                           wrf_cu_cur_state_0_port, ZN => n118);
   U80 : NAND3_X1 port map( A1 => n155, A2 => n83, A3 => 
                           wrf_cu_cur_state_0_port, ZN => n156);
   U81 : INV_X1 port map( A => OP(1), ZN => n155);
   U82 : NOR3_X1 port map( A1 => n32, A2 => n34, A3 => n151, ZN => n152);
   U83 : INV_X1 port map( A => n86, ZN => n122);
   U84 : NOR2_X1 port map( A1 => n138, A2 => n127, ZN => n86);
   U85 : AND4_X1 port map( A1 => n39, A2 => n38, A3 => n40, A4 => n157, ZN => 
                           n127);
   U86 : NAND3_X1 port map( A1 => TRNSF_CPLT_ACK, A2 => n119, A3 => 
                           wrf_cu_cur_state_0_port, ZN => n138);
   U87 : MUX2_X1 port map( A => wrf_cu_cur_state_1_port, B => n119, S => 
                           wrf_cu_cur_state_0_port, Z => N66);
   U88 : INV_X1 port map( A => STATE_0_port, ZN => n119);
   U89 : NAND2_X1 port map( A1 => n84, A2 => n83, ZN => STATE_0_port);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_WRF_DATA_W8_N_WIN3_N_REG_PER_WIN5_N_GLOBAL_REG5.all;

entity WRF_DATA_W8_N_WIN3_N_REG_PER_WIN5_N_GLOBAL_REG5 is

   port( CLK, RESET, ENABLE, RD1_EN, RD2_EN, WR_EN : in std_logic;  WADDR, 
         RADDR1, RADDR2 : in std_logic_vector (4 downto 0);  DIN : in 
         std_logic_vector (7 downto 0);  DOUT1, DOUT2 : out std_logic_vector (7
         downto 0);  TRNSF_CPLT_ACK : in std_logic;  OP : in wrf_op;  STATE : 
         out wrf_state;  CWP, SWP : out std_logic_vector (5 downto 0));

end WRF_DATA_W8_N_WIN3_N_REG_PER_WIN5_N_GLOBAL_REG5;

architecture SYN_Behavioural of WRF_DATA_W8_N_WIN3_N_REG_PER_WIN5_N_GLOBAL_REG5
   is

   component RF_ADDR_W6_DATA_W8
      port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
            ADD_RD2 : in std_logic_vector (5 downto 0);  DATAIN : in 
            std_logic_vector (7 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (7 downto 0));
   end component;
   
   component ADDR_DEC_N_GLOBAL_REG5_N_REG_PER_WIN5_N_WIN3_1
      port( VIRT_ADDR : in std_logic_vector (4 downto 0);  CWP : in 
            std_logic_vector (5 downto 0);  PHY_ADDR : out std_logic_vector (5 
            downto 0));
   end component;
   
   component ADDR_DEC_N_GLOBAL_REG5_N_REG_PER_WIN5_N_WIN3_2
      port( VIRT_ADDR : in std_logic_vector (4 downto 0);  CWP : in 
            std_logic_vector (5 downto 0);  PHY_ADDR : out std_logic_vector (5 
            downto 0));
   end component;
   
   component ADDR_DEC_N_GLOBAL_REG5_N_REG_PER_WIN5_N_WIN3_0
      port( VIRT_ADDR : in std_logic_vector (4 downto 0);  CWP : in 
            std_logic_vector (5 downto 0);  PHY_ADDR : out std_logic_vector (5 
            downto 0));
   end component;
   
   component WRF_CU_N_GLOBAL_REG5_N_REG_PER_WIN5_N_WIN3
      port( CLK, RESET, TRNSF_CPLT_ACK : in std_logic;  OP : in 
            std_logic_vector (0 to 1);  STATE : out std_logic_vector (0 to 1); 
            CWP, SWP : out std_logic_vector (5 downto 0));
   end component;
   
   signal OP_1_port, OP_0_port, STATE_1_port, STATE_0_port, CWP_5_port, 
      CWP_4_port, CWP_3_port, CWP_2_port, CWP_1_port, SWP_5_port, SWP_4_port, 
      SWP_3_port, SWP_2_port, SWP_1_port, waddr_phys_5_port, waddr_phys_4_port,
      waddr_phys_3_port, waddr_phys_2_port, waddr_phys_1_port, 
      waddr_phys_0_port, raddr1_phys_5_port, raddr1_phys_4_port, 
      raddr1_phys_3_port, raddr1_phys_2_port, raddr1_phys_1_port, 
      raddr1_phys_0_port, raddr2_phys_5_port, raddr2_phys_4_port, 
      raddr2_phys_3_port, raddr2_phys_2_port, raddr2_phys_1_port, 
      raddr2_phys_0_port, SWP_0_port, n_1294, n_1295, n_1296, n_1297 : 
      std_logic;
   
   signal STATE_pin : std_logic_vector (0 to 1);

begin
   (OP_1_port, OP_0_port) <= wrf_op_to_std_logic_vector(OP);
   STATE <= std_logic_vector_to_wrf_state((STATE_1_port, STATE_0_port));
   CWP <= ( CWP_5_port, CWP_4_port, CWP_3_port, CWP_2_port, CWP_1_port, 
      SWP_0_port );
   SWP <= ( SWP_5_port, SWP_4_port, SWP_3_port, SWP_2_port, SWP_1_port, 
      SWP_0_port );
   
   ( STATE_1_port, STATE_0_port ) <= STATE_pin;
   U_WRF_CU : WRF_CU_N_GLOBAL_REG5_N_REG_PER_WIN5_N_WIN3 port map( CLK => CLK, 
      RESET => RESET, TRNSF_CPLT_ACK => TRNSF_CPLT_ACK, OP(0) => OP_1_port, 
      OP(1) => OP_0_port, STATE => STATE_pin, CWP(5) => n_1294, CWP(4) => 
      CWP_4_port, CWP(3) => CWP_3_port, CWP(2) => CWP_2_port, CWP(1) => 
      CWP_1_port, CWP(0) => n_1295, SWP(5) => n_1296, SWP(4) => SWP_4_port, 
      SWP(3) => SWP_3_port, SWP(2) => SWP_2_port, SWP(1) => SWP_1_port, SWP(0) 
      => n_1297);
   U_ADDR_DEC_WADDR : ADDR_DEC_N_GLOBAL_REG5_N_REG_PER_WIN5_N_WIN3_0 port map( 
                           VIRT_ADDR(4) => WADDR(4), VIRT_ADDR(3) => WADDR(3), 
                           VIRT_ADDR(2) => WADDR(2), VIRT_ADDR(1) => WADDR(1), 
                           VIRT_ADDR(0) => WADDR(0), CWP(5) => CWP_5_port, 
                           CWP(4) => CWP_4_port, CWP(3) => CWP_3_port, CWP(2) 
                           => CWP_2_port, CWP(1) => CWP_1_port, CWP(0) => 
                           SWP_0_port, PHY_ADDR(5) => waddr_phys_5_port, 
                           PHY_ADDR(4) => waddr_phys_4_port, PHY_ADDR(3) => 
                           waddr_phys_3_port, PHY_ADDR(2) => waddr_phys_2_port,
                           PHY_ADDR(1) => waddr_phys_1_port, PHY_ADDR(0) => 
                           waddr_phys_0_port);
   U_ADDR_DEC_RADDR1 : ADDR_DEC_N_GLOBAL_REG5_N_REG_PER_WIN5_N_WIN3_2 port map(
                           VIRT_ADDR(4) => RADDR1(4), VIRT_ADDR(3) => RADDR1(3)
                           , VIRT_ADDR(2) => RADDR1(2), VIRT_ADDR(1) => 
                           RADDR1(1), VIRT_ADDR(0) => RADDR1(0), CWP(5) => 
                           CWP_5_port, CWP(4) => CWP_4_port, CWP(3) => 
                           CWP_3_port, CWP(2) => CWP_2_port, CWP(1) => 
                           CWP_1_port, CWP(0) => SWP_0_port, PHY_ADDR(5) => 
                           raddr1_phys_5_port, PHY_ADDR(4) => 
                           raddr1_phys_4_port, PHY_ADDR(3) => 
                           raddr1_phys_3_port, PHY_ADDR(2) => 
                           raddr1_phys_2_port, PHY_ADDR(1) => 
                           raddr1_phys_1_port, PHY_ADDR(0) => 
                           raddr1_phys_0_port);
   U_ADDR_DEC_RADDR2 : ADDR_DEC_N_GLOBAL_REG5_N_REG_PER_WIN5_N_WIN3_1 port map(
                           VIRT_ADDR(4) => RADDR2(4), VIRT_ADDR(3) => RADDR2(3)
                           , VIRT_ADDR(2) => RADDR2(2), VIRT_ADDR(1) => 
                           RADDR2(1), VIRT_ADDR(0) => RADDR2(0), CWP(5) => 
                           CWP_5_port, CWP(4) => CWP_4_port, CWP(3) => 
                           CWP_3_port, CWP(2) => CWP_2_port, CWP(1) => 
                           CWP_1_port, CWP(0) => SWP_0_port, PHY_ADDR(5) => 
                           raddr2_phys_5_port, PHY_ADDR(4) => 
                           raddr2_phys_4_port, PHY_ADDR(3) => 
                           raddr2_phys_3_port, PHY_ADDR(2) => 
                           raddr2_phys_2_port, PHY_ADDR(1) => 
                           raddr2_phys_1_port, PHY_ADDR(0) => 
                           raddr2_phys_0_port);
   U_RF : RF_ADDR_W6_DATA_W8 port map( CLK => CLK, RESET => RESET, ENABLE => 
                           ENABLE, RD1 => RD1_EN, RD2 => RD2_EN, WR => WR_EN, 
                           ADD_WR(5) => waddr_phys_5_port, ADD_WR(4) => 
                           waddr_phys_4_port, ADD_WR(3) => waddr_phys_3_port, 
                           ADD_WR(2) => waddr_phys_2_port, ADD_WR(1) => 
                           waddr_phys_1_port, ADD_WR(0) => waddr_phys_0_port, 
                           ADD_RD1(5) => raddr1_phys_5_port, ADD_RD1(4) => 
                           raddr1_phys_4_port, ADD_RD1(3) => raddr1_phys_3_port
                           , ADD_RD1(2) => raddr1_phys_2_port, ADD_RD1(1) => 
                           raddr1_phys_1_port, ADD_RD1(0) => raddr1_phys_0_port
                           , ADD_RD2(5) => raddr2_phys_5_port, ADD_RD2(4) => 
                           raddr2_phys_4_port, ADD_RD2(3) => raddr2_phys_3_port
                           , ADD_RD2(2) => raddr2_phys_2_port, ADD_RD2(1) => 
                           raddr2_phys_1_port, ADD_RD2(0) => raddr2_phys_0_port
                           , DATAIN(7) => DIN(7), DATAIN(6) => DIN(6), 
                           DATAIN(5) => DIN(5), DATAIN(4) => DIN(4), DATAIN(3) 
                           => DIN(3), DATAIN(2) => DIN(2), DATAIN(1) => DIN(1),
                           DATAIN(0) => DIN(0), OUT1(7) => DOUT1(7), OUT1(6) =>
                           DOUT1(6), OUT1(5) => DOUT1(5), OUT1(4) => DOUT1(4), 
                           OUT1(3) => DOUT1(3), OUT1(2) => DOUT1(2), OUT1(1) =>
                           DOUT1(1), OUT1(0) => DOUT1(0), OUT2(7) => DOUT2(7), 
                           OUT2(6) => DOUT2(6), OUT2(5) => DOUT2(5), OUT2(4) =>
                           DOUT2(4), OUT2(3) => DOUT2(3), OUT2(2) => DOUT2(2), 
                           OUT2(1) => DOUT2(1), OUT2(0) => DOUT2(0));
   SWP_0_port <= '0';
   SWP_5_port <= '0';
   CWP_5_port <= '0';

end SYN_Behavioural;
