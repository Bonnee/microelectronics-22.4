LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_unsigned.ALL;

ENTITY TBSUM_GENERATOR IS
END TBSUM_GENERATOR;

ARCHITECTURE TEST OF TBSUM_GENERATOR IS
	CONSTANT BIT_PER_BLOCK : INTEGER := 3;
	CONSTANT BLOCKS : INTEGER := 2;

	COMPONENT SUM_GENERATOR IS
		GENERIC (
			NBIT_PER_BLOCK : INTEGER;
			NBLOCKS : INTEGER);
		PORT (
			A : IN STD_LOGIC_VECTOR((NBIT_PER_BLOCK * NBLOCKS) - 1 DOWNTO 0);
			B : IN STD_LOGIC_VECTOR((NBIT_PER_BLOCK * NBLOCKS) - 1 DOWNTO 0);
			Ci : IN STD_LOGIC_VECTOR(NBLOCKS - 1 DOWNTO 0);
			S : OUT STD_LOGIC_VECTOR((NBIT_PER_BLOCK * NBLOCKS) - 1 DOWNTO 0));
	END COMPONENT;

	SIGNAL A : STD_LOGIC_VECTOR((BIT_PER_BLOCK * BLOCKS) - 1 DOWNTO 0);
	SIGNAL B : STD_LOGIC_VECTOR((BIT_PER_BLOCK * BLOCKS) - 1 DOWNTO 0);
	SIGNAL Ci : STD_LOGIC_VECTOR(BLOCKS - 1 DOWNTO 0);
	SIGNAL S : STD_LOGIC_VECTOR((BIT_PER_BLOCK * BLOCKS) - 1 DOWNTO 0);

BEGIN

	SUM_GEN : SUM_GENERATOR
	GENERIC MAP(NBIT_PER_BLOCK => BIT_PER_BLOCK, NBLOCKS => BLOCKS)
	PORT MAP(A => A, B => B, Ci => Ci, S => S);

	A <= "000000", "000001" AFTER 0.5 ns, "000010" AFTER 1 ns, "111110" AFTER 1.5 ns, "111111" AFTER 2 ns;
	B <= "000000", "000000" AFTER 0.5 ns, "111010" AFTER 1 ns, "000001" AFTER 1.5 ns, "000001" AFTER 2 ns;
	Ci <= "00",  "00"   AFTER 0.5 ns, "01"   AFTER 1 ns, "10"   AFTER 1.5 ns, "11"   AFTER 2 ns;

END TEST;

CONFIGURATION SUM_GENERATORTEST OF TBSUM_GENERATOR IS
	FOR TEST
		FOR ALL : SUM_GENERATOR
			USE CONFIGURATION WORK.CFG_SUM_GENERATOR_STRUCTURAL;
		END FOR;
	END FOR;
END SUM_GENERATORTEST;
