PACKAGE CONSTANTS IS
   CONSTANT NumBit : INTEGER := 4;
END CONSTANTS;