
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_BOOTHMUL_NBIT32_1 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_BOOTHMUL_NBIT32_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity RCA_NBIT64_16_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_NBIT64_16_DW01_add_0;

architecture SYN_rpl of RCA_NBIT64_16_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_63_port, carry_62_port, carry_61_port, carry_60_port, 
      carry_59_port, carry_58_port, carry_57_port, carry_56_port, carry_55_port
      , carry_54_port, carry_53_port, carry_52_port, carry_51_port, 
      carry_50_port, carry_49_port, carry_48_port, carry_47_port, carry_46_port
      , carry_45_port, carry_44_port, carry_43_port, carry_42_port, 
      carry_41_port, carry_40_port, carry_39_port, carry_38_port, carry_37_port
      , carry_36_port, carry_35_port, carry_34_port, carry_33_port, 
      carry_32_port, carry_31_port, carry_30_port, carry_29_port, carry_28_port
      , carry_27_port, carry_26_port, carry_25_port, carry_24_port, 
      carry_23_port, carry_22_port, carry_21_port, carry_20_port, carry_19_port
      , carry_18_port, carry_17_port, carry_16_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_10_port
      , carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1_61 : FA_X1 port map( A => A(61), B => B(61), CI => carry_61_port, CO => 
                           carry_62_port, S => SUM(61));
   U1_60 : FA_X1 port map( A => A(60), B => B(60), CI => carry_60_port, CO => 
                           carry_61_port, S => SUM(60));
   U1_59 : FA_X1 port map( A => A(59), B => B(59), CI => carry_59_port, CO => 
                           carry_60_port, S => SUM(59));
   U1_58 : FA_X1 port map( A => A(58), B => B(58), CI => carry_58_port, CO => 
                           carry_59_port, S => SUM(58));
   U1_57 : FA_X1 port map( A => A(57), B => B(57), CI => carry_57_port, CO => 
                           carry_58_port, S => SUM(57));
   U1_56 : FA_X1 port map( A => A(56), B => B(56), CI => carry_56_port, CO => 
                           carry_57_port, S => SUM(56));
   U1_55 : FA_X1 port map( A => A(55), B => B(55), CI => carry_55_port, CO => 
                           carry_56_port, S => SUM(55));
   U1_54 : FA_X1 port map( A => A(54), B => B(54), CI => carry_54_port, CO => 
                           carry_55_port, S => SUM(54));
   U1_53 : FA_X1 port map( A => A(53), B => B(53), CI => carry_53_port, CO => 
                           carry_54_port, S => SUM(53));
   U1_52 : FA_X1 port map( A => A(52), B => B(52), CI => carry_52_port, CO => 
                           carry_53_port, S => SUM(52));
   U1_51 : FA_X1 port map( A => A(51), B => B(51), CI => carry_51_port, CO => 
                           carry_52_port, S => SUM(51));
   U1_50 : FA_X1 port map( A => A(50), B => B(50), CI => carry_50_port, CO => 
                           carry_51_port, S => SUM(50));
   U1_49 : FA_X1 port map( A => A(49), B => B(49), CI => carry_49_port, CO => 
                           carry_50_port, S => SUM(49));
   U1_48 : FA_X1 port map( A => A(48), B => B(48), CI => carry_48_port, CO => 
                           carry_49_port, S => SUM(48));
   U1_47 : FA_X1 port map( A => A(47), B => B(47), CI => carry_47_port, CO => 
                           carry_48_port, S => SUM(47));
   U1_46 : FA_X1 port map( A => A(46), B => B(46), CI => carry_46_port, CO => 
                           carry_47_port, S => SUM(46));
   U1_45 : FA_X1 port map( A => A(45), B => B(45), CI => carry_45_port, CO => 
                           carry_46_port, S => SUM(45));
   U1_44 : FA_X1 port map( A => A(44), B => B(44), CI => carry_44_port, CO => 
                           carry_45_port, S => SUM(44));
   U1_43 : FA_X1 port map( A => A(43), B => B(43), CI => carry_43_port, CO => 
                           carry_44_port, S => SUM(43));
   U1_42 : FA_X1 port map( A => A(42), B => B(42), CI => carry_42_port, CO => 
                           carry_43_port, S => SUM(42));
   U1_41 : FA_X1 port map( A => A(41), B => B(41), CI => carry_41_port, CO => 
                           carry_42_port, S => SUM(41));
   U1_40 : FA_X1 port map( A => A(40), B => B(40), CI => carry_40_port, CO => 
                           carry_41_port, S => SUM(40));
   U1_39 : FA_X1 port map( A => A(39), B => B(39), CI => carry_39_port, CO => 
                           carry_40_port, S => SUM(39));
   U1_38 : FA_X1 port map( A => A(38), B => B(38), CI => carry_38_port, CO => 
                           carry_39_port, S => SUM(38));
   U1_37 : FA_X1 port map( A => A(37), B => B(37), CI => carry_37_port, CO => 
                           carry_38_port, S => SUM(37));
   U1_36 : FA_X1 port map( A => A(36), B => B(36), CI => carry_36_port, CO => 
                           carry_37_port, S => SUM(36));
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => carry_35_port, CO => 
                           carry_36_port, S => SUM(35));
   U1_34 : FA_X1 port map( A => A(34), B => B(34), CI => carry_34_port, CO => 
                           carry_35_port, S => SUM(34));
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => carry_32_port, CO => 
                           carry_33_port, S => SUM(32));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity RCA_NBIT64_17_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_NBIT64_17_DW01_add_0;

architecture SYN_rpl of RCA_NBIT64_17_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_63_port, carry_62_port, carry_61_port, carry_60_port, 
      carry_59_port, carry_58_port, carry_57_port, carry_56_port, carry_55_port
      , carry_54_port, carry_53_port, carry_52_port, carry_51_port, 
      carry_50_port, carry_49_port, carry_48_port, carry_47_port, carry_46_port
      , carry_45_port, carry_44_port, carry_43_port, carry_42_port, 
      carry_41_port, carry_40_port, carry_39_port, carry_38_port, carry_37_port
      , carry_36_port, carry_35_port, carry_34_port, carry_33_port, 
      carry_32_port, carry_31_port, carry_30_port, carry_29_port, carry_28_port
      , carry_27_port, carry_26_port, carry_25_port, carry_24_port, 
      carry_23_port, carry_22_port, carry_21_port, carry_20_port, carry_19_port
      , carry_18_port, carry_17_port, carry_16_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_10_port
      , carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1_61 : FA_X1 port map( A => A(61), B => B(61), CI => carry_61_port, CO => 
                           carry_62_port, S => SUM(61));
   U1_60 : FA_X1 port map( A => A(60), B => B(60), CI => carry_60_port, CO => 
                           carry_61_port, S => SUM(60));
   U1_59 : FA_X1 port map( A => A(59), B => B(59), CI => carry_59_port, CO => 
                           carry_60_port, S => SUM(59));
   U1_58 : FA_X1 port map( A => A(58), B => B(58), CI => carry_58_port, CO => 
                           carry_59_port, S => SUM(58));
   U1_57 : FA_X1 port map( A => A(57), B => B(57), CI => carry_57_port, CO => 
                           carry_58_port, S => SUM(57));
   U1_56 : FA_X1 port map( A => A(56), B => B(56), CI => carry_56_port, CO => 
                           carry_57_port, S => SUM(56));
   U1_55 : FA_X1 port map( A => A(55), B => B(55), CI => carry_55_port, CO => 
                           carry_56_port, S => SUM(55));
   U1_54 : FA_X1 port map( A => A(54), B => B(54), CI => carry_54_port, CO => 
                           carry_55_port, S => SUM(54));
   U1_53 : FA_X1 port map( A => A(53), B => B(53), CI => carry_53_port, CO => 
                           carry_54_port, S => SUM(53));
   U1_52 : FA_X1 port map( A => A(52), B => B(52), CI => carry_52_port, CO => 
                           carry_53_port, S => SUM(52));
   U1_51 : FA_X1 port map( A => A(51), B => B(51), CI => carry_51_port, CO => 
                           carry_52_port, S => SUM(51));
   U1_50 : FA_X1 port map( A => A(50), B => B(50), CI => carry_50_port, CO => 
                           carry_51_port, S => SUM(50));
   U1_49 : FA_X1 port map( A => A(49), B => B(49), CI => carry_49_port, CO => 
                           carry_50_port, S => SUM(49));
   U1_48 : FA_X1 port map( A => A(48), B => B(48), CI => carry_48_port, CO => 
                           carry_49_port, S => SUM(48));
   U1_47 : FA_X1 port map( A => A(47), B => B(47), CI => carry_47_port, CO => 
                           carry_48_port, S => SUM(47));
   U1_46 : FA_X1 port map( A => A(46), B => B(46), CI => carry_46_port, CO => 
                           carry_47_port, S => SUM(46));
   U1_45 : FA_X1 port map( A => A(45), B => B(45), CI => carry_45_port, CO => 
                           carry_46_port, S => SUM(45));
   U1_44 : FA_X1 port map( A => A(44), B => B(44), CI => carry_44_port, CO => 
                           carry_45_port, S => SUM(44));
   U1_43 : FA_X1 port map( A => A(43), B => B(43), CI => carry_43_port, CO => 
                           carry_44_port, S => SUM(43));
   U1_42 : FA_X1 port map( A => A(42), B => B(42), CI => carry_42_port, CO => 
                           carry_43_port, S => SUM(42));
   U1_41 : FA_X1 port map( A => A(41), B => B(41), CI => carry_41_port, CO => 
                           carry_42_port, S => SUM(41));
   U1_40 : FA_X1 port map( A => A(40), B => B(40), CI => carry_40_port, CO => 
                           carry_41_port, S => SUM(40));
   U1_39 : FA_X1 port map( A => A(39), B => B(39), CI => carry_39_port, CO => 
                           carry_40_port, S => SUM(39));
   U1_38 : FA_X1 port map( A => A(38), B => B(38), CI => carry_38_port, CO => 
                           carry_39_port, S => SUM(38));
   U1_37 : FA_X1 port map( A => A(37), B => B(37), CI => carry_37_port, CO => 
                           carry_38_port, S => SUM(37));
   U1_36 : FA_X1 port map( A => A(36), B => B(36), CI => carry_36_port, CO => 
                           carry_37_port, S => SUM(36));
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => carry_35_port, CO => 
                           carry_36_port, S => SUM(35));
   U1_34 : FA_X1 port map( A => A(34), B => B(34), CI => carry_34_port, CO => 
                           carry_35_port, S => SUM(34));
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => carry_32_port, CO => 
                           carry_33_port, S => SUM(32));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity RCA_NBIT64_18_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_NBIT64_18_DW01_add_0;

architecture SYN_rpl of RCA_NBIT64_18_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_63_port, carry_62_port, carry_61_port, carry_60_port, 
      carry_59_port, carry_58_port, carry_57_port, carry_56_port, carry_55_port
      , carry_54_port, carry_53_port, carry_52_port, carry_51_port, 
      carry_50_port, carry_49_port, carry_48_port, carry_47_port, carry_46_port
      , carry_45_port, carry_44_port, carry_43_port, carry_42_port, 
      carry_41_port, carry_40_port, carry_39_port, carry_38_port, carry_37_port
      , carry_36_port, carry_35_port, carry_34_port, carry_33_port, 
      carry_32_port, carry_31_port, carry_30_port, carry_29_port, carry_28_port
      , carry_27_port, carry_26_port, carry_25_port, carry_24_port, 
      carry_23_port, carry_22_port, carry_21_port, carry_20_port, carry_19_port
      , carry_18_port, carry_17_port, carry_16_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_10_port
      , carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1_61 : FA_X1 port map( A => A(61), B => B(61), CI => carry_61_port, CO => 
                           carry_62_port, S => SUM(61));
   U1_60 : FA_X1 port map( A => A(60), B => B(60), CI => carry_60_port, CO => 
                           carry_61_port, S => SUM(60));
   U1_59 : FA_X1 port map( A => A(59), B => B(59), CI => carry_59_port, CO => 
                           carry_60_port, S => SUM(59));
   U1_58 : FA_X1 port map( A => A(58), B => B(58), CI => carry_58_port, CO => 
                           carry_59_port, S => SUM(58));
   U1_57 : FA_X1 port map( A => A(57), B => B(57), CI => carry_57_port, CO => 
                           carry_58_port, S => SUM(57));
   U1_56 : FA_X1 port map( A => A(56), B => B(56), CI => carry_56_port, CO => 
                           carry_57_port, S => SUM(56));
   U1_55 : FA_X1 port map( A => A(55), B => B(55), CI => carry_55_port, CO => 
                           carry_56_port, S => SUM(55));
   U1_54 : FA_X1 port map( A => A(54), B => B(54), CI => carry_54_port, CO => 
                           carry_55_port, S => SUM(54));
   U1_53 : FA_X1 port map( A => A(53), B => B(53), CI => carry_53_port, CO => 
                           carry_54_port, S => SUM(53));
   U1_52 : FA_X1 port map( A => A(52), B => B(52), CI => carry_52_port, CO => 
                           carry_53_port, S => SUM(52));
   U1_51 : FA_X1 port map( A => A(51), B => B(51), CI => carry_51_port, CO => 
                           carry_52_port, S => SUM(51));
   U1_50 : FA_X1 port map( A => A(50), B => B(50), CI => carry_50_port, CO => 
                           carry_51_port, S => SUM(50));
   U1_49 : FA_X1 port map( A => A(49), B => B(49), CI => carry_49_port, CO => 
                           carry_50_port, S => SUM(49));
   U1_48 : FA_X1 port map( A => A(48), B => B(48), CI => carry_48_port, CO => 
                           carry_49_port, S => SUM(48));
   U1_47 : FA_X1 port map( A => A(47), B => B(47), CI => carry_47_port, CO => 
                           carry_48_port, S => SUM(47));
   U1_46 : FA_X1 port map( A => A(46), B => B(46), CI => carry_46_port, CO => 
                           carry_47_port, S => SUM(46));
   U1_45 : FA_X1 port map( A => A(45), B => B(45), CI => carry_45_port, CO => 
                           carry_46_port, S => SUM(45));
   U1_44 : FA_X1 port map( A => A(44), B => B(44), CI => carry_44_port, CO => 
                           carry_45_port, S => SUM(44));
   U1_43 : FA_X1 port map( A => A(43), B => B(43), CI => carry_43_port, CO => 
                           carry_44_port, S => SUM(43));
   U1_42 : FA_X1 port map( A => A(42), B => B(42), CI => carry_42_port, CO => 
                           carry_43_port, S => SUM(42));
   U1_41 : FA_X1 port map( A => A(41), B => B(41), CI => carry_41_port, CO => 
                           carry_42_port, S => SUM(41));
   U1_40 : FA_X1 port map( A => A(40), B => B(40), CI => carry_40_port, CO => 
                           carry_41_port, S => SUM(40));
   U1_39 : FA_X1 port map( A => A(39), B => B(39), CI => carry_39_port, CO => 
                           carry_40_port, S => SUM(39));
   U1_38 : FA_X1 port map( A => A(38), B => B(38), CI => carry_38_port, CO => 
                           carry_39_port, S => SUM(38));
   U1_37 : FA_X1 port map( A => A(37), B => B(37), CI => carry_37_port, CO => 
                           carry_38_port, S => SUM(37));
   U1_36 : FA_X1 port map( A => A(36), B => B(36), CI => carry_36_port, CO => 
                           carry_37_port, S => SUM(36));
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => carry_35_port, CO => 
                           carry_36_port, S => SUM(35));
   U1_34 : FA_X1 port map( A => A(34), B => B(34), CI => carry_34_port, CO => 
                           carry_35_port, S => SUM(34));
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => carry_32_port, CO => 
                           carry_33_port, S => SUM(32));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity RCA_NBIT64_19_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_NBIT64_19_DW01_add_0;

architecture SYN_rpl of RCA_NBIT64_19_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_63_port, carry_62_port, carry_61_port, carry_60_port, 
      carry_59_port, carry_58_port, carry_57_port, carry_56_port, carry_55_port
      , carry_54_port, carry_53_port, carry_52_port, carry_51_port, 
      carry_50_port, carry_49_port, carry_48_port, carry_47_port, carry_46_port
      , carry_45_port, carry_44_port, carry_43_port, carry_42_port, 
      carry_41_port, carry_40_port, carry_39_port, carry_38_port, carry_37_port
      , carry_36_port, carry_35_port, carry_34_port, carry_33_port, 
      carry_32_port, carry_31_port, carry_30_port, carry_29_port, carry_28_port
      , carry_27_port, carry_26_port, carry_25_port, carry_24_port, 
      carry_23_port, carry_22_port, carry_21_port, carry_20_port, carry_19_port
      , carry_18_port, carry_17_port, carry_16_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_10_port
      , carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1_61 : FA_X1 port map( A => A(61), B => B(61), CI => carry_61_port, CO => 
                           carry_62_port, S => SUM(61));
   U1_60 : FA_X1 port map( A => A(60), B => B(60), CI => carry_60_port, CO => 
                           carry_61_port, S => SUM(60));
   U1_59 : FA_X1 port map( A => A(59), B => B(59), CI => carry_59_port, CO => 
                           carry_60_port, S => SUM(59));
   U1_58 : FA_X1 port map( A => A(58), B => B(58), CI => carry_58_port, CO => 
                           carry_59_port, S => SUM(58));
   U1_57 : FA_X1 port map( A => A(57), B => B(57), CI => carry_57_port, CO => 
                           carry_58_port, S => SUM(57));
   U1_56 : FA_X1 port map( A => A(56), B => B(56), CI => carry_56_port, CO => 
                           carry_57_port, S => SUM(56));
   U1_55 : FA_X1 port map( A => A(55), B => B(55), CI => carry_55_port, CO => 
                           carry_56_port, S => SUM(55));
   U1_54 : FA_X1 port map( A => A(54), B => B(54), CI => carry_54_port, CO => 
                           carry_55_port, S => SUM(54));
   U1_53 : FA_X1 port map( A => A(53), B => B(53), CI => carry_53_port, CO => 
                           carry_54_port, S => SUM(53));
   U1_52 : FA_X1 port map( A => A(52), B => B(52), CI => carry_52_port, CO => 
                           carry_53_port, S => SUM(52));
   U1_51 : FA_X1 port map( A => A(51), B => B(51), CI => carry_51_port, CO => 
                           carry_52_port, S => SUM(51));
   U1_50 : FA_X1 port map( A => A(50), B => B(50), CI => carry_50_port, CO => 
                           carry_51_port, S => SUM(50));
   U1_49 : FA_X1 port map( A => A(49), B => B(49), CI => carry_49_port, CO => 
                           carry_50_port, S => SUM(49));
   U1_48 : FA_X1 port map( A => A(48), B => B(48), CI => carry_48_port, CO => 
                           carry_49_port, S => SUM(48));
   U1_47 : FA_X1 port map( A => A(47), B => B(47), CI => carry_47_port, CO => 
                           carry_48_port, S => SUM(47));
   U1_46 : FA_X1 port map( A => A(46), B => B(46), CI => carry_46_port, CO => 
                           carry_47_port, S => SUM(46));
   U1_45 : FA_X1 port map( A => A(45), B => B(45), CI => carry_45_port, CO => 
                           carry_46_port, S => SUM(45));
   U1_44 : FA_X1 port map( A => A(44), B => B(44), CI => carry_44_port, CO => 
                           carry_45_port, S => SUM(44));
   U1_43 : FA_X1 port map( A => A(43), B => B(43), CI => carry_43_port, CO => 
                           carry_44_port, S => SUM(43));
   U1_42 : FA_X1 port map( A => A(42), B => B(42), CI => carry_42_port, CO => 
                           carry_43_port, S => SUM(42));
   U1_41 : FA_X1 port map( A => A(41), B => B(41), CI => carry_41_port, CO => 
                           carry_42_port, S => SUM(41));
   U1_40 : FA_X1 port map( A => A(40), B => B(40), CI => carry_40_port, CO => 
                           carry_41_port, S => SUM(40));
   U1_39 : FA_X1 port map( A => A(39), B => B(39), CI => carry_39_port, CO => 
                           carry_40_port, S => SUM(39));
   U1_38 : FA_X1 port map( A => A(38), B => B(38), CI => carry_38_port, CO => 
                           carry_39_port, S => SUM(38));
   U1_37 : FA_X1 port map( A => A(37), B => B(37), CI => carry_37_port, CO => 
                           carry_38_port, S => SUM(37));
   U1_36 : FA_X1 port map( A => A(36), B => B(36), CI => carry_36_port, CO => 
                           carry_37_port, S => SUM(36));
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => carry_35_port, CO => 
                           carry_36_port, S => SUM(35));
   U1_34 : FA_X1 port map( A => A(34), B => B(34), CI => carry_34_port, CO => 
                           carry_35_port, S => SUM(34));
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => carry_32_port, CO => 
                           carry_33_port, S => SUM(32));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity RCA_NBIT64_20_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_NBIT64_20_DW01_add_0;

architecture SYN_rpl of RCA_NBIT64_20_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_63_port, carry_62_port, carry_61_port, carry_60_port, 
      carry_59_port, carry_58_port, carry_57_port, carry_56_port, carry_55_port
      , carry_54_port, carry_53_port, carry_52_port, carry_51_port, 
      carry_50_port, carry_49_port, carry_48_port, carry_47_port, carry_46_port
      , carry_45_port, carry_44_port, carry_43_port, carry_42_port, 
      carry_41_port, carry_40_port, carry_39_port, carry_38_port, carry_37_port
      , carry_36_port, carry_35_port, carry_34_port, carry_33_port, 
      carry_32_port, carry_31_port, carry_30_port, carry_29_port, carry_28_port
      , carry_27_port, carry_26_port, carry_25_port, carry_24_port, 
      carry_23_port, carry_22_port, carry_21_port, carry_20_port, carry_19_port
      , carry_18_port, carry_17_port, carry_16_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_10_port
      , carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1_61 : FA_X1 port map( A => A(61), B => B(61), CI => carry_61_port, CO => 
                           carry_62_port, S => SUM(61));
   U1_60 : FA_X1 port map( A => A(60), B => B(60), CI => carry_60_port, CO => 
                           carry_61_port, S => SUM(60));
   U1_59 : FA_X1 port map( A => A(59), B => B(59), CI => carry_59_port, CO => 
                           carry_60_port, S => SUM(59));
   U1_58 : FA_X1 port map( A => A(58), B => B(58), CI => carry_58_port, CO => 
                           carry_59_port, S => SUM(58));
   U1_57 : FA_X1 port map( A => A(57), B => B(57), CI => carry_57_port, CO => 
                           carry_58_port, S => SUM(57));
   U1_56 : FA_X1 port map( A => A(56), B => B(56), CI => carry_56_port, CO => 
                           carry_57_port, S => SUM(56));
   U1_55 : FA_X1 port map( A => A(55), B => B(55), CI => carry_55_port, CO => 
                           carry_56_port, S => SUM(55));
   U1_54 : FA_X1 port map( A => A(54), B => B(54), CI => carry_54_port, CO => 
                           carry_55_port, S => SUM(54));
   U1_53 : FA_X1 port map( A => A(53), B => B(53), CI => carry_53_port, CO => 
                           carry_54_port, S => SUM(53));
   U1_52 : FA_X1 port map( A => A(52), B => B(52), CI => carry_52_port, CO => 
                           carry_53_port, S => SUM(52));
   U1_51 : FA_X1 port map( A => A(51), B => B(51), CI => carry_51_port, CO => 
                           carry_52_port, S => SUM(51));
   U1_50 : FA_X1 port map( A => A(50), B => B(50), CI => carry_50_port, CO => 
                           carry_51_port, S => SUM(50));
   U1_49 : FA_X1 port map( A => A(49), B => B(49), CI => carry_49_port, CO => 
                           carry_50_port, S => SUM(49));
   U1_48 : FA_X1 port map( A => A(48), B => B(48), CI => carry_48_port, CO => 
                           carry_49_port, S => SUM(48));
   U1_47 : FA_X1 port map( A => A(47), B => B(47), CI => carry_47_port, CO => 
                           carry_48_port, S => SUM(47));
   U1_46 : FA_X1 port map( A => A(46), B => B(46), CI => carry_46_port, CO => 
                           carry_47_port, S => SUM(46));
   U1_45 : FA_X1 port map( A => A(45), B => B(45), CI => carry_45_port, CO => 
                           carry_46_port, S => SUM(45));
   U1_44 : FA_X1 port map( A => A(44), B => B(44), CI => carry_44_port, CO => 
                           carry_45_port, S => SUM(44));
   U1_43 : FA_X1 port map( A => A(43), B => B(43), CI => carry_43_port, CO => 
                           carry_44_port, S => SUM(43));
   U1_42 : FA_X1 port map( A => A(42), B => B(42), CI => carry_42_port, CO => 
                           carry_43_port, S => SUM(42));
   U1_41 : FA_X1 port map( A => A(41), B => B(41), CI => carry_41_port, CO => 
                           carry_42_port, S => SUM(41));
   U1_40 : FA_X1 port map( A => A(40), B => B(40), CI => carry_40_port, CO => 
                           carry_41_port, S => SUM(40));
   U1_39 : FA_X1 port map( A => A(39), B => B(39), CI => carry_39_port, CO => 
                           carry_40_port, S => SUM(39));
   U1_38 : FA_X1 port map( A => A(38), B => B(38), CI => carry_38_port, CO => 
                           carry_39_port, S => SUM(38));
   U1_37 : FA_X1 port map( A => A(37), B => B(37), CI => carry_37_port, CO => 
                           carry_38_port, S => SUM(37));
   U1_36 : FA_X1 port map( A => A(36), B => B(36), CI => carry_36_port, CO => 
                           carry_37_port, S => SUM(36));
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => carry_35_port, CO => 
                           carry_36_port, S => SUM(35));
   U1_34 : FA_X1 port map( A => A(34), B => B(34), CI => carry_34_port, CO => 
                           carry_35_port, S => SUM(34));
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => carry_32_port, CO => 
                           carry_33_port, S => SUM(32));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity RCA_NBIT64_21_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_NBIT64_21_DW01_add_0;

architecture SYN_rpl of RCA_NBIT64_21_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_63_port, carry_62_port, carry_61_port, carry_60_port, 
      carry_59_port, carry_58_port, carry_57_port, carry_56_port, carry_55_port
      , carry_54_port, carry_53_port, carry_52_port, carry_51_port, 
      carry_50_port, carry_49_port, carry_48_port, carry_47_port, carry_46_port
      , carry_45_port, carry_44_port, carry_43_port, carry_42_port, 
      carry_41_port, carry_40_port, carry_39_port, carry_38_port, carry_37_port
      , carry_36_port, carry_35_port, carry_34_port, carry_33_port, 
      carry_32_port, carry_31_port, carry_30_port, carry_29_port, carry_28_port
      , carry_27_port, carry_26_port, carry_25_port, carry_24_port, 
      carry_23_port, carry_22_port, carry_21_port, carry_20_port, carry_19_port
      , carry_18_port, carry_17_port, carry_16_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_10_port
      , carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1_61 : FA_X1 port map( A => A(61), B => B(61), CI => carry_61_port, CO => 
                           carry_62_port, S => SUM(61));
   U1_60 : FA_X1 port map( A => A(60), B => B(60), CI => carry_60_port, CO => 
                           carry_61_port, S => SUM(60));
   U1_59 : FA_X1 port map( A => A(59), B => B(59), CI => carry_59_port, CO => 
                           carry_60_port, S => SUM(59));
   U1_58 : FA_X1 port map( A => A(58), B => B(58), CI => carry_58_port, CO => 
                           carry_59_port, S => SUM(58));
   U1_57 : FA_X1 port map( A => A(57), B => B(57), CI => carry_57_port, CO => 
                           carry_58_port, S => SUM(57));
   U1_56 : FA_X1 port map( A => A(56), B => B(56), CI => carry_56_port, CO => 
                           carry_57_port, S => SUM(56));
   U1_55 : FA_X1 port map( A => A(55), B => B(55), CI => carry_55_port, CO => 
                           carry_56_port, S => SUM(55));
   U1_54 : FA_X1 port map( A => A(54), B => B(54), CI => carry_54_port, CO => 
                           carry_55_port, S => SUM(54));
   U1_53 : FA_X1 port map( A => A(53), B => B(53), CI => carry_53_port, CO => 
                           carry_54_port, S => SUM(53));
   U1_52 : FA_X1 port map( A => A(52), B => B(52), CI => carry_52_port, CO => 
                           carry_53_port, S => SUM(52));
   U1_51 : FA_X1 port map( A => A(51), B => B(51), CI => carry_51_port, CO => 
                           carry_52_port, S => SUM(51));
   U1_50 : FA_X1 port map( A => A(50), B => B(50), CI => carry_50_port, CO => 
                           carry_51_port, S => SUM(50));
   U1_49 : FA_X1 port map( A => A(49), B => B(49), CI => carry_49_port, CO => 
                           carry_50_port, S => SUM(49));
   U1_48 : FA_X1 port map( A => A(48), B => B(48), CI => carry_48_port, CO => 
                           carry_49_port, S => SUM(48));
   U1_47 : FA_X1 port map( A => A(47), B => B(47), CI => carry_47_port, CO => 
                           carry_48_port, S => SUM(47));
   U1_46 : FA_X1 port map( A => A(46), B => B(46), CI => carry_46_port, CO => 
                           carry_47_port, S => SUM(46));
   U1_45 : FA_X1 port map( A => A(45), B => B(45), CI => carry_45_port, CO => 
                           carry_46_port, S => SUM(45));
   U1_44 : FA_X1 port map( A => A(44), B => B(44), CI => carry_44_port, CO => 
                           carry_45_port, S => SUM(44));
   U1_43 : FA_X1 port map( A => A(43), B => B(43), CI => carry_43_port, CO => 
                           carry_44_port, S => SUM(43));
   U1_42 : FA_X1 port map( A => A(42), B => B(42), CI => carry_42_port, CO => 
                           carry_43_port, S => SUM(42));
   U1_41 : FA_X1 port map( A => A(41), B => B(41), CI => carry_41_port, CO => 
                           carry_42_port, S => SUM(41));
   U1_40 : FA_X1 port map( A => A(40), B => B(40), CI => carry_40_port, CO => 
                           carry_41_port, S => SUM(40));
   U1_39 : FA_X1 port map( A => A(39), B => B(39), CI => carry_39_port, CO => 
                           carry_40_port, S => SUM(39));
   U1_38 : FA_X1 port map( A => A(38), B => B(38), CI => carry_38_port, CO => 
                           carry_39_port, S => SUM(38));
   U1_37 : FA_X1 port map( A => A(37), B => B(37), CI => carry_37_port, CO => 
                           carry_38_port, S => SUM(37));
   U1_36 : FA_X1 port map( A => A(36), B => B(36), CI => carry_36_port, CO => 
                           carry_37_port, S => SUM(36));
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => carry_35_port, CO => 
                           carry_36_port, S => SUM(35));
   U1_34 : FA_X1 port map( A => A(34), B => B(34), CI => carry_34_port, CO => 
                           carry_35_port, S => SUM(34));
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => carry_32_port, CO => 
                           carry_33_port, S => SUM(32));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity RCA_NBIT64_22_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_NBIT64_22_DW01_add_0;

architecture SYN_rpl of RCA_NBIT64_22_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_63_port, carry_62_port, carry_61_port, carry_60_port, 
      carry_59_port, carry_58_port, carry_57_port, carry_56_port, carry_55_port
      , carry_54_port, carry_53_port, carry_52_port, carry_51_port, 
      carry_50_port, carry_49_port, carry_48_port, carry_47_port, carry_46_port
      , carry_45_port, carry_44_port, carry_43_port, carry_42_port, 
      carry_41_port, carry_40_port, carry_39_port, carry_38_port, carry_37_port
      , carry_36_port, carry_35_port, carry_34_port, carry_33_port, 
      carry_32_port, carry_31_port, carry_30_port, carry_29_port, carry_28_port
      , carry_27_port, carry_26_port, carry_25_port, carry_24_port, 
      carry_23_port, carry_22_port, carry_21_port, carry_20_port, carry_19_port
      , carry_18_port, carry_17_port, carry_16_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_10_port
      , carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1_61 : FA_X1 port map( A => A(61), B => B(61), CI => carry_61_port, CO => 
                           carry_62_port, S => SUM(61));
   U1_60 : FA_X1 port map( A => A(60), B => B(60), CI => carry_60_port, CO => 
                           carry_61_port, S => SUM(60));
   U1_59 : FA_X1 port map( A => A(59), B => B(59), CI => carry_59_port, CO => 
                           carry_60_port, S => SUM(59));
   U1_58 : FA_X1 port map( A => A(58), B => B(58), CI => carry_58_port, CO => 
                           carry_59_port, S => SUM(58));
   U1_57 : FA_X1 port map( A => A(57), B => B(57), CI => carry_57_port, CO => 
                           carry_58_port, S => SUM(57));
   U1_56 : FA_X1 port map( A => A(56), B => B(56), CI => carry_56_port, CO => 
                           carry_57_port, S => SUM(56));
   U1_55 : FA_X1 port map( A => A(55), B => B(55), CI => carry_55_port, CO => 
                           carry_56_port, S => SUM(55));
   U1_54 : FA_X1 port map( A => A(54), B => B(54), CI => carry_54_port, CO => 
                           carry_55_port, S => SUM(54));
   U1_53 : FA_X1 port map( A => A(53), B => B(53), CI => carry_53_port, CO => 
                           carry_54_port, S => SUM(53));
   U1_52 : FA_X1 port map( A => A(52), B => B(52), CI => carry_52_port, CO => 
                           carry_53_port, S => SUM(52));
   U1_51 : FA_X1 port map( A => A(51), B => B(51), CI => carry_51_port, CO => 
                           carry_52_port, S => SUM(51));
   U1_50 : FA_X1 port map( A => A(50), B => B(50), CI => carry_50_port, CO => 
                           carry_51_port, S => SUM(50));
   U1_49 : FA_X1 port map( A => A(49), B => B(49), CI => carry_49_port, CO => 
                           carry_50_port, S => SUM(49));
   U1_48 : FA_X1 port map( A => A(48), B => B(48), CI => carry_48_port, CO => 
                           carry_49_port, S => SUM(48));
   U1_47 : FA_X1 port map( A => A(47), B => B(47), CI => carry_47_port, CO => 
                           carry_48_port, S => SUM(47));
   U1_46 : FA_X1 port map( A => A(46), B => B(46), CI => carry_46_port, CO => 
                           carry_47_port, S => SUM(46));
   U1_45 : FA_X1 port map( A => A(45), B => B(45), CI => carry_45_port, CO => 
                           carry_46_port, S => SUM(45));
   U1_44 : FA_X1 port map( A => A(44), B => B(44), CI => carry_44_port, CO => 
                           carry_45_port, S => SUM(44));
   U1_43 : FA_X1 port map( A => A(43), B => B(43), CI => carry_43_port, CO => 
                           carry_44_port, S => SUM(43));
   U1_42 : FA_X1 port map( A => A(42), B => B(42), CI => carry_42_port, CO => 
                           carry_43_port, S => SUM(42));
   U1_41 : FA_X1 port map( A => A(41), B => B(41), CI => carry_41_port, CO => 
                           carry_42_port, S => SUM(41));
   U1_40 : FA_X1 port map( A => A(40), B => B(40), CI => carry_40_port, CO => 
                           carry_41_port, S => SUM(40));
   U1_39 : FA_X1 port map( A => A(39), B => B(39), CI => carry_39_port, CO => 
                           carry_40_port, S => SUM(39));
   U1_38 : FA_X1 port map( A => A(38), B => B(38), CI => carry_38_port, CO => 
                           carry_39_port, S => SUM(38));
   U1_37 : FA_X1 port map( A => A(37), B => B(37), CI => carry_37_port, CO => 
                           carry_38_port, S => SUM(37));
   U1_36 : FA_X1 port map( A => A(36), B => B(36), CI => carry_36_port, CO => 
                           carry_37_port, S => SUM(36));
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => carry_35_port, CO => 
                           carry_36_port, S => SUM(35));
   U1_34 : FA_X1 port map( A => A(34), B => B(34), CI => carry_34_port, CO => 
                           carry_35_port, S => SUM(34));
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => carry_32_port, CO => 
                           carry_33_port, S => SUM(32));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity RCA_NBIT64_23_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_NBIT64_23_DW01_add_0;

architecture SYN_rpl of RCA_NBIT64_23_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_63_port, carry_62_port, carry_61_port, carry_60_port, 
      carry_59_port, carry_58_port, carry_57_port, carry_56_port, carry_55_port
      , carry_54_port, carry_53_port, carry_52_port, carry_51_port, 
      carry_50_port, carry_49_port, carry_48_port, carry_47_port, carry_46_port
      , carry_45_port, carry_44_port, carry_43_port, carry_42_port, 
      carry_41_port, carry_40_port, carry_39_port, carry_38_port, carry_37_port
      , carry_36_port, carry_35_port, carry_34_port, carry_33_port, 
      carry_32_port, carry_31_port, carry_30_port, carry_29_port, carry_28_port
      , carry_27_port, carry_26_port, carry_25_port, carry_24_port, 
      carry_23_port, carry_22_port, carry_21_port, carry_20_port, carry_19_port
      , carry_18_port, carry_17_port, carry_16_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_10_port
      , carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1_61 : FA_X1 port map( A => A(61), B => B(61), CI => carry_61_port, CO => 
                           carry_62_port, S => SUM(61));
   U1_60 : FA_X1 port map( A => A(60), B => B(60), CI => carry_60_port, CO => 
                           carry_61_port, S => SUM(60));
   U1_59 : FA_X1 port map( A => A(59), B => B(59), CI => carry_59_port, CO => 
                           carry_60_port, S => SUM(59));
   U1_58 : FA_X1 port map( A => A(58), B => B(58), CI => carry_58_port, CO => 
                           carry_59_port, S => SUM(58));
   U1_57 : FA_X1 port map( A => A(57), B => B(57), CI => carry_57_port, CO => 
                           carry_58_port, S => SUM(57));
   U1_56 : FA_X1 port map( A => A(56), B => B(56), CI => carry_56_port, CO => 
                           carry_57_port, S => SUM(56));
   U1_55 : FA_X1 port map( A => A(55), B => B(55), CI => carry_55_port, CO => 
                           carry_56_port, S => SUM(55));
   U1_54 : FA_X1 port map( A => A(54), B => B(54), CI => carry_54_port, CO => 
                           carry_55_port, S => SUM(54));
   U1_53 : FA_X1 port map( A => A(53), B => B(53), CI => carry_53_port, CO => 
                           carry_54_port, S => SUM(53));
   U1_52 : FA_X1 port map( A => A(52), B => B(52), CI => carry_52_port, CO => 
                           carry_53_port, S => SUM(52));
   U1_51 : FA_X1 port map( A => A(51), B => B(51), CI => carry_51_port, CO => 
                           carry_52_port, S => SUM(51));
   U1_50 : FA_X1 port map( A => A(50), B => B(50), CI => carry_50_port, CO => 
                           carry_51_port, S => SUM(50));
   U1_49 : FA_X1 port map( A => A(49), B => B(49), CI => carry_49_port, CO => 
                           carry_50_port, S => SUM(49));
   U1_48 : FA_X1 port map( A => A(48), B => B(48), CI => carry_48_port, CO => 
                           carry_49_port, S => SUM(48));
   U1_47 : FA_X1 port map( A => A(47), B => B(47), CI => carry_47_port, CO => 
                           carry_48_port, S => SUM(47));
   U1_46 : FA_X1 port map( A => A(46), B => B(46), CI => carry_46_port, CO => 
                           carry_47_port, S => SUM(46));
   U1_45 : FA_X1 port map( A => A(45), B => B(45), CI => carry_45_port, CO => 
                           carry_46_port, S => SUM(45));
   U1_44 : FA_X1 port map( A => A(44), B => B(44), CI => carry_44_port, CO => 
                           carry_45_port, S => SUM(44));
   U1_43 : FA_X1 port map( A => A(43), B => B(43), CI => carry_43_port, CO => 
                           carry_44_port, S => SUM(43));
   U1_42 : FA_X1 port map( A => A(42), B => B(42), CI => carry_42_port, CO => 
                           carry_43_port, S => SUM(42));
   U1_41 : FA_X1 port map( A => A(41), B => B(41), CI => carry_41_port, CO => 
                           carry_42_port, S => SUM(41));
   U1_40 : FA_X1 port map( A => A(40), B => B(40), CI => carry_40_port, CO => 
                           carry_41_port, S => SUM(40));
   U1_39 : FA_X1 port map( A => A(39), B => B(39), CI => carry_39_port, CO => 
                           carry_40_port, S => SUM(39));
   U1_38 : FA_X1 port map( A => A(38), B => B(38), CI => carry_38_port, CO => 
                           carry_39_port, S => SUM(38));
   U1_37 : FA_X1 port map( A => A(37), B => B(37), CI => carry_37_port, CO => 
                           carry_38_port, S => SUM(37));
   U1_36 : FA_X1 port map( A => A(36), B => B(36), CI => carry_36_port, CO => 
                           carry_37_port, S => SUM(36));
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => carry_35_port, CO => 
                           carry_36_port, S => SUM(35));
   U1_34 : FA_X1 port map( A => A(34), B => B(34), CI => carry_34_port, CO => 
                           carry_35_port, S => SUM(34));
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => carry_32_port, CO => 
                           carry_33_port, S => SUM(32));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity RCA_NBIT64_24_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_NBIT64_24_DW01_add_0;

architecture SYN_rpl of RCA_NBIT64_24_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_63_port, carry_62_port, carry_61_port, carry_60_port, 
      carry_59_port, carry_58_port, carry_57_port, carry_56_port, carry_55_port
      , carry_54_port, carry_53_port, carry_52_port, carry_51_port, 
      carry_50_port, carry_49_port, carry_48_port, carry_47_port, carry_46_port
      , carry_45_port, carry_44_port, carry_43_port, carry_42_port, 
      carry_41_port, carry_40_port, carry_39_port, carry_38_port, carry_37_port
      , carry_36_port, carry_35_port, carry_34_port, carry_33_port, 
      carry_32_port, carry_31_port, carry_30_port, carry_29_port, carry_28_port
      , carry_27_port, carry_26_port, carry_25_port, carry_24_port, 
      carry_23_port, carry_22_port, carry_21_port, carry_20_port, carry_19_port
      , carry_18_port, carry_17_port, carry_16_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_10_port
      , carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1_61 : FA_X1 port map( A => A(61), B => B(61), CI => carry_61_port, CO => 
                           carry_62_port, S => SUM(61));
   U1_60 : FA_X1 port map( A => A(60), B => B(60), CI => carry_60_port, CO => 
                           carry_61_port, S => SUM(60));
   U1_59 : FA_X1 port map( A => A(59), B => B(59), CI => carry_59_port, CO => 
                           carry_60_port, S => SUM(59));
   U1_58 : FA_X1 port map( A => A(58), B => B(58), CI => carry_58_port, CO => 
                           carry_59_port, S => SUM(58));
   U1_57 : FA_X1 port map( A => A(57), B => B(57), CI => carry_57_port, CO => 
                           carry_58_port, S => SUM(57));
   U1_56 : FA_X1 port map( A => A(56), B => B(56), CI => carry_56_port, CO => 
                           carry_57_port, S => SUM(56));
   U1_55 : FA_X1 port map( A => A(55), B => B(55), CI => carry_55_port, CO => 
                           carry_56_port, S => SUM(55));
   U1_54 : FA_X1 port map( A => A(54), B => B(54), CI => carry_54_port, CO => 
                           carry_55_port, S => SUM(54));
   U1_53 : FA_X1 port map( A => A(53), B => B(53), CI => carry_53_port, CO => 
                           carry_54_port, S => SUM(53));
   U1_52 : FA_X1 port map( A => A(52), B => B(52), CI => carry_52_port, CO => 
                           carry_53_port, S => SUM(52));
   U1_51 : FA_X1 port map( A => A(51), B => B(51), CI => carry_51_port, CO => 
                           carry_52_port, S => SUM(51));
   U1_50 : FA_X1 port map( A => A(50), B => B(50), CI => carry_50_port, CO => 
                           carry_51_port, S => SUM(50));
   U1_49 : FA_X1 port map( A => A(49), B => B(49), CI => carry_49_port, CO => 
                           carry_50_port, S => SUM(49));
   U1_48 : FA_X1 port map( A => A(48), B => B(48), CI => carry_48_port, CO => 
                           carry_49_port, S => SUM(48));
   U1_47 : FA_X1 port map( A => A(47), B => B(47), CI => carry_47_port, CO => 
                           carry_48_port, S => SUM(47));
   U1_46 : FA_X1 port map( A => A(46), B => B(46), CI => carry_46_port, CO => 
                           carry_47_port, S => SUM(46));
   U1_45 : FA_X1 port map( A => A(45), B => B(45), CI => carry_45_port, CO => 
                           carry_46_port, S => SUM(45));
   U1_44 : FA_X1 port map( A => A(44), B => B(44), CI => carry_44_port, CO => 
                           carry_45_port, S => SUM(44));
   U1_43 : FA_X1 port map( A => A(43), B => B(43), CI => carry_43_port, CO => 
                           carry_44_port, S => SUM(43));
   U1_42 : FA_X1 port map( A => A(42), B => B(42), CI => carry_42_port, CO => 
                           carry_43_port, S => SUM(42));
   U1_41 : FA_X1 port map( A => A(41), B => B(41), CI => carry_41_port, CO => 
                           carry_42_port, S => SUM(41));
   U1_40 : FA_X1 port map( A => A(40), B => B(40), CI => carry_40_port, CO => 
                           carry_41_port, S => SUM(40));
   U1_39 : FA_X1 port map( A => A(39), B => B(39), CI => carry_39_port, CO => 
                           carry_40_port, S => SUM(39));
   U1_38 : FA_X1 port map( A => A(38), B => B(38), CI => carry_38_port, CO => 
                           carry_39_port, S => SUM(38));
   U1_37 : FA_X1 port map( A => A(37), B => B(37), CI => carry_37_port, CO => 
                           carry_38_port, S => SUM(37));
   U1_36 : FA_X1 port map( A => A(36), B => B(36), CI => carry_36_port, CO => 
                           carry_37_port, S => SUM(36));
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => carry_35_port, CO => 
                           carry_36_port, S => SUM(35));
   U1_34 : FA_X1 port map( A => A(34), B => B(34), CI => carry_34_port, CO => 
                           carry_35_port, S => SUM(34));
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => carry_32_port, CO => 
                           carry_33_port, S => SUM(32));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity RCA_NBIT64_25_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_NBIT64_25_DW01_add_0;

architecture SYN_rpl of RCA_NBIT64_25_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_63_port, carry_62_port, carry_61_port, carry_60_port, 
      carry_59_port, carry_58_port, carry_57_port, carry_56_port, carry_55_port
      , carry_54_port, carry_53_port, carry_52_port, carry_51_port, 
      carry_50_port, carry_49_port, carry_48_port, carry_47_port, carry_46_port
      , carry_45_port, carry_44_port, carry_43_port, carry_42_port, 
      carry_41_port, carry_40_port, carry_39_port, carry_38_port, carry_37_port
      , carry_36_port, carry_35_port, carry_34_port, carry_33_port, 
      carry_32_port, carry_31_port, carry_30_port, carry_29_port, carry_28_port
      , carry_27_port, carry_26_port, carry_25_port, carry_24_port, 
      carry_23_port, carry_22_port, carry_21_port, carry_20_port, carry_19_port
      , carry_18_port, carry_17_port, carry_16_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_10_port
      , carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1_61 : FA_X1 port map( A => A(61), B => B(61), CI => carry_61_port, CO => 
                           carry_62_port, S => SUM(61));
   U1_60 : FA_X1 port map( A => A(60), B => B(60), CI => carry_60_port, CO => 
                           carry_61_port, S => SUM(60));
   U1_59 : FA_X1 port map( A => A(59), B => B(59), CI => carry_59_port, CO => 
                           carry_60_port, S => SUM(59));
   U1_58 : FA_X1 port map( A => A(58), B => B(58), CI => carry_58_port, CO => 
                           carry_59_port, S => SUM(58));
   U1_57 : FA_X1 port map( A => A(57), B => B(57), CI => carry_57_port, CO => 
                           carry_58_port, S => SUM(57));
   U1_56 : FA_X1 port map( A => A(56), B => B(56), CI => carry_56_port, CO => 
                           carry_57_port, S => SUM(56));
   U1_55 : FA_X1 port map( A => A(55), B => B(55), CI => carry_55_port, CO => 
                           carry_56_port, S => SUM(55));
   U1_54 : FA_X1 port map( A => A(54), B => B(54), CI => carry_54_port, CO => 
                           carry_55_port, S => SUM(54));
   U1_53 : FA_X1 port map( A => A(53), B => B(53), CI => carry_53_port, CO => 
                           carry_54_port, S => SUM(53));
   U1_52 : FA_X1 port map( A => A(52), B => B(52), CI => carry_52_port, CO => 
                           carry_53_port, S => SUM(52));
   U1_51 : FA_X1 port map( A => A(51), B => B(51), CI => carry_51_port, CO => 
                           carry_52_port, S => SUM(51));
   U1_50 : FA_X1 port map( A => A(50), B => B(50), CI => carry_50_port, CO => 
                           carry_51_port, S => SUM(50));
   U1_49 : FA_X1 port map( A => A(49), B => B(49), CI => carry_49_port, CO => 
                           carry_50_port, S => SUM(49));
   U1_48 : FA_X1 port map( A => A(48), B => B(48), CI => carry_48_port, CO => 
                           carry_49_port, S => SUM(48));
   U1_47 : FA_X1 port map( A => A(47), B => B(47), CI => carry_47_port, CO => 
                           carry_48_port, S => SUM(47));
   U1_46 : FA_X1 port map( A => A(46), B => B(46), CI => carry_46_port, CO => 
                           carry_47_port, S => SUM(46));
   U1_45 : FA_X1 port map( A => A(45), B => B(45), CI => carry_45_port, CO => 
                           carry_46_port, S => SUM(45));
   U1_44 : FA_X1 port map( A => A(44), B => B(44), CI => carry_44_port, CO => 
                           carry_45_port, S => SUM(44));
   U1_43 : FA_X1 port map( A => A(43), B => B(43), CI => carry_43_port, CO => 
                           carry_44_port, S => SUM(43));
   U1_42 : FA_X1 port map( A => A(42), B => B(42), CI => carry_42_port, CO => 
                           carry_43_port, S => SUM(42));
   U1_41 : FA_X1 port map( A => A(41), B => B(41), CI => carry_41_port, CO => 
                           carry_42_port, S => SUM(41));
   U1_40 : FA_X1 port map( A => A(40), B => B(40), CI => carry_40_port, CO => 
                           carry_41_port, S => SUM(40));
   U1_39 : FA_X1 port map( A => A(39), B => B(39), CI => carry_39_port, CO => 
                           carry_40_port, S => SUM(39));
   U1_38 : FA_X1 port map( A => A(38), B => B(38), CI => carry_38_port, CO => 
                           carry_39_port, S => SUM(38));
   U1_37 : FA_X1 port map( A => A(37), B => B(37), CI => carry_37_port, CO => 
                           carry_38_port, S => SUM(37));
   U1_36 : FA_X1 port map( A => A(36), B => B(36), CI => carry_36_port, CO => 
                           carry_37_port, S => SUM(36));
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => carry_35_port, CO => 
                           carry_36_port, S => SUM(35));
   U1_34 : FA_X1 port map( A => A(34), B => B(34), CI => carry_34_port, CO => 
                           carry_35_port, S => SUM(34));
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => carry_32_port, CO => 
                           carry_33_port, S => SUM(32));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity RCA_NBIT64_26_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_NBIT64_26_DW01_add_0;

architecture SYN_rpl of RCA_NBIT64_26_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_63_port, carry_62_port, carry_61_port, carry_60_port, 
      carry_59_port, carry_58_port, carry_57_port, carry_56_port, carry_55_port
      , carry_54_port, carry_53_port, carry_52_port, carry_51_port, 
      carry_50_port, carry_49_port, carry_48_port, carry_47_port, carry_46_port
      , carry_45_port, carry_44_port, carry_43_port, carry_42_port, 
      carry_41_port, carry_40_port, carry_39_port, carry_38_port, carry_37_port
      , carry_36_port, carry_35_port, carry_34_port, carry_33_port, 
      carry_32_port, carry_31_port, carry_30_port, carry_29_port, carry_28_port
      , carry_27_port, carry_26_port, carry_25_port, carry_24_port, 
      carry_23_port, carry_22_port, carry_21_port, carry_20_port, carry_19_port
      , carry_18_port, carry_17_port, carry_16_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_10_port
      , carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1_61 : FA_X1 port map( A => A(61), B => B(61), CI => carry_61_port, CO => 
                           carry_62_port, S => SUM(61));
   U1_60 : FA_X1 port map( A => A(60), B => B(60), CI => carry_60_port, CO => 
                           carry_61_port, S => SUM(60));
   U1_59 : FA_X1 port map( A => A(59), B => B(59), CI => carry_59_port, CO => 
                           carry_60_port, S => SUM(59));
   U1_58 : FA_X1 port map( A => A(58), B => B(58), CI => carry_58_port, CO => 
                           carry_59_port, S => SUM(58));
   U1_57 : FA_X1 port map( A => A(57), B => B(57), CI => carry_57_port, CO => 
                           carry_58_port, S => SUM(57));
   U1_56 : FA_X1 port map( A => A(56), B => B(56), CI => carry_56_port, CO => 
                           carry_57_port, S => SUM(56));
   U1_55 : FA_X1 port map( A => A(55), B => B(55), CI => carry_55_port, CO => 
                           carry_56_port, S => SUM(55));
   U1_54 : FA_X1 port map( A => A(54), B => B(54), CI => carry_54_port, CO => 
                           carry_55_port, S => SUM(54));
   U1_53 : FA_X1 port map( A => A(53), B => B(53), CI => carry_53_port, CO => 
                           carry_54_port, S => SUM(53));
   U1_52 : FA_X1 port map( A => A(52), B => B(52), CI => carry_52_port, CO => 
                           carry_53_port, S => SUM(52));
   U1_51 : FA_X1 port map( A => A(51), B => B(51), CI => carry_51_port, CO => 
                           carry_52_port, S => SUM(51));
   U1_50 : FA_X1 port map( A => A(50), B => B(50), CI => carry_50_port, CO => 
                           carry_51_port, S => SUM(50));
   U1_49 : FA_X1 port map( A => A(49), B => B(49), CI => carry_49_port, CO => 
                           carry_50_port, S => SUM(49));
   U1_48 : FA_X1 port map( A => A(48), B => B(48), CI => carry_48_port, CO => 
                           carry_49_port, S => SUM(48));
   U1_47 : FA_X1 port map( A => A(47), B => B(47), CI => carry_47_port, CO => 
                           carry_48_port, S => SUM(47));
   U1_46 : FA_X1 port map( A => A(46), B => B(46), CI => carry_46_port, CO => 
                           carry_47_port, S => SUM(46));
   U1_45 : FA_X1 port map( A => A(45), B => B(45), CI => carry_45_port, CO => 
                           carry_46_port, S => SUM(45));
   U1_44 : FA_X1 port map( A => A(44), B => B(44), CI => carry_44_port, CO => 
                           carry_45_port, S => SUM(44));
   U1_43 : FA_X1 port map( A => A(43), B => B(43), CI => carry_43_port, CO => 
                           carry_44_port, S => SUM(43));
   U1_42 : FA_X1 port map( A => A(42), B => B(42), CI => carry_42_port, CO => 
                           carry_43_port, S => SUM(42));
   U1_41 : FA_X1 port map( A => A(41), B => B(41), CI => carry_41_port, CO => 
                           carry_42_port, S => SUM(41));
   U1_40 : FA_X1 port map( A => A(40), B => B(40), CI => carry_40_port, CO => 
                           carry_41_port, S => SUM(40));
   U1_39 : FA_X1 port map( A => A(39), B => B(39), CI => carry_39_port, CO => 
                           carry_40_port, S => SUM(39));
   U1_38 : FA_X1 port map( A => A(38), B => B(38), CI => carry_38_port, CO => 
                           carry_39_port, S => SUM(38));
   U1_37 : FA_X1 port map( A => A(37), B => B(37), CI => carry_37_port, CO => 
                           carry_38_port, S => SUM(37));
   U1_36 : FA_X1 port map( A => A(36), B => B(36), CI => carry_36_port, CO => 
                           carry_37_port, S => SUM(36));
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => carry_35_port, CO => 
                           carry_36_port, S => SUM(35));
   U1_34 : FA_X1 port map( A => A(34), B => B(34), CI => carry_34_port, CO => 
                           carry_35_port, S => SUM(34));
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => carry_32_port, CO => 
                           carry_33_port, S => SUM(32));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity RCA_NBIT64_27_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_NBIT64_27_DW01_add_0;

architecture SYN_rpl of RCA_NBIT64_27_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_63_port, carry_62_port, carry_61_port, carry_60_port, 
      carry_59_port, carry_58_port, carry_57_port, carry_56_port, carry_55_port
      , carry_54_port, carry_53_port, carry_52_port, carry_51_port, 
      carry_50_port, carry_49_port, carry_48_port, carry_47_port, carry_46_port
      , carry_45_port, carry_44_port, carry_43_port, carry_42_port, 
      carry_41_port, carry_40_port, carry_39_port, carry_38_port, carry_37_port
      , carry_36_port, carry_35_port, carry_34_port, carry_33_port, 
      carry_32_port, carry_31_port, carry_30_port, carry_29_port, carry_28_port
      , carry_27_port, carry_26_port, carry_25_port, carry_24_port, 
      carry_23_port, carry_22_port, carry_21_port, carry_20_port, carry_19_port
      , carry_18_port, carry_17_port, carry_16_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_10_port
      , carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1_61 : FA_X1 port map( A => A(61), B => B(61), CI => carry_61_port, CO => 
                           carry_62_port, S => SUM(61));
   U1_60 : FA_X1 port map( A => A(60), B => B(60), CI => carry_60_port, CO => 
                           carry_61_port, S => SUM(60));
   U1_59 : FA_X1 port map( A => A(59), B => B(59), CI => carry_59_port, CO => 
                           carry_60_port, S => SUM(59));
   U1_58 : FA_X1 port map( A => A(58), B => B(58), CI => carry_58_port, CO => 
                           carry_59_port, S => SUM(58));
   U1_57 : FA_X1 port map( A => A(57), B => B(57), CI => carry_57_port, CO => 
                           carry_58_port, S => SUM(57));
   U1_56 : FA_X1 port map( A => A(56), B => B(56), CI => carry_56_port, CO => 
                           carry_57_port, S => SUM(56));
   U1_55 : FA_X1 port map( A => A(55), B => B(55), CI => carry_55_port, CO => 
                           carry_56_port, S => SUM(55));
   U1_54 : FA_X1 port map( A => A(54), B => B(54), CI => carry_54_port, CO => 
                           carry_55_port, S => SUM(54));
   U1_53 : FA_X1 port map( A => A(53), B => B(53), CI => carry_53_port, CO => 
                           carry_54_port, S => SUM(53));
   U1_52 : FA_X1 port map( A => A(52), B => B(52), CI => carry_52_port, CO => 
                           carry_53_port, S => SUM(52));
   U1_51 : FA_X1 port map( A => A(51), B => B(51), CI => carry_51_port, CO => 
                           carry_52_port, S => SUM(51));
   U1_50 : FA_X1 port map( A => A(50), B => B(50), CI => carry_50_port, CO => 
                           carry_51_port, S => SUM(50));
   U1_49 : FA_X1 port map( A => A(49), B => B(49), CI => carry_49_port, CO => 
                           carry_50_port, S => SUM(49));
   U1_48 : FA_X1 port map( A => A(48), B => B(48), CI => carry_48_port, CO => 
                           carry_49_port, S => SUM(48));
   U1_47 : FA_X1 port map( A => A(47), B => B(47), CI => carry_47_port, CO => 
                           carry_48_port, S => SUM(47));
   U1_46 : FA_X1 port map( A => A(46), B => B(46), CI => carry_46_port, CO => 
                           carry_47_port, S => SUM(46));
   U1_45 : FA_X1 port map( A => A(45), B => B(45), CI => carry_45_port, CO => 
                           carry_46_port, S => SUM(45));
   U1_44 : FA_X1 port map( A => A(44), B => B(44), CI => carry_44_port, CO => 
                           carry_45_port, S => SUM(44));
   U1_43 : FA_X1 port map( A => A(43), B => B(43), CI => carry_43_port, CO => 
                           carry_44_port, S => SUM(43));
   U1_42 : FA_X1 port map( A => A(42), B => B(42), CI => carry_42_port, CO => 
                           carry_43_port, S => SUM(42));
   U1_41 : FA_X1 port map( A => A(41), B => B(41), CI => carry_41_port, CO => 
                           carry_42_port, S => SUM(41));
   U1_40 : FA_X1 port map( A => A(40), B => B(40), CI => carry_40_port, CO => 
                           carry_41_port, S => SUM(40));
   U1_39 : FA_X1 port map( A => A(39), B => B(39), CI => carry_39_port, CO => 
                           carry_40_port, S => SUM(39));
   U1_38 : FA_X1 port map( A => A(38), B => B(38), CI => carry_38_port, CO => 
                           carry_39_port, S => SUM(38));
   U1_37 : FA_X1 port map( A => A(37), B => B(37), CI => carry_37_port, CO => 
                           carry_38_port, S => SUM(37));
   U1_36 : FA_X1 port map( A => A(36), B => B(36), CI => carry_36_port, CO => 
                           carry_37_port, S => SUM(36));
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => carry_35_port, CO => 
                           carry_36_port, S => SUM(35));
   U1_34 : FA_X1 port map( A => A(34), B => B(34), CI => carry_34_port, CO => 
                           carry_35_port, S => SUM(34));
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => carry_32_port, CO => 
                           carry_33_port, S => SUM(32));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity RCA_NBIT64_28_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_NBIT64_28_DW01_add_0;

architecture SYN_rpl of RCA_NBIT64_28_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_63_port, carry_62_port, carry_61_port, carry_60_port, 
      carry_59_port, carry_58_port, carry_57_port, carry_56_port, carry_55_port
      , carry_54_port, carry_53_port, carry_52_port, carry_51_port, 
      carry_50_port, carry_49_port, carry_48_port, carry_47_port, carry_46_port
      , carry_45_port, carry_44_port, carry_43_port, carry_42_port, 
      carry_41_port, carry_40_port, carry_39_port, carry_38_port, carry_37_port
      , carry_36_port, carry_35_port, carry_34_port, carry_33_port, 
      carry_32_port, carry_31_port, carry_30_port, carry_29_port, carry_28_port
      , carry_27_port, carry_26_port, carry_25_port, carry_24_port, 
      carry_23_port, carry_22_port, carry_21_port, carry_20_port, carry_19_port
      , carry_18_port, carry_17_port, carry_16_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_10_port
      , carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1_61 : FA_X1 port map( A => A(61), B => B(61), CI => carry_61_port, CO => 
                           carry_62_port, S => SUM(61));
   U1_60 : FA_X1 port map( A => A(60), B => B(60), CI => carry_60_port, CO => 
                           carry_61_port, S => SUM(60));
   U1_59 : FA_X1 port map( A => A(59), B => B(59), CI => carry_59_port, CO => 
                           carry_60_port, S => SUM(59));
   U1_58 : FA_X1 port map( A => A(58), B => B(58), CI => carry_58_port, CO => 
                           carry_59_port, S => SUM(58));
   U1_57 : FA_X1 port map( A => A(57), B => B(57), CI => carry_57_port, CO => 
                           carry_58_port, S => SUM(57));
   U1_56 : FA_X1 port map( A => A(56), B => B(56), CI => carry_56_port, CO => 
                           carry_57_port, S => SUM(56));
   U1_55 : FA_X1 port map( A => A(55), B => B(55), CI => carry_55_port, CO => 
                           carry_56_port, S => SUM(55));
   U1_54 : FA_X1 port map( A => A(54), B => B(54), CI => carry_54_port, CO => 
                           carry_55_port, S => SUM(54));
   U1_53 : FA_X1 port map( A => A(53), B => B(53), CI => carry_53_port, CO => 
                           carry_54_port, S => SUM(53));
   U1_52 : FA_X1 port map( A => A(52), B => B(52), CI => carry_52_port, CO => 
                           carry_53_port, S => SUM(52));
   U1_51 : FA_X1 port map( A => A(51), B => B(51), CI => carry_51_port, CO => 
                           carry_52_port, S => SUM(51));
   U1_50 : FA_X1 port map( A => A(50), B => B(50), CI => carry_50_port, CO => 
                           carry_51_port, S => SUM(50));
   U1_49 : FA_X1 port map( A => A(49), B => B(49), CI => carry_49_port, CO => 
                           carry_50_port, S => SUM(49));
   U1_48 : FA_X1 port map( A => A(48), B => B(48), CI => carry_48_port, CO => 
                           carry_49_port, S => SUM(48));
   U1_47 : FA_X1 port map( A => A(47), B => B(47), CI => carry_47_port, CO => 
                           carry_48_port, S => SUM(47));
   U1_46 : FA_X1 port map( A => A(46), B => B(46), CI => carry_46_port, CO => 
                           carry_47_port, S => SUM(46));
   U1_45 : FA_X1 port map( A => A(45), B => B(45), CI => carry_45_port, CO => 
                           carry_46_port, S => SUM(45));
   U1_44 : FA_X1 port map( A => A(44), B => B(44), CI => carry_44_port, CO => 
                           carry_45_port, S => SUM(44));
   U1_43 : FA_X1 port map( A => A(43), B => B(43), CI => carry_43_port, CO => 
                           carry_44_port, S => SUM(43));
   U1_42 : FA_X1 port map( A => A(42), B => B(42), CI => carry_42_port, CO => 
                           carry_43_port, S => SUM(42));
   U1_41 : FA_X1 port map( A => A(41), B => B(41), CI => carry_41_port, CO => 
                           carry_42_port, S => SUM(41));
   U1_40 : FA_X1 port map( A => A(40), B => B(40), CI => carry_40_port, CO => 
                           carry_41_port, S => SUM(40));
   U1_39 : FA_X1 port map( A => A(39), B => B(39), CI => carry_39_port, CO => 
                           carry_40_port, S => SUM(39));
   U1_38 : FA_X1 port map( A => A(38), B => B(38), CI => carry_38_port, CO => 
                           carry_39_port, S => SUM(38));
   U1_37 : FA_X1 port map( A => A(37), B => B(37), CI => carry_37_port, CO => 
                           carry_38_port, S => SUM(37));
   U1_36 : FA_X1 port map( A => A(36), B => B(36), CI => carry_36_port, CO => 
                           carry_37_port, S => SUM(36));
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => carry_35_port, CO => 
                           carry_36_port, S => SUM(35));
   U1_34 : FA_X1 port map( A => A(34), B => B(34), CI => carry_34_port, CO => 
                           carry_35_port, S => SUM(34));
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => carry_32_port, CO => 
                           carry_33_port, S => SUM(32));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity RCA_NBIT64_29_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_NBIT64_29_DW01_add_0;

architecture SYN_rpl of RCA_NBIT64_29_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_63_port, carry_62_port, carry_61_port, carry_60_port, 
      carry_59_port, carry_58_port, carry_57_port, carry_56_port, carry_55_port
      , carry_54_port, carry_53_port, carry_52_port, carry_51_port, 
      carry_50_port, carry_49_port, carry_48_port, carry_47_port, carry_46_port
      , carry_45_port, carry_44_port, carry_43_port, carry_42_port, 
      carry_41_port, carry_40_port, carry_39_port, carry_38_port, carry_37_port
      , carry_36_port, carry_35_port, carry_34_port, carry_33_port, 
      carry_32_port, carry_31_port, carry_30_port, carry_29_port, carry_28_port
      , carry_27_port, carry_26_port, carry_25_port, carry_24_port, 
      carry_23_port, carry_22_port, carry_21_port, carry_20_port, carry_19_port
      , carry_18_port, carry_17_port, carry_16_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_10_port
      , carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1_61 : FA_X1 port map( A => A(61), B => B(61), CI => carry_61_port, CO => 
                           carry_62_port, S => SUM(61));
   U1_60 : FA_X1 port map( A => A(60), B => B(60), CI => carry_60_port, CO => 
                           carry_61_port, S => SUM(60));
   U1_59 : FA_X1 port map( A => A(59), B => B(59), CI => carry_59_port, CO => 
                           carry_60_port, S => SUM(59));
   U1_58 : FA_X1 port map( A => A(58), B => B(58), CI => carry_58_port, CO => 
                           carry_59_port, S => SUM(58));
   U1_57 : FA_X1 port map( A => A(57), B => B(57), CI => carry_57_port, CO => 
                           carry_58_port, S => SUM(57));
   U1_56 : FA_X1 port map( A => A(56), B => B(56), CI => carry_56_port, CO => 
                           carry_57_port, S => SUM(56));
   U1_55 : FA_X1 port map( A => A(55), B => B(55), CI => carry_55_port, CO => 
                           carry_56_port, S => SUM(55));
   U1_54 : FA_X1 port map( A => A(54), B => B(54), CI => carry_54_port, CO => 
                           carry_55_port, S => SUM(54));
   U1_53 : FA_X1 port map( A => A(53), B => B(53), CI => carry_53_port, CO => 
                           carry_54_port, S => SUM(53));
   U1_52 : FA_X1 port map( A => A(52), B => B(52), CI => carry_52_port, CO => 
                           carry_53_port, S => SUM(52));
   U1_51 : FA_X1 port map( A => A(51), B => B(51), CI => carry_51_port, CO => 
                           carry_52_port, S => SUM(51));
   U1_50 : FA_X1 port map( A => A(50), B => B(50), CI => carry_50_port, CO => 
                           carry_51_port, S => SUM(50));
   U1_49 : FA_X1 port map( A => A(49), B => B(49), CI => carry_49_port, CO => 
                           carry_50_port, S => SUM(49));
   U1_48 : FA_X1 port map( A => A(48), B => B(48), CI => carry_48_port, CO => 
                           carry_49_port, S => SUM(48));
   U1_47 : FA_X1 port map( A => A(47), B => B(47), CI => carry_47_port, CO => 
                           carry_48_port, S => SUM(47));
   U1_46 : FA_X1 port map( A => A(46), B => B(46), CI => carry_46_port, CO => 
                           carry_47_port, S => SUM(46));
   U1_45 : FA_X1 port map( A => A(45), B => B(45), CI => carry_45_port, CO => 
                           carry_46_port, S => SUM(45));
   U1_44 : FA_X1 port map( A => A(44), B => B(44), CI => carry_44_port, CO => 
                           carry_45_port, S => SUM(44));
   U1_43 : FA_X1 port map( A => A(43), B => B(43), CI => carry_43_port, CO => 
                           carry_44_port, S => SUM(43));
   U1_42 : FA_X1 port map( A => A(42), B => B(42), CI => carry_42_port, CO => 
                           carry_43_port, S => SUM(42));
   U1_41 : FA_X1 port map( A => A(41), B => B(41), CI => carry_41_port, CO => 
                           carry_42_port, S => SUM(41));
   U1_40 : FA_X1 port map( A => A(40), B => B(40), CI => carry_40_port, CO => 
                           carry_41_port, S => SUM(40));
   U1_39 : FA_X1 port map( A => A(39), B => B(39), CI => carry_39_port, CO => 
                           carry_40_port, S => SUM(39));
   U1_38 : FA_X1 port map( A => A(38), B => B(38), CI => carry_38_port, CO => 
                           carry_39_port, S => SUM(38));
   U1_37 : FA_X1 port map( A => A(37), B => B(37), CI => carry_37_port, CO => 
                           carry_38_port, S => SUM(37));
   U1_36 : FA_X1 port map( A => A(36), B => B(36), CI => carry_36_port, CO => 
                           carry_37_port, S => SUM(36));
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => carry_35_port, CO => 
                           carry_36_port, S => SUM(35));
   U1_34 : FA_X1 port map( A => A(34), B => B(34), CI => carry_34_port, CO => 
                           carry_35_port, S => SUM(34));
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => carry_32_port, CO => 
                           carry_33_port, S => SUM(32));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity RCA_NBIT64_15_DW01_add_0 is

   port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (64 downto 0);  CO : out std_logic);

end RCA_NBIT64_15_DW01_add_0;

architecture SYN_rpl of RCA_NBIT64_15_DW01_add_0 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_63_port, carry_62_port, carry_61_port, carry_60_port, 
      carry_59_port, carry_58_port, carry_57_port, carry_56_port, carry_55_port
      , carry_54_port, carry_53_port, carry_52_port, carry_51_port, 
      carry_50_port, carry_49_port, carry_48_port, carry_47_port, carry_46_port
      , carry_45_port, carry_44_port, carry_43_port, carry_42_port, 
      carry_41_port, carry_40_port, carry_39_port, carry_38_port, carry_37_port
      , carry_36_port, carry_35_port, carry_34_port, carry_33_port, 
      carry_32_port, carry_31_port, carry_30_port, carry_29_port, carry_28_port
      , carry_27_port, carry_26_port, carry_25_port, carry_24_port, 
      carry_23_port, carry_22_port, carry_21_port, carry_20_port, carry_19_port
      , carry_18_port, carry_17_port, carry_16_port, carry_15_port, 
      carry_14_port, carry_13_port, carry_12_port, carry_11_port, carry_10_port
      , carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   U1_63 : FA_X1 port map( A => A(63), B => B(63), CI => carry_63_port, CO => 
                           SUM(64), S => SUM(63));
   U1_62 : FA_X1 port map( A => A(62), B => B(62), CI => carry_62_port, CO => 
                           carry_63_port, S => SUM(62));
   U1_61 : FA_X1 port map( A => A(61), B => B(61), CI => carry_61_port, CO => 
                           carry_62_port, S => SUM(61));
   U1_60 : FA_X1 port map( A => A(60), B => B(60), CI => carry_60_port, CO => 
                           carry_61_port, S => SUM(60));
   U1_59 : FA_X1 port map( A => A(59), B => B(59), CI => carry_59_port, CO => 
                           carry_60_port, S => SUM(59));
   U1_58 : FA_X1 port map( A => A(58), B => B(58), CI => carry_58_port, CO => 
                           carry_59_port, S => SUM(58));
   U1_57 : FA_X1 port map( A => A(57), B => B(57), CI => carry_57_port, CO => 
                           carry_58_port, S => SUM(57));
   U1_56 : FA_X1 port map( A => A(56), B => B(56), CI => carry_56_port, CO => 
                           carry_57_port, S => SUM(56));
   U1_55 : FA_X1 port map( A => A(55), B => B(55), CI => carry_55_port, CO => 
                           carry_56_port, S => SUM(55));
   U1_54 : FA_X1 port map( A => A(54), B => B(54), CI => carry_54_port, CO => 
                           carry_55_port, S => SUM(54));
   U1_53 : FA_X1 port map( A => A(53), B => B(53), CI => carry_53_port, CO => 
                           carry_54_port, S => SUM(53));
   U1_52 : FA_X1 port map( A => A(52), B => B(52), CI => carry_52_port, CO => 
                           carry_53_port, S => SUM(52));
   U1_51 : FA_X1 port map( A => A(51), B => B(51), CI => carry_51_port, CO => 
                           carry_52_port, S => SUM(51));
   U1_50 : FA_X1 port map( A => A(50), B => B(50), CI => carry_50_port, CO => 
                           carry_51_port, S => SUM(50));
   U1_49 : FA_X1 port map( A => A(49), B => B(49), CI => carry_49_port, CO => 
                           carry_50_port, S => SUM(49));
   U1_48 : FA_X1 port map( A => A(48), B => B(48), CI => carry_48_port, CO => 
                           carry_49_port, S => SUM(48));
   U1_47 : FA_X1 port map( A => A(47), B => B(47), CI => carry_47_port, CO => 
                           carry_48_port, S => SUM(47));
   U1_46 : FA_X1 port map( A => A(46), B => B(46), CI => carry_46_port, CO => 
                           carry_47_port, S => SUM(46));
   U1_45 : FA_X1 port map( A => A(45), B => B(45), CI => carry_45_port, CO => 
                           carry_46_port, S => SUM(45));
   U1_44 : FA_X1 port map( A => A(44), B => B(44), CI => carry_44_port, CO => 
                           carry_45_port, S => SUM(44));
   U1_43 : FA_X1 port map( A => A(43), B => B(43), CI => carry_43_port, CO => 
                           carry_44_port, S => SUM(43));
   U1_42 : FA_X1 port map( A => A(42), B => B(42), CI => carry_42_port, CO => 
                           carry_43_port, S => SUM(42));
   U1_41 : FA_X1 port map( A => A(41), B => B(41), CI => carry_41_port, CO => 
                           carry_42_port, S => SUM(41));
   U1_40 : FA_X1 port map( A => A(40), B => B(40), CI => carry_40_port, CO => 
                           carry_41_port, S => SUM(40));
   U1_39 : FA_X1 port map( A => A(39), B => B(39), CI => carry_39_port, CO => 
                           carry_40_port, S => SUM(39));
   U1_38 : FA_X1 port map( A => A(38), B => B(38), CI => carry_38_port, CO => 
                           carry_39_port, S => SUM(38));
   U1_37 : FA_X1 port map( A => A(37), B => B(37), CI => carry_37_port, CO => 
                           carry_38_port, S => SUM(37));
   U1_36 : FA_X1 port map( A => A(36), B => B(36), CI => carry_36_port, CO => 
                           carry_37_port, S => SUM(36));
   U1_35 : FA_X1 port map( A => A(35), B => B(35), CI => carry_35_port, CO => 
                           carry_36_port, S => SUM(35));
   U1_34 : FA_X1 port map( A => A(34), B => B(34), CI => carry_34_port, CO => 
                           carry_35_port, S => SUM(34));
   U1_33 : FA_X1 port map( A => A(33), B => B(33), CI => carry_33_port, CO => 
                           carry_34_port, S => SUM(33));
   U1_32 : FA_X1 port map( A => A(32), B => B(32), CI => carry_32_port, CO => 
                           carry_33_port, S => SUM(32));
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           carry_32_port, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1_0 : FA_X1 port map( A => A(0), B => B(0), CI => CI, CO => carry_1_port, S
                           => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity BOOTHMUL_NBIT32_1_DW01_sub_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end BOOTHMUL_NBIT32_1_DW01_sub_0;

architecture SYN_rpl of BOOTHMUL_NBIT32_1_DW01_sub_0 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal DIFF_1_port, DIFF_2_port, DIFF_3_port, DIFF_4_port, DIFF_5_port, 
      DIFF_6_port, DIFF_7_port, DIFF_9_port, DIFF_10_port, DIFF_11_port, 
      DIFF_12_port, DIFF_13_port, DIFF_14_port, DIFF_15_port, DIFF_16_port, 
      DIFF_17_port, DIFF_18_port, DIFF_19_port, DIFF_20_port, DIFF_21_port, 
      DIFF_22_port, DIFF_23_port, DIFF_24_port, DIFF_25_port, DIFF_26_port, 
      DIFF_27_port, DIFF_28_port, DIFF_29_port, DIFF_30_port, DIFF_8_port, n96,
      n97, n98, n99, n101, n102, n103, n104, n105, n106, n107, n108, n110, n111
      , n112, n114, n115, n116, n118, n119, n120, n122, n123, n94, DIFF_31_port
      , n100, n109, n113, n117, n121, n124, n125, n126 : std_logic;

begin
   DIFF <= ( DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, 
      DIFF_2_port, DIFF_1_port, B(0) );
   
   U42 : XOR2_X1 port map( A => n97, B => B(9), Z => DIFF_9_port);
   U43 : XOR2_X1 port map( A => n99, B => B(7), Z => DIFF_7_port);
   U45 : XOR2_X1 port map( A => n101, B => B(5), Z => DIFF_5_port);
   U46 : XOR2_X1 port map( A => n103, B => B(3), Z => DIFF_3_port);
   U47 : XOR2_X1 port map( A => n96, B => B(30), Z => DIFF_30_port);
   U48 : XOR2_X1 port map( A => n106, B => B(27), Z => DIFF_27_port);
   U50 : XOR2_X1 port map( A => n108, B => B(25), Z => DIFF_25_port);
   U51 : XOR2_X1 port map( A => n110, B => B(23), Z => DIFF_23_port);
   U53 : XOR2_X1 port map( A => n112, B => B(21), Z => DIFF_21_port);
   U54 : XOR2_X1 port map( A => B(1), B => B(0), Z => DIFF_1_port);
   U55 : XOR2_X1 port map( A => n114, B => B(19), Z => DIFF_19_port);
   U57 : XOR2_X1 port map( A => n116, B => B(17), Z => DIFF_17_port);
   U58 : XOR2_X1 port map( A => n118, B => B(15), Z => DIFF_15_port);
   U60 : XOR2_X1 port map( A => n120, B => B(13), Z => DIFF_13_port);
   U61 : XOR2_X1 port map( A => n122, B => B(11), Z => DIFF_11_port);
   U1 : XOR2_X1 port map( A => n100, B => B(31), Z => n94);
   U2 : INV_X2 port map( A => n94, ZN => DIFF_31_port);
   U3 : NOR2_X1 port map( A1 => n96, A2 => B(30), ZN => n100);
   U4 : NOR3_X1 port map( A1 => B(27), A2 => B(28), A3 => n106, ZN => n104);
   U5 : NAND2_X1 port map( A1 => n104, A2 => n126, ZN => n96);
   U6 : INV_X1 port map( A => B(29), ZN => n126);
   U7 : OR3_X1 port map( A1 => B(25), A2 => B(26), A3 => n108, ZN => n106);
   U8 : OR3_X1 port map( A1 => B(1), A2 => B(2), A3 => B(0), ZN => n103);
   U9 : OR3_X1 port map( A1 => B(5), A2 => B(6), A3 => n101, ZN => n99);
   U10 : OR3_X1 port map( A1 => B(10), A2 => B(9), A3 => n97, ZN => n122);
   U11 : OR3_X1 port map( A1 => B(13), A2 => B(14), A3 => n120, ZN => n118);
   U12 : OR3_X1 port map( A1 => B(17), A2 => B(18), A3 => n116, ZN => n114);
   U13 : OR3_X1 port map( A1 => B(21), A2 => B(22), A3 => n112, ZN => n110);
   U14 : OR3_X1 port map( A1 => B(3), A2 => B(4), A3 => n103, ZN => n101);
   U15 : OR3_X1 port map( A1 => B(7), A2 => B(8), A3 => n99, ZN => n97);
   U16 : OR3_X1 port map( A1 => B(11), A2 => B(12), A3 => n122, ZN => n120);
   U17 : OR3_X1 port map( A1 => B(15), A2 => B(16), A3 => n118, ZN => n116);
   U18 : OR3_X1 port map( A1 => B(19), A2 => B(20), A3 => n114, ZN => n112);
   U19 : OR3_X1 port map( A1 => B(23), A2 => B(24), A3 => n110, ZN => n108);
   U20 : XNOR2_X1 port map( A => n104, B => B(29), ZN => DIFF_29_port);
   U21 : XNOR2_X1 port map( A => n109, B => B(6), ZN => DIFF_6_port);
   U22 : NOR2_X1 port map( A1 => n101, A2 => B(5), ZN => n109);
   U23 : XNOR2_X1 port map( A => n113, B => B(10), ZN => DIFF_10_port);
   U24 : NOR2_X1 port map( A1 => n97, A2 => B(9), ZN => n113);
   U25 : XNOR2_X1 port map( A => n117, B => B(14), ZN => DIFF_14_port);
   U26 : NOR2_X1 port map( A1 => n120, A2 => B(13), ZN => n117);
   U27 : XNOR2_X1 port map( A => n121, B => B(18), ZN => DIFF_18_port);
   U28 : NOR2_X1 port map( A1 => n116, A2 => B(17), ZN => n121);
   U29 : XNOR2_X1 port map( A => n124, B => B(22), ZN => DIFF_22_port);
   U30 : NOR2_X1 port map( A1 => n112, A2 => B(21), ZN => n124);
   U31 : XNOR2_X1 port map( A => n125, B => B(26), ZN => DIFF_26_port);
   U32 : NOR2_X1 port map( A1 => n108, A2 => B(25), ZN => n125);
   U33 : XNOR2_X1 port map( A => B(2), B => n105, ZN => DIFF_2_port);
   U34 : NOR2_X1 port map( A1 => B(0), A2 => B(1), ZN => n105);
   U35 : XNOR2_X1 port map( A => B(4), B => n102, ZN => DIFF_4_port);
   U36 : NOR2_X1 port map( A1 => B(3), A2 => n103, ZN => n102);
   U37 : XNOR2_X1 port map( A => B(12), B => n123, ZN => DIFF_12_port);
   U38 : NOR2_X1 port map( A1 => B(11), A2 => n122, ZN => n123);
   U39 : XNOR2_X1 port map( A => B(16), B => n119, ZN => DIFF_16_port);
   U40 : NOR2_X1 port map( A1 => B(15), A2 => n118, ZN => n119);
   U41 : XNOR2_X1 port map( A => B(20), B => n115, ZN => DIFF_20_port);
   U44 : NOR2_X1 port map( A1 => B(19), A2 => n114, ZN => n115);
   U49 : XNOR2_X1 port map( A => B(24), B => n111, ZN => DIFF_24_port);
   U52 : NOR2_X1 port map( A1 => B(23), A2 => n110, ZN => n111);
   U56 : XNOR2_X1 port map( A => B(28), B => n107, ZN => DIFF_28_port);
   U59 : NOR2_X1 port map( A1 => B(27), A2 => n106, ZN => n107);
   U62 : XNOR2_X1 port map( A => B(8), B => n98, ZN => DIFF_8_port);
   U63 : NOR2_X1 port map( A1 => B(7), A2 => n99, ZN => n98);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity RCA_NBIT64_16 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_16;

architecture SYN_BEHAVIORAL of RCA_NBIT64_16 is

   component RCA_NBIT64_16_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1079 : std_logic;

begin
   
   n1 <= '0';
   add_1_root_add_81_2 : RCA_NBIT64_16_DW01_add_0 port map( A(64) => n1, A(63) 
                           => A(63), A(62) => A(62), A(61) => A(61), A(60) => 
                           A(60), A(59) => A(59), A(58) => A(58), A(57) => 
                           A(57), A(56) => A(56), A(55) => A(55), A(54) => 
                           A(54), A(53) => A(53), A(52) => A(52), A(51) => 
                           A(51), A(50) => A(50), A(49) => A(49), A(48) => 
                           A(48), A(47) => A(47), A(46) => A(46), A(45) => 
                           A(45), A(44) => A(44), A(43) => A(43), A(42) => 
                           A(42), A(41) => A(41), A(40) => A(40), A(39) => 
                           A(39), A(38) => A(38), A(37) => A(37), A(36) => 
                           A(36), A(35) => A(35), A(34) => A(34), A(33) => 
                           A(33), A(32) => A(32), A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(64) => n1, B(63) => B(63), 
                           B(62) => B(62), B(61) => B(61), B(60) => B(60), 
                           B(59) => B(59), B(58) => B(58), B(57) => B(57), 
                           B(56) => B(56), B(55) => B(55), B(54) => B(54), 
                           B(53) => B(53), B(52) => B(52), B(51) => B(51), 
                           B(50) => B(50), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, SUM(63)
                           => S(63), SUM(62) => S(62), SUM(61) => S(61), 
                           SUM(60) => S(60), SUM(59) => S(59), SUM(58) => S(58)
                           , SUM(57) => S(57), SUM(56) => S(56), SUM(55) => 
                           S(55), SUM(54) => S(54), SUM(53) => S(53), SUM(52) 
                           => S(52), SUM(51) => S(51), SUM(50) => S(50), 
                           SUM(49) => S(49), SUM(48) => S(48), SUM(47) => S(47)
                           , SUM(46) => S(46), SUM(45) => S(45), SUM(44) => 
                           S(44), SUM(43) => S(43), SUM(42) => S(42), SUM(41) 
                           => S(41), SUM(40) => S(40), SUM(39) => S(39), 
                           SUM(38) => S(38), SUM(37) => S(37), SUM(36) => S(36)
                           , SUM(35) => S(35), SUM(34) => S(34), SUM(33) => 
                           S(33), SUM(32) => S(32), SUM(31) => S(31), SUM(30) 
                           => S(30), SUM(29) => S(29), SUM(28) => S(28), 
                           SUM(27) => S(27), SUM(26) => S(26), SUM(25) => S(25)
                           , SUM(24) => S(24), SUM(23) => S(23), SUM(22) => 
                           S(22), SUM(21) => S(21), SUM(20) => S(20), SUM(19) 
                           => S(19), SUM(18) => S(18), SUM(17) => S(17), 
                           SUM(16) => S(16), SUM(15) => S(15), SUM(14) => S(14)
                           , SUM(13) => S(13), SUM(12) => S(12), SUM(11) => 
                           S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) => 
                           S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5)
                           , SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1079);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity RCA_NBIT64_17 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_17;

architecture SYN_BEHAVIORAL of RCA_NBIT64_17 is

   component RCA_NBIT64_17_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1080 : std_logic;

begin
   
   n1 <= '0';
   add_1_root_add_81_2 : RCA_NBIT64_17_DW01_add_0 port map( A(64) => n1, A(63) 
                           => A(63), A(62) => A(62), A(61) => A(61), A(60) => 
                           A(60), A(59) => A(59), A(58) => A(58), A(57) => 
                           A(57), A(56) => A(56), A(55) => A(55), A(54) => 
                           A(54), A(53) => A(53), A(52) => A(52), A(51) => 
                           A(51), A(50) => A(50), A(49) => A(49), A(48) => 
                           A(48), A(47) => A(47), A(46) => A(46), A(45) => 
                           A(45), A(44) => A(44), A(43) => A(43), A(42) => 
                           A(42), A(41) => A(41), A(40) => A(40), A(39) => 
                           A(39), A(38) => A(38), A(37) => A(37), A(36) => 
                           A(36), A(35) => A(35), A(34) => A(34), A(33) => 
                           A(33), A(32) => A(32), A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(64) => n1, B(63) => B(63), 
                           B(62) => B(62), B(61) => B(61), B(60) => B(60), 
                           B(59) => B(59), B(58) => B(58), B(57) => B(57), 
                           B(56) => B(56), B(55) => B(55), B(54) => B(54), 
                           B(53) => B(53), B(52) => B(52), B(51) => B(51), 
                           B(50) => B(50), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, SUM(63)
                           => S(63), SUM(62) => S(62), SUM(61) => S(61), 
                           SUM(60) => S(60), SUM(59) => S(59), SUM(58) => S(58)
                           , SUM(57) => S(57), SUM(56) => S(56), SUM(55) => 
                           S(55), SUM(54) => S(54), SUM(53) => S(53), SUM(52) 
                           => S(52), SUM(51) => S(51), SUM(50) => S(50), 
                           SUM(49) => S(49), SUM(48) => S(48), SUM(47) => S(47)
                           , SUM(46) => S(46), SUM(45) => S(45), SUM(44) => 
                           S(44), SUM(43) => S(43), SUM(42) => S(42), SUM(41) 
                           => S(41), SUM(40) => S(40), SUM(39) => S(39), 
                           SUM(38) => S(38), SUM(37) => S(37), SUM(36) => S(36)
                           , SUM(35) => S(35), SUM(34) => S(34), SUM(33) => 
                           S(33), SUM(32) => S(32), SUM(31) => S(31), SUM(30) 
                           => S(30), SUM(29) => S(29), SUM(28) => S(28), 
                           SUM(27) => S(27), SUM(26) => S(26), SUM(25) => S(25)
                           , SUM(24) => S(24), SUM(23) => S(23), SUM(22) => 
                           S(22), SUM(21) => S(21), SUM(20) => S(20), SUM(19) 
                           => S(19), SUM(18) => S(18), SUM(17) => S(17), 
                           SUM(16) => S(16), SUM(15) => S(15), SUM(14) => S(14)
                           , SUM(13) => S(13), SUM(12) => S(12), SUM(11) => 
                           S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) => 
                           S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5)
                           , SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1080);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity RCA_NBIT64_18 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_18;

architecture SYN_BEHAVIORAL of RCA_NBIT64_18 is

   component RCA_NBIT64_18_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1081 : std_logic;

begin
   
   n1 <= '0';
   add_1_root_add_81_2 : RCA_NBIT64_18_DW01_add_0 port map( A(64) => n1, A(63) 
                           => A(63), A(62) => A(62), A(61) => A(61), A(60) => 
                           A(60), A(59) => A(59), A(58) => A(58), A(57) => 
                           A(57), A(56) => A(56), A(55) => A(55), A(54) => 
                           A(54), A(53) => A(53), A(52) => A(52), A(51) => 
                           A(51), A(50) => A(50), A(49) => A(49), A(48) => 
                           A(48), A(47) => A(47), A(46) => A(46), A(45) => 
                           A(45), A(44) => A(44), A(43) => A(43), A(42) => 
                           A(42), A(41) => A(41), A(40) => A(40), A(39) => 
                           A(39), A(38) => A(38), A(37) => A(37), A(36) => 
                           A(36), A(35) => A(35), A(34) => A(34), A(33) => 
                           A(33), A(32) => A(32), A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(64) => n1, B(63) => B(63), 
                           B(62) => B(62), B(61) => B(61), B(60) => B(60), 
                           B(59) => B(59), B(58) => B(58), B(57) => B(57), 
                           B(56) => B(56), B(55) => B(55), B(54) => B(54), 
                           B(53) => B(53), B(52) => B(52), B(51) => B(51), 
                           B(50) => B(50), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, SUM(63)
                           => S(63), SUM(62) => S(62), SUM(61) => S(61), 
                           SUM(60) => S(60), SUM(59) => S(59), SUM(58) => S(58)
                           , SUM(57) => S(57), SUM(56) => S(56), SUM(55) => 
                           S(55), SUM(54) => S(54), SUM(53) => S(53), SUM(52) 
                           => S(52), SUM(51) => S(51), SUM(50) => S(50), 
                           SUM(49) => S(49), SUM(48) => S(48), SUM(47) => S(47)
                           , SUM(46) => S(46), SUM(45) => S(45), SUM(44) => 
                           S(44), SUM(43) => S(43), SUM(42) => S(42), SUM(41) 
                           => S(41), SUM(40) => S(40), SUM(39) => S(39), 
                           SUM(38) => S(38), SUM(37) => S(37), SUM(36) => S(36)
                           , SUM(35) => S(35), SUM(34) => S(34), SUM(33) => 
                           S(33), SUM(32) => S(32), SUM(31) => S(31), SUM(30) 
                           => S(30), SUM(29) => S(29), SUM(28) => S(28), 
                           SUM(27) => S(27), SUM(26) => S(26), SUM(25) => S(25)
                           , SUM(24) => S(24), SUM(23) => S(23), SUM(22) => 
                           S(22), SUM(21) => S(21), SUM(20) => S(20), SUM(19) 
                           => S(19), SUM(18) => S(18), SUM(17) => S(17), 
                           SUM(16) => S(16), SUM(15) => S(15), SUM(14) => S(14)
                           , SUM(13) => S(13), SUM(12) => S(12), SUM(11) => 
                           S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) => 
                           S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5)
                           , SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1081);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity RCA_NBIT64_19 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_19;

architecture SYN_BEHAVIORAL of RCA_NBIT64_19 is

   component RCA_NBIT64_19_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1082 : std_logic;

begin
   
   n1 <= '0';
   add_1_root_add_81_2 : RCA_NBIT64_19_DW01_add_0 port map( A(64) => n1, A(63) 
                           => A(63), A(62) => A(62), A(61) => A(61), A(60) => 
                           A(60), A(59) => A(59), A(58) => A(58), A(57) => 
                           A(57), A(56) => A(56), A(55) => A(55), A(54) => 
                           A(54), A(53) => A(53), A(52) => A(52), A(51) => 
                           A(51), A(50) => A(50), A(49) => A(49), A(48) => 
                           A(48), A(47) => A(47), A(46) => A(46), A(45) => 
                           A(45), A(44) => A(44), A(43) => A(43), A(42) => 
                           A(42), A(41) => A(41), A(40) => A(40), A(39) => 
                           A(39), A(38) => A(38), A(37) => A(37), A(36) => 
                           A(36), A(35) => A(35), A(34) => A(34), A(33) => 
                           A(33), A(32) => A(32), A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(64) => n1, B(63) => B(63), 
                           B(62) => B(62), B(61) => B(61), B(60) => B(60), 
                           B(59) => B(59), B(58) => B(58), B(57) => B(57), 
                           B(56) => B(56), B(55) => B(55), B(54) => B(54), 
                           B(53) => B(53), B(52) => B(52), B(51) => B(51), 
                           B(50) => B(50), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, SUM(63)
                           => S(63), SUM(62) => S(62), SUM(61) => S(61), 
                           SUM(60) => S(60), SUM(59) => S(59), SUM(58) => S(58)
                           , SUM(57) => S(57), SUM(56) => S(56), SUM(55) => 
                           S(55), SUM(54) => S(54), SUM(53) => S(53), SUM(52) 
                           => S(52), SUM(51) => S(51), SUM(50) => S(50), 
                           SUM(49) => S(49), SUM(48) => S(48), SUM(47) => S(47)
                           , SUM(46) => S(46), SUM(45) => S(45), SUM(44) => 
                           S(44), SUM(43) => S(43), SUM(42) => S(42), SUM(41) 
                           => S(41), SUM(40) => S(40), SUM(39) => S(39), 
                           SUM(38) => S(38), SUM(37) => S(37), SUM(36) => S(36)
                           , SUM(35) => S(35), SUM(34) => S(34), SUM(33) => 
                           S(33), SUM(32) => S(32), SUM(31) => S(31), SUM(30) 
                           => S(30), SUM(29) => S(29), SUM(28) => S(28), 
                           SUM(27) => S(27), SUM(26) => S(26), SUM(25) => S(25)
                           , SUM(24) => S(24), SUM(23) => S(23), SUM(22) => 
                           S(22), SUM(21) => S(21), SUM(20) => S(20), SUM(19) 
                           => S(19), SUM(18) => S(18), SUM(17) => S(17), 
                           SUM(16) => S(16), SUM(15) => S(15), SUM(14) => S(14)
                           , SUM(13) => S(13), SUM(12) => S(12), SUM(11) => 
                           S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) => 
                           S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5)
                           , SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1082);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity RCA_NBIT64_20 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_20;

architecture SYN_BEHAVIORAL of RCA_NBIT64_20 is

   component RCA_NBIT64_20_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1083 : std_logic;

begin
   
   n1 <= '0';
   add_1_root_add_81_2 : RCA_NBIT64_20_DW01_add_0 port map( A(64) => n1, A(63) 
                           => A(63), A(62) => A(62), A(61) => A(61), A(60) => 
                           A(60), A(59) => A(59), A(58) => A(58), A(57) => 
                           A(57), A(56) => A(56), A(55) => A(55), A(54) => 
                           A(54), A(53) => A(53), A(52) => A(52), A(51) => 
                           A(51), A(50) => A(50), A(49) => A(49), A(48) => 
                           A(48), A(47) => A(47), A(46) => A(46), A(45) => 
                           A(45), A(44) => A(44), A(43) => A(43), A(42) => 
                           A(42), A(41) => A(41), A(40) => A(40), A(39) => 
                           A(39), A(38) => A(38), A(37) => A(37), A(36) => 
                           A(36), A(35) => A(35), A(34) => A(34), A(33) => 
                           A(33), A(32) => A(32), A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(64) => n1, B(63) => B(63), 
                           B(62) => B(62), B(61) => B(61), B(60) => B(60), 
                           B(59) => B(59), B(58) => B(58), B(57) => B(57), 
                           B(56) => B(56), B(55) => B(55), B(54) => B(54), 
                           B(53) => B(53), B(52) => B(52), B(51) => B(51), 
                           B(50) => B(50), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, SUM(63)
                           => S(63), SUM(62) => S(62), SUM(61) => S(61), 
                           SUM(60) => S(60), SUM(59) => S(59), SUM(58) => S(58)
                           , SUM(57) => S(57), SUM(56) => S(56), SUM(55) => 
                           S(55), SUM(54) => S(54), SUM(53) => S(53), SUM(52) 
                           => S(52), SUM(51) => S(51), SUM(50) => S(50), 
                           SUM(49) => S(49), SUM(48) => S(48), SUM(47) => S(47)
                           , SUM(46) => S(46), SUM(45) => S(45), SUM(44) => 
                           S(44), SUM(43) => S(43), SUM(42) => S(42), SUM(41) 
                           => S(41), SUM(40) => S(40), SUM(39) => S(39), 
                           SUM(38) => S(38), SUM(37) => S(37), SUM(36) => S(36)
                           , SUM(35) => S(35), SUM(34) => S(34), SUM(33) => 
                           S(33), SUM(32) => S(32), SUM(31) => S(31), SUM(30) 
                           => S(30), SUM(29) => S(29), SUM(28) => S(28), 
                           SUM(27) => S(27), SUM(26) => S(26), SUM(25) => S(25)
                           , SUM(24) => S(24), SUM(23) => S(23), SUM(22) => 
                           S(22), SUM(21) => S(21), SUM(20) => S(20), SUM(19) 
                           => S(19), SUM(18) => S(18), SUM(17) => S(17), 
                           SUM(16) => S(16), SUM(15) => S(15), SUM(14) => S(14)
                           , SUM(13) => S(13), SUM(12) => S(12), SUM(11) => 
                           S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) => 
                           S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5)
                           , SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1083);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity RCA_NBIT64_21 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_21;

architecture SYN_BEHAVIORAL of RCA_NBIT64_21 is

   component RCA_NBIT64_21_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1084 : std_logic;

begin
   
   n1 <= '0';
   add_1_root_add_81_2 : RCA_NBIT64_21_DW01_add_0 port map( A(64) => n1, A(63) 
                           => A(63), A(62) => A(62), A(61) => A(61), A(60) => 
                           A(60), A(59) => A(59), A(58) => A(58), A(57) => 
                           A(57), A(56) => A(56), A(55) => A(55), A(54) => 
                           A(54), A(53) => A(53), A(52) => A(52), A(51) => 
                           A(51), A(50) => A(50), A(49) => A(49), A(48) => 
                           A(48), A(47) => A(47), A(46) => A(46), A(45) => 
                           A(45), A(44) => A(44), A(43) => A(43), A(42) => 
                           A(42), A(41) => A(41), A(40) => A(40), A(39) => 
                           A(39), A(38) => A(38), A(37) => A(37), A(36) => 
                           A(36), A(35) => A(35), A(34) => A(34), A(33) => 
                           A(33), A(32) => A(32), A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(64) => n1, B(63) => B(63), 
                           B(62) => B(62), B(61) => B(61), B(60) => B(60), 
                           B(59) => B(59), B(58) => B(58), B(57) => B(57), 
                           B(56) => B(56), B(55) => B(55), B(54) => B(54), 
                           B(53) => B(53), B(52) => B(52), B(51) => B(51), 
                           B(50) => B(50), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, SUM(63)
                           => S(63), SUM(62) => S(62), SUM(61) => S(61), 
                           SUM(60) => S(60), SUM(59) => S(59), SUM(58) => S(58)
                           , SUM(57) => S(57), SUM(56) => S(56), SUM(55) => 
                           S(55), SUM(54) => S(54), SUM(53) => S(53), SUM(52) 
                           => S(52), SUM(51) => S(51), SUM(50) => S(50), 
                           SUM(49) => S(49), SUM(48) => S(48), SUM(47) => S(47)
                           , SUM(46) => S(46), SUM(45) => S(45), SUM(44) => 
                           S(44), SUM(43) => S(43), SUM(42) => S(42), SUM(41) 
                           => S(41), SUM(40) => S(40), SUM(39) => S(39), 
                           SUM(38) => S(38), SUM(37) => S(37), SUM(36) => S(36)
                           , SUM(35) => S(35), SUM(34) => S(34), SUM(33) => 
                           S(33), SUM(32) => S(32), SUM(31) => S(31), SUM(30) 
                           => S(30), SUM(29) => S(29), SUM(28) => S(28), 
                           SUM(27) => S(27), SUM(26) => S(26), SUM(25) => S(25)
                           , SUM(24) => S(24), SUM(23) => S(23), SUM(22) => 
                           S(22), SUM(21) => S(21), SUM(20) => S(20), SUM(19) 
                           => S(19), SUM(18) => S(18), SUM(17) => S(17), 
                           SUM(16) => S(16), SUM(15) => S(15), SUM(14) => S(14)
                           , SUM(13) => S(13), SUM(12) => S(12), SUM(11) => 
                           S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) => 
                           S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5)
                           , SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1084);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity RCA_NBIT64_22 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_22;

architecture SYN_BEHAVIORAL of RCA_NBIT64_22 is

   component RCA_NBIT64_22_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1085 : std_logic;

begin
   
   n1 <= '0';
   add_1_root_add_81_2 : RCA_NBIT64_22_DW01_add_0 port map( A(64) => n1, A(63) 
                           => A(63), A(62) => A(62), A(61) => A(61), A(60) => 
                           A(60), A(59) => A(59), A(58) => A(58), A(57) => 
                           A(57), A(56) => A(56), A(55) => A(55), A(54) => 
                           A(54), A(53) => A(53), A(52) => A(52), A(51) => 
                           A(51), A(50) => A(50), A(49) => A(49), A(48) => 
                           A(48), A(47) => A(47), A(46) => A(46), A(45) => 
                           A(45), A(44) => A(44), A(43) => A(43), A(42) => 
                           A(42), A(41) => A(41), A(40) => A(40), A(39) => 
                           A(39), A(38) => A(38), A(37) => A(37), A(36) => 
                           A(36), A(35) => A(35), A(34) => A(34), A(33) => 
                           A(33), A(32) => A(32), A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(64) => n1, B(63) => B(63), 
                           B(62) => B(62), B(61) => B(61), B(60) => B(60), 
                           B(59) => B(59), B(58) => B(58), B(57) => B(57), 
                           B(56) => B(56), B(55) => B(55), B(54) => B(54), 
                           B(53) => B(53), B(52) => B(52), B(51) => B(51), 
                           B(50) => B(50), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, SUM(63)
                           => S(63), SUM(62) => S(62), SUM(61) => S(61), 
                           SUM(60) => S(60), SUM(59) => S(59), SUM(58) => S(58)
                           , SUM(57) => S(57), SUM(56) => S(56), SUM(55) => 
                           S(55), SUM(54) => S(54), SUM(53) => S(53), SUM(52) 
                           => S(52), SUM(51) => S(51), SUM(50) => S(50), 
                           SUM(49) => S(49), SUM(48) => S(48), SUM(47) => S(47)
                           , SUM(46) => S(46), SUM(45) => S(45), SUM(44) => 
                           S(44), SUM(43) => S(43), SUM(42) => S(42), SUM(41) 
                           => S(41), SUM(40) => S(40), SUM(39) => S(39), 
                           SUM(38) => S(38), SUM(37) => S(37), SUM(36) => S(36)
                           , SUM(35) => S(35), SUM(34) => S(34), SUM(33) => 
                           S(33), SUM(32) => S(32), SUM(31) => S(31), SUM(30) 
                           => S(30), SUM(29) => S(29), SUM(28) => S(28), 
                           SUM(27) => S(27), SUM(26) => S(26), SUM(25) => S(25)
                           , SUM(24) => S(24), SUM(23) => S(23), SUM(22) => 
                           S(22), SUM(21) => S(21), SUM(20) => S(20), SUM(19) 
                           => S(19), SUM(18) => S(18), SUM(17) => S(17), 
                           SUM(16) => S(16), SUM(15) => S(15), SUM(14) => S(14)
                           , SUM(13) => S(13), SUM(12) => S(12), SUM(11) => 
                           S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) => 
                           S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5)
                           , SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1085);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity RCA_NBIT64_23 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_23;

architecture SYN_BEHAVIORAL of RCA_NBIT64_23 is

   component RCA_NBIT64_23_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1086 : std_logic;

begin
   
   n1 <= '0';
   add_1_root_add_81_2 : RCA_NBIT64_23_DW01_add_0 port map( A(64) => n1, A(63) 
                           => A(63), A(62) => A(62), A(61) => A(61), A(60) => 
                           A(60), A(59) => A(59), A(58) => A(58), A(57) => 
                           A(57), A(56) => A(56), A(55) => A(55), A(54) => 
                           A(54), A(53) => A(53), A(52) => A(52), A(51) => 
                           A(51), A(50) => A(50), A(49) => A(49), A(48) => 
                           A(48), A(47) => A(47), A(46) => A(46), A(45) => 
                           A(45), A(44) => A(44), A(43) => A(43), A(42) => 
                           A(42), A(41) => A(41), A(40) => A(40), A(39) => 
                           A(39), A(38) => A(38), A(37) => A(37), A(36) => 
                           A(36), A(35) => A(35), A(34) => A(34), A(33) => 
                           A(33), A(32) => A(32), A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(64) => n1, B(63) => B(63), 
                           B(62) => B(62), B(61) => B(61), B(60) => B(60), 
                           B(59) => B(59), B(58) => B(58), B(57) => B(57), 
                           B(56) => B(56), B(55) => B(55), B(54) => B(54), 
                           B(53) => B(53), B(52) => B(52), B(51) => B(51), 
                           B(50) => B(50), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, SUM(63)
                           => S(63), SUM(62) => S(62), SUM(61) => S(61), 
                           SUM(60) => S(60), SUM(59) => S(59), SUM(58) => S(58)
                           , SUM(57) => S(57), SUM(56) => S(56), SUM(55) => 
                           S(55), SUM(54) => S(54), SUM(53) => S(53), SUM(52) 
                           => S(52), SUM(51) => S(51), SUM(50) => S(50), 
                           SUM(49) => S(49), SUM(48) => S(48), SUM(47) => S(47)
                           , SUM(46) => S(46), SUM(45) => S(45), SUM(44) => 
                           S(44), SUM(43) => S(43), SUM(42) => S(42), SUM(41) 
                           => S(41), SUM(40) => S(40), SUM(39) => S(39), 
                           SUM(38) => S(38), SUM(37) => S(37), SUM(36) => S(36)
                           , SUM(35) => S(35), SUM(34) => S(34), SUM(33) => 
                           S(33), SUM(32) => S(32), SUM(31) => S(31), SUM(30) 
                           => S(30), SUM(29) => S(29), SUM(28) => S(28), 
                           SUM(27) => S(27), SUM(26) => S(26), SUM(25) => S(25)
                           , SUM(24) => S(24), SUM(23) => S(23), SUM(22) => 
                           S(22), SUM(21) => S(21), SUM(20) => S(20), SUM(19) 
                           => S(19), SUM(18) => S(18), SUM(17) => S(17), 
                           SUM(16) => S(16), SUM(15) => S(15), SUM(14) => S(14)
                           , SUM(13) => S(13), SUM(12) => S(12), SUM(11) => 
                           S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) => 
                           S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5)
                           , SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1086);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity RCA_NBIT64_24 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_24;

architecture SYN_BEHAVIORAL of RCA_NBIT64_24 is

   component RCA_NBIT64_24_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1087 : std_logic;

begin
   
   n1 <= '0';
   add_1_root_add_81_2 : RCA_NBIT64_24_DW01_add_0 port map( A(64) => n1, A(63) 
                           => A(63), A(62) => A(62), A(61) => A(61), A(60) => 
                           A(60), A(59) => A(59), A(58) => A(58), A(57) => 
                           A(57), A(56) => A(56), A(55) => A(55), A(54) => 
                           A(54), A(53) => A(53), A(52) => A(52), A(51) => 
                           A(51), A(50) => A(50), A(49) => A(49), A(48) => 
                           A(48), A(47) => A(47), A(46) => A(46), A(45) => 
                           A(45), A(44) => A(44), A(43) => A(43), A(42) => 
                           A(42), A(41) => A(41), A(40) => A(40), A(39) => 
                           A(39), A(38) => A(38), A(37) => A(37), A(36) => 
                           A(36), A(35) => A(35), A(34) => A(34), A(33) => 
                           A(33), A(32) => A(32), A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(64) => n1, B(63) => B(63), 
                           B(62) => B(62), B(61) => B(61), B(60) => B(60), 
                           B(59) => B(59), B(58) => B(58), B(57) => B(57), 
                           B(56) => B(56), B(55) => B(55), B(54) => B(54), 
                           B(53) => B(53), B(52) => B(52), B(51) => B(51), 
                           B(50) => B(50), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, SUM(63)
                           => S(63), SUM(62) => S(62), SUM(61) => S(61), 
                           SUM(60) => S(60), SUM(59) => S(59), SUM(58) => S(58)
                           , SUM(57) => S(57), SUM(56) => S(56), SUM(55) => 
                           S(55), SUM(54) => S(54), SUM(53) => S(53), SUM(52) 
                           => S(52), SUM(51) => S(51), SUM(50) => S(50), 
                           SUM(49) => S(49), SUM(48) => S(48), SUM(47) => S(47)
                           , SUM(46) => S(46), SUM(45) => S(45), SUM(44) => 
                           S(44), SUM(43) => S(43), SUM(42) => S(42), SUM(41) 
                           => S(41), SUM(40) => S(40), SUM(39) => S(39), 
                           SUM(38) => S(38), SUM(37) => S(37), SUM(36) => S(36)
                           , SUM(35) => S(35), SUM(34) => S(34), SUM(33) => 
                           S(33), SUM(32) => S(32), SUM(31) => S(31), SUM(30) 
                           => S(30), SUM(29) => S(29), SUM(28) => S(28), 
                           SUM(27) => S(27), SUM(26) => S(26), SUM(25) => S(25)
                           , SUM(24) => S(24), SUM(23) => S(23), SUM(22) => 
                           S(22), SUM(21) => S(21), SUM(20) => S(20), SUM(19) 
                           => S(19), SUM(18) => S(18), SUM(17) => S(17), 
                           SUM(16) => S(16), SUM(15) => S(15), SUM(14) => S(14)
                           , SUM(13) => S(13), SUM(12) => S(12), SUM(11) => 
                           S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) => 
                           S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5)
                           , SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1087);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity RCA_NBIT64_25 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_25;

architecture SYN_BEHAVIORAL of RCA_NBIT64_25 is

   component RCA_NBIT64_25_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1088 : std_logic;

begin
   
   n1 <= '0';
   add_1_root_add_81_2 : RCA_NBIT64_25_DW01_add_0 port map( A(64) => n1, A(63) 
                           => A(63), A(62) => A(62), A(61) => A(61), A(60) => 
                           A(60), A(59) => A(59), A(58) => A(58), A(57) => 
                           A(57), A(56) => A(56), A(55) => A(55), A(54) => 
                           A(54), A(53) => A(53), A(52) => A(52), A(51) => 
                           A(51), A(50) => A(50), A(49) => A(49), A(48) => 
                           A(48), A(47) => A(47), A(46) => A(46), A(45) => 
                           A(45), A(44) => A(44), A(43) => A(43), A(42) => 
                           A(42), A(41) => A(41), A(40) => A(40), A(39) => 
                           A(39), A(38) => A(38), A(37) => A(37), A(36) => 
                           A(36), A(35) => A(35), A(34) => A(34), A(33) => 
                           A(33), A(32) => A(32), A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(64) => n1, B(63) => B(63), 
                           B(62) => B(62), B(61) => B(61), B(60) => B(60), 
                           B(59) => B(59), B(58) => B(58), B(57) => B(57), 
                           B(56) => B(56), B(55) => B(55), B(54) => B(54), 
                           B(53) => B(53), B(52) => B(52), B(51) => B(51), 
                           B(50) => B(50), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, SUM(63)
                           => S(63), SUM(62) => S(62), SUM(61) => S(61), 
                           SUM(60) => S(60), SUM(59) => S(59), SUM(58) => S(58)
                           , SUM(57) => S(57), SUM(56) => S(56), SUM(55) => 
                           S(55), SUM(54) => S(54), SUM(53) => S(53), SUM(52) 
                           => S(52), SUM(51) => S(51), SUM(50) => S(50), 
                           SUM(49) => S(49), SUM(48) => S(48), SUM(47) => S(47)
                           , SUM(46) => S(46), SUM(45) => S(45), SUM(44) => 
                           S(44), SUM(43) => S(43), SUM(42) => S(42), SUM(41) 
                           => S(41), SUM(40) => S(40), SUM(39) => S(39), 
                           SUM(38) => S(38), SUM(37) => S(37), SUM(36) => S(36)
                           , SUM(35) => S(35), SUM(34) => S(34), SUM(33) => 
                           S(33), SUM(32) => S(32), SUM(31) => S(31), SUM(30) 
                           => S(30), SUM(29) => S(29), SUM(28) => S(28), 
                           SUM(27) => S(27), SUM(26) => S(26), SUM(25) => S(25)
                           , SUM(24) => S(24), SUM(23) => S(23), SUM(22) => 
                           S(22), SUM(21) => S(21), SUM(20) => S(20), SUM(19) 
                           => S(19), SUM(18) => S(18), SUM(17) => S(17), 
                           SUM(16) => S(16), SUM(15) => S(15), SUM(14) => S(14)
                           , SUM(13) => S(13), SUM(12) => S(12), SUM(11) => 
                           S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) => 
                           S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5)
                           , SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1088);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity RCA_NBIT64_26 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_26;

architecture SYN_BEHAVIORAL of RCA_NBIT64_26 is

   component RCA_NBIT64_26_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1089 : std_logic;

begin
   
   n1 <= '0';
   add_1_root_add_81_2 : RCA_NBIT64_26_DW01_add_0 port map( A(64) => n1, A(63) 
                           => A(63), A(62) => A(62), A(61) => A(61), A(60) => 
                           A(60), A(59) => A(59), A(58) => A(58), A(57) => 
                           A(57), A(56) => A(56), A(55) => A(55), A(54) => 
                           A(54), A(53) => A(53), A(52) => A(52), A(51) => 
                           A(51), A(50) => A(50), A(49) => A(49), A(48) => 
                           A(48), A(47) => A(47), A(46) => A(46), A(45) => 
                           A(45), A(44) => A(44), A(43) => A(43), A(42) => 
                           A(42), A(41) => A(41), A(40) => A(40), A(39) => 
                           A(39), A(38) => A(38), A(37) => A(37), A(36) => 
                           A(36), A(35) => A(35), A(34) => A(34), A(33) => 
                           A(33), A(32) => A(32), A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(64) => n1, B(63) => B(63), 
                           B(62) => B(62), B(61) => B(61), B(60) => B(60), 
                           B(59) => B(59), B(58) => B(58), B(57) => B(57), 
                           B(56) => B(56), B(55) => B(55), B(54) => B(54), 
                           B(53) => B(53), B(52) => B(52), B(51) => B(51), 
                           B(50) => B(50), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, SUM(63)
                           => S(63), SUM(62) => S(62), SUM(61) => S(61), 
                           SUM(60) => S(60), SUM(59) => S(59), SUM(58) => S(58)
                           , SUM(57) => S(57), SUM(56) => S(56), SUM(55) => 
                           S(55), SUM(54) => S(54), SUM(53) => S(53), SUM(52) 
                           => S(52), SUM(51) => S(51), SUM(50) => S(50), 
                           SUM(49) => S(49), SUM(48) => S(48), SUM(47) => S(47)
                           , SUM(46) => S(46), SUM(45) => S(45), SUM(44) => 
                           S(44), SUM(43) => S(43), SUM(42) => S(42), SUM(41) 
                           => S(41), SUM(40) => S(40), SUM(39) => S(39), 
                           SUM(38) => S(38), SUM(37) => S(37), SUM(36) => S(36)
                           , SUM(35) => S(35), SUM(34) => S(34), SUM(33) => 
                           S(33), SUM(32) => S(32), SUM(31) => S(31), SUM(30) 
                           => S(30), SUM(29) => S(29), SUM(28) => S(28), 
                           SUM(27) => S(27), SUM(26) => S(26), SUM(25) => S(25)
                           , SUM(24) => S(24), SUM(23) => S(23), SUM(22) => 
                           S(22), SUM(21) => S(21), SUM(20) => S(20), SUM(19) 
                           => S(19), SUM(18) => S(18), SUM(17) => S(17), 
                           SUM(16) => S(16), SUM(15) => S(15), SUM(14) => S(14)
                           , SUM(13) => S(13), SUM(12) => S(12), SUM(11) => 
                           S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) => 
                           S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5)
                           , SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1089);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity RCA_NBIT64_27 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_27;

architecture SYN_BEHAVIORAL of RCA_NBIT64_27 is

   component RCA_NBIT64_27_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1090 : std_logic;

begin
   
   n1 <= '0';
   add_1_root_add_81_2 : RCA_NBIT64_27_DW01_add_0 port map( A(64) => n1, A(63) 
                           => A(63), A(62) => A(62), A(61) => A(61), A(60) => 
                           A(60), A(59) => A(59), A(58) => A(58), A(57) => 
                           A(57), A(56) => A(56), A(55) => A(55), A(54) => 
                           A(54), A(53) => A(53), A(52) => A(52), A(51) => 
                           A(51), A(50) => A(50), A(49) => A(49), A(48) => 
                           A(48), A(47) => A(47), A(46) => A(46), A(45) => 
                           A(45), A(44) => A(44), A(43) => A(43), A(42) => 
                           A(42), A(41) => A(41), A(40) => A(40), A(39) => 
                           A(39), A(38) => A(38), A(37) => A(37), A(36) => 
                           A(36), A(35) => A(35), A(34) => A(34), A(33) => 
                           A(33), A(32) => A(32), A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(64) => n1, B(63) => B(63), 
                           B(62) => B(62), B(61) => B(61), B(60) => B(60), 
                           B(59) => B(59), B(58) => B(58), B(57) => B(57), 
                           B(56) => B(56), B(55) => B(55), B(54) => B(54), 
                           B(53) => B(53), B(52) => B(52), B(51) => B(51), 
                           B(50) => B(50), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, SUM(63)
                           => S(63), SUM(62) => S(62), SUM(61) => S(61), 
                           SUM(60) => S(60), SUM(59) => S(59), SUM(58) => S(58)
                           , SUM(57) => S(57), SUM(56) => S(56), SUM(55) => 
                           S(55), SUM(54) => S(54), SUM(53) => S(53), SUM(52) 
                           => S(52), SUM(51) => S(51), SUM(50) => S(50), 
                           SUM(49) => S(49), SUM(48) => S(48), SUM(47) => S(47)
                           , SUM(46) => S(46), SUM(45) => S(45), SUM(44) => 
                           S(44), SUM(43) => S(43), SUM(42) => S(42), SUM(41) 
                           => S(41), SUM(40) => S(40), SUM(39) => S(39), 
                           SUM(38) => S(38), SUM(37) => S(37), SUM(36) => S(36)
                           , SUM(35) => S(35), SUM(34) => S(34), SUM(33) => 
                           S(33), SUM(32) => S(32), SUM(31) => S(31), SUM(30) 
                           => S(30), SUM(29) => S(29), SUM(28) => S(28), 
                           SUM(27) => S(27), SUM(26) => S(26), SUM(25) => S(25)
                           , SUM(24) => S(24), SUM(23) => S(23), SUM(22) => 
                           S(22), SUM(21) => S(21), SUM(20) => S(20), SUM(19) 
                           => S(19), SUM(18) => S(18), SUM(17) => S(17), 
                           SUM(16) => S(16), SUM(15) => S(15), SUM(14) => S(14)
                           , SUM(13) => S(13), SUM(12) => S(12), SUM(11) => 
                           S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) => 
                           S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5)
                           , SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1090);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity RCA_NBIT64_28 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_28;

architecture SYN_BEHAVIORAL of RCA_NBIT64_28 is

   component RCA_NBIT64_28_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1091 : std_logic;

begin
   
   n1 <= '0';
   add_1_root_add_81_2 : RCA_NBIT64_28_DW01_add_0 port map( A(64) => n1, A(63) 
                           => A(63), A(62) => A(62), A(61) => A(61), A(60) => 
                           A(60), A(59) => A(59), A(58) => A(58), A(57) => 
                           A(57), A(56) => A(56), A(55) => A(55), A(54) => 
                           A(54), A(53) => A(53), A(52) => A(52), A(51) => 
                           A(51), A(50) => A(50), A(49) => A(49), A(48) => 
                           A(48), A(47) => A(47), A(46) => A(46), A(45) => 
                           A(45), A(44) => A(44), A(43) => A(43), A(42) => 
                           A(42), A(41) => A(41), A(40) => A(40), A(39) => 
                           A(39), A(38) => A(38), A(37) => A(37), A(36) => 
                           A(36), A(35) => A(35), A(34) => A(34), A(33) => 
                           A(33), A(32) => A(32), A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(64) => n1, B(63) => B(63), 
                           B(62) => B(62), B(61) => B(61), B(60) => B(60), 
                           B(59) => B(59), B(58) => B(58), B(57) => B(57), 
                           B(56) => B(56), B(55) => B(55), B(54) => B(54), 
                           B(53) => B(53), B(52) => B(52), B(51) => B(51), 
                           B(50) => B(50), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, SUM(63)
                           => S(63), SUM(62) => S(62), SUM(61) => S(61), 
                           SUM(60) => S(60), SUM(59) => S(59), SUM(58) => S(58)
                           , SUM(57) => S(57), SUM(56) => S(56), SUM(55) => 
                           S(55), SUM(54) => S(54), SUM(53) => S(53), SUM(52) 
                           => S(52), SUM(51) => S(51), SUM(50) => S(50), 
                           SUM(49) => S(49), SUM(48) => S(48), SUM(47) => S(47)
                           , SUM(46) => S(46), SUM(45) => S(45), SUM(44) => 
                           S(44), SUM(43) => S(43), SUM(42) => S(42), SUM(41) 
                           => S(41), SUM(40) => S(40), SUM(39) => S(39), 
                           SUM(38) => S(38), SUM(37) => S(37), SUM(36) => S(36)
                           , SUM(35) => S(35), SUM(34) => S(34), SUM(33) => 
                           S(33), SUM(32) => S(32), SUM(31) => S(31), SUM(30) 
                           => S(30), SUM(29) => S(29), SUM(28) => S(28), 
                           SUM(27) => S(27), SUM(26) => S(26), SUM(25) => S(25)
                           , SUM(24) => S(24), SUM(23) => S(23), SUM(22) => 
                           S(22), SUM(21) => S(21), SUM(20) => S(20), SUM(19) 
                           => S(19), SUM(18) => S(18), SUM(17) => S(17), 
                           SUM(16) => S(16), SUM(15) => S(15), SUM(14) => S(14)
                           , SUM(13) => S(13), SUM(12) => S(12), SUM(11) => 
                           S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) => 
                           S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5)
                           , SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1091);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity RCA_NBIT64_29 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_29;

architecture SYN_BEHAVIORAL of RCA_NBIT64_29 is

   component RCA_NBIT64_29_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n_1092 : std_logic;

begin
   
   n1 <= '0';
   add_1_root_add_81_2 : RCA_NBIT64_29_DW01_add_0 port map( A(64) => n1, A(63) 
                           => A(63), A(62) => A(62), A(61) => A(61), A(60) => 
                           A(60), A(59) => A(59), A(58) => A(58), A(57) => 
                           A(57), A(56) => A(56), A(55) => A(55), A(54) => 
                           A(54), A(53) => A(53), A(52) => A(52), A(51) => 
                           A(51), A(50) => A(50), A(49) => A(49), A(48) => 
                           A(48), A(47) => A(47), A(46) => A(46), A(45) => 
                           A(45), A(44) => A(44), A(43) => A(43), A(42) => 
                           A(42), A(41) => A(41), A(40) => A(40), A(39) => 
                           A(39), A(38) => A(38), A(37) => A(37), A(36) => 
                           A(36), A(35) => A(35), A(34) => A(34), A(33) => 
                           A(33), A(32) => A(32), A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(64) => n1, B(63) => B(63), 
                           B(62) => B(62), B(61) => B(61), B(60) => B(60), 
                           B(59) => B(59), B(58) => B(58), B(57) => B(57), 
                           B(56) => B(56), B(55) => B(55), B(54) => B(54), 
                           B(53) => B(53), B(52) => B(52), B(51) => B(51), 
                           B(50) => B(50), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, SUM(63)
                           => S(63), SUM(62) => S(62), SUM(61) => S(61), 
                           SUM(60) => S(60), SUM(59) => S(59), SUM(58) => S(58)
                           , SUM(57) => S(57), SUM(56) => S(56), SUM(55) => 
                           S(55), SUM(54) => S(54), SUM(53) => S(53), SUM(52) 
                           => S(52), SUM(51) => S(51), SUM(50) => S(50), 
                           SUM(49) => S(49), SUM(48) => S(48), SUM(47) => S(47)
                           , SUM(46) => S(46), SUM(45) => S(45), SUM(44) => 
                           S(44), SUM(43) => S(43), SUM(42) => S(42), SUM(41) 
                           => S(41), SUM(40) => S(40), SUM(39) => S(39), 
                           SUM(38) => S(38), SUM(37) => S(37), SUM(36) => S(36)
                           , SUM(35) => S(35), SUM(34) => S(34), SUM(33) => 
                           S(33), SUM(32) => S(32), SUM(31) => S(31), SUM(30) 
                           => S(30), SUM(29) => S(29), SUM(28) => S(28), 
                           SUM(27) => S(27), SUM(26) => S(26), SUM(25) => S(25)
                           , SUM(24) => S(24), SUM(23) => S(23), SUM(22) => 
                           S(22), SUM(21) => S(21), SUM(20) => S(20), SUM(19) 
                           => S(19), SUM(18) => S(18), SUM(17) => S(17), 
                           SUM(16) => S(16), SUM(15) => S(15), SUM(14) => S(14)
                           , SUM(13) => S(13), SUM(12) => S(12), SUM(11) => 
                           S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) => 
                           S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5)
                           , SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1092);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity RCA_NBIT64_15 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_NBIT64_15;

architecture SYN_BEHAVIORAL of RCA_NBIT64_15 is

   component RCA_NBIT64_15_DW01_add_0
      port( A, B : in std_logic_vector (64 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (64 downto 0);  CO : out std_logic);
   end component;
   
   signal n2, n_1093 : std_logic;

begin
   
   n2 <= '0';
   add_1_root_add_81_2 : RCA_NBIT64_15_DW01_add_0 port map( A(64) => n2, A(63) 
                           => A(63), A(62) => A(62), A(61) => A(61), A(60) => 
                           A(60), A(59) => A(59), A(58) => A(58), A(57) => 
                           A(57), A(56) => A(56), A(55) => A(55), A(54) => 
                           A(54), A(53) => A(53), A(52) => A(52), A(51) => 
                           A(51), A(50) => A(50), A(49) => A(49), A(48) => 
                           A(48), A(47) => A(47), A(46) => A(46), A(45) => 
                           A(45), A(44) => A(44), A(43) => A(43), A(42) => 
                           A(42), A(41) => A(41), A(40) => A(40), A(39) => 
                           A(39), A(38) => A(38), A(37) => A(37), A(36) => 
                           A(36), A(35) => A(35), A(34) => A(34), A(33) => 
                           A(33), A(32) => A(32), A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(64) => n2, B(63) => B(63), 
                           B(62) => B(62), B(61) => B(61), B(60) => B(60), 
                           B(59) => B(59), B(58) => B(58), B(57) => B(57), 
                           B(56) => B(56), B(55) => B(55), B(54) => B(54), 
                           B(53) => B(53), B(52) => B(52), B(51) => B(51), 
                           B(50) => B(50), B(49) => B(49), B(48) => B(48), 
                           B(47) => B(47), B(46) => B(46), B(45) => B(45), 
                           B(44) => B(44), B(43) => B(43), B(42) => B(42), 
                           B(41) => B(41), B(40) => B(40), B(39) => B(39), 
                           B(38) => B(38), B(37) => B(37), B(36) => B(36), 
                           B(35) => B(35), B(34) => B(34), B(33) => B(33), 
                           B(32) => B(32), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), CI => Ci, SUM(64) => Co, SUM(63)
                           => S(63), SUM(62) => S(62), SUM(61) => S(61), 
                           SUM(60) => S(60), SUM(59) => S(59), SUM(58) => S(58)
                           , SUM(57) => S(57), SUM(56) => S(56), SUM(55) => 
                           S(55), SUM(54) => S(54), SUM(53) => S(53), SUM(52) 
                           => S(52), SUM(51) => S(51), SUM(50) => S(50), 
                           SUM(49) => S(49), SUM(48) => S(48), SUM(47) => S(47)
                           , SUM(46) => S(46), SUM(45) => S(45), SUM(44) => 
                           S(44), SUM(43) => S(43), SUM(42) => S(42), SUM(41) 
                           => S(41), SUM(40) => S(40), SUM(39) => S(39), 
                           SUM(38) => S(38), SUM(37) => S(37), SUM(36) => S(36)
                           , SUM(35) => S(35), SUM(34) => S(34), SUM(33) => 
                           S(33), SUM(32) => S(32), SUM(31) => S(31), SUM(30) 
                           => S(30), SUM(29) => S(29), SUM(28) => S(28), 
                           SUM(27) => S(27), SUM(26) => S(26), SUM(25) => S(25)
                           , SUM(24) => S(24), SUM(23) => S(23), SUM(22) => 
                           S(22), SUM(21) => S(21), SUM(20) => S(20), SUM(19) 
                           => S(19), SUM(18) => S(18), SUM(17) => S(17), 
                           SUM(16) => S(16), SUM(15) => S(15), SUM(14) => S(14)
                           , SUM(13) => S(13), SUM(12) => S(12), SUM(11) => 
                           S(11), SUM(10) => S(10), SUM(9) => S(9), SUM(8) => 
                           S(8), SUM(7) => S(7), SUM(6) => S(6), SUM(5) => S(5)
                           , SUM(4) => S(4), SUM(3) => S(3), SUM(2) => S(2), 
                           SUM(1) => S(1), SUM(0) => S(0), CO => n_1093);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity BOOTHENC_NBIT64_i30 is

   port( A, A_n, A_ns, A_s, B : in std_logic_vector (63 downto 0);  O, A_so, 
         A_nso : out std_logic_vector (63 downto 0));

end BOOTHENC_NBIT64_i30;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT64_i30 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, O_63_port, O_62_port, O_61_port, O_60_port, O_59_port,
      O_58_port, O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, 
      O_52_port, O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, 
      O_46_port, O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, 
      O_40_port, O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, 
      O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, 
      O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, 
      O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, 
      O_16_port, O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, 
      O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, 
      O_3_port, O_2_port, O_1_port, n391, n392, n393, n394, n395, n396, n397, 
      n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, 
      n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, 
      n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, 
      n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, 
      n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, 
      n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, 
      n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, 
      n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, 
      n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, 
      n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, 
      n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, 
      n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, 
      n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, 
      n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, 
      n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, 
      n578, n579, n580, n581, n582, n583, n584, n585 : std_logic;

begin
   O <= ( O_63_port, O_62_port, O_61_port, O_60_port, O_59_port, O_58_port, 
      O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, O_52_port, 
      O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, O_46_port, 
      O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, O_40_port, 
      O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, 
      O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, 
      O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, 
      O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, O_16_port, 
      O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, O_10_port, 
      O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, O_3_port, 
      O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(61), A_s(60), A_s(59), A_s(58), A_s(57), A_s(56), A_s(55), 
      A_s(54), A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), 
      A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), 
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   A_nso <= ( A_s(61), A_s(60), A_s(59), A_s(58), A_s(57), A_s(56), A_s(55), 
      A_s(54), A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), 
      A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), 
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : AND3_X1 port map( A1 => B(30), A2 => n585, A3 => B(29), ZN => n391);
   U3 : INV_X4 port map( A => n391, ZN => n392);
   U4 : INV_X4 port map( A => n552, ZN => n398);
   U5 : OR3_X4 port map( A1 => B(29), A2 => B(30), A3 => n585, ZN => n393);
   U6 : INV_X4 port map( A => n553, ZN => n397);
   U7 : OAI221_X1 port map( B1 => n393, B2 => n394, C1 => n392, C2 => n395, A 
                           => n396, ZN => O_9_port);
   U8 : AOI22_X1 port map( A1 => A_ns(8), A2 => n397, B1 => A_s(8), B2 => n398,
                           ZN => n396);
   U9 : INV_X1 port map( A => A_s(7), ZN => n395);
   U10 : INV_X1 port map( A => A_ns(7), ZN => n394);
   U11 : OAI221_X1 port map( B1 => n393, B2 => n399, C1 => n392, C2 => n400, A 
                           => n401, ZN => O_8_port);
   U12 : AOI22_X1 port map( A1 => A_ns(7), A2 => n397, B1 => A_s(7), B2 => n398
                           , ZN => n401);
   U13 : INV_X1 port map( A => A_s(6), ZN => n400);
   U14 : INV_X1 port map( A => A_ns(6), ZN => n399);
   U15 : OAI221_X1 port map( B1 => n393, B2 => n402, C1 => n392, C2 => n403, A 
                           => n404, ZN => O_7_port);
   U16 : AOI22_X1 port map( A1 => A_ns(6), A2 => n397, B1 => A_s(6), B2 => n398
                           , ZN => n404);
   U17 : INV_X1 port map( A => A_s(5), ZN => n403);
   U18 : INV_X1 port map( A => A_ns(5), ZN => n402);
   U19 : OAI221_X1 port map( B1 => n393, B2 => n405, C1 => n392, C2 => n406, A 
                           => n407, ZN => O_6_port);
   U20 : AOI22_X1 port map( A1 => A_ns(5), A2 => n397, B1 => A_s(5), B2 => n398
                           , ZN => n407);
   U21 : INV_X1 port map( A => A_s(4), ZN => n406);
   U22 : INV_X1 port map( A => A_ns(4), ZN => n405);
   U23 : OAI221_X1 port map( B1 => n393, B2 => n408, C1 => n392, C2 => n409, A 
                           => n410, ZN => O_63_port);
   U24 : AOI22_X1 port map( A1 => A_ns(62), A2 => n397, B1 => A_s(62), B2 => 
                           n398, ZN => n410);
   U25 : INV_X1 port map( A => A_s(61), ZN => n409);
   U26 : INV_X1 port map( A => A_ns(61), ZN => n408);
   U27 : OAI221_X1 port map( B1 => n393, B2 => n411, C1 => n392, C2 => n412, A 
                           => n413, ZN => O_62_port);
   U28 : AOI22_X1 port map( A1 => A_ns(61), A2 => n397, B1 => A_s(61), B2 => 
                           n398, ZN => n413);
   U29 : INV_X1 port map( A => A_s(60), ZN => n412);
   U30 : INV_X1 port map( A => A_ns(60), ZN => n411);
   U31 : OAI221_X1 port map( B1 => n393, B2 => n414, C1 => n392, C2 => n415, A 
                           => n416, ZN => O_61_port);
   U32 : AOI22_X1 port map( A1 => A_ns(60), A2 => n397, B1 => A_s(60), B2 => 
                           n398, ZN => n416);
   U33 : INV_X1 port map( A => A_s(59), ZN => n415);
   U34 : INV_X1 port map( A => A_ns(59), ZN => n414);
   U35 : OAI221_X1 port map( B1 => n393, B2 => n417, C1 => n392, C2 => n418, A 
                           => n419, ZN => O_60_port);
   U36 : AOI22_X1 port map( A1 => A_ns(59), A2 => n397, B1 => A_s(59), B2 => 
                           n398, ZN => n419);
   U37 : INV_X1 port map( A => A_s(58), ZN => n418);
   U38 : INV_X1 port map( A => A_ns(58), ZN => n417);
   U39 : OAI221_X1 port map( B1 => n393, B2 => n420, C1 => n392, C2 => n421, A 
                           => n422, ZN => O_5_port);
   U40 : AOI22_X1 port map( A1 => A_ns(4), A2 => n397, B1 => A_s(4), B2 => n398
                           , ZN => n422);
   U41 : INV_X1 port map( A => A_s(3), ZN => n421);
   U42 : INV_X1 port map( A => A_ns(3), ZN => n420);
   U43 : OAI221_X1 port map( B1 => n393, B2 => n423, C1 => n392, C2 => n424, A 
                           => n425, ZN => O_59_port);
   U44 : AOI22_X1 port map( A1 => A_ns(58), A2 => n397, B1 => A_s(58), B2 => 
                           n398, ZN => n425);
   U45 : INV_X1 port map( A => A_s(57), ZN => n424);
   U46 : INV_X1 port map( A => A_ns(57), ZN => n423);
   U47 : OAI221_X1 port map( B1 => n393, B2 => n426, C1 => n392, C2 => n427, A 
                           => n428, ZN => O_58_port);
   U48 : AOI22_X1 port map( A1 => A_ns(57), A2 => n397, B1 => A_s(57), B2 => 
                           n398, ZN => n428);
   U49 : INV_X1 port map( A => A_s(56), ZN => n427);
   U50 : INV_X1 port map( A => A_ns(56), ZN => n426);
   U51 : OAI221_X1 port map( B1 => n393, B2 => n429, C1 => n392, C2 => n430, A 
                           => n431, ZN => O_57_port);
   U52 : AOI22_X1 port map( A1 => A_ns(56), A2 => n397, B1 => A_s(56), B2 => 
                           n398, ZN => n431);
   U53 : INV_X1 port map( A => A_s(55), ZN => n430);
   U54 : INV_X1 port map( A => A_ns(55), ZN => n429);
   U55 : OAI221_X1 port map( B1 => n393, B2 => n432, C1 => n392, C2 => n433, A 
                           => n434, ZN => O_56_port);
   U56 : AOI22_X1 port map( A1 => A_ns(55), A2 => n397, B1 => A_s(55), B2 => 
                           n398, ZN => n434);
   U57 : INV_X1 port map( A => A_s(54), ZN => n433);
   U58 : INV_X1 port map( A => A_ns(54), ZN => n432);
   U59 : OAI221_X1 port map( B1 => n393, B2 => n435, C1 => n392, C2 => n436, A 
                           => n437, ZN => O_55_port);
   U60 : AOI22_X1 port map( A1 => A_ns(54), A2 => n397, B1 => A_s(54), B2 => 
                           n398, ZN => n437);
   U61 : INV_X1 port map( A => A_s(53), ZN => n436);
   U62 : INV_X1 port map( A => A_ns(53), ZN => n435);
   U63 : OAI221_X1 port map( B1 => n393, B2 => n438, C1 => n392, C2 => n439, A 
                           => n440, ZN => O_54_port);
   U64 : AOI22_X1 port map( A1 => A_ns(53), A2 => n397, B1 => A_s(53), B2 => 
                           n398, ZN => n440);
   U65 : INV_X1 port map( A => A_s(52), ZN => n439);
   U66 : INV_X1 port map( A => A_ns(52), ZN => n438);
   U67 : OAI221_X1 port map( B1 => n393, B2 => n441, C1 => n392, C2 => n442, A 
                           => n443, ZN => O_53_port);
   U68 : AOI22_X1 port map( A1 => A_ns(52), A2 => n397, B1 => A_s(52), B2 => 
                           n398, ZN => n443);
   U69 : INV_X1 port map( A => A_s(51), ZN => n442);
   U70 : INV_X1 port map( A => A_ns(51), ZN => n441);
   U71 : OAI221_X1 port map( B1 => n393, B2 => n444, C1 => n392, C2 => n445, A 
                           => n446, ZN => O_52_port);
   U72 : AOI22_X1 port map( A1 => A_ns(51), A2 => n397, B1 => A_s(51), B2 => 
                           n398, ZN => n446);
   U73 : INV_X1 port map( A => A_s(50), ZN => n445);
   U74 : INV_X1 port map( A => A_ns(50), ZN => n444);
   U75 : OAI221_X1 port map( B1 => n393, B2 => n447, C1 => n392, C2 => n448, A 
                           => n449, ZN => O_51_port);
   U76 : AOI22_X1 port map( A1 => A_ns(50), A2 => n397, B1 => A_s(50), B2 => 
                           n398, ZN => n449);
   U77 : INV_X1 port map( A => A_s(49), ZN => n448);
   U78 : INV_X1 port map( A => A_ns(49), ZN => n447);
   U79 : OAI221_X1 port map( B1 => n393, B2 => n450, C1 => n392, C2 => n451, A 
                           => n452, ZN => O_50_port);
   U80 : AOI22_X1 port map( A1 => A_ns(49), A2 => n397, B1 => A_s(49), B2 => 
                           n398, ZN => n452);
   U81 : INV_X1 port map( A => A_s(48), ZN => n451);
   U82 : INV_X1 port map( A => A_ns(48), ZN => n450);
   U83 : OAI221_X1 port map( B1 => n393, B2 => n453, C1 => n392, C2 => n454, A 
                           => n455, ZN => O_4_port);
   U84 : AOI22_X1 port map( A1 => A_ns(3), A2 => n397, B1 => A_s(3), B2 => n398
                           , ZN => n455);
   U85 : INV_X1 port map( A => A_s(2), ZN => n454);
   U86 : INV_X1 port map( A => A_ns(2), ZN => n453);
   U87 : OAI221_X1 port map( B1 => n393, B2 => n456, C1 => n392, C2 => n457, A 
                           => n458, ZN => O_49_port);
   U88 : AOI22_X1 port map( A1 => A_ns(48), A2 => n397, B1 => A_s(48), B2 => 
                           n398, ZN => n458);
   U89 : INV_X1 port map( A => A_s(47), ZN => n457);
   U90 : INV_X1 port map( A => A_ns(47), ZN => n456);
   U91 : OAI221_X1 port map( B1 => n393, B2 => n459, C1 => n392, C2 => n460, A 
                           => n461, ZN => O_48_port);
   U92 : AOI22_X1 port map( A1 => A_ns(47), A2 => n397, B1 => A_s(47), B2 => 
                           n398, ZN => n461);
   U93 : INV_X1 port map( A => A_s(46), ZN => n460);
   U94 : INV_X1 port map( A => A_ns(46), ZN => n459);
   U95 : OAI221_X1 port map( B1 => n393, B2 => n462, C1 => n392, C2 => n463, A 
                           => n464, ZN => O_47_port);
   U96 : AOI22_X1 port map( A1 => A_ns(46), A2 => n397, B1 => A_s(46), B2 => 
                           n398, ZN => n464);
   U97 : INV_X1 port map( A => A_s(45), ZN => n463);
   U98 : INV_X1 port map( A => A_ns(45), ZN => n462);
   U99 : OAI221_X1 port map( B1 => n393, B2 => n465, C1 => n392, C2 => n466, A 
                           => n467, ZN => O_46_port);
   U100 : AOI22_X1 port map( A1 => A_ns(45), A2 => n397, B1 => A_s(45), B2 => 
                           n398, ZN => n467);
   U101 : INV_X1 port map( A => A_s(44), ZN => n466);
   U102 : INV_X1 port map( A => A_ns(44), ZN => n465);
   U103 : OAI221_X1 port map( B1 => n393, B2 => n468, C1 => n392, C2 => n469, A
                           => n470, ZN => O_45_port);
   U104 : AOI22_X1 port map( A1 => A_ns(44), A2 => n397, B1 => A_s(44), B2 => 
                           n398, ZN => n470);
   U105 : INV_X1 port map( A => A_s(43), ZN => n469);
   U106 : INV_X1 port map( A => A_ns(43), ZN => n468);
   U107 : OAI221_X1 port map( B1 => n393, B2 => n471, C1 => n392, C2 => n472, A
                           => n473, ZN => O_44_port);
   U108 : AOI22_X1 port map( A1 => A_ns(43), A2 => n397, B1 => A_s(43), B2 => 
                           n398, ZN => n473);
   U109 : INV_X1 port map( A => A_s(42), ZN => n472);
   U110 : INV_X1 port map( A => A_ns(42), ZN => n471);
   U111 : OAI221_X1 port map( B1 => n393, B2 => n474, C1 => n392, C2 => n475, A
                           => n476, ZN => O_43_port);
   U112 : AOI22_X1 port map( A1 => A_ns(42), A2 => n397, B1 => A_s(42), B2 => 
                           n398, ZN => n476);
   U113 : INV_X1 port map( A => A_s(41), ZN => n475);
   U114 : INV_X1 port map( A => A_ns(41), ZN => n474);
   U115 : OAI221_X1 port map( B1 => n393, B2 => n477, C1 => n392, C2 => n478, A
                           => n479, ZN => O_42_port);
   U116 : AOI22_X1 port map( A1 => A_ns(41), A2 => n397, B1 => A_s(41), B2 => 
                           n398, ZN => n479);
   U117 : INV_X1 port map( A => A_s(40), ZN => n478);
   U118 : INV_X1 port map( A => A_ns(40), ZN => n477);
   U119 : OAI221_X1 port map( B1 => n393, B2 => n480, C1 => n392, C2 => n481, A
                           => n482, ZN => O_41_port);
   U120 : AOI22_X1 port map( A1 => A_ns(40), A2 => n397, B1 => A_s(40), B2 => 
                           n398, ZN => n482);
   U121 : INV_X1 port map( A => A_s(39), ZN => n481);
   U122 : INV_X1 port map( A => A_ns(39), ZN => n480);
   U123 : OAI221_X1 port map( B1 => n393, B2 => n483, C1 => n392, C2 => n484, A
                           => n485, ZN => O_40_port);
   U124 : AOI22_X1 port map( A1 => A_ns(39), A2 => n397, B1 => A_s(39), B2 => 
                           n398, ZN => n485);
   U125 : INV_X1 port map( A => A_s(38), ZN => n484);
   U126 : INV_X1 port map( A => A_ns(38), ZN => n483);
   U127 : OAI221_X1 port map( B1 => n393, B2 => n486, C1 => n392, C2 => n487, A
                           => n488, ZN => O_3_port);
   U128 : AOI22_X1 port map( A1 => A_ns(2), A2 => n397, B1 => A_s(2), B2 => 
                           n398, ZN => n488);
   U129 : INV_X1 port map( A => A_s(1), ZN => n487);
   U130 : INV_X1 port map( A => A_ns(1), ZN => n486);
   U131 : OAI221_X1 port map( B1 => n393, B2 => n489, C1 => n392, C2 => n490, A
                           => n491, ZN => O_39_port);
   U132 : AOI22_X1 port map( A1 => A_ns(38), A2 => n397, B1 => A_s(38), B2 => 
                           n398, ZN => n491);
   U133 : INV_X1 port map( A => A_s(37), ZN => n490);
   U134 : INV_X1 port map( A => A_ns(37), ZN => n489);
   U135 : OAI221_X1 port map( B1 => n393, B2 => n492, C1 => n392, C2 => n493, A
                           => n494, ZN => O_38_port);
   U136 : AOI22_X1 port map( A1 => A_ns(37), A2 => n397, B1 => A_s(37), B2 => 
                           n398, ZN => n494);
   U137 : INV_X1 port map( A => A_s(36), ZN => n493);
   U138 : INV_X1 port map( A => A_ns(36), ZN => n492);
   U139 : OAI221_X1 port map( B1 => n393, B2 => n495, C1 => n392, C2 => n496, A
                           => n497, ZN => O_37_port);
   U140 : AOI22_X1 port map( A1 => A_ns(36), A2 => n397, B1 => A_s(36), B2 => 
                           n398, ZN => n497);
   U141 : INV_X1 port map( A => A_s(35), ZN => n496);
   U142 : INV_X1 port map( A => A_ns(35), ZN => n495);
   U143 : OAI221_X1 port map( B1 => n393, B2 => n498, C1 => n392, C2 => n499, A
                           => n500, ZN => O_36_port);
   U144 : AOI22_X1 port map( A1 => A_ns(35), A2 => n397, B1 => A_s(35), B2 => 
                           n398, ZN => n500);
   U145 : INV_X1 port map( A => A_s(34), ZN => n499);
   U146 : INV_X1 port map( A => A_ns(34), ZN => n498);
   U147 : OAI221_X1 port map( B1 => n393, B2 => n501, C1 => n392, C2 => n502, A
                           => n503, ZN => O_35_port);
   U148 : AOI22_X1 port map( A1 => A_ns(34), A2 => n397, B1 => A_s(34), B2 => 
                           n398, ZN => n503);
   U149 : INV_X1 port map( A => A_s(33), ZN => n502);
   U150 : INV_X1 port map( A => A_ns(33), ZN => n501);
   U151 : OAI221_X1 port map( B1 => n393, B2 => n504, C1 => n392, C2 => n505, A
                           => n506, ZN => O_34_port);
   U152 : AOI22_X1 port map( A1 => A_ns(33), A2 => n397, B1 => A_s(33), B2 => 
                           n398, ZN => n506);
   U153 : INV_X1 port map( A => A_s(32), ZN => n505);
   U154 : INV_X1 port map( A => A_ns(32), ZN => n504);
   U155 : OAI221_X1 port map( B1 => n393, B2 => n507, C1 => n392, C2 => n508, A
                           => n509, ZN => O_33_port);
   U156 : AOI22_X1 port map( A1 => A_ns(32), A2 => n397, B1 => A_s(32), B2 => 
                           n398, ZN => n509);
   U157 : INV_X1 port map( A => A_s(31), ZN => n508);
   U158 : INV_X1 port map( A => A_ns(31), ZN => n507);
   U159 : OAI221_X1 port map( B1 => n393, B2 => n510, C1 => n392, C2 => n511, A
                           => n512, ZN => O_32_port);
   U160 : AOI22_X1 port map( A1 => A_ns(31), A2 => n397, B1 => A_s(31), B2 => 
                           n398, ZN => n512);
   U161 : INV_X1 port map( A => A_s(30), ZN => n511);
   U162 : INV_X1 port map( A => A_ns(30), ZN => n510);
   U163 : OAI221_X1 port map( B1 => n393, B2 => n513, C1 => n392, C2 => n514, A
                           => n515, ZN => O_31_port);
   U164 : AOI22_X1 port map( A1 => A_ns(30), A2 => n397, B1 => A_s(30), B2 => 
                           n398, ZN => n515);
   U165 : INV_X1 port map( A => A_s(29), ZN => n514);
   U166 : INV_X1 port map( A => A_ns(29), ZN => n513);
   U167 : OAI221_X1 port map( B1 => n393, B2 => n516, C1 => n392, C2 => n517, A
                           => n518, ZN => O_30_port);
   U168 : AOI22_X1 port map( A1 => A_ns(29), A2 => n397, B1 => A_s(29), B2 => 
                           n398, ZN => n518);
   U169 : INV_X1 port map( A => A_s(28), ZN => n517);
   U170 : INV_X1 port map( A => A_ns(28), ZN => n516);
   U171 : OAI221_X1 port map( B1 => n393, B2 => n519, C1 => n392, C2 => n520, A
                           => n521, ZN => O_2_port);
   U172 : AOI22_X1 port map( A1 => A_ns(1), A2 => n397, B1 => A_s(1), B2 => 
                           n398, ZN => n521);
   U173 : OAI221_X1 port map( B1 => n393, B2 => n522, C1 => n392, C2 => n523, A
                           => n524, ZN => O_29_port);
   U174 : AOI22_X1 port map( A1 => A_ns(28), A2 => n397, B1 => A_s(28), B2 => 
                           n398, ZN => n524);
   U175 : INV_X1 port map( A => A_s(27), ZN => n523);
   U176 : INV_X1 port map( A => A_ns(27), ZN => n522);
   U177 : OAI221_X1 port map( B1 => n393, B2 => n525, C1 => n392, C2 => n526, A
                           => n527, ZN => O_28_port);
   U178 : AOI22_X1 port map( A1 => A_ns(27), A2 => n397, B1 => A_s(27), B2 => 
                           n398, ZN => n527);
   U179 : INV_X1 port map( A => A_s(26), ZN => n526);
   U180 : INV_X1 port map( A => A_ns(26), ZN => n525);
   U181 : OAI221_X1 port map( B1 => n393, B2 => n528, C1 => n392, C2 => n529, A
                           => n530, ZN => O_27_port);
   U182 : AOI22_X1 port map( A1 => A_ns(26), A2 => n397, B1 => A_s(26), B2 => 
                           n398, ZN => n530);
   U183 : INV_X1 port map( A => A_s(25), ZN => n529);
   U184 : INV_X1 port map( A => A_ns(25), ZN => n528);
   U185 : OAI221_X1 port map( B1 => n393, B2 => n531, C1 => n392, C2 => n532, A
                           => n533, ZN => O_26_port);
   U186 : AOI22_X1 port map( A1 => A_ns(25), A2 => n397, B1 => A_s(25), B2 => 
                           n398, ZN => n533);
   U187 : INV_X1 port map( A => A_s(24), ZN => n532);
   U188 : INV_X1 port map( A => A_ns(24), ZN => n531);
   U189 : OAI221_X1 port map( B1 => n393, B2 => n534, C1 => n392, C2 => n535, A
                           => n536, ZN => O_25_port);
   U190 : AOI22_X1 port map( A1 => A_ns(24), A2 => n397, B1 => A_s(24), B2 => 
                           n398, ZN => n536);
   U191 : INV_X1 port map( A => A_s(23), ZN => n535);
   U192 : INV_X1 port map( A => A_ns(23), ZN => n534);
   U193 : OAI221_X1 port map( B1 => n393, B2 => n537, C1 => n392, C2 => n538, A
                           => n539, ZN => O_24_port);
   U194 : AOI22_X1 port map( A1 => A_ns(23), A2 => n397, B1 => A_s(23), B2 => 
                           n398, ZN => n539);
   U195 : INV_X1 port map( A => A_s(22), ZN => n538);
   U196 : INV_X1 port map( A => A_ns(22), ZN => n537);
   U197 : OAI221_X1 port map( B1 => n393, B2 => n540, C1 => n392, C2 => n541, A
                           => n542, ZN => O_23_port);
   U198 : AOI22_X1 port map( A1 => A_ns(22), A2 => n397, B1 => A_s(22), B2 => 
                           n398, ZN => n542);
   U199 : INV_X1 port map( A => A_s(21), ZN => n541);
   U200 : INV_X1 port map( A => A_ns(21), ZN => n540);
   U201 : OAI221_X1 port map( B1 => n393, B2 => n543, C1 => n392, C2 => n544, A
                           => n545, ZN => O_22_port);
   U202 : AOI22_X1 port map( A1 => A_ns(21), A2 => n397, B1 => A_s(21), B2 => 
                           n398, ZN => n545);
   U203 : INV_X1 port map( A => A_s(20), ZN => n544);
   U204 : INV_X1 port map( A => A_ns(20), ZN => n543);
   U205 : OAI221_X1 port map( B1 => n393, B2 => n546, C1 => n392, C2 => n547, A
                           => n548, ZN => O_21_port);
   U206 : AOI22_X1 port map( A1 => A_ns(20), A2 => n397, B1 => A_s(20), B2 => 
                           n398, ZN => n548);
   U207 : INV_X1 port map( A => A_s(19), ZN => n547);
   U208 : INV_X1 port map( A => A_ns(19), ZN => n546);
   U209 : OAI221_X1 port map( B1 => n393, B2 => n549, C1 => n392, C2 => n550, A
                           => n551, ZN => O_20_port);
   U210 : AOI22_X1 port map( A1 => A_ns(19), A2 => n397, B1 => A_s(19), B2 => 
                           n398, ZN => n551);
   U211 : INV_X1 port map( A => A_s(18), ZN => n550);
   U212 : INV_X1 port map( A => A_ns(18), ZN => n549);
   U213 : OAI22_X1 port map( A1 => n552, A2 => n520, B1 => n553, B2 => n519, ZN
                           => O_1_port);
   U214 : INV_X1 port map( A => A_ns(0), ZN => n519);
   U215 : INV_X1 port map( A => A_s(0), ZN => n520);
   U216 : OAI221_X1 port map( B1 => n393, B2 => n554, C1 => n392, C2 => n555, A
                           => n556, ZN => O_19_port);
   U217 : AOI22_X1 port map( A1 => A_ns(18), A2 => n397, B1 => A_s(18), B2 => 
                           n398, ZN => n556);
   U218 : INV_X1 port map( A => A_s(17), ZN => n555);
   U219 : INV_X1 port map( A => A_ns(17), ZN => n554);
   U220 : OAI221_X1 port map( B1 => n393, B2 => n557, C1 => n392, C2 => n558, A
                           => n559, ZN => O_18_port);
   U221 : AOI22_X1 port map( A1 => A_ns(17), A2 => n397, B1 => A_s(17), B2 => 
                           n398, ZN => n559);
   U222 : INV_X1 port map( A => A_s(16), ZN => n558);
   U223 : INV_X1 port map( A => A_ns(16), ZN => n557);
   U224 : OAI221_X1 port map( B1 => n393, B2 => n560, C1 => n392, C2 => n561, A
                           => n562, ZN => O_17_port);
   U225 : AOI22_X1 port map( A1 => A_ns(16), A2 => n397, B1 => A_s(16), B2 => 
                           n398, ZN => n562);
   U226 : INV_X1 port map( A => A_s(15), ZN => n561);
   U227 : INV_X1 port map( A => A_ns(15), ZN => n560);
   U228 : OAI221_X1 port map( B1 => n393, B2 => n563, C1 => n392, C2 => n564, A
                           => n565, ZN => O_16_port);
   U229 : AOI22_X1 port map( A1 => A_ns(15), A2 => n397, B1 => A_s(15), B2 => 
                           n398, ZN => n565);
   U230 : INV_X1 port map( A => A_s(14), ZN => n564);
   U231 : INV_X1 port map( A => A_ns(14), ZN => n563);
   U232 : OAI221_X1 port map( B1 => n393, B2 => n566, C1 => n392, C2 => n567, A
                           => n568, ZN => O_15_port);
   U233 : AOI22_X1 port map( A1 => A_ns(14), A2 => n397, B1 => A_s(14), B2 => 
                           n398, ZN => n568);
   U234 : INV_X1 port map( A => A_s(13), ZN => n567);
   U235 : INV_X1 port map( A => A_ns(13), ZN => n566);
   U236 : OAI221_X1 port map( B1 => n393, B2 => n569, C1 => n392, C2 => n570, A
                           => n571, ZN => O_14_port);
   U237 : AOI22_X1 port map( A1 => A_ns(13), A2 => n397, B1 => A_s(13), B2 => 
                           n398, ZN => n571);
   U238 : INV_X1 port map( A => A_s(12), ZN => n570);
   U239 : INV_X1 port map( A => A_ns(12), ZN => n569);
   U240 : OAI221_X1 port map( B1 => n393, B2 => n572, C1 => n392, C2 => n573, A
                           => n574, ZN => O_13_port);
   U241 : AOI22_X1 port map( A1 => A_ns(12), A2 => n397, B1 => A_s(12), B2 => 
                           n398, ZN => n574);
   U242 : INV_X1 port map( A => A_s(11), ZN => n573);
   U243 : INV_X1 port map( A => A_ns(11), ZN => n572);
   U244 : OAI221_X1 port map( B1 => n393, B2 => n575, C1 => n392, C2 => n576, A
                           => n577, ZN => O_12_port);
   U245 : AOI22_X1 port map( A1 => A_ns(11), A2 => n397, B1 => A_s(11), B2 => 
                           n398, ZN => n577);
   U246 : INV_X1 port map( A => A_s(10), ZN => n576);
   U247 : INV_X1 port map( A => A_ns(10), ZN => n575);
   U248 : OAI221_X1 port map( B1 => n393, B2 => n578, C1 => n392, C2 => n579, A
                           => n580, ZN => O_11_port);
   U249 : AOI22_X1 port map( A1 => A_ns(10), A2 => n397, B1 => A_s(10), B2 => 
                           n398, ZN => n580);
   U250 : INV_X1 port map( A => A_s(9), ZN => n579);
   U251 : INV_X1 port map( A => A_ns(9), ZN => n578);
   U252 : OAI221_X1 port map( B1 => n581, B2 => n393, C1 => n582, C2 => n392, A
                           => n583, ZN => O_10_port);
   U253 : AOI22_X1 port map( A1 => A_ns(9), A2 => n397, B1 => A_s(9), B2 => 
                           n398, ZN => n583);
   U254 : NAND2_X1 port map( A1 => n584, A2 => n552, ZN => n553);
   U255 : NAND2_X1 port map( A1 => n584, A2 => n585, ZN => n552);
   U256 : XOR2_X1 port map( A => B(29), B => B(30), Z => n584);
   U257 : INV_X1 port map( A => A_s(8), ZN => n582);
   U258 : INV_X1 port map( A => B(31), ZN => n585);
   U259 : INV_X1 port map( A => A_ns(8), ZN => n581);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity BOOTHENC_NBIT64_i28 is

   port( A, A_n, A_ns, A_s, B : in std_logic_vector (63 downto 0);  O, A_so, 
         A_nso : out std_logic_vector (63 downto 0));

end BOOTHENC_NBIT64_i28;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT64_i28 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, O_63_port, O_62_port, O_61_port, O_60_port, O_59_port,
      O_58_port, O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, 
      O_52_port, O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, 
      O_46_port, O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, 
      O_40_port, O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, 
      O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, 
      O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, 
      O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, 
      O_16_port, O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, 
      O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, 
      O_3_port, O_2_port, O_1_port, n391, n392, n393, n394, n395, n396, n397, 
      n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, 
      n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, 
      n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, 
      n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, 
      n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, 
      n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, 
      n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, 
      n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, 
      n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, 
      n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, 
      n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, 
      n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, 
      n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, 
      n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, 
      n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, 
      n578, n579, n580, n581, n582, n583, n584, n585 : std_logic;

begin
   O <= ( O_63_port, O_62_port, O_61_port, O_60_port, O_59_port, O_58_port, 
      O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, O_52_port, 
      O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, O_46_port, 
      O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, O_40_port, 
      O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, 
      O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, 
      O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, 
      O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, O_16_port, 
      O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, O_10_port, 
      O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, O_3_port, 
      O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(61), A_s(60), A_s(59), A_s(58), A_s(57), A_s(56), A_s(55), 
      A_s(54), A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), 
      A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), 
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   A_nso <= ( A_s(61), A_s(60), A_s(59), A_s(58), A_s(57), A_s(56), A_s(55), 
      A_s(54), A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), 
      A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), 
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : AND3_X1 port map( A1 => B(28), A2 => n585, A3 => B(27), ZN => n391);
   U3 : INV_X4 port map( A => n391, ZN => n392);
   U4 : INV_X4 port map( A => n552, ZN => n398);
   U5 : OR3_X4 port map( A1 => B(27), A2 => B(28), A3 => n585, ZN => n393);
   U6 : INV_X4 port map( A => n553, ZN => n397);
   U7 : OAI221_X1 port map( B1 => n393, B2 => n394, C1 => n392, C2 => n395, A 
                           => n396, ZN => O_9_port);
   U8 : AOI22_X1 port map( A1 => A_ns(8), A2 => n397, B1 => A_s(8), B2 => n398,
                           ZN => n396);
   U9 : INV_X1 port map( A => A_s(7), ZN => n395);
   U10 : INV_X1 port map( A => A_ns(7), ZN => n394);
   U11 : OAI221_X1 port map( B1 => n393, B2 => n399, C1 => n392, C2 => n400, A 
                           => n401, ZN => O_8_port);
   U12 : AOI22_X1 port map( A1 => A_ns(7), A2 => n397, B1 => A_s(7), B2 => n398
                           , ZN => n401);
   U13 : INV_X1 port map( A => A_s(6), ZN => n400);
   U14 : INV_X1 port map( A => A_ns(6), ZN => n399);
   U15 : OAI221_X1 port map( B1 => n393, B2 => n402, C1 => n392, C2 => n403, A 
                           => n404, ZN => O_7_port);
   U16 : AOI22_X1 port map( A1 => A_ns(6), A2 => n397, B1 => A_s(6), B2 => n398
                           , ZN => n404);
   U17 : INV_X1 port map( A => A_s(5), ZN => n403);
   U18 : INV_X1 port map( A => A_ns(5), ZN => n402);
   U19 : OAI221_X1 port map( B1 => n393, B2 => n405, C1 => n392, C2 => n406, A 
                           => n407, ZN => O_6_port);
   U20 : AOI22_X1 port map( A1 => A_ns(5), A2 => n397, B1 => A_s(5), B2 => n398
                           , ZN => n407);
   U21 : INV_X1 port map( A => A_s(4), ZN => n406);
   U22 : INV_X1 port map( A => A_ns(4), ZN => n405);
   U23 : OAI221_X1 port map( B1 => n393, B2 => n408, C1 => n392, C2 => n409, A 
                           => n410, ZN => O_63_port);
   U24 : AOI22_X1 port map( A1 => A_ns(62), A2 => n397, B1 => A_s(62), B2 => 
                           n398, ZN => n410);
   U25 : INV_X1 port map( A => A_s(61), ZN => n409);
   U26 : INV_X1 port map( A => A_ns(61), ZN => n408);
   U27 : OAI221_X1 port map( B1 => n393, B2 => n411, C1 => n392, C2 => n412, A 
                           => n413, ZN => O_62_port);
   U28 : AOI22_X1 port map( A1 => A_ns(61), A2 => n397, B1 => A_s(61), B2 => 
                           n398, ZN => n413);
   U29 : INV_X1 port map( A => A_s(60), ZN => n412);
   U30 : INV_X1 port map( A => A_ns(60), ZN => n411);
   U31 : OAI221_X1 port map( B1 => n393, B2 => n414, C1 => n392, C2 => n415, A 
                           => n416, ZN => O_61_port);
   U32 : AOI22_X1 port map( A1 => A_ns(60), A2 => n397, B1 => A_s(60), B2 => 
                           n398, ZN => n416);
   U33 : INV_X1 port map( A => A_s(59), ZN => n415);
   U34 : INV_X1 port map( A => A_ns(59), ZN => n414);
   U35 : OAI221_X1 port map( B1 => n393, B2 => n417, C1 => n392, C2 => n418, A 
                           => n419, ZN => O_60_port);
   U36 : AOI22_X1 port map( A1 => A_ns(59), A2 => n397, B1 => A_s(59), B2 => 
                           n398, ZN => n419);
   U37 : INV_X1 port map( A => A_s(58), ZN => n418);
   U38 : INV_X1 port map( A => A_ns(58), ZN => n417);
   U39 : OAI221_X1 port map( B1 => n393, B2 => n420, C1 => n392, C2 => n421, A 
                           => n422, ZN => O_5_port);
   U40 : AOI22_X1 port map( A1 => A_ns(4), A2 => n397, B1 => A_s(4), B2 => n398
                           , ZN => n422);
   U41 : INV_X1 port map( A => A_s(3), ZN => n421);
   U42 : INV_X1 port map( A => A_ns(3), ZN => n420);
   U43 : OAI221_X1 port map( B1 => n393, B2 => n423, C1 => n392, C2 => n424, A 
                           => n425, ZN => O_59_port);
   U44 : AOI22_X1 port map( A1 => A_ns(58), A2 => n397, B1 => A_s(58), B2 => 
                           n398, ZN => n425);
   U45 : INV_X1 port map( A => A_s(57), ZN => n424);
   U46 : INV_X1 port map( A => A_ns(57), ZN => n423);
   U47 : OAI221_X1 port map( B1 => n393, B2 => n426, C1 => n392, C2 => n427, A 
                           => n428, ZN => O_58_port);
   U48 : AOI22_X1 port map( A1 => A_ns(57), A2 => n397, B1 => A_s(57), B2 => 
                           n398, ZN => n428);
   U49 : INV_X1 port map( A => A_s(56), ZN => n427);
   U50 : INV_X1 port map( A => A_ns(56), ZN => n426);
   U51 : OAI221_X1 port map( B1 => n393, B2 => n429, C1 => n392, C2 => n430, A 
                           => n431, ZN => O_57_port);
   U52 : AOI22_X1 port map( A1 => A_ns(56), A2 => n397, B1 => A_s(56), B2 => 
                           n398, ZN => n431);
   U53 : INV_X1 port map( A => A_s(55), ZN => n430);
   U54 : INV_X1 port map( A => A_ns(55), ZN => n429);
   U55 : OAI221_X1 port map( B1 => n393, B2 => n432, C1 => n392, C2 => n433, A 
                           => n434, ZN => O_56_port);
   U56 : AOI22_X1 port map( A1 => A_ns(55), A2 => n397, B1 => A_s(55), B2 => 
                           n398, ZN => n434);
   U57 : INV_X1 port map( A => A_s(54), ZN => n433);
   U58 : INV_X1 port map( A => A_ns(54), ZN => n432);
   U59 : OAI221_X1 port map( B1 => n393, B2 => n435, C1 => n392, C2 => n436, A 
                           => n437, ZN => O_55_port);
   U60 : AOI22_X1 port map( A1 => A_ns(54), A2 => n397, B1 => A_s(54), B2 => 
                           n398, ZN => n437);
   U61 : INV_X1 port map( A => A_s(53), ZN => n436);
   U62 : INV_X1 port map( A => A_ns(53), ZN => n435);
   U63 : OAI221_X1 port map( B1 => n393, B2 => n438, C1 => n392, C2 => n439, A 
                           => n440, ZN => O_54_port);
   U64 : AOI22_X1 port map( A1 => A_ns(53), A2 => n397, B1 => A_s(53), B2 => 
                           n398, ZN => n440);
   U65 : INV_X1 port map( A => A_s(52), ZN => n439);
   U66 : INV_X1 port map( A => A_ns(52), ZN => n438);
   U67 : OAI221_X1 port map( B1 => n393, B2 => n441, C1 => n392, C2 => n442, A 
                           => n443, ZN => O_53_port);
   U68 : AOI22_X1 port map( A1 => A_ns(52), A2 => n397, B1 => A_s(52), B2 => 
                           n398, ZN => n443);
   U69 : INV_X1 port map( A => A_s(51), ZN => n442);
   U70 : INV_X1 port map( A => A_ns(51), ZN => n441);
   U71 : OAI221_X1 port map( B1 => n393, B2 => n444, C1 => n392, C2 => n445, A 
                           => n446, ZN => O_52_port);
   U72 : AOI22_X1 port map( A1 => A_ns(51), A2 => n397, B1 => A_s(51), B2 => 
                           n398, ZN => n446);
   U73 : INV_X1 port map( A => A_s(50), ZN => n445);
   U74 : INV_X1 port map( A => A_ns(50), ZN => n444);
   U75 : OAI221_X1 port map( B1 => n393, B2 => n447, C1 => n392, C2 => n448, A 
                           => n449, ZN => O_51_port);
   U76 : AOI22_X1 port map( A1 => A_ns(50), A2 => n397, B1 => A_s(50), B2 => 
                           n398, ZN => n449);
   U77 : INV_X1 port map( A => A_s(49), ZN => n448);
   U78 : INV_X1 port map( A => A_ns(49), ZN => n447);
   U79 : OAI221_X1 port map( B1 => n393, B2 => n450, C1 => n392, C2 => n451, A 
                           => n452, ZN => O_50_port);
   U80 : AOI22_X1 port map( A1 => A_ns(49), A2 => n397, B1 => A_s(49), B2 => 
                           n398, ZN => n452);
   U81 : INV_X1 port map( A => A_s(48), ZN => n451);
   U82 : INV_X1 port map( A => A_ns(48), ZN => n450);
   U83 : OAI221_X1 port map( B1 => n393, B2 => n453, C1 => n392, C2 => n454, A 
                           => n455, ZN => O_4_port);
   U84 : AOI22_X1 port map( A1 => A_ns(3), A2 => n397, B1 => A_s(3), B2 => n398
                           , ZN => n455);
   U85 : INV_X1 port map( A => A_s(2), ZN => n454);
   U86 : INV_X1 port map( A => A_ns(2), ZN => n453);
   U87 : OAI221_X1 port map( B1 => n393, B2 => n456, C1 => n392, C2 => n457, A 
                           => n458, ZN => O_49_port);
   U88 : AOI22_X1 port map( A1 => A_ns(48), A2 => n397, B1 => A_s(48), B2 => 
                           n398, ZN => n458);
   U89 : INV_X1 port map( A => A_s(47), ZN => n457);
   U90 : INV_X1 port map( A => A_ns(47), ZN => n456);
   U91 : OAI221_X1 port map( B1 => n393, B2 => n459, C1 => n392, C2 => n460, A 
                           => n461, ZN => O_48_port);
   U92 : AOI22_X1 port map( A1 => A_ns(47), A2 => n397, B1 => A_s(47), B2 => 
                           n398, ZN => n461);
   U93 : INV_X1 port map( A => A_s(46), ZN => n460);
   U94 : INV_X1 port map( A => A_ns(46), ZN => n459);
   U95 : OAI221_X1 port map( B1 => n393, B2 => n462, C1 => n392, C2 => n463, A 
                           => n464, ZN => O_47_port);
   U96 : AOI22_X1 port map( A1 => A_ns(46), A2 => n397, B1 => A_s(46), B2 => 
                           n398, ZN => n464);
   U97 : INV_X1 port map( A => A_s(45), ZN => n463);
   U98 : INV_X1 port map( A => A_ns(45), ZN => n462);
   U99 : OAI221_X1 port map( B1 => n393, B2 => n465, C1 => n392, C2 => n466, A 
                           => n467, ZN => O_46_port);
   U100 : AOI22_X1 port map( A1 => A_ns(45), A2 => n397, B1 => A_s(45), B2 => 
                           n398, ZN => n467);
   U101 : INV_X1 port map( A => A_s(44), ZN => n466);
   U102 : INV_X1 port map( A => A_ns(44), ZN => n465);
   U103 : OAI221_X1 port map( B1 => n393, B2 => n468, C1 => n392, C2 => n469, A
                           => n470, ZN => O_45_port);
   U104 : AOI22_X1 port map( A1 => A_ns(44), A2 => n397, B1 => A_s(44), B2 => 
                           n398, ZN => n470);
   U105 : INV_X1 port map( A => A_s(43), ZN => n469);
   U106 : INV_X1 port map( A => A_ns(43), ZN => n468);
   U107 : OAI221_X1 port map( B1 => n393, B2 => n471, C1 => n392, C2 => n472, A
                           => n473, ZN => O_44_port);
   U108 : AOI22_X1 port map( A1 => A_ns(43), A2 => n397, B1 => A_s(43), B2 => 
                           n398, ZN => n473);
   U109 : INV_X1 port map( A => A_s(42), ZN => n472);
   U110 : INV_X1 port map( A => A_ns(42), ZN => n471);
   U111 : OAI221_X1 port map( B1 => n393, B2 => n474, C1 => n392, C2 => n475, A
                           => n476, ZN => O_43_port);
   U112 : AOI22_X1 port map( A1 => A_ns(42), A2 => n397, B1 => A_s(42), B2 => 
                           n398, ZN => n476);
   U113 : INV_X1 port map( A => A_s(41), ZN => n475);
   U114 : INV_X1 port map( A => A_ns(41), ZN => n474);
   U115 : OAI221_X1 port map( B1 => n393, B2 => n477, C1 => n392, C2 => n478, A
                           => n479, ZN => O_42_port);
   U116 : AOI22_X1 port map( A1 => A_ns(41), A2 => n397, B1 => A_s(41), B2 => 
                           n398, ZN => n479);
   U117 : INV_X1 port map( A => A_s(40), ZN => n478);
   U118 : INV_X1 port map( A => A_ns(40), ZN => n477);
   U119 : OAI221_X1 port map( B1 => n393, B2 => n480, C1 => n392, C2 => n481, A
                           => n482, ZN => O_41_port);
   U120 : AOI22_X1 port map( A1 => A_ns(40), A2 => n397, B1 => A_s(40), B2 => 
                           n398, ZN => n482);
   U121 : INV_X1 port map( A => A_s(39), ZN => n481);
   U122 : INV_X1 port map( A => A_ns(39), ZN => n480);
   U123 : OAI221_X1 port map( B1 => n393, B2 => n483, C1 => n392, C2 => n484, A
                           => n485, ZN => O_40_port);
   U124 : AOI22_X1 port map( A1 => A_ns(39), A2 => n397, B1 => A_s(39), B2 => 
                           n398, ZN => n485);
   U125 : INV_X1 port map( A => A_s(38), ZN => n484);
   U126 : INV_X1 port map( A => A_ns(38), ZN => n483);
   U127 : OAI221_X1 port map( B1 => n393, B2 => n486, C1 => n392, C2 => n487, A
                           => n488, ZN => O_3_port);
   U128 : AOI22_X1 port map( A1 => A_ns(2), A2 => n397, B1 => A_s(2), B2 => 
                           n398, ZN => n488);
   U129 : INV_X1 port map( A => A_s(1), ZN => n487);
   U130 : INV_X1 port map( A => A_ns(1), ZN => n486);
   U131 : OAI221_X1 port map( B1 => n393, B2 => n489, C1 => n392, C2 => n490, A
                           => n491, ZN => O_39_port);
   U132 : AOI22_X1 port map( A1 => A_ns(38), A2 => n397, B1 => A_s(38), B2 => 
                           n398, ZN => n491);
   U133 : INV_X1 port map( A => A_s(37), ZN => n490);
   U134 : INV_X1 port map( A => A_ns(37), ZN => n489);
   U135 : OAI221_X1 port map( B1 => n393, B2 => n492, C1 => n392, C2 => n493, A
                           => n494, ZN => O_38_port);
   U136 : AOI22_X1 port map( A1 => A_ns(37), A2 => n397, B1 => A_s(37), B2 => 
                           n398, ZN => n494);
   U137 : INV_X1 port map( A => A_s(36), ZN => n493);
   U138 : INV_X1 port map( A => A_ns(36), ZN => n492);
   U139 : OAI221_X1 port map( B1 => n393, B2 => n495, C1 => n392, C2 => n496, A
                           => n497, ZN => O_37_port);
   U140 : AOI22_X1 port map( A1 => A_ns(36), A2 => n397, B1 => A_s(36), B2 => 
                           n398, ZN => n497);
   U141 : INV_X1 port map( A => A_s(35), ZN => n496);
   U142 : INV_X1 port map( A => A_ns(35), ZN => n495);
   U143 : OAI221_X1 port map( B1 => n393, B2 => n498, C1 => n392, C2 => n499, A
                           => n500, ZN => O_36_port);
   U144 : AOI22_X1 port map( A1 => A_ns(35), A2 => n397, B1 => A_s(35), B2 => 
                           n398, ZN => n500);
   U145 : INV_X1 port map( A => A_s(34), ZN => n499);
   U146 : INV_X1 port map( A => A_ns(34), ZN => n498);
   U147 : OAI221_X1 port map( B1 => n393, B2 => n501, C1 => n392, C2 => n502, A
                           => n503, ZN => O_35_port);
   U148 : AOI22_X1 port map( A1 => A_ns(34), A2 => n397, B1 => A_s(34), B2 => 
                           n398, ZN => n503);
   U149 : INV_X1 port map( A => A_s(33), ZN => n502);
   U150 : INV_X1 port map( A => A_ns(33), ZN => n501);
   U151 : OAI221_X1 port map( B1 => n393, B2 => n504, C1 => n392, C2 => n505, A
                           => n506, ZN => O_34_port);
   U152 : AOI22_X1 port map( A1 => A_ns(33), A2 => n397, B1 => A_s(33), B2 => 
                           n398, ZN => n506);
   U153 : INV_X1 port map( A => A_s(32), ZN => n505);
   U154 : INV_X1 port map( A => A_ns(32), ZN => n504);
   U155 : OAI221_X1 port map( B1 => n393, B2 => n507, C1 => n392, C2 => n508, A
                           => n509, ZN => O_33_port);
   U156 : AOI22_X1 port map( A1 => A_ns(32), A2 => n397, B1 => A_s(32), B2 => 
                           n398, ZN => n509);
   U157 : INV_X1 port map( A => A_s(31), ZN => n508);
   U158 : INV_X1 port map( A => A_ns(31), ZN => n507);
   U159 : OAI221_X1 port map( B1 => n393, B2 => n510, C1 => n392, C2 => n511, A
                           => n512, ZN => O_32_port);
   U160 : AOI22_X1 port map( A1 => A_ns(31), A2 => n397, B1 => A_s(31), B2 => 
                           n398, ZN => n512);
   U161 : INV_X1 port map( A => A_s(30), ZN => n511);
   U162 : INV_X1 port map( A => A_ns(30), ZN => n510);
   U163 : OAI221_X1 port map( B1 => n393, B2 => n513, C1 => n392, C2 => n514, A
                           => n515, ZN => O_31_port);
   U164 : AOI22_X1 port map( A1 => A_ns(30), A2 => n397, B1 => A_s(30), B2 => 
                           n398, ZN => n515);
   U165 : INV_X1 port map( A => A_s(29), ZN => n514);
   U166 : INV_X1 port map( A => A_ns(29), ZN => n513);
   U167 : OAI221_X1 port map( B1 => n393, B2 => n516, C1 => n392, C2 => n517, A
                           => n518, ZN => O_30_port);
   U168 : AOI22_X1 port map( A1 => A_ns(29), A2 => n397, B1 => A_s(29), B2 => 
                           n398, ZN => n518);
   U169 : INV_X1 port map( A => A_s(28), ZN => n517);
   U170 : INV_X1 port map( A => A_ns(28), ZN => n516);
   U171 : OAI221_X1 port map( B1 => n393, B2 => n519, C1 => n392, C2 => n520, A
                           => n521, ZN => O_2_port);
   U172 : AOI22_X1 port map( A1 => A_ns(1), A2 => n397, B1 => A_s(1), B2 => 
                           n398, ZN => n521);
   U173 : OAI221_X1 port map( B1 => n393, B2 => n522, C1 => n392, C2 => n523, A
                           => n524, ZN => O_29_port);
   U174 : AOI22_X1 port map( A1 => A_ns(28), A2 => n397, B1 => A_s(28), B2 => 
                           n398, ZN => n524);
   U175 : INV_X1 port map( A => A_s(27), ZN => n523);
   U176 : INV_X1 port map( A => A_ns(27), ZN => n522);
   U177 : OAI221_X1 port map( B1 => n393, B2 => n525, C1 => n392, C2 => n526, A
                           => n527, ZN => O_28_port);
   U178 : AOI22_X1 port map( A1 => A_ns(27), A2 => n397, B1 => A_s(27), B2 => 
                           n398, ZN => n527);
   U179 : INV_X1 port map( A => A_s(26), ZN => n526);
   U180 : INV_X1 port map( A => A_ns(26), ZN => n525);
   U181 : OAI221_X1 port map( B1 => n393, B2 => n528, C1 => n392, C2 => n529, A
                           => n530, ZN => O_27_port);
   U182 : AOI22_X1 port map( A1 => A_ns(26), A2 => n397, B1 => A_s(26), B2 => 
                           n398, ZN => n530);
   U183 : INV_X1 port map( A => A_s(25), ZN => n529);
   U184 : INV_X1 port map( A => A_ns(25), ZN => n528);
   U185 : OAI221_X1 port map( B1 => n393, B2 => n531, C1 => n392, C2 => n532, A
                           => n533, ZN => O_26_port);
   U186 : AOI22_X1 port map( A1 => A_ns(25), A2 => n397, B1 => A_s(25), B2 => 
                           n398, ZN => n533);
   U187 : INV_X1 port map( A => A_s(24), ZN => n532);
   U188 : INV_X1 port map( A => A_ns(24), ZN => n531);
   U189 : OAI221_X1 port map( B1 => n393, B2 => n534, C1 => n392, C2 => n535, A
                           => n536, ZN => O_25_port);
   U190 : AOI22_X1 port map( A1 => A_ns(24), A2 => n397, B1 => A_s(24), B2 => 
                           n398, ZN => n536);
   U191 : INV_X1 port map( A => A_s(23), ZN => n535);
   U192 : INV_X1 port map( A => A_ns(23), ZN => n534);
   U193 : OAI221_X1 port map( B1 => n393, B2 => n537, C1 => n392, C2 => n538, A
                           => n539, ZN => O_24_port);
   U194 : AOI22_X1 port map( A1 => A_ns(23), A2 => n397, B1 => A_s(23), B2 => 
                           n398, ZN => n539);
   U195 : INV_X1 port map( A => A_s(22), ZN => n538);
   U196 : INV_X1 port map( A => A_ns(22), ZN => n537);
   U197 : OAI221_X1 port map( B1 => n393, B2 => n540, C1 => n392, C2 => n541, A
                           => n542, ZN => O_23_port);
   U198 : AOI22_X1 port map( A1 => A_ns(22), A2 => n397, B1 => A_s(22), B2 => 
                           n398, ZN => n542);
   U199 : INV_X1 port map( A => A_s(21), ZN => n541);
   U200 : INV_X1 port map( A => A_ns(21), ZN => n540);
   U201 : OAI221_X1 port map( B1 => n393, B2 => n543, C1 => n392, C2 => n544, A
                           => n545, ZN => O_22_port);
   U202 : AOI22_X1 port map( A1 => A_ns(21), A2 => n397, B1 => A_s(21), B2 => 
                           n398, ZN => n545);
   U203 : INV_X1 port map( A => A_s(20), ZN => n544);
   U204 : INV_X1 port map( A => A_ns(20), ZN => n543);
   U205 : OAI221_X1 port map( B1 => n393, B2 => n546, C1 => n392, C2 => n547, A
                           => n548, ZN => O_21_port);
   U206 : AOI22_X1 port map( A1 => A_ns(20), A2 => n397, B1 => A_s(20), B2 => 
                           n398, ZN => n548);
   U207 : INV_X1 port map( A => A_s(19), ZN => n547);
   U208 : INV_X1 port map( A => A_ns(19), ZN => n546);
   U209 : OAI221_X1 port map( B1 => n393, B2 => n549, C1 => n392, C2 => n550, A
                           => n551, ZN => O_20_port);
   U210 : AOI22_X1 port map( A1 => A_ns(19), A2 => n397, B1 => A_s(19), B2 => 
                           n398, ZN => n551);
   U211 : INV_X1 port map( A => A_s(18), ZN => n550);
   U212 : INV_X1 port map( A => A_ns(18), ZN => n549);
   U213 : OAI22_X1 port map( A1 => n552, A2 => n520, B1 => n553, B2 => n519, ZN
                           => O_1_port);
   U214 : INV_X1 port map( A => A_ns(0), ZN => n519);
   U215 : INV_X1 port map( A => A_s(0), ZN => n520);
   U216 : OAI221_X1 port map( B1 => n393, B2 => n554, C1 => n392, C2 => n555, A
                           => n556, ZN => O_19_port);
   U217 : AOI22_X1 port map( A1 => A_ns(18), A2 => n397, B1 => A_s(18), B2 => 
                           n398, ZN => n556);
   U218 : INV_X1 port map( A => A_s(17), ZN => n555);
   U219 : INV_X1 port map( A => A_ns(17), ZN => n554);
   U220 : OAI221_X1 port map( B1 => n393, B2 => n557, C1 => n392, C2 => n558, A
                           => n559, ZN => O_18_port);
   U221 : AOI22_X1 port map( A1 => A_ns(17), A2 => n397, B1 => A_s(17), B2 => 
                           n398, ZN => n559);
   U222 : INV_X1 port map( A => A_s(16), ZN => n558);
   U223 : INV_X1 port map( A => A_ns(16), ZN => n557);
   U224 : OAI221_X1 port map( B1 => n393, B2 => n560, C1 => n392, C2 => n561, A
                           => n562, ZN => O_17_port);
   U225 : AOI22_X1 port map( A1 => A_ns(16), A2 => n397, B1 => A_s(16), B2 => 
                           n398, ZN => n562);
   U226 : INV_X1 port map( A => A_s(15), ZN => n561);
   U227 : INV_X1 port map( A => A_ns(15), ZN => n560);
   U228 : OAI221_X1 port map( B1 => n393, B2 => n563, C1 => n392, C2 => n564, A
                           => n565, ZN => O_16_port);
   U229 : AOI22_X1 port map( A1 => A_ns(15), A2 => n397, B1 => A_s(15), B2 => 
                           n398, ZN => n565);
   U230 : INV_X1 port map( A => A_s(14), ZN => n564);
   U231 : INV_X1 port map( A => A_ns(14), ZN => n563);
   U232 : OAI221_X1 port map( B1 => n393, B2 => n566, C1 => n392, C2 => n567, A
                           => n568, ZN => O_15_port);
   U233 : AOI22_X1 port map( A1 => A_ns(14), A2 => n397, B1 => A_s(14), B2 => 
                           n398, ZN => n568);
   U234 : INV_X1 port map( A => A_s(13), ZN => n567);
   U235 : INV_X1 port map( A => A_ns(13), ZN => n566);
   U236 : OAI221_X1 port map( B1 => n393, B2 => n569, C1 => n392, C2 => n570, A
                           => n571, ZN => O_14_port);
   U237 : AOI22_X1 port map( A1 => A_ns(13), A2 => n397, B1 => A_s(13), B2 => 
                           n398, ZN => n571);
   U238 : INV_X1 port map( A => A_s(12), ZN => n570);
   U239 : INV_X1 port map( A => A_ns(12), ZN => n569);
   U240 : OAI221_X1 port map( B1 => n393, B2 => n572, C1 => n392, C2 => n573, A
                           => n574, ZN => O_13_port);
   U241 : AOI22_X1 port map( A1 => A_ns(12), A2 => n397, B1 => A_s(12), B2 => 
                           n398, ZN => n574);
   U242 : INV_X1 port map( A => A_s(11), ZN => n573);
   U243 : INV_X1 port map( A => A_ns(11), ZN => n572);
   U244 : OAI221_X1 port map( B1 => n393, B2 => n575, C1 => n392, C2 => n576, A
                           => n577, ZN => O_12_port);
   U245 : AOI22_X1 port map( A1 => A_ns(11), A2 => n397, B1 => A_s(11), B2 => 
                           n398, ZN => n577);
   U246 : INV_X1 port map( A => A_s(10), ZN => n576);
   U247 : INV_X1 port map( A => A_ns(10), ZN => n575);
   U248 : OAI221_X1 port map( B1 => n393, B2 => n578, C1 => n392, C2 => n579, A
                           => n580, ZN => O_11_port);
   U249 : AOI22_X1 port map( A1 => A_ns(10), A2 => n397, B1 => A_s(10), B2 => 
                           n398, ZN => n580);
   U250 : INV_X1 port map( A => A_s(9), ZN => n579);
   U251 : INV_X1 port map( A => A_ns(9), ZN => n578);
   U252 : OAI221_X1 port map( B1 => n581, B2 => n393, C1 => n582, C2 => n392, A
                           => n583, ZN => O_10_port);
   U253 : AOI22_X1 port map( A1 => A_ns(9), A2 => n397, B1 => A_s(9), B2 => 
                           n398, ZN => n583);
   U254 : NAND2_X1 port map( A1 => n584, A2 => n552, ZN => n553);
   U255 : NAND2_X1 port map( A1 => n584, A2 => n585, ZN => n552);
   U256 : XOR2_X1 port map( A => B(27), B => B(28), Z => n584);
   U257 : INV_X1 port map( A => A_s(8), ZN => n582);
   U258 : INV_X1 port map( A => B(29), ZN => n585);
   U259 : INV_X1 port map( A => A_ns(8), ZN => n581);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity BOOTHENC_NBIT64_i26 is

   port( A, A_n, A_ns, A_s, B : in std_logic_vector (63 downto 0);  O, A_so, 
         A_nso : out std_logic_vector (63 downto 0));

end BOOTHENC_NBIT64_i26;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT64_i26 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, O_63_port, O_62_port, O_61_port, O_60_port, O_59_port,
      O_58_port, O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, 
      O_52_port, O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, 
      O_46_port, O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, 
      O_40_port, O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, 
      O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, 
      O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, 
      O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, 
      O_16_port, O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, 
      O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, 
      O_3_port, O_2_port, O_1_port, n391, n392, n393, n394, n395, n396, n397, 
      n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, 
      n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, 
      n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, 
      n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, 
      n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, 
      n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, 
      n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, 
      n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, 
      n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, 
      n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, 
      n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, 
      n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, 
      n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, 
      n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, 
      n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, 
      n578, n579, n580, n581, n582, n583, n584, n585 : std_logic;

begin
   O <= ( O_63_port, O_62_port, O_61_port, O_60_port, O_59_port, O_58_port, 
      O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, O_52_port, 
      O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, O_46_port, 
      O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, O_40_port, 
      O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, 
      O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, 
      O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, 
      O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, O_16_port, 
      O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, O_10_port, 
      O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, O_3_port, 
      O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(61), A_s(60), A_s(59), A_s(58), A_s(57), A_s(56), A_s(55), 
      A_s(54), A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), 
      A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), 
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   A_nso <= ( A_s(61), A_s(60), A_s(59), A_s(58), A_s(57), A_s(56), A_s(55), 
      A_s(54), A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), 
      A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), 
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : AND3_X1 port map( A1 => B(26), A2 => n585, A3 => B(25), ZN => n391);
   U3 : INV_X4 port map( A => n391, ZN => n392);
   U4 : INV_X4 port map( A => n552, ZN => n398);
   U5 : OR3_X4 port map( A1 => B(25), A2 => B(26), A3 => n585, ZN => n393);
   U6 : INV_X4 port map( A => n553, ZN => n397);
   U7 : OAI221_X1 port map( B1 => n393, B2 => n394, C1 => n392, C2 => n395, A 
                           => n396, ZN => O_9_port);
   U8 : AOI22_X1 port map( A1 => A_ns(8), A2 => n397, B1 => A_s(8), B2 => n398,
                           ZN => n396);
   U9 : INV_X1 port map( A => A_s(7), ZN => n395);
   U10 : INV_X1 port map( A => A_ns(7), ZN => n394);
   U11 : OAI221_X1 port map( B1 => n393, B2 => n399, C1 => n392, C2 => n400, A 
                           => n401, ZN => O_8_port);
   U12 : AOI22_X1 port map( A1 => A_ns(7), A2 => n397, B1 => A_s(7), B2 => n398
                           , ZN => n401);
   U13 : INV_X1 port map( A => A_s(6), ZN => n400);
   U14 : INV_X1 port map( A => A_ns(6), ZN => n399);
   U15 : OAI221_X1 port map( B1 => n393, B2 => n402, C1 => n392, C2 => n403, A 
                           => n404, ZN => O_7_port);
   U16 : AOI22_X1 port map( A1 => A_ns(6), A2 => n397, B1 => A_s(6), B2 => n398
                           , ZN => n404);
   U17 : INV_X1 port map( A => A_s(5), ZN => n403);
   U18 : INV_X1 port map( A => A_ns(5), ZN => n402);
   U19 : OAI221_X1 port map( B1 => n393, B2 => n405, C1 => n392, C2 => n406, A 
                           => n407, ZN => O_6_port);
   U20 : AOI22_X1 port map( A1 => A_ns(5), A2 => n397, B1 => A_s(5), B2 => n398
                           , ZN => n407);
   U21 : INV_X1 port map( A => A_s(4), ZN => n406);
   U22 : INV_X1 port map( A => A_ns(4), ZN => n405);
   U23 : OAI221_X1 port map( B1 => n393, B2 => n408, C1 => n392, C2 => n409, A 
                           => n410, ZN => O_63_port);
   U24 : AOI22_X1 port map( A1 => A_ns(62), A2 => n397, B1 => A_s(62), B2 => 
                           n398, ZN => n410);
   U25 : INV_X1 port map( A => A_s(61), ZN => n409);
   U26 : INV_X1 port map( A => A_ns(61), ZN => n408);
   U27 : OAI221_X1 port map( B1 => n393, B2 => n411, C1 => n392, C2 => n412, A 
                           => n413, ZN => O_62_port);
   U28 : AOI22_X1 port map( A1 => A_ns(61), A2 => n397, B1 => A_s(61), B2 => 
                           n398, ZN => n413);
   U29 : INV_X1 port map( A => A_s(60), ZN => n412);
   U30 : INV_X1 port map( A => A_ns(60), ZN => n411);
   U31 : OAI221_X1 port map( B1 => n393, B2 => n414, C1 => n392, C2 => n415, A 
                           => n416, ZN => O_61_port);
   U32 : AOI22_X1 port map( A1 => A_ns(60), A2 => n397, B1 => A_s(60), B2 => 
                           n398, ZN => n416);
   U33 : INV_X1 port map( A => A_s(59), ZN => n415);
   U34 : INV_X1 port map( A => A_ns(59), ZN => n414);
   U35 : OAI221_X1 port map( B1 => n393, B2 => n417, C1 => n392, C2 => n418, A 
                           => n419, ZN => O_60_port);
   U36 : AOI22_X1 port map( A1 => A_ns(59), A2 => n397, B1 => A_s(59), B2 => 
                           n398, ZN => n419);
   U37 : INV_X1 port map( A => A_s(58), ZN => n418);
   U38 : INV_X1 port map( A => A_ns(58), ZN => n417);
   U39 : OAI221_X1 port map( B1 => n393, B2 => n420, C1 => n392, C2 => n421, A 
                           => n422, ZN => O_5_port);
   U40 : AOI22_X1 port map( A1 => A_ns(4), A2 => n397, B1 => A_s(4), B2 => n398
                           , ZN => n422);
   U41 : INV_X1 port map( A => A_s(3), ZN => n421);
   U42 : INV_X1 port map( A => A_ns(3), ZN => n420);
   U43 : OAI221_X1 port map( B1 => n393, B2 => n423, C1 => n392, C2 => n424, A 
                           => n425, ZN => O_59_port);
   U44 : AOI22_X1 port map( A1 => A_ns(58), A2 => n397, B1 => A_s(58), B2 => 
                           n398, ZN => n425);
   U45 : INV_X1 port map( A => A_s(57), ZN => n424);
   U46 : INV_X1 port map( A => A_ns(57), ZN => n423);
   U47 : OAI221_X1 port map( B1 => n393, B2 => n426, C1 => n392, C2 => n427, A 
                           => n428, ZN => O_58_port);
   U48 : AOI22_X1 port map( A1 => A_ns(57), A2 => n397, B1 => A_s(57), B2 => 
                           n398, ZN => n428);
   U49 : INV_X1 port map( A => A_s(56), ZN => n427);
   U50 : INV_X1 port map( A => A_ns(56), ZN => n426);
   U51 : OAI221_X1 port map( B1 => n393, B2 => n429, C1 => n392, C2 => n430, A 
                           => n431, ZN => O_57_port);
   U52 : AOI22_X1 port map( A1 => A_ns(56), A2 => n397, B1 => A_s(56), B2 => 
                           n398, ZN => n431);
   U53 : INV_X1 port map( A => A_s(55), ZN => n430);
   U54 : INV_X1 port map( A => A_ns(55), ZN => n429);
   U55 : OAI221_X1 port map( B1 => n393, B2 => n432, C1 => n392, C2 => n433, A 
                           => n434, ZN => O_56_port);
   U56 : AOI22_X1 port map( A1 => A_ns(55), A2 => n397, B1 => A_s(55), B2 => 
                           n398, ZN => n434);
   U57 : INV_X1 port map( A => A_s(54), ZN => n433);
   U58 : INV_X1 port map( A => A_ns(54), ZN => n432);
   U59 : OAI221_X1 port map( B1 => n393, B2 => n435, C1 => n392, C2 => n436, A 
                           => n437, ZN => O_55_port);
   U60 : AOI22_X1 port map( A1 => A_ns(54), A2 => n397, B1 => A_s(54), B2 => 
                           n398, ZN => n437);
   U61 : INV_X1 port map( A => A_s(53), ZN => n436);
   U62 : INV_X1 port map( A => A_ns(53), ZN => n435);
   U63 : OAI221_X1 port map( B1 => n393, B2 => n438, C1 => n392, C2 => n439, A 
                           => n440, ZN => O_54_port);
   U64 : AOI22_X1 port map( A1 => A_ns(53), A2 => n397, B1 => A_s(53), B2 => 
                           n398, ZN => n440);
   U65 : INV_X1 port map( A => A_s(52), ZN => n439);
   U66 : INV_X1 port map( A => A_ns(52), ZN => n438);
   U67 : OAI221_X1 port map( B1 => n393, B2 => n441, C1 => n392, C2 => n442, A 
                           => n443, ZN => O_53_port);
   U68 : AOI22_X1 port map( A1 => A_ns(52), A2 => n397, B1 => A_s(52), B2 => 
                           n398, ZN => n443);
   U69 : INV_X1 port map( A => A_s(51), ZN => n442);
   U70 : INV_X1 port map( A => A_ns(51), ZN => n441);
   U71 : OAI221_X1 port map( B1 => n393, B2 => n444, C1 => n392, C2 => n445, A 
                           => n446, ZN => O_52_port);
   U72 : AOI22_X1 port map( A1 => A_ns(51), A2 => n397, B1 => A_s(51), B2 => 
                           n398, ZN => n446);
   U73 : INV_X1 port map( A => A_s(50), ZN => n445);
   U74 : INV_X1 port map( A => A_ns(50), ZN => n444);
   U75 : OAI221_X1 port map( B1 => n393, B2 => n447, C1 => n392, C2 => n448, A 
                           => n449, ZN => O_51_port);
   U76 : AOI22_X1 port map( A1 => A_ns(50), A2 => n397, B1 => A_s(50), B2 => 
                           n398, ZN => n449);
   U77 : INV_X1 port map( A => A_s(49), ZN => n448);
   U78 : INV_X1 port map( A => A_ns(49), ZN => n447);
   U79 : OAI221_X1 port map( B1 => n393, B2 => n450, C1 => n392, C2 => n451, A 
                           => n452, ZN => O_50_port);
   U80 : AOI22_X1 port map( A1 => A_ns(49), A2 => n397, B1 => A_s(49), B2 => 
                           n398, ZN => n452);
   U81 : INV_X1 port map( A => A_s(48), ZN => n451);
   U82 : INV_X1 port map( A => A_ns(48), ZN => n450);
   U83 : OAI221_X1 port map( B1 => n393, B2 => n453, C1 => n392, C2 => n454, A 
                           => n455, ZN => O_4_port);
   U84 : AOI22_X1 port map( A1 => A_ns(3), A2 => n397, B1 => A_s(3), B2 => n398
                           , ZN => n455);
   U85 : INV_X1 port map( A => A_s(2), ZN => n454);
   U86 : INV_X1 port map( A => A_ns(2), ZN => n453);
   U87 : OAI221_X1 port map( B1 => n393, B2 => n456, C1 => n392, C2 => n457, A 
                           => n458, ZN => O_49_port);
   U88 : AOI22_X1 port map( A1 => A_ns(48), A2 => n397, B1 => A_s(48), B2 => 
                           n398, ZN => n458);
   U89 : INV_X1 port map( A => A_s(47), ZN => n457);
   U90 : INV_X1 port map( A => A_ns(47), ZN => n456);
   U91 : OAI221_X1 port map( B1 => n393, B2 => n459, C1 => n392, C2 => n460, A 
                           => n461, ZN => O_48_port);
   U92 : AOI22_X1 port map( A1 => A_ns(47), A2 => n397, B1 => A_s(47), B2 => 
                           n398, ZN => n461);
   U93 : INV_X1 port map( A => A_s(46), ZN => n460);
   U94 : INV_X1 port map( A => A_ns(46), ZN => n459);
   U95 : OAI221_X1 port map( B1 => n393, B2 => n462, C1 => n392, C2 => n463, A 
                           => n464, ZN => O_47_port);
   U96 : AOI22_X1 port map( A1 => A_ns(46), A2 => n397, B1 => A_s(46), B2 => 
                           n398, ZN => n464);
   U97 : INV_X1 port map( A => A_s(45), ZN => n463);
   U98 : INV_X1 port map( A => A_ns(45), ZN => n462);
   U99 : OAI221_X1 port map( B1 => n393, B2 => n465, C1 => n392, C2 => n466, A 
                           => n467, ZN => O_46_port);
   U100 : AOI22_X1 port map( A1 => A_ns(45), A2 => n397, B1 => A_s(45), B2 => 
                           n398, ZN => n467);
   U101 : INV_X1 port map( A => A_s(44), ZN => n466);
   U102 : INV_X1 port map( A => A_ns(44), ZN => n465);
   U103 : OAI221_X1 port map( B1 => n393, B2 => n468, C1 => n392, C2 => n469, A
                           => n470, ZN => O_45_port);
   U104 : AOI22_X1 port map( A1 => A_ns(44), A2 => n397, B1 => A_s(44), B2 => 
                           n398, ZN => n470);
   U105 : INV_X1 port map( A => A_s(43), ZN => n469);
   U106 : INV_X1 port map( A => A_ns(43), ZN => n468);
   U107 : OAI221_X1 port map( B1 => n393, B2 => n471, C1 => n392, C2 => n472, A
                           => n473, ZN => O_44_port);
   U108 : AOI22_X1 port map( A1 => A_ns(43), A2 => n397, B1 => A_s(43), B2 => 
                           n398, ZN => n473);
   U109 : INV_X1 port map( A => A_s(42), ZN => n472);
   U110 : INV_X1 port map( A => A_ns(42), ZN => n471);
   U111 : OAI221_X1 port map( B1 => n393, B2 => n474, C1 => n392, C2 => n475, A
                           => n476, ZN => O_43_port);
   U112 : AOI22_X1 port map( A1 => A_ns(42), A2 => n397, B1 => A_s(42), B2 => 
                           n398, ZN => n476);
   U113 : INV_X1 port map( A => A_s(41), ZN => n475);
   U114 : INV_X1 port map( A => A_ns(41), ZN => n474);
   U115 : OAI221_X1 port map( B1 => n393, B2 => n477, C1 => n392, C2 => n478, A
                           => n479, ZN => O_42_port);
   U116 : AOI22_X1 port map( A1 => A_ns(41), A2 => n397, B1 => A_s(41), B2 => 
                           n398, ZN => n479);
   U117 : INV_X1 port map( A => A_s(40), ZN => n478);
   U118 : INV_X1 port map( A => A_ns(40), ZN => n477);
   U119 : OAI221_X1 port map( B1 => n393, B2 => n480, C1 => n392, C2 => n481, A
                           => n482, ZN => O_41_port);
   U120 : AOI22_X1 port map( A1 => A_ns(40), A2 => n397, B1 => A_s(40), B2 => 
                           n398, ZN => n482);
   U121 : INV_X1 port map( A => A_s(39), ZN => n481);
   U122 : INV_X1 port map( A => A_ns(39), ZN => n480);
   U123 : OAI221_X1 port map( B1 => n393, B2 => n483, C1 => n392, C2 => n484, A
                           => n485, ZN => O_40_port);
   U124 : AOI22_X1 port map( A1 => A_ns(39), A2 => n397, B1 => A_s(39), B2 => 
                           n398, ZN => n485);
   U125 : INV_X1 port map( A => A_s(38), ZN => n484);
   U126 : INV_X1 port map( A => A_ns(38), ZN => n483);
   U127 : OAI221_X1 port map( B1 => n393, B2 => n486, C1 => n392, C2 => n487, A
                           => n488, ZN => O_3_port);
   U128 : AOI22_X1 port map( A1 => A_ns(2), A2 => n397, B1 => A_s(2), B2 => 
                           n398, ZN => n488);
   U129 : INV_X1 port map( A => A_s(1), ZN => n487);
   U130 : INV_X1 port map( A => A_ns(1), ZN => n486);
   U131 : OAI221_X1 port map( B1 => n393, B2 => n489, C1 => n392, C2 => n490, A
                           => n491, ZN => O_39_port);
   U132 : AOI22_X1 port map( A1 => A_ns(38), A2 => n397, B1 => A_s(38), B2 => 
                           n398, ZN => n491);
   U133 : INV_X1 port map( A => A_s(37), ZN => n490);
   U134 : INV_X1 port map( A => A_ns(37), ZN => n489);
   U135 : OAI221_X1 port map( B1 => n393, B2 => n492, C1 => n392, C2 => n493, A
                           => n494, ZN => O_38_port);
   U136 : AOI22_X1 port map( A1 => A_ns(37), A2 => n397, B1 => A_s(37), B2 => 
                           n398, ZN => n494);
   U137 : INV_X1 port map( A => A_s(36), ZN => n493);
   U138 : INV_X1 port map( A => A_ns(36), ZN => n492);
   U139 : OAI221_X1 port map( B1 => n393, B2 => n495, C1 => n392, C2 => n496, A
                           => n497, ZN => O_37_port);
   U140 : AOI22_X1 port map( A1 => A_ns(36), A2 => n397, B1 => A_s(36), B2 => 
                           n398, ZN => n497);
   U141 : INV_X1 port map( A => A_s(35), ZN => n496);
   U142 : INV_X1 port map( A => A_ns(35), ZN => n495);
   U143 : OAI221_X1 port map( B1 => n393, B2 => n498, C1 => n392, C2 => n499, A
                           => n500, ZN => O_36_port);
   U144 : AOI22_X1 port map( A1 => A_ns(35), A2 => n397, B1 => A_s(35), B2 => 
                           n398, ZN => n500);
   U145 : INV_X1 port map( A => A_s(34), ZN => n499);
   U146 : INV_X1 port map( A => A_ns(34), ZN => n498);
   U147 : OAI221_X1 port map( B1 => n393, B2 => n501, C1 => n392, C2 => n502, A
                           => n503, ZN => O_35_port);
   U148 : AOI22_X1 port map( A1 => A_ns(34), A2 => n397, B1 => A_s(34), B2 => 
                           n398, ZN => n503);
   U149 : INV_X1 port map( A => A_s(33), ZN => n502);
   U150 : INV_X1 port map( A => A_ns(33), ZN => n501);
   U151 : OAI221_X1 port map( B1 => n393, B2 => n504, C1 => n392, C2 => n505, A
                           => n506, ZN => O_34_port);
   U152 : AOI22_X1 port map( A1 => A_ns(33), A2 => n397, B1 => A_s(33), B2 => 
                           n398, ZN => n506);
   U153 : INV_X1 port map( A => A_s(32), ZN => n505);
   U154 : INV_X1 port map( A => A_ns(32), ZN => n504);
   U155 : OAI221_X1 port map( B1 => n393, B2 => n507, C1 => n392, C2 => n508, A
                           => n509, ZN => O_33_port);
   U156 : AOI22_X1 port map( A1 => A_ns(32), A2 => n397, B1 => A_s(32), B2 => 
                           n398, ZN => n509);
   U157 : INV_X1 port map( A => A_s(31), ZN => n508);
   U158 : INV_X1 port map( A => A_ns(31), ZN => n507);
   U159 : OAI221_X1 port map( B1 => n393, B2 => n510, C1 => n392, C2 => n511, A
                           => n512, ZN => O_32_port);
   U160 : AOI22_X1 port map( A1 => A_ns(31), A2 => n397, B1 => A_s(31), B2 => 
                           n398, ZN => n512);
   U161 : INV_X1 port map( A => A_s(30), ZN => n511);
   U162 : INV_X1 port map( A => A_ns(30), ZN => n510);
   U163 : OAI221_X1 port map( B1 => n393, B2 => n513, C1 => n392, C2 => n514, A
                           => n515, ZN => O_31_port);
   U164 : AOI22_X1 port map( A1 => A_ns(30), A2 => n397, B1 => A_s(30), B2 => 
                           n398, ZN => n515);
   U165 : INV_X1 port map( A => A_s(29), ZN => n514);
   U166 : INV_X1 port map( A => A_ns(29), ZN => n513);
   U167 : OAI221_X1 port map( B1 => n393, B2 => n516, C1 => n392, C2 => n517, A
                           => n518, ZN => O_30_port);
   U168 : AOI22_X1 port map( A1 => A_ns(29), A2 => n397, B1 => A_s(29), B2 => 
                           n398, ZN => n518);
   U169 : INV_X1 port map( A => A_s(28), ZN => n517);
   U170 : INV_X1 port map( A => A_ns(28), ZN => n516);
   U171 : OAI221_X1 port map( B1 => n393, B2 => n519, C1 => n392, C2 => n520, A
                           => n521, ZN => O_2_port);
   U172 : AOI22_X1 port map( A1 => A_ns(1), A2 => n397, B1 => A_s(1), B2 => 
                           n398, ZN => n521);
   U173 : OAI221_X1 port map( B1 => n393, B2 => n522, C1 => n392, C2 => n523, A
                           => n524, ZN => O_29_port);
   U174 : AOI22_X1 port map( A1 => A_ns(28), A2 => n397, B1 => A_s(28), B2 => 
                           n398, ZN => n524);
   U175 : INV_X1 port map( A => A_s(27), ZN => n523);
   U176 : INV_X1 port map( A => A_ns(27), ZN => n522);
   U177 : OAI221_X1 port map( B1 => n393, B2 => n525, C1 => n392, C2 => n526, A
                           => n527, ZN => O_28_port);
   U178 : AOI22_X1 port map( A1 => A_ns(27), A2 => n397, B1 => A_s(27), B2 => 
                           n398, ZN => n527);
   U179 : INV_X1 port map( A => A_s(26), ZN => n526);
   U180 : INV_X1 port map( A => A_ns(26), ZN => n525);
   U181 : OAI221_X1 port map( B1 => n393, B2 => n528, C1 => n392, C2 => n529, A
                           => n530, ZN => O_27_port);
   U182 : AOI22_X1 port map( A1 => A_ns(26), A2 => n397, B1 => A_s(26), B2 => 
                           n398, ZN => n530);
   U183 : INV_X1 port map( A => A_s(25), ZN => n529);
   U184 : INV_X1 port map( A => A_ns(25), ZN => n528);
   U185 : OAI221_X1 port map( B1 => n393, B2 => n531, C1 => n392, C2 => n532, A
                           => n533, ZN => O_26_port);
   U186 : AOI22_X1 port map( A1 => A_ns(25), A2 => n397, B1 => A_s(25), B2 => 
                           n398, ZN => n533);
   U187 : INV_X1 port map( A => A_s(24), ZN => n532);
   U188 : INV_X1 port map( A => A_ns(24), ZN => n531);
   U189 : OAI221_X1 port map( B1 => n393, B2 => n534, C1 => n392, C2 => n535, A
                           => n536, ZN => O_25_port);
   U190 : AOI22_X1 port map( A1 => A_ns(24), A2 => n397, B1 => A_s(24), B2 => 
                           n398, ZN => n536);
   U191 : INV_X1 port map( A => A_s(23), ZN => n535);
   U192 : INV_X1 port map( A => A_ns(23), ZN => n534);
   U193 : OAI221_X1 port map( B1 => n393, B2 => n537, C1 => n392, C2 => n538, A
                           => n539, ZN => O_24_port);
   U194 : AOI22_X1 port map( A1 => A_ns(23), A2 => n397, B1 => A_s(23), B2 => 
                           n398, ZN => n539);
   U195 : INV_X1 port map( A => A_s(22), ZN => n538);
   U196 : INV_X1 port map( A => A_ns(22), ZN => n537);
   U197 : OAI221_X1 port map( B1 => n393, B2 => n540, C1 => n392, C2 => n541, A
                           => n542, ZN => O_23_port);
   U198 : AOI22_X1 port map( A1 => A_ns(22), A2 => n397, B1 => A_s(22), B2 => 
                           n398, ZN => n542);
   U199 : INV_X1 port map( A => A_s(21), ZN => n541);
   U200 : INV_X1 port map( A => A_ns(21), ZN => n540);
   U201 : OAI221_X1 port map( B1 => n393, B2 => n543, C1 => n392, C2 => n544, A
                           => n545, ZN => O_22_port);
   U202 : AOI22_X1 port map( A1 => A_ns(21), A2 => n397, B1 => A_s(21), B2 => 
                           n398, ZN => n545);
   U203 : INV_X1 port map( A => A_s(20), ZN => n544);
   U204 : INV_X1 port map( A => A_ns(20), ZN => n543);
   U205 : OAI221_X1 port map( B1 => n393, B2 => n546, C1 => n392, C2 => n547, A
                           => n548, ZN => O_21_port);
   U206 : AOI22_X1 port map( A1 => A_ns(20), A2 => n397, B1 => A_s(20), B2 => 
                           n398, ZN => n548);
   U207 : INV_X1 port map( A => A_s(19), ZN => n547);
   U208 : INV_X1 port map( A => A_ns(19), ZN => n546);
   U209 : OAI221_X1 port map( B1 => n393, B2 => n549, C1 => n392, C2 => n550, A
                           => n551, ZN => O_20_port);
   U210 : AOI22_X1 port map( A1 => A_ns(19), A2 => n397, B1 => A_s(19), B2 => 
                           n398, ZN => n551);
   U211 : INV_X1 port map( A => A_s(18), ZN => n550);
   U212 : INV_X1 port map( A => A_ns(18), ZN => n549);
   U213 : OAI22_X1 port map( A1 => n552, A2 => n520, B1 => n553, B2 => n519, ZN
                           => O_1_port);
   U214 : INV_X1 port map( A => A_ns(0), ZN => n519);
   U215 : INV_X1 port map( A => A_s(0), ZN => n520);
   U216 : OAI221_X1 port map( B1 => n393, B2 => n554, C1 => n392, C2 => n555, A
                           => n556, ZN => O_19_port);
   U217 : AOI22_X1 port map( A1 => A_ns(18), A2 => n397, B1 => A_s(18), B2 => 
                           n398, ZN => n556);
   U218 : INV_X1 port map( A => A_s(17), ZN => n555);
   U219 : INV_X1 port map( A => A_ns(17), ZN => n554);
   U220 : OAI221_X1 port map( B1 => n393, B2 => n557, C1 => n392, C2 => n558, A
                           => n559, ZN => O_18_port);
   U221 : AOI22_X1 port map( A1 => A_ns(17), A2 => n397, B1 => A_s(17), B2 => 
                           n398, ZN => n559);
   U222 : INV_X1 port map( A => A_s(16), ZN => n558);
   U223 : INV_X1 port map( A => A_ns(16), ZN => n557);
   U224 : OAI221_X1 port map( B1 => n393, B2 => n560, C1 => n392, C2 => n561, A
                           => n562, ZN => O_17_port);
   U225 : AOI22_X1 port map( A1 => A_ns(16), A2 => n397, B1 => A_s(16), B2 => 
                           n398, ZN => n562);
   U226 : INV_X1 port map( A => A_s(15), ZN => n561);
   U227 : INV_X1 port map( A => A_ns(15), ZN => n560);
   U228 : OAI221_X1 port map( B1 => n393, B2 => n563, C1 => n392, C2 => n564, A
                           => n565, ZN => O_16_port);
   U229 : AOI22_X1 port map( A1 => A_ns(15), A2 => n397, B1 => A_s(15), B2 => 
                           n398, ZN => n565);
   U230 : INV_X1 port map( A => A_s(14), ZN => n564);
   U231 : INV_X1 port map( A => A_ns(14), ZN => n563);
   U232 : OAI221_X1 port map( B1 => n393, B2 => n566, C1 => n392, C2 => n567, A
                           => n568, ZN => O_15_port);
   U233 : AOI22_X1 port map( A1 => A_ns(14), A2 => n397, B1 => A_s(14), B2 => 
                           n398, ZN => n568);
   U234 : INV_X1 port map( A => A_s(13), ZN => n567);
   U235 : INV_X1 port map( A => A_ns(13), ZN => n566);
   U236 : OAI221_X1 port map( B1 => n393, B2 => n569, C1 => n392, C2 => n570, A
                           => n571, ZN => O_14_port);
   U237 : AOI22_X1 port map( A1 => A_ns(13), A2 => n397, B1 => A_s(13), B2 => 
                           n398, ZN => n571);
   U238 : INV_X1 port map( A => A_s(12), ZN => n570);
   U239 : INV_X1 port map( A => A_ns(12), ZN => n569);
   U240 : OAI221_X1 port map( B1 => n393, B2 => n572, C1 => n392, C2 => n573, A
                           => n574, ZN => O_13_port);
   U241 : AOI22_X1 port map( A1 => A_ns(12), A2 => n397, B1 => A_s(12), B2 => 
                           n398, ZN => n574);
   U242 : INV_X1 port map( A => A_s(11), ZN => n573);
   U243 : INV_X1 port map( A => A_ns(11), ZN => n572);
   U244 : OAI221_X1 port map( B1 => n393, B2 => n575, C1 => n392, C2 => n576, A
                           => n577, ZN => O_12_port);
   U245 : AOI22_X1 port map( A1 => A_ns(11), A2 => n397, B1 => A_s(11), B2 => 
                           n398, ZN => n577);
   U246 : INV_X1 port map( A => A_s(10), ZN => n576);
   U247 : INV_X1 port map( A => A_ns(10), ZN => n575);
   U248 : OAI221_X1 port map( B1 => n393, B2 => n578, C1 => n392, C2 => n579, A
                           => n580, ZN => O_11_port);
   U249 : AOI22_X1 port map( A1 => A_ns(10), A2 => n397, B1 => A_s(10), B2 => 
                           n398, ZN => n580);
   U250 : INV_X1 port map( A => A_s(9), ZN => n579);
   U251 : INV_X1 port map( A => A_ns(9), ZN => n578);
   U252 : OAI221_X1 port map( B1 => n581, B2 => n393, C1 => n582, C2 => n392, A
                           => n583, ZN => O_10_port);
   U253 : AOI22_X1 port map( A1 => A_ns(9), A2 => n397, B1 => A_s(9), B2 => 
                           n398, ZN => n583);
   U254 : NAND2_X1 port map( A1 => n584, A2 => n552, ZN => n553);
   U255 : NAND2_X1 port map( A1 => n584, A2 => n585, ZN => n552);
   U256 : XOR2_X1 port map( A => B(25), B => B(26), Z => n584);
   U257 : INV_X1 port map( A => A_s(8), ZN => n582);
   U258 : INV_X1 port map( A => B(27), ZN => n585);
   U259 : INV_X1 port map( A => A_ns(8), ZN => n581);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity BOOTHENC_NBIT64_i24 is

   port( A, A_n, A_ns, A_s, B : in std_logic_vector (63 downto 0);  O, A_so, 
         A_nso : out std_logic_vector (63 downto 0));

end BOOTHENC_NBIT64_i24;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT64_i24 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, O_63_port, O_62_port, O_61_port, O_60_port, O_59_port,
      O_58_port, O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, 
      O_52_port, O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, 
      O_46_port, O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, 
      O_40_port, O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, 
      O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, 
      O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, 
      O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, 
      O_16_port, O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, 
      O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, 
      O_3_port, O_2_port, O_1_port, n391, n392, n393, n394, n395, n396, n397, 
      n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, 
      n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, 
      n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, 
      n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, 
      n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, 
      n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, 
      n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, 
      n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, 
      n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, 
      n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, 
      n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, 
      n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, 
      n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, 
      n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, 
      n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, 
      n578, n579, n580, n581, n582, n583, n584, n585 : std_logic;

begin
   O <= ( O_63_port, O_62_port, O_61_port, O_60_port, O_59_port, O_58_port, 
      O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, O_52_port, 
      O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, O_46_port, 
      O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, O_40_port, 
      O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, 
      O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, 
      O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, 
      O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, O_16_port, 
      O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, O_10_port, 
      O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, O_3_port, 
      O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(61), A_s(60), A_s(59), A_s(58), A_s(57), A_s(56), A_s(55), 
      A_s(54), A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), 
      A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), 
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   A_nso <= ( A_s(61), A_s(60), A_s(59), A_s(58), A_s(57), A_s(56), A_s(55), 
      A_s(54), A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), 
      A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), 
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : AND3_X1 port map( A1 => B(24), A2 => n585, A3 => B(23), ZN => n391);
   U3 : INV_X4 port map( A => n391, ZN => n392);
   U4 : INV_X4 port map( A => n552, ZN => n398);
   U5 : OR3_X4 port map( A1 => B(23), A2 => B(24), A3 => n585, ZN => n393);
   U6 : INV_X4 port map( A => n553, ZN => n397);
   U7 : OAI221_X1 port map( B1 => n393, B2 => n394, C1 => n392, C2 => n395, A 
                           => n396, ZN => O_9_port);
   U8 : AOI22_X1 port map( A1 => A_ns(8), A2 => n397, B1 => A_s(8), B2 => n398,
                           ZN => n396);
   U9 : INV_X1 port map( A => A_s(7), ZN => n395);
   U10 : INV_X1 port map( A => A_ns(7), ZN => n394);
   U11 : OAI221_X1 port map( B1 => n393, B2 => n399, C1 => n392, C2 => n400, A 
                           => n401, ZN => O_8_port);
   U12 : AOI22_X1 port map( A1 => A_ns(7), A2 => n397, B1 => A_s(7), B2 => n398
                           , ZN => n401);
   U13 : INV_X1 port map( A => A_s(6), ZN => n400);
   U14 : INV_X1 port map( A => A_ns(6), ZN => n399);
   U15 : OAI221_X1 port map( B1 => n393, B2 => n402, C1 => n392, C2 => n403, A 
                           => n404, ZN => O_7_port);
   U16 : AOI22_X1 port map( A1 => A_ns(6), A2 => n397, B1 => A_s(6), B2 => n398
                           , ZN => n404);
   U17 : INV_X1 port map( A => A_s(5), ZN => n403);
   U18 : INV_X1 port map( A => A_ns(5), ZN => n402);
   U19 : OAI221_X1 port map( B1 => n393, B2 => n405, C1 => n392, C2 => n406, A 
                           => n407, ZN => O_6_port);
   U20 : AOI22_X1 port map( A1 => A_ns(5), A2 => n397, B1 => A_s(5), B2 => n398
                           , ZN => n407);
   U21 : INV_X1 port map( A => A_s(4), ZN => n406);
   U22 : INV_X1 port map( A => A_ns(4), ZN => n405);
   U23 : OAI221_X1 port map( B1 => n393, B2 => n408, C1 => n392, C2 => n409, A 
                           => n410, ZN => O_63_port);
   U24 : AOI22_X1 port map( A1 => A_ns(62), A2 => n397, B1 => A_s(62), B2 => 
                           n398, ZN => n410);
   U25 : INV_X1 port map( A => A_s(61), ZN => n409);
   U26 : INV_X1 port map( A => A_ns(61), ZN => n408);
   U27 : OAI221_X1 port map( B1 => n393, B2 => n411, C1 => n392, C2 => n412, A 
                           => n413, ZN => O_62_port);
   U28 : AOI22_X1 port map( A1 => A_ns(61), A2 => n397, B1 => A_s(61), B2 => 
                           n398, ZN => n413);
   U29 : INV_X1 port map( A => A_s(60), ZN => n412);
   U30 : INV_X1 port map( A => A_ns(60), ZN => n411);
   U31 : OAI221_X1 port map( B1 => n393, B2 => n414, C1 => n392, C2 => n415, A 
                           => n416, ZN => O_61_port);
   U32 : AOI22_X1 port map( A1 => A_ns(60), A2 => n397, B1 => A_s(60), B2 => 
                           n398, ZN => n416);
   U33 : INV_X1 port map( A => A_s(59), ZN => n415);
   U34 : INV_X1 port map( A => A_ns(59), ZN => n414);
   U35 : OAI221_X1 port map( B1 => n393, B2 => n417, C1 => n392, C2 => n418, A 
                           => n419, ZN => O_60_port);
   U36 : AOI22_X1 port map( A1 => A_ns(59), A2 => n397, B1 => A_s(59), B2 => 
                           n398, ZN => n419);
   U37 : INV_X1 port map( A => A_s(58), ZN => n418);
   U38 : INV_X1 port map( A => A_ns(58), ZN => n417);
   U39 : OAI221_X1 port map( B1 => n393, B2 => n420, C1 => n392, C2 => n421, A 
                           => n422, ZN => O_5_port);
   U40 : AOI22_X1 port map( A1 => A_ns(4), A2 => n397, B1 => A_s(4), B2 => n398
                           , ZN => n422);
   U41 : INV_X1 port map( A => A_s(3), ZN => n421);
   U42 : INV_X1 port map( A => A_ns(3), ZN => n420);
   U43 : OAI221_X1 port map( B1 => n393, B2 => n423, C1 => n392, C2 => n424, A 
                           => n425, ZN => O_59_port);
   U44 : AOI22_X1 port map( A1 => A_ns(58), A2 => n397, B1 => A_s(58), B2 => 
                           n398, ZN => n425);
   U45 : INV_X1 port map( A => A_s(57), ZN => n424);
   U46 : INV_X1 port map( A => A_ns(57), ZN => n423);
   U47 : OAI221_X1 port map( B1 => n393, B2 => n426, C1 => n392, C2 => n427, A 
                           => n428, ZN => O_58_port);
   U48 : AOI22_X1 port map( A1 => A_ns(57), A2 => n397, B1 => A_s(57), B2 => 
                           n398, ZN => n428);
   U49 : INV_X1 port map( A => A_s(56), ZN => n427);
   U50 : INV_X1 port map( A => A_ns(56), ZN => n426);
   U51 : OAI221_X1 port map( B1 => n393, B2 => n429, C1 => n392, C2 => n430, A 
                           => n431, ZN => O_57_port);
   U52 : AOI22_X1 port map( A1 => A_ns(56), A2 => n397, B1 => A_s(56), B2 => 
                           n398, ZN => n431);
   U53 : INV_X1 port map( A => A_s(55), ZN => n430);
   U54 : INV_X1 port map( A => A_ns(55), ZN => n429);
   U55 : OAI221_X1 port map( B1 => n393, B2 => n432, C1 => n392, C2 => n433, A 
                           => n434, ZN => O_56_port);
   U56 : AOI22_X1 port map( A1 => A_ns(55), A2 => n397, B1 => A_s(55), B2 => 
                           n398, ZN => n434);
   U57 : INV_X1 port map( A => A_s(54), ZN => n433);
   U58 : INV_X1 port map( A => A_ns(54), ZN => n432);
   U59 : OAI221_X1 port map( B1 => n393, B2 => n435, C1 => n392, C2 => n436, A 
                           => n437, ZN => O_55_port);
   U60 : AOI22_X1 port map( A1 => A_ns(54), A2 => n397, B1 => A_s(54), B2 => 
                           n398, ZN => n437);
   U61 : INV_X1 port map( A => A_s(53), ZN => n436);
   U62 : INV_X1 port map( A => A_ns(53), ZN => n435);
   U63 : OAI221_X1 port map( B1 => n393, B2 => n438, C1 => n392, C2 => n439, A 
                           => n440, ZN => O_54_port);
   U64 : AOI22_X1 port map( A1 => A_ns(53), A2 => n397, B1 => A_s(53), B2 => 
                           n398, ZN => n440);
   U65 : INV_X1 port map( A => A_s(52), ZN => n439);
   U66 : INV_X1 port map( A => A_ns(52), ZN => n438);
   U67 : OAI221_X1 port map( B1 => n393, B2 => n441, C1 => n392, C2 => n442, A 
                           => n443, ZN => O_53_port);
   U68 : AOI22_X1 port map( A1 => A_ns(52), A2 => n397, B1 => A_s(52), B2 => 
                           n398, ZN => n443);
   U69 : INV_X1 port map( A => A_s(51), ZN => n442);
   U70 : INV_X1 port map( A => A_ns(51), ZN => n441);
   U71 : OAI221_X1 port map( B1 => n393, B2 => n444, C1 => n392, C2 => n445, A 
                           => n446, ZN => O_52_port);
   U72 : AOI22_X1 port map( A1 => A_ns(51), A2 => n397, B1 => A_s(51), B2 => 
                           n398, ZN => n446);
   U73 : INV_X1 port map( A => A_s(50), ZN => n445);
   U74 : INV_X1 port map( A => A_ns(50), ZN => n444);
   U75 : OAI221_X1 port map( B1 => n393, B2 => n447, C1 => n392, C2 => n448, A 
                           => n449, ZN => O_51_port);
   U76 : AOI22_X1 port map( A1 => A_ns(50), A2 => n397, B1 => A_s(50), B2 => 
                           n398, ZN => n449);
   U77 : INV_X1 port map( A => A_s(49), ZN => n448);
   U78 : INV_X1 port map( A => A_ns(49), ZN => n447);
   U79 : OAI221_X1 port map( B1 => n393, B2 => n450, C1 => n392, C2 => n451, A 
                           => n452, ZN => O_50_port);
   U80 : AOI22_X1 port map( A1 => A_ns(49), A2 => n397, B1 => A_s(49), B2 => 
                           n398, ZN => n452);
   U81 : INV_X1 port map( A => A_s(48), ZN => n451);
   U82 : INV_X1 port map( A => A_ns(48), ZN => n450);
   U83 : OAI221_X1 port map( B1 => n393, B2 => n453, C1 => n392, C2 => n454, A 
                           => n455, ZN => O_4_port);
   U84 : AOI22_X1 port map( A1 => A_ns(3), A2 => n397, B1 => A_s(3), B2 => n398
                           , ZN => n455);
   U85 : INV_X1 port map( A => A_s(2), ZN => n454);
   U86 : INV_X1 port map( A => A_ns(2), ZN => n453);
   U87 : OAI221_X1 port map( B1 => n393, B2 => n456, C1 => n392, C2 => n457, A 
                           => n458, ZN => O_49_port);
   U88 : AOI22_X1 port map( A1 => A_ns(48), A2 => n397, B1 => A_s(48), B2 => 
                           n398, ZN => n458);
   U89 : INV_X1 port map( A => A_s(47), ZN => n457);
   U90 : INV_X1 port map( A => A_ns(47), ZN => n456);
   U91 : OAI221_X1 port map( B1 => n393, B2 => n459, C1 => n392, C2 => n460, A 
                           => n461, ZN => O_48_port);
   U92 : AOI22_X1 port map( A1 => A_ns(47), A2 => n397, B1 => A_s(47), B2 => 
                           n398, ZN => n461);
   U93 : INV_X1 port map( A => A_s(46), ZN => n460);
   U94 : INV_X1 port map( A => A_ns(46), ZN => n459);
   U95 : OAI221_X1 port map( B1 => n393, B2 => n462, C1 => n392, C2 => n463, A 
                           => n464, ZN => O_47_port);
   U96 : AOI22_X1 port map( A1 => A_ns(46), A2 => n397, B1 => A_s(46), B2 => 
                           n398, ZN => n464);
   U97 : INV_X1 port map( A => A_s(45), ZN => n463);
   U98 : INV_X1 port map( A => A_ns(45), ZN => n462);
   U99 : OAI221_X1 port map( B1 => n393, B2 => n465, C1 => n392, C2 => n466, A 
                           => n467, ZN => O_46_port);
   U100 : AOI22_X1 port map( A1 => A_ns(45), A2 => n397, B1 => A_s(45), B2 => 
                           n398, ZN => n467);
   U101 : INV_X1 port map( A => A_s(44), ZN => n466);
   U102 : INV_X1 port map( A => A_ns(44), ZN => n465);
   U103 : OAI221_X1 port map( B1 => n393, B2 => n468, C1 => n392, C2 => n469, A
                           => n470, ZN => O_45_port);
   U104 : AOI22_X1 port map( A1 => A_ns(44), A2 => n397, B1 => A_s(44), B2 => 
                           n398, ZN => n470);
   U105 : INV_X1 port map( A => A_s(43), ZN => n469);
   U106 : INV_X1 port map( A => A_ns(43), ZN => n468);
   U107 : OAI221_X1 port map( B1 => n393, B2 => n471, C1 => n392, C2 => n472, A
                           => n473, ZN => O_44_port);
   U108 : AOI22_X1 port map( A1 => A_ns(43), A2 => n397, B1 => A_s(43), B2 => 
                           n398, ZN => n473);
   U109 : INV_X1 port map( A => A_s(42), ZN => n472);
   U110 : INV_X1 port map( A => A_ns(42), ZN => n471);
   U111 : OAI221_X1 port map( B1 => n393, B2 => n474, C1 => n392, C2 => n475, A
                           => n476, ZN => O_43_port);
   U112 : AOI22_X1 port map( A1 => A_ns(42), A2 => n397, B1 => A_s(42), B2 => 
                           n398, ZN => n476);
   U113 : INV_X1 port map( A => A_s(41), ZN => n475);
   U114 : INV_X1 port map( A => A_ns(41), ZN => n474);
   U115 : OAI221_X1 port map( B1 => n393, B2 => n477, C1 => n392, C2 => n478, A
                           => n479, ZN => O_42_port);
   U116 : AOI22_X1 port map( A1 => A_ns(41), A2 => n397, B1 => A_s(41), B2 => 
                           n398, ZN => n479);
   U117 : INV_X1 port map( A => A_s(40), ZN => n478);
   U118 : INV_X1 port map( A => A_ns(40), ZN => n477);
   U119 : OAI221_X1 port map( B1 => n393, B2 => n480, C1 => n392, C2 => n481, A
                           => n482, ZN => O_41_port);
   U120 : AOI22_X1 port map( A1 => A_ns(40), A2 => n397, B1 => A_s(40), B2 => 
                           n398, ZN => n482);
   U121 : INV_X1 port map( A => A_s(39), ZN => n481);
   U122 : INV_X1 port map( A => A_ns(39), ZN => n480);
   U123 : OAI221_X1 port map( B1 => n393, B2 => n483, C1 => n392, C2 => n484, A
                           => n485, ZN => O_40_port);
   U124 : AOI22_X1 port map( A1 => A_ns(39), A2 => n397, B1 => A_s(39), B2 => 
                           n398, ZN => n485);
   U125 : INV_X1 port map( A => A_s(38), ZN => n484);
   U126 : INV_X1 port map( A => A_ns(38), ZN => n483);
   U127 : OAI221_X1 port map( B1 => n393, B2 => n486, C1 => n392, C2 => n487, A
                           => n488, ZN => O_3_port);
   U128 : AOI22_X1 port map( A1 => A_ns(2), A2 => n397, B1 => A_s(2), B2 => 
                           n398, ZN => n488);
   U129 : INV_X1 port map( A => A_s(1), ZN => n487);
   U130 : INV_X1 port map( A => A_ns(1), ZN => n486);
   U131 : OAI221_X1 port map( B1 => n393, B2 => n489, C1 => n392, C2 => n490, A
                           => n491, ZN => O_39_port);
   U132 : AOI22_X1 port map( A1 => A_ns(38), A2 => n397, B1 => A_s(38), B2 => 
                           n398, ZN => n491);
   U133 : INV_X1 port map( A => A_s(37), ZN => n490);
   U134 : INV_X1 port map( A => A_ns(37), ZN => n489);
   U135 : OAI221_X1 port map( B1 => n393, B2 => n492, C1 => n392, C2 => n493, A
                           => n494, ZN => O_38_port);
   U136 : AOI22_X1 port map( A1 => A_ns(37), A2 => n397, B1 => A_s(37), B2 => 
                           n398, ZN => n494);
   U137 : INV_X1 port map( A => A_s(36), ZN => n493);
   U138 : INV_X1 port map( A => A_ns(36), ZN => n492);
   U139 : OAI221_X1 port map( B1 => n393, B2 => n495, C1 => n392, C2 => n496, A
                           => n497, ZN => O_37_port);
   U140 : AOI22_X1 port map( A1 => A_ns(36), A2 => n397, B1 => A_s(36), B2 => 
                           n398, ZN => n497);
   U141 : INV_X1 port map( A => A_s(35), ZN => n496);
   U142 : INV_X1 port map( A => A_ns(35), ZN => n495);
   U143 : OAI221_X1 port map( B1 => n393, B2 => n498, C1 => n392, C2 => n499, A
                           => n500, ZN => O_36_port);
   U144 : AOI22_X1 port map( A1 => A_ns(35), A2 => n397, B1 => A_s(35), B2 => 
                           n398, ZN => n500);
   U145 : INV_X1 port map( A => A_s(34), ZN => n499);
   U146 : INV_X1 port map( A => A_ns(34), ZN => n498);
   U147 : OAI221_X1 port map( B1 => n393, B2 => n501, C1 => n392, C2 => n502, A
                           => n503, ZN => O_35_port);
   U148 : AOI22_X1 port map( A1 => A_ns(34), A2 => n397, B1 => A_s(34), B2 => 
                           n398, ZN => n503);
   U149 : INV_X1 port map( A => A_s(33), ZN => n502);
   U150 : INV_X1 port map( A => A_ns(33), ZN => n501);
   U151 : OAI221_X1 port map( B1 => n393, B2 => n504, C1 => n392, C2 => n505, A
                           => n506, ZN => O_34_port);
   U152 : AOI22_X1 port map( A1 => A_ns(33), A2 => n397, B1 => A_s(33), B2 => 
                           n398, ZN => n506);
   U153 : INV_X1 port map( A => A_s(32), ZN => n505);
   U154 : INV_X1 port map( A => A_ns(32), ZN => n504);
   U155 : OAI221_X1 port map( B1 => n393, B2 => n507, C1 => n392, C2 => n508, A
                           => n509, ZN => O_33_port);
   U156 : AOI22_X1 port map( A1 => A_ns(32), A2 => n397, B1 => A_s(32), B2 => 
                           n398, ZN => n509);
   U157 : INV_X1 port map( A => A_s(31), ZN => n508);
   U158 : INV_X1 port map( A => A_ns(31), ZN => n507);
   U159 : OAI221_X1 port map( B1 => n393, B2 => n510, C1 => n392, C2 => n511, A
                           => n512, ZN => O_32_port);
   U160 : AOI22_X1 port map( A1 => A_ns(31), A2 => n397, B1 => A_s(31), B2 => 
                           n398, ZN => n512);
   U161 : INV_X1 port map( A => A_s(30), ZN => n511);
   U162 : INV_X1 port map( A => A_ns(30), ZN => n510);
   U163 : OAI221_X1 port map( B1 => n393, B2 => n513, C1 => n392, C2 => n514, A
                           => n515, ZN => O_31_port);
   U164 : AOI22_X1 port map( A1 => A_ns(30), A2 => n397, B1 => A_s(30), B2 => 
                           n398, ZN => n515);
   U165 : INV_X1 port map( A => A_s(29), ZN => n514);
   U166 : INV_X1 port map( A => A_ns(29), ZN => n513);
   U167 : OAI221_X1 port map( B1 => n393, B2 => n516, C1 => n392, C2 => n517, A
                           => n518, ZN => O_30_port);
   U168 : AOI22_X1 port map( A1 => A_ns(29), A2 => n397, B1 => A_s(29), B2 => 
                           n398, ZN => n518);
   U169 : INV_X1 port map( A => A_s(28), ZN => n517);
   U170 : INV_X1 port map( A => A_ns(28), ZN => n516);
   U171 : OAI221_X1 port map( B1 => n393, B2 => n519, C1 => n392, C2 => n520, A
                           => n521, ZN => O_2_port);
   U172 : AOI22_X1 port map( A1 => A_ns(1), A2 => n397, B1 => A_s(1), B2 => 
                           n398, ZN => n521);
   U173 : OAI221_X1 port map( B1 => n393, B2 => n522, C1 => n392, C2 => n523, A
                           => n524, ZN => O_29_port);
   U174 : AOI22_X1 port map( A1 => A_ns(28), A2 => n397, B1 => A_s(28), B2 => 
                           n398, ZN => n524);
   U175 : INV_X1 port map( A => A_s(27), ZN => n523);
   U176 : INV_X1 port map( A => A_ns(27), ZN => n522);
   U177 : OAI221_X1 port map( B1 => n393, B2 => n525, C1 => n392, C2 => n526, A
                           => n527, ZN => O_28_port);
   U178 : AOI22_X1 port map( A1 => A_ns(27), A2 => n397, B1 => A_s(27), B2 => 
                           n398, ZN => n527);
   U179 : INV_X1 port map( A => A_s(26), ZN => n526);
   U180 : INV_X1 port map( A => A_ns(26), ZN => n525);
   U181 : OAI221_X1 port map( B1 => n393, B2 => n528, C1 => n392, C2 => n529, A
                           => n530, ZN => O_27_port);
   U182 : AOI22_X1 port map( A1 => A_ns(26), A2 => n397, B1 => A_s(26), B2 => 
                           n398, ZN => n530);
   U183 : INV_X1 port map( A => A_s(25), ZN => n529);
   U184 : INV_X1 port map( A => A_ns(25), ZN => n528);
   U185 : OAI221_X1 port map( B1 => n393, B2 => n531, C1 => n392, C2 => n532, A
                           => n533, ZN => O_26_port);
   U186 : AOI22_X1 port map( A1 => A_ns(25), A2 => n397, B1 => A_s(25), B2 => 
                           n398, ZN => n533);
   U187 : INV_X1 port map( A => A_s(24), ZN => n532);
   U188 : INV_X1 port map( A => A_ns(24), ZN => n531);
   U189 : OAI221_X1 port map( B1 => n393, B2 => n534, C1 => n392, C2 => n535, A
                           => n536, ZN => O_25_port);
   U190 : AOI22_X1 port map( A1 => A_ns(24), A2 => n397, B1 => A_s(24), B2 => 
                           n398, ZN => n536);
   U191 : INV_X1 port map( A => A_s(23), ZN => n535);
   U192 : INV_X1 port map( A => A_ns(23), ZN => n534);
   U193 : OAI221_X1 port map( B1 => n393, B2 => n537, C1 => n392, C2 => n538, A
                           => n539, ZN => O_24_port);
   U194 : AOI22_X1 port map( A1 => A_ns(23), A2 => n397, B1 => A_s(23), B2 => 
                           n398, ZN => n539);
   U195 : INV_X1 port map( A => A_s(22), ZN => n538);
   U196 : INV_X1 port map( A => A_ns(22), ZN => n537);
   U197 : OAI221_X1 port map( B1 => n393, B2 => n540, C1 => n392, C2 => n541, A
                           => n542, ZN => O_23_port);
   U198 : AOI22_X1 port map( A1 => A_ns(22), A2 => n397, B1 => A_s(22), B2 => 
                           n398, ZN => n542);
   U199 : INV_X1 port map( A => A_s(21), ZN => n541);
   U200 : INV_X1 port map( A => A_ns(21), ZN => n540);
   U201 : OAI221_X1 port map( B1 => n393, B2 => n543, C1 => n392, C2 => n544, A
                           => n545, ZN => O_22_port);
   U202 : AOI22_X1 port map( A1 => A_ns(21), A2 => n397, B1 => A_s(21), B2 => 
                           n398, ZN => n545);
   U203 : INV_X1 port map( A => A_s(20), ZN => n544);
   U204 : INV_X1 port map( A => A_ns(20), ZN => n543);
   U205 : OAI221_X1 port map( B1 => n393, B2 => n546, C1 => n392, C2 => n547, A
                           => n548, ZN => O_21_port);
   U206 : AOI22_X1 port map( A1 => A_ns(20), A2 => n397, B1 => A_s(20), B2 => 
                           n398, ZN => n548);
   U207 : INV_X1 port map( A => A_s(19), ZN => n547);
   U208 : INV_X1 port map( A => A_ns(19), ZN => n546);
   U209 : OAI221_X1 port map( B1 => n393, B2 => n549, C1 => n392, C2 => n550, A
                           => n551, ZN => O_20_port);
   U210 : AOI22_X1 port map( A1 => A_ns(19), A2 => n397, B1 => A_s(19), B2 => 
                           n398, ZN => n551);
   U211 : INV_X1 port map( A => A_s(18), ZN => n550);
   U212 : INV_X1 port map( A => A_ns(18), ZN => n549);
   U213 : OAI22_X1 port map( A1 => n552, A2 => n520, B1 => n553, B2 => n519, ZN
                           => O_1_port);
   U214 : INV_X1 port map( A => A_ns(0), ZN => n519);
   U215 : INV_X1 port map( A => A_s(0), ZN => n520);
   U216 : OAI221_X1 port map( B1 => n393, B2 => n554, C1 => n392, C2 => n555, A
                           => n556, ZN => O_19_port);
   U217 : AOI22_X1 port map( A1 => A_ns(18), A2 => n397, B1 => A_s(18), B2 => 
                           n398, ZN => n556);
   U218 : INV_X1 port map( A => A_s(17), ZN => n555);
   U219 : INV_X1 port map( A => A_ns(17), ZN => n554);
   U220 : OAI221_X1 port map( B1 => n393, B2 => n557, C1 => n392, C2 => n558, A
                           => n559, ZN => O_18_port);
   U221 : AOI22_X1 port map( A1 => A_ns(17), A2 => n397, B1 => A_s(17), B2 => 
                           n398, ZN => n559);
   U222 : INV_X1 port map( A => A_s(16), ZN => n558);
   U223 : INV_X1 port map( A => A_ns(16), ZN => n557);
   U224 : OAI221_X1 port map( B1 => n393, B2 => n560, C1 => n392, C2 => n561, A
                           => n562, ZN => O_17_port);
   U225 : AOI22_X1 port map( A1 => A_ns(16), A2 => n397, B1 => A_s(16), B2 => 
                           n398, ZN => n562);
   U226 : INV_X1 port map( A => A_s(15), ZN => n561);
   U227 : INV_X1 port map( A => A_ns(15), ZN => n560);
   U228 : OAI221_X1 port map( B1 => n393, B2 => n563, C1 => n392, C2 => n564, A
                           => n565, ZN => O_16_port);
   U229 : AOI22_X1 port map( A1 => A_ns(15), A2 => n397, B1 => A_s(15), B2 => 
                           n398, ZN => n565);
   U230 : INV_X1 port map( A => A_s(14), ZN => n564);
   U231 : INV_X1 port map( A => A_ns(14), ZN => n563);
   U232 : OAI221_X1 port map( B1 => n393, B2 => n566, C1 => n392, C2 => n567, A
                           => n568, ZN => O_15_port);
   U233 : AOI22_X1 port map( A1 => A_ns(14), A2 => n397, B1 => A_s(14), B2 => 
                           n398, ZN => n568);
   U234 : INV_X1 port map( A => A_s(13), ZN => n567);
   U235 : INV_X1 port map( A => A_ns(13), ZN => n566);
   U236 : OAI221_X1 port map( B1 => n393, B2 => n569, C1 => n392, C2 => n570, A
                           => n571, ZN => O_14_port);
   U237 : AOI22_X1 port map( A1 => A_ns(13), A2 => n397, B1 => A_s(13), B2 => 
                           n398, ZN => n571);
   U238 : INV_X1 port map( A => A_s(12), ZN => n570);
   U239 : INV_X1 port map( A => A_ns(12), ZN => n569);
   U240 : OAI221_X1 port map( B1 => n393, B2 => n572, C1 => n392, C2 => n573, A
                           => n574, ZN => O_13_port);
   U241 : AOI22_X1 port map( A1 => A_ns(12), A2 => n397, B1 => A_s(12), B2 => 
                           n398, ZN => n574);
   U242 : INV_X1 port map( A => A_s(11), ZN => n573);
   U243 : INV_X1 port map( A => A_ns(11), ZN => n572);
   U244 : OAI221_X1 port map( B1 => n393, B2 => n575, C1 => n392, C2 => n576, A
                           => n577, ZN => O_12_port);
   U245 : AOI22_X1 port map( A1 => A_ns(11), A2 => n397, B1 => A_s(11), B2 => 
                           n398, ZN => n577);
   U246 : INV_X1 port map( A => A_s(10), ZN => n576);
   U247 : INV_X1 port map( A => A_ns(10), ZN => n575);
   U248 : OAI221_X1 port map( B1 => n393, B2 => n578, C1 => n392, C2 => n579, A
                           => n580, ZN => O_11_port);
   U249 : AOI22_X1 port map( A1 => A_ns(10), A2 => n397, B1 => A_s(10), B2 => 
                           n398, ZN => n580);
   U250 : INV_X1 port map( A => A_s(9), ZN => n579);
   U251 : INV_X1 port map( A => A_ns(9), ZN => n578);
   U252 : OAI221_X1 port map( B1 => n581, B2 => n393, C1 => n582, C2 => n392, A
                           => n583, ZN => O_10_port);
   U253 : AOI22_X1 port map( A1 => A_ns(9), A2 => n397, B1 => A_s(9), B2 => 
                           n398, ZN => n583);
   U254 : NAND2_X1 port map( A1 => n584, A2 => n552, ZN => n553);
   U255 : NAND2_X1 port map( A1 => n584, A2 => n585, ZN => n552);
   U256 : XOR2_X1 port map( A => B(23), B => B(24), Z => n584);
   U257 : INV_X1 port map( A => A_s(8), ZN => n582);
   U258 : INV_X1 port map( A => B(25), ZN => n585);
   U259 : INV_X1 port map( A => A_ns(8), ZN => n581);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity BOOTHENC_NBIT64_i22 is

   port( A, A_n, A_ns, A_s, B : in std_logic_vector (63 downto 0);  O, A_so, 
         A_nso : out std_logic_vector (63 downto 0));

end BOOTHENC_NBIT64_i22;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT64_i22 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, O_63_port, O_62_port, O_61_port, O_60_port, O_59_port,
      O_58_port, O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, 
      O_52_port, O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, 
      O_46_port, O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, 
      O_40_port, O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, 
      O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, 
      O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, 
      O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, 
      O_16_port, O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, 
      O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, 
      O_3_port, O_2_port, O_1_port, n391, n392, n393, n394, n395, n396, n397, 
      n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, 
      n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, 
      n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, 
      n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, 
      n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, 
      n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, 
      n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, 
      n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, 
      n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, 
      n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, 
      n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, 
      n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, 
      n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, 
      n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, 
      n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, 
      n578, n579, n580, n581, n582, n583, n584, n585 : std_logic;

begin
   O <= ( O_63_port, O_62_port, O_61_port, O_60_port, O_59_port, O_58_port, 
      O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, O_52_port, 
      O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, O_46_port, 
      O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, O_40_port, 
      O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, 
      O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, 
      O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, 
      O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, O_16_port, 
      O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, O_10_port, 
      O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, O_3_port, 
      O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(61), A_s(60), A_s(59), A_s(58), A_s(57), A_s(56), A_s(55), 
      A_s(54), A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), 
      A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), 
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   A_nso <= ( A_s(61), A_s(60), A_s(59), A_s(58), A_s(57), A_s(56), A_s(55), 
      A_s(54), A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), 
      A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), 
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : AND3_X1 port map( A1 => B(22), A2 => n585, A3 => B(21), ZN => n391);
   U3 : INV_X4 port map( A => n391, ZN => n392);
   U4 : INV_X4 port map( A => n552, ZN => n398);
   U5 : OR3_X4 port map( A1 => B(21), A2 => B(22), A3 => n585, ZN => n393);
   U6 : INV_X4 port map( A => n553, ZN => n397);
   U7 : OAI221_X1 port map( B1 => n393, B2 => n394, C1 => n392, C2 => n395, A 
                           => n396, ZN => O_9_port);
   U8 : AOI22_X1 port map( A1 => A_ns(8), A2 => n397, B1 => A_s(8), B2 => n398,
                           ZN => n396);
   U9 : INV_X1 port map( A => A_s(7), ZN => n395);
   U10 : INV_X1 port map( A => A_ns(7), ZN => n394);
   U11 : OAI221_X1 port map( B1 => n393, B2 => n399, C1 => n392, C2 => n400, A 
                           => n401, ZN => O_8_port);
   U12 : AOI22_X1 port map( A1 => A_ns(7), A2 => n397, B1 => A_s(7), B2 => n398
                           , ZN => n401);
   U13 : INV_X1 port map( A => A_s(6), ZN => n400);
   U14 : INV_X1 port map( A => A_ns(6), ZN => n399);
   U15 : OAI221_X1 port map( B1 => n393, B2 => n402, C1 => n392, C2 => n403, A 
                           => n404, ZN => O_7_port);
   U16 : AOI22_X1 port map( A1 => A_ns(6), A2 => n397, B1 => A_s(6), B2 => n398
                           , ZN => n404);
   U17 : INV_X1 port map( A => A_s(5), ZN => n403);
   U18 : INV_X1 port map( A => A_ns(5), ZN => n402);
   U19 : OAI221_X1 port map( B1 => n393, B2 => n405, C1 => n392, C2 => n406, A 
                           => n407, ZN => O_6_port);
   U20 : AOI22_X1 port map( A1 => A_ns(5), A2 => n397, B1 => A_s(5), B2 => n398
                           , ZN => n407);
   U21 : INV_X1 port map( A => A_s(4), ZN => n406);
   U22 : INV_X1 port map( A => A_ns(4), ZN => n405);
   U23 : OAI221_X1 port map( B1 => n393, B2 => n408, C1 => n392, C2 => n409, A 
                           => n410, ZN => O_63_port);
   U24 : AOI22_X1 port map( A1 => A_ns(62), A2 => n397, B1 => A_s(62), B2 => 
                           n398, ZN => n410);
   U25 : INV_X1 port map( A => A_s(61), ZN => n409);
   U26 : INV_X1 port map( A => A_ns(61), ZN => n408);
   U27 : OAI221_X1 port map( B1 => n393, B2 => n411, C1 => n392, C2 => n412, A 
                           => n413, ZN => O_62_port);
   U28 : AOI22_X1 port map( A1 => A_ns(61), A2 => n397, B1 => A_s(61), B2 => 
                           n398, ZN => n413);
   U29 : INV_X1 port map( A => A_s(60), ZN => n412);
   U30 : INV_X1 port map( A => A_ns(60), ZN => n411);
   U31 : OAI221_X1 port map( B1 => n393, B2 => n414, C1 => n392, C2 => n415, A 
                           => n416, ZN => O_61_port);
   U32 : AOI22_X1 port map( A1 => A_ns(60), A2 => n397, B1 => A_s(60), B2 => 
                           n398, ZN => n416);
   U33 : INV_X1 port map( A => A_s(59), ZN => n415);
   U34 : INV_X1 port map( A => A_ns(59), ZN => n414);
   U35 : OAI221_X1 port map( B1 => n393, B2 => n417, C1 => n392, C2 => n418, A 
                           => n419, ZN => O_60_port);
   U36 : AOI22_X1 port map( A1 => A_ns(59), A2 => n397, B1 => A_s(59), B2 => 
                           n398, ZN => n419);
   U37 : INV_X1 port map( A => A_s(58), ZN => n418);
   U38 : INV_X1 port map( A => A_ns(58), ZN => n417);
   U39 : OAI221_X1 port map( B1 => n393, B2 => n420, C1 => n392, C2 => n421, A 
                           => n422, ZN => O_5_port);
   U40 : AOI22_X1 port map( A1 => A_ns(4), A2 => n397, B1 => A_s(4), B2 => n398
                           , ZN => n422);
   U41 : INV_X1 port map( A => A_s(3), ZN => n421);
   U42 : INV_X1 port map( A => A_ns(3), ZN => n420);
   U43 : OAI221_X1 port map( B1 => n393, B2 => n423, C1 => n392, C2 => n424, A 
                           => n425, ZN => O_59_port);
   U44 : AOI22_X1 port map( A1 => A_ns(58), A2 => n397, B1 => A_s(58), B2 => 
                           n398, ZN => n425);
   U45 : INV_X1 port map( A => A_s(57), ZN => n424);
   U46 : INV_X1 port map( A => A_ns(57), ZN => n423);
   U47 : OAI221_X1 port map( B1 => n393, B2 => n426, C1 => n392, C2 => n427, A 
                           => n428, ZN => O_58_port);
   U48 : AOI22_X1 port map( A1 => A_ns(57), A2 => n397, B1 => A_s(57), B2 => 
                           n398, ZN => n428);
   U49 : INV_X1 port map( A => A_s(56), ZN => n427);
   U50 : INV_X1 port map( A => A_ns(56), ZN => n426);
   U51 : OAI221_X1 port map( B1 => n393, B2 => n429, C1 => n392, C2 => n430, A 
                           => n431, ZN => O_57_port);
   U52 : AOI22_X1 port map( A1 => A_ns(56), A2 => n397, B1 => A_s(56), B2 => 
                           n398, ZN => n431);
   U53 : INV_X1 port map( A => A_s(55), ZN => n430);
   U54 : INV_X1 port map( A => A_ns(55), ZN => n429);
   U55 : OAI221_X1 port map( B1 => n393, B2 => n432, C1 => n392, C2 => n433, A 
                           => n434, ZN => O_56_port);
   U56 : AOI22_X1 port map( A1 => A_ns(55), A2 => n397, B1 => A_s(55), B2 => 
                           n398, ZN => n434);
   U57 : INV_X1 port map( A => A_s(54), ZN => n433);
   U58 : INV_X1 port map( A => A_ns(54), ZN => n432);
   U59 : OAI221_X1 port map( B1 => n393, B2 => n435, C1 => n392, C2 => n436, A 
                           => n437, ZN => O_55_port);
   U60 : AOI22_X1 port map( A1 => A_ns(54), A2 => n397, B1 => A_s(54), B2 => 
                           n398, ZN => n437);
   U61 : INV_X1 port map( A => A_s(53), ZN => n436);
   U62 : INV_X1 port map( A => A_ns(53), ZN => n435);
   U63 : OAI221_X1 port map( B1 => n393, B2 => n438, C1 => n392, C2 => n439, A 
                           => n440, ZN => O_54_port);
   U64 : AOI22_X1 port map( A1 => A_ns(53), A2 => n397, B1 => A_s(53), B2 => 
                           n398, ZN => n440);
   U65 : INV_X1 port map( A => A_s(52), ZN => n439);
   U66 : INV_X1 port map( A => A_ns(52), ZN => n438);
   U67 : OAI221_X1 port map( B1 => n393, B2 => n441, C1 => n392, C2 => n442, A 
                           => n443, ZN => O_53_port);
   U68 : AOI22_X1 port map( A1 => A_ns(52), A2 => n397, B1 => A_s(52), B2 => 
                           n398, ZN => n443);
   U69 : INV_X1 port map( A => A_s(51), ZN => n442);
   U70 : INV_X1 port map( A => A_ns(51), ZN => n441);
   U71 : OAI221_X1 port map( B1 => n393, B2 => n444, C1 => n392, C2 => n445, A 
                           => n446, ZN => O_52_port);
   U72 : AOI22_X1 port map( A1 => A_ns(51), A2 => n397, B1 => A_s(51), B2 => 
                           n398, ZN => n446);
   U73 : INV_X1 port map( A => A_s(50), ZN => n445);
   U74 : INV_X1 port map( A => A_ns(50), ZN => n444);
   U75 : OAI221_X1 port map( B1 => n393, B2 => n447, C1 => n392, C2 => n448, A 
                           => n449, ZN => O_51_port);
   U76 : AOI22_X1 port map( A1 => A_ns(50), A2 => n397, B1 => A_s(50), B2 => 
                           n398, ZN => n449);
   U77 : INV_X1 port map( A => A_s(49), ZN => n448);
   U78 : INV_X1 port map( A => A_ns(49), ZN => n447);
   U79 : OAI221_X1 port map( B1 => n393, B2 => n450, C1 => n392, C2 => n451, A 
                           => n452, ZN => O_50_port);
   U80 : AOI22_X1 port map( A1 => A_ns(49), A2 => n397, B1 => A_s(49), B2 => 
                           n398, ZN => n452);
   U81 : INV_X1 port map( A => A_s(48), ZN => n451);
   U82 : INV_X1 port map( A => A_ns(48), ZN => n450);
   U83 : OAI221_X1 port map( B1 => n393, B2 => n453, C1 => n392, C2 => n454, A 
                           => n455, ZN => O_4_port);
   U84 : AOI22_X1 port map( A1 => A_ns(3), A2 => n397, B1 => A_s(3), B2 => n398
                           , ZN => n455);
   U85 : INV_X1 port map( A => A_s(2), ZN => n454);
   U86 : INV_X1 port map( A => A_ns(2), ZN => n453);
   U87 : OAI221_X1 port map( B1 => n393, B2 => n456, C1 => n392, C2 => n457, A 
                           => n458, ZN => O_49_port);
   U88 : AOI22_X1 port map( A1 => A_ns(48), A2 => n397, B1 => A_s(48), B2 => 
                           n398, ZN => n458);
   U89 : INV_X1 port map( A => A_s(47), ZN => n457);
   U90 : INV_X1 port map( A => A_ns(47), ZN => n456);
   U91 : OAI221_X1 port map( B1 => n393, B2 => n459, C1 => n392, C2 => n460, A 
                           => n461, ZN => O_48_port);
   U92 : AOI22_X1 port map( A1 => A_ns(47), A2 => n397, B1 => A_s(47), B2 => 
                           n398, ZN => n461);
   U93 : INV_X1 port map( A => A_s(46), ZN => n460);
   U94 : INV_X1 port map( A => A_ns(46), ZN => n459);
   U95 : OAI221_X1 port map( B1 => n393, B2 => n462, C1 => n392, C2 => n463, A 
                           => n464, ZN => O_47_port);
   U96 : AOI22_X1 port map( A1 => A_ns(46), A2 => n397, B1 => A_s(46), B2 => 
                           n398, ZN => n464);
   U97 : INV_X1 port map( A => A_s(45), ZN => n463);
   U98 : INV_X1 port map( A => A_ns(45), ZN => n462);
   U99 : OAI221_X1 port map( B1 => n393, B2 => n465, C1 => n392, C2 => n466, A 
                           => n467, ZN => O_46_port);
   U100 : AOI22_X1 port map( A1 => A_ns(45), A2 => n397, B1 => A_s(45), B2 => 
                           n398, ZN => n467);
   U101 : INV_X1 port map( A => A_s(44), ZN => n466);
   U102 : INV_X1 port map( A => A_ns(44), ZN => n465);
   U103 : OAI221_X1 port map( B1 => n393, B2 => n468, C1 => n392, C2 => n469, A
                           => n470, ZN => O_45_port);
   U104 : AOI22_X1 port map( A1 => A_ns(44), A2 => n397, B1 => A_s(44), B2 => 
                           n398, ZN => n470);
   U105 : INV_X1 port map( A => A_s(43), ZN => n469);
   U106 : INV_X1 port map( A => A_ns(43), ZN => n468);
   U107 : OAI221_X1 port map( B1 => n393, B2 => n471, C1 => n392, C2 => n472, A
                           => n473, ZN => O_44_port);
   U108 : AOI22_X1 port map( A1 => A_ns(43), A2 => n397, B1 => A_s(43), B2 => 
                           n398, ZN => n473);
   U109 : INV_X1 port map( A => A_s(42), ZN => n472);
   U110 : INV_X1 port map( A => A_ns(42), ZN => n471);
   U111 : OAI221_X1 port map( B1 => n393, B2 => n474, C1 => n392, C2 => n475, A
                           => n476, ZN => O_43_port);
   U112 : AOI22_X1 port map( A1 => A_ns(42), A2 => n397, B1 => A_s(42), B2 => 
                           n398, ZN => n476);
   U113 : INV_X1 port map( A => A_s(41), ZN => n475);
   U114 : INV_X1 port map( A => A_ns(41), ZN => n474);
   U115 : OAI221_X1 port map( B1 => n393, B2 => n477, C1 => n392, C2 => n478, A
                           => n479, ZN => O_42_port);
   U116 : AOI22_X1 port map( A1 => A_ns(41), A2 => n397, B1 => A_s(41), B2 => 
                           n398, ZN => n479);
   U117 : INV_X1 port map( A => A_s(40), ZN => n478);
   U118 : INV_X1 port map( A => A_ns(40), ZN => n477);
   U119 : OAI221_X1 port map( B1 => n393, B2 => n480, C1 => n392, C2 => n481, A
                           => n482, ZN => O_41_port);
   U120 : AOI22_X1 port map( A1 => A_ns(40), A2 => n397, B1 => A_s(40), B2 => 
                           n398, ZN => n482);
   U121 : INV_X1 port map( A => A_s(39), ZN => n481);
   U122 : INV_X1 port map( A => A_ns(39), ZN => n480);
   U123 : OAI221_X1 port map( B1 => n393, B2 => n483, C1 => n392, C2 => n484, A
                           => n485, ZN => O_40_port);
   U124 : AOI22_X1 port map( A1 => A_ns(39), A2 => n397, B1 => A_s(39), B2 => 
                           n398, ZN => n485);
   U125 : INV_X1 port map( A => A_s(38), ZN => n484);
   U126 : INV_X1 port map( A => A_ns(38), ZN => n483);
   U127 : OAI221_X1 port map( B1 => n393, B2 => n486, C1 => n392, C2 => n487, A
                           => n488, ZN => O_3_port);
   U128 : AOI22_X1 port map( A1 => A_ns(2), A2 => n397, B1 => A_s(2), B2 => 
                           n398, ZN => n488);
   U129 : INV_X1 port map( A => A_s(1), ZN => n487);
   U130 : INV_X1 port map( A => A_ns(1), ZN => n486);
   U131 : OAI221_X1 port map( B1 => n393, B2 => n489, C1 => n392, C2 => n490, A
                           => n491, ZN => O_39_port);
   U132 : AOI22_X1 port map( A1 => A_ns(38), A2 => n397, B1 => A_s(38), B2 => 
                           n398, ZN => n491);
   U133 : INV_X1 port map( A => A_s(37), ZN => n490);
   U134 : INV_X1 port map( A => A_ns(37), ZN => n489);
   U135 : OAI221_X1 port map( B1 => n393, B2 => n492, C1 => n392, C2 => n493, A
                           => n494, ZN => O_38_port);
   U136 : AOI22_X1 port map( A1 => A_ns(37), A2 => n397, B1 => A_s(37), B2 => 
                           n398, ZN => n494);
   U137 : INV_X1 port map( A => A_s(36), ZN => n493);
   U138 : INV_X1 port map( A => A_ns(36), ZN => n492);
   U139 : OAI221_X1 port map( B1 => n393, B2 => n495, C1 => n392, C2 => n496, A
                           => n497, ZN => O_37_port);
   U140 : AOI22_X1 port map( A1 => A_ns(36), A2 => n397, B1 => A_s(36), B2 => 
                           n398, ZN => n497);
   U141 : INV_X1 port map( A => A_s(35), ZN => n496);
   U142 : INV_X1 port map( A => A_ns(35), ZN => n495);
   U143 : OAI221_X1 port map( B1 => n393, B2 => n498, C1 => n392, C2 => n499, A
                           => n500, ZN => O_36_port);
   U144 : AOI22_X1 port map( A1 => A_ns(35), A2 => n397, B1 => A_s(35), B2 => 
                           n398, ZN => n500);
   U145 : INV_X1 port map( A => A_s(34), ZN => n499);
   U146 : INV_X1 port map( A => A_ns(34), ZN => n498);
   U147 : OAI221_X1 port map( B1 => n393, B2 => n501, C1 => n392, C2 => n502, A
                           => n503, ZN => O_35_port);
   U148 : AOI22_X1 port map( A1 => A_ns(34), A2 => n397, B1 => A_s(34), B2 => 
                           n398, ZN => n503);
   U149 : INV_X1 port map( A => A_s(33), ZN => n502);
   U150 : INV_X1 port map( A => A_ns(33), ZN => n501);
   U151 : OAI221_X1 port map( B1 => n393, B2 => n504, C1 => n392, C2 => n505, A
                           => n506, ZN => O_34_port);
   U152 : AOI22_X1 port map( A1 => A_ns(33), A2 => n397, B1 => A_s(33), B2 => 
                           n398, ZN => n506);
   U153 : INV_X1 port map( A => A_s(32), ZN => n505);
   U154 : INV_X1 port map( A => A_ns(32), ZN => n504);
   U155 : OAI221_X1 port map( B1 => n393, B2 => n507, C1 => n392, C2 => n508, A
                           => n509, ZN => O_33_port);
   U156 : AOI22_X1 port map( A1 => A_ns(32), A2 => n397, B1 => A_s(32), B2 => 
                           n398, ZN => n509);
   U157 : INV_X1 port map( A => A_s(31), ZN => n508);
   U158 : INV_X1 port map( A => A_ns(31), ZN => n507);
   U159 : OAI221_X1 port map( B1 => n393, B2 => n510, C1 => n392, C2 => n511, A
                           => n512, ZN => O_32_port);
   U160 : AOI22_X1 port map( A1 => A_ns(31), A2 => n397, B1 => A_s(31), B2 => 
                           n398, ZN => n512);
   U161 : INV_X1 port map( A => A_s(30), ZN => n511);
   U162 : INV_X1 port map( A => A_ns(30), ZN => n510);
   U163 : OAI221_X1 port map( B1 => n393, B2 => n513, C1 => n392, C2 => n514, A
                           => n515, ZN => O_31_port);
   U164 : AOI22_X1 port map( A1 => A_ns(30), A2 => n397, B1 => A_s(30), B2 => 
                           n398, ZN => n515);
   U165 : INV_X1 port map( A => A_s(29), ZN => n514);
   U166 : INV_X1 port map( A => A_ns(29), ZN => n513);
   U167 : OAI221_X1 port map( B1 => n393, B2 => n516, C1 => n392, C2 => n517, A
                           => n518, ZN => O_30_port);
   U168 : AOI22_X1 port map( A1 => A_ns(29), A2 => n397, B1 => A_s(29), B2 => 
                           n398, ZN => n518);
   U169 : INV_X1 port map( A => A_s(28), ZN => n517);
   U170 : INV_X1 port map( A => A_ns(28), ZN => n516);
   U171 : OAI221_X1 port map( B1 => n393, B2 => n519, C1 => n392, C2 => n520, A
                           => n521, ZN => O_2_port);
   U172 : AOI22_X1 port map( A1 => A_ns(1), A2 => n397, B1 => A_s(1), B2 => 
                           n398, ZN => n521);
   U173 : OAI221_X1 port map( B1 => n393, B2 => n522, C1 => n392, C2 => n523, A
                           => n524, ZN => O_29_port);
   U174 : AOI22_X1 port map( A1 => A_ns(28), A2 => n397, B1 => A_s(28), B2 => 
                           n398, ZN => n524);
   U175 : INV_X1 port map( A => A_s(27), ZN => n523);
   U176 : INV_X1 port map( A => A_ns(27), ZN => n522);
   U177 : OAI221_X1 port map( B1 => n393, B2 => n525, C1 => n392, C2 => n526, A
                           => n527, ZN => O_28_port);
   U178 : AOI22_X1 port map( A1 => A_ns(27), A2 => n397, B1 => A_s(27), B2 => 
                           n398, ZN => n527);
   U179 : INV_X1 port map( A => A_s(26), ZN => n526);
   U180 : INV_X1 port map( A => A_ns(26), ZN => n525);
   U181 : OAI221_X1 port map( B1 => n393, B2 => n528, C1 => n392, C2 => n529, A
                           => n530, ZN => O_27_port);
   U182 : AOI22_X1 port map( A1 => A_ns(26), A2 => n397, B1 => A_s(26), B2 => 
                           n398, ZN => n530);
   U183 : INV_X1 port map( A => A_s(25), ZN => n529);
   U184 : INV_X1 port map( A => A_ns(25), ZN => n528);
   U185 : OAI221_X1 port map( B1 => n393, B2 => n531, C1 => n392, C2 => n532, A
                           => n533, ZN => O_26_port);
   U186 : AOI22_X1 port map( A1 => A_ns(25), A2 => n397, B1 => A_s(25), B2 => 
                           n398, ZN => n533);
   U187 : INV_X1 port map( A => A_s(24), ZN => n532);
   U188 : INV_X1 port map( A => A_ns(24), ZN => n531);
   U189 : OAI221_X1 port map( B1 => n393, B2 => n534, C1 => n392, C2 => n535, A
                           => n536, ZN => O_25_port);
   U190 : AOI22_X1 port map( A1 => A_ns(24), A2 => n397, B1 => A_s(24), B2 => 
                           n398, ZN => n536);
   U191 : INV_X1 port map( A => A_s(23), ZN => n535);
   U192 : INV_X1 port map( A => A_ns(23), ZN => n534);
   U193 : OAI221_X1 port map( B1 => n393, B2 => n537, C1 => n392, C2 => n538, A
                           => n539, ZN => O_24_port);
   U194 : AOI22_X1 port map( A1 => A_ns(23), A2 => n397, B1 => A_s(23), B2 => 
                           n398, ZN => n539);
   U195 : INV_X1 port map( A => A_s(22), ZN => n538);
   U196 : INV_X1 port map( A => A_ns(22), ZN => n537);
   U197 : OAI221_X1 port map( B1 => n393, B2 => n540, C1 => n392, C2 => n541, A
                           => n542, ZN => O_23_port);
   U198 : AOI22_X1 port map( A1 => A_ns(22), A2 => n397, B1 => A_s(22), B2 => 
                           n398, ZN => n542);
   U199 : INV_X1 port map( A => A_s(21), ZN => n541);
   U200 : INV_X1 port map( A => A_ns(21), ZN => n540);
   U201 : OAI221_X1 port map( B1 => n393, B2 => n543, C1 => n392, C2 => n544, A
                           => n545, ZN => O_22_port);
   U202 : AOI22_X1 port map( A1 => A_ns(21), A2 => n397, B1 => A_s(21), B2 => 
                           n398, ZN => n545);
   U203 : INV_X1 port map( A => A_s(20), ZN => n544);
   U204 : INV_X1 port map( A => A_ns(20), ZN => n543);
   U205 : OAI221_X1 port map( B1 => n393, B2 => n546, C1 => n392, C2 => n547, A
                           => n548, ZN => O_21_port);
   U206 : AOI22_X1 port map( A1 => A_ns(20), A2 => n397, B1 => A_s(20), B2 => 
                           n398, ZN => n548);
   U207 : INV_X1 port map( A => A_s(19), ZN => n547);
   U208 : INV_X1 port map( A => A_ns(19), ZN => n546);
   U209 : OAI221_X1 port map( B1 => n393, B2 => n549, C1 => n392, C2 => n550, A
                           => n551, ZN => O_20_port);
   U210 : AOI22_X1 port map( A1 => A_ns(19), A2 => n397, B1 => A_s(19), B2 => 
                           n398, ZN => n551);
   U211 : INV_X1 port map( A => A_s(18), ZN => n550);
   U212 : INV_X1 port map( A => A_ns(18), ZN => n549);
   U213 : OAI22_X1 port map( A1 => n552, A2 => n520, B1 => n553, B2 => n519, ZN
                           => O_1_port);
   U214 : INV_X1 port map( A => A_ns(0), ZN => n519);
   U215 : INV_X1 port map( A => A_s(0), ZN => n520);
   U216 : OAI221_X1 port map( B1 => n393, B2 => n554, C1 => n392, C2 => n555, A
                           => n556, ZN => O_19_port);
   U217 : AOI22_X1 port map( A1 => A_ns(18), A2 => n397, B1 => A_s(18), B2 => 
                           n398, ZN => n556);
   U218 : INV_X1 port map( A => A_s(17), ZN => n555);
   U219 : INV_X1 port map( A => A_ns(17), ZN => n554);
   U220 : OAI221_X1 port map( B1 => n393, B2 => n557, C1 => n392, C2 => n558, A
                           => n559, ZN => O_18_port);
   U221 : AOI22_X1 port map( A1 => A_ns(17), A2 => n397, B1 => A_s(17), B2 => 
                           n398, ZN => n559);
   U222 : INV_X1 port map( A => A_s(16), ZN => n558);
   U223 : INV_X1 port map( A => A_ns(16), ZN => n557);
   U224 : OAI221_X1 port map( B1 => n393, B2 => n560, C1 => n392, C2 => n561, A
                           => n562, ZN => O_17_port);
   U225 : AOI22_X1 port map( A1 => A_ns(16), A2 => n397, B1 => A_s(16), B2 => 
                           n398, ZN => n562);
   U226 : INV_X1 port map( A => A_s(15), ZN => n561);
   U227 : INV_X1 port map( A => A_ns(15), ZN => n560);
   U228 : OAI221_X1 port map( B1 => n393, B2 => n563, C1 => n392, C2 => n564, A
                           => n565, ZN => O_16_port);
   U229 : AOI22_X1 port map( A1 => A_ns(15), A2 => n397, B1 => A_s(15), B2 => 
                           n398, ZN => n565);
   U230 : INV_X1 port map( A => A_s(14), ZN => n564);
   U231 : INV_X1 port map( A => A_ns(14), ZN => n563);
   U232 : OAI221_X1 port map( B1 => n393, B2 => n566, C1 => n392, C2 => n567, A
                           => n568, ZN => O_15_port);
   U233 : AOI22_X1 port map( A1 => A_ns(14), A2 => n397, B1 => A_s(14), B2 => 
                           n398, ZN => n568);
   U234 : INV_X1 port map( A => A_s(13), ZN => n567);
   U235 : INV_X1 port map( A => A_ns(13), ZN => n566);
   U236 : OAI221_X1 port map( B1 => n393, B2 => n569, C1 => n392, C2 => n570, A
                           => n571, ZN => O_14_port);
   U237 : AOI22_X1 port map( A1 => A_ns(13), A2 => n397, B1 => A_s(13), B2 => 
                           n398, ZN => n571);
   U238 : INV_X1 port map( A => A_s(12), ZN => n570);
   U239 : INV_X1 port map( A => A_ns(12), ZN => n569);
   U240 : OAI221_X1 port map( B1 => n393, B2 => n572, C1 => n392, C2 => n573, A
                           => n574, ZN => O_13_port);
   U241 : AOI22_X1 port map( A1 => A_ns(12), A2 => n397, B1 => A_s(12), B2 => 
                           n398, ZN => n574);
   U242 : INV_X1 port map( A => A_s(11), ZN => n573);
   U243 : INV_X1 port map( A => A_ns(11), ZN => n572);
   U244 : OAI221_X1 port map( B1 => n393, B2 => n575, C1 => n392, C2 => n576, A
                           => n577, ZN => O_12_port);
   U245 : AOI22_X1 port map( A1 => A_ns(11), A2 => n397, B1 => A_s(11), B2 => 
                           n398, ZN => n577);
   U246 : INV_X1 port map( A => A_s(10), ZN => n576);
   U247 : INV_X1 port map( A => A_ns(10), ZN => n575);
   U248 : OAI221_X1 port map( B1 => n393, B2 => n578, C1 => n392, C2 => n579, A
                           => n580, ZN => O_11_port);
   U249 : AOI22_X1 port map( A1 => A_ns(10), A2 => n397, B1 => A_s(10), B2 => 
                           n398, ZN => n580);
   U250 : INV_X1 port map( A => A_s(9), ZN => n579);
   U251 : INV_X1 port map( A => A_ns(9), ZN => n578);
   U252 : OAI221_X1 port map( B1 => n581, B2 => n393, C1 => n582, C2 => n392, A
                           => n583, ZN => O_10_port);
   U253 : AOI22_X1 port map( A1 => A_ns(9), A2 => n397, B1 => A_s(9), B2 => 
                           n398, ZN => n583);
   U254 : NAND2_X1 port map( A1 => n584, A2 => n552, ZN => n553);
   U255 : NAND2_X1 port map( A1 => n584, A2 => n585, ZN => n552);
   U256 : XOR2_X1 port map( A => B(21), B => B(22), Z => n584);
   U257 : INV_X1 port map( A => A_s(8), ZN => n582);
   U258 : INV_X1 port map( A => B(23), ZN => n585);
   U259 : INV_X1 port map( A => A_ns(8), ZN => n581);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity BOOTHENC_NBIT64_i20 is

   port( A, A_n, A_ns, A_s, B : in std_logic_vector (63 downto 0);  O, A_so, 
         A_nso : out std_logic_vector (63 downto 0));

end BOOTHENC_NBIT64_i20;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT64_i20 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, O_63_port, O_62_port, O_61_port, O_60_port, O_59_port,
      O_58_port, O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, 
      O_52_port, O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, 
      O_46_port, O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, 
      O_40_port, O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, 
      O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, 
      O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, 
      O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, 
      O_16_port, O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, 
      O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, 
      O_3_port, O_2_port, O_1_port, n391, n392, n393, n394, n395, n396, n397, 
      n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, 
      n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, 
      n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, 
      n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, 
      n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, 
      n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, 
      n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, 
      n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, 
      n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, 
      n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, 
      n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, 
      n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, 
      n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, 
      n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, 
      n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, 
      n578, n579, n580, n581, n582, n583, n584, n585 : std_logic;

begin
   O <= ( O_63_port, O_62_port, O_61_port, O_60_port, O_59_port, O_58_port, 
      O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, O_52_port, 
      O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, O_46_port, 
      O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, O_40_port, 
      O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, 
      O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, 
      O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, 
      O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, O_16_port, 
      O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, O_10_port, 
      O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, O_3_port, 
      O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(61), A_s(60), A_s(59), A_s(58), A_s(57), A_s(56), A_s(55), 
      A_s(54), A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), 
      A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), 
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   A_nso <= ( A_s(61), A_s(60), A_s(59), A_s(58), A_s(57), A_s(56), A_s(55), 
      A_s(54), A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), 
      A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), 
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : AND3_X1 port map( A1 => B(20), A2 => n585, A3 => B(19), ZN => n391);
   U3 : INV_X4 port map( A => n391, ZN => n392);
   U4 : INV_X4 port map( A => n552, ZN => n398);
   U5 : OR3_X4 port map( A1 => B(19), A2 => B(20), A3 => n585, ZN => n393);
   U6 : INV_X4 port map( A => n553, ZN => n397);
   U7 : OAI221_X1 port map( B1 => n393, B2 => n394, C1 => n392, C2 => n395, A 
                           => n396, ZN => O_9_port);
   U8 : AOI22_X1 port map( A1 => A_ns(8), A2 => n397, B1 => A_s(8), B2 => n398,
                           ZN => n396);
   U9 : INV_X1 port map( A => A_s(7), ZN => n395);
   U10 : INV_X1 port map( A => A_ns(7), ZN => n394);
   U11 : OAI221_X1 port map( B1 => n393, B2 => n399, C1 => n392, C2 => n400, A 
                           => n401, ZN => O_8_port);
   U12 : AOI22_X1 port map( A1 => A_ns(7), A2 => n397, B1 => A_s(7), B2 => n398
                           , ZN => n401);
   U13 : INV_X1 port map( A => A_s(6), ZN => n400);
   U14 : INV_X1 port map( A => A_ns(6), ZN => n399);
   U15 : OAI221_X1 port map( B1 => n393, B2 => n402, C1 => n392, C2 => n403, A 
                           => n404, ZN => O_7_port);
   U16 : AOI22_X1 port map( A1 => A_ns(6), A2 => n397, B1 => A_s(6), B2 => n398
                           , ZN => n404);
   U17 : INV_X1 port map( A => A_s(5), ZN => n403);
   U18 : INV_X1 port map( A => A_ns(5), ZN => n402);
   U19 : OAI221_X1 port map( B1 => n393, B2 => n405, C1 => n392, C2 => n406, A 
                           => n407, ZN => O_6_port);
   U20 : AOI22_X1 port map( A1 => A_ns(5), A2 => n397, B1 => A_s(5), B2 => n398
                           , ZN => n407);
   U21 : INV_X1 port map( A => A_s(4), ZN => n406);
   U22 : INV_X1 port map( A => A_ns(4), ZN => n405);
   U23 : OAI221_X1 port map( B1 => n393, B2 => n408, C1 => n392, C2 => n409, A 
                           => n410, ZN => O_63_port);
   U24 : AOI22_X1 port map( A1 => A_ns(62), A2 => n397, B1 => A_s(62), B2 => 
                           n398, ZN => n410);
   U25 : INV_X1 port map( A => A_s(61), ZN => n409);
   U26 : INV_X1 port map( A => A_ns(61), ZN => n408);
   U27 : OAI221_X1 port map( B1 => n393, B2 => n411, C1 => n392, C2 => n412, A 
                           => n413, ZN => O_62_port);
   U28 : AOI22_X1 port map( A1 => A_ns(61), A2 => n397, B1 => A_s(61), B2 => 
                           n398, ZN => n413);
   U29 : INV_X1 port map( A => A_s(60), ZN => n412);
   U30 : INV_X1 port map( A => A_ns(60), ZN => n411);
   U31 : OAI221_X1 port map( B1 => n393, B2 => n414, C1 => n392, C2 => n415, A 
                           => n416, ZN => O_61_port);
   U32 : AOI22_X1 port map( A1 => A_ns(60), A2 => n397, B1 => A_s(60), B2 => 
                           n398, ZN => n416);
   U33 : INV_X1 port map( A => A_s(59), ZN => n415);
   U34 : INV_X1 port map( A => A_ns(59), ZN => n414);
   U35 : OAI221_X1 port map( B1 => n393, B2 => n417, C1 => n392, C2 => n418, A 
                           => n419, ZN => O_60_port);
   U36 : AOI22_X1 port map( A1 => A_ns(59), A2 => n397, B1 => A_s(59), B2 => 
                           n398, ZN => n419);
   U37 : INV_X1 port map( A => A_s(58), ZN => n418);
   U38 : INV_X1 port map( A => A_ns(58), ZN => n417);
   U39 : OAI221_X1 port map( B1 => n393, B2 => n420, C1 => n392, C2 => n421, A 
                           => n422, ZN => O_5_port);
   U40 : AOI22_X1 port map( A1 => A_ns(4), A2 => n397, B1 => A_s(4), B2 => n398
                           , ZN => n422);
   U41 : INV_X1 port map( A => A_s(3), ZN => n421);
   U42 : INV_X1 port map( A => A_ns(3), ZN => n420);
   U43 : OAI221_X1 port map( B1 => n393, B2 => n423, C1 => n392, C2 => n424, A 
                           => n425, ZN => O_59_port);
   U44 : AOI22_X1 port map( A1 => A_ns(58), A2 => n397, B1 => A_s(58), B2 => 
                           n398, ZN => n425);
   U45 : INV_X1 port map( A => A_s(57), ZN => n424);
   U46 : INV_X1 port map( A => A_ns(57), ZN => n423);
   U47 : OAI221_X1 port map( B1 => n393, B2 => n426, C1 => n392, C2 => n427, A 
                           => n428, ZN => O_58_port);
   U48 : AOI22_X1 port map( A1 => A_ns(57), A2 => n397, B1 => A_s(57), B2 => 
                           n398, ZN => n428);
   U49 : INV_X1 port map( A => A_s(56), ZN => n427);
   U50 : INV_X1 port map( A => A_ns(56), ZN => n426);
   U51 : OAI221_X1 port map( B1 => n393, B2 => n429, C1 => n392, C2 => n430, A 
                           => n431, ZN => O_57_port);
   U52 : AOI22_X1 port map( A1 => A_ns(56), A2 => n397, B1 => A_s(56), B2 => 
                           n398, ZN => n431);
   U53 : INV_X1 port map( A => A_s(55), ZN => n430);
   U54 : INV_X1 port map( A => A_ns(55), ZN => n429);
   U55 : OAI221_X1 port map( B1 => n393, B2 => n432, C1 => n392, C2 => n433, A 
                           => n434, ZN => O_56_port);
   U56 : AOI22_X1 port map( A1 => A_ns(55), A2 => n397, B1 => A_s(55), B2 => 
                           n398, ZN => n434);
   U57 : INV_X1 port map( A => A_s(54), ZN => n433);
   U58 : INV_X1 port map( A => A_ns(54), ZN => n432);
   U59 : OAI221_X1 port map( B1 => n393, B2 => n435, C1 => n392, C2 => n436, A 
                           => n437, ZN => O_55_port);
   U60 : AOI22_X1 port map( A1 => A_ns(54), A2 => n397, B1 => A_s(54), B2 => 
                           n398, ZN => n437);
   U61 : INV_X1 port map( A => A_s(53), ZN => n436);
   U62 : INV_X1 port map( A => A_ns(53), ZN => n435);
   U63 : OAI221_X1 port map( B1 => n393, B2 => n438, C1 => n392, C2 => n439, A 
                           => n440, ZN => O_54_port);
   U64 : AOI22_X1 port map( A1 => A_ns(53), A2 => n397, B1 => A_s(53), B2 => 
                           n398, ZN => n440);
   U65 : INV_X1 port map( A => A_s(52), ZN => n439);
   U66 : INV_X1 port map( A => A_ns(52), ZN => n438);
   U67 : OAI221_X1 port map( B1 => n393, B2 => n441, C1 => n392, C2 => n442, A 
                           => n443, ZN => O_53_port);
   U68 : AOI22_X1 port map( A1 => A_ns(52), A2 => n397, B1 => A_s(52), B2 => 
                           n398, ZN => n443);
   U69 : INV_X1 port map( A => A_s(51), ZN => n442);
   U70 : INV_X1 port map( A => A_ns(51), ZN => n441);
   U71 : OAI221_X1 port map( B1 => n393, B2 => n444, C1 => n392, C2 => n445, A 
                           => n446, ZN => O_52_port);
   U72 : AOI22_X1 port map( A1 => A_ns(51), A2 => n397, B1 => A_s(51), B2 => 
                           n398, ZN => n446);
   U73 : INV_X1 port map( A => A_s(50), ZN => n445);
   U74 : INV_X1 port map( A => A_ns(50), ZN => n444);
   U75 : OAI221_X1 port map( B1 => n393, B2 => n447, C1 => n392, C2 => n448, A 
                           => n449, ZN => O_51_port);
   U76 : AOI22_X1 port map( A1 => A_ns(50), A2 => n397, B1 => A_s(50), B2 => 
                           n398, ZN => n449);
   U77 : INV_X1 port map( A => A_s(49), ZN => n448);
   U78 : INV_X1 port map( A => A_ns(49), ZN => n447);
   U79 : OAI221_X1 port map( B1 => n393, B2 => n450, C1 => n392, C2 => n451, A 
                           => n452, ZN => O_50_port);
   U80 : AOI22_X1 port map( A1 => A_ns(49), A2 => n397, B1 => A_s(49), B2 => 
                           n398, ZN => n452);
   U81 : INV_X1 port map( A => A_s(48), ZN => n451);
   U82 : INV_X1 port map( A => A_ns(48), ZN => n450);
   U83 : OAI221_X1 port map( B1 => n393, B2 => n453, C1 => n392, C2 => n454, A 
                           => n455, ZN => O_4_port);
   U84 : AOI22_X1 port map( A1 => A_ns(3), A2 => n397, B1 => A_s(3), B2 => n398
                           , ZN => n455);
   U85 : INV_X1 port map( A => A_s(2), ZN => n454);
   U86 : INV_X1 port map( A => A_ns(2), ZN => n453);
   U87 : OAI221_X1 port map( B1 => n393, B2 => n456, C1 => n392, C2 => n457, A 
                           => n458, ZN => O_49_port);
   U88 : AOI22_X1 port map( A1 => A_ns(48), A2 => n397, B1 => A_s(48), B2 => 
                           n398, ZN => n458);
   U89 : INV_X1 port map( A => A_s(47), ZN => n457);
   U90 : INV_X1 port map( A => A_ns(47), ZN => n456);
   U91 : OAI221_X1 port map( B1 => n393, B2 => n459, C1 => n392, C2 => n460, A 
                           => n461, ZN => O_48_port);
   U92 : AOI22_X1 port map( A1 => A_ns(47), A2 => n397, B1 => A_s(47), B2 => 
                           n398, ZN => n461);
   U93 : INV_X1 port map( A => A_s(46), ZN => n460);
   U94 : INV_X1 port map( A => A_ns(46), ZN => n459);
   U95 : OAI221_X1 port map( B1 => n393, B2 => n462, C1 => n392, C2 => n463, A 
                           => n464, ZN => O_47_port);
   U96 : AOI22_X1 port map( A1 => A_ns(46), A2 => n397, B1 => A_s(46), B2 => 
                           n398, ZN => n464);
   U97 : INV_X1 port map( A => A_s(45), ZN => n463);
   U98 : INV_X1 port map( A => A_ns(45), ZN => n462);
   U99 : OAI221_X1 port map( B1 => n393, B2 => n465, C1 => n392, C2 => n466, A 
                           => n467, ZN => O_46_port);
   U100 : AOI22_X1 port map( A1 => A_ns(45), A2 => n397, B1 => A_s(45), B2 => 
                           n398, ZN => n467);
   U101 : INV_X1 port map( A => A_s(44), ZN => n466);
   U102 : INV_X1 port map( A => A_ns(44), ZN => n465);
   U103 : OAI221_X1 port map( B1 => n393, B2 => n468, C1 => n392, C2 => n469, A
                           => n470, ZN => O_45_port);
   U104 : AOI22_X1 port map( A1 => A_ns(44), A2 => n397, B1 => A_s(44), B2 => 
                           n398, ZN => n470);
   U105 : INV_X1 port map( A => A_s(43), ZN => n469);
   U106 : INV_X1 port map( A => A_ns(43), ZN => n468);
   U107 : OAI221_X1 port map( B1 => n393, B2 => n471, C1 => n392, C2 => n472, A
                           => n473, ZN => O_44_port);
   U108 : AOI22_X1 port map( A1 => A_ns(43), A2 => n397, B1 => A_s(43), B2 => 
                           n398, ZN => n473);
   U109 : INV_X1 port map( A => A_s(42), ZN => n472);
   U110 : INV_X1 port map( A => A_ns(42), ZN => n471);
   U111 : OAI221_X1 port map( B1 => n393, B2 => n474, C1 => n392, C2 => n475, A
                           => n476, ZN => O_43_port);
   U112 : AOI22_X1 port map( A1 => A_ns(42), A2 => n397, B1 => A_s(42), B2 => 
                           n398, ZN => n476);
   U113 : INV_X1 port map( A => A_s(41), ZN => n475);
   U114 : INV_X1 port map( A => A_ns(41), ZN => n474);
   U115 : OAI221_X1 port map( B1 => n393, B2 => n477, C1 => n392, C2 => n478, A
                           => n479, ZN => O_42_port);
   U116 : AOI22_X1 port map( A1 => A_ns(41), A2 => n397, B1 => A_s(41), B2 => 
                           n398, ZN => n479);
   U117 : INV_X1 port map( A => A_s(40), ZN => n478);
   U118 : INV_X1 port map( A => A_ns(40), ZN => n477);
   U119 : OAI221_X1 port map( B1 => n393, B2 => n480, C1 => n392, C2 => n481, A
                           => n482, ZN => O_41_port);
   U120 : AOI22_X1 port map( A1 => A_ns(40), A2 => n397, B1 => A_s(40), B2 => 
                           n398, ZN => n482);
   U121 : INV_X1 port map( A => A_s(39), ZN => n481);
   U122 : INV_X1 port map( A => A_ns(39), ZN => n480);
   U123 : OAI221_X1 port map( B1 => n393, B2 => n483, C1 => n392, C2 => n484, A
                           => n485, ZN => O_40_port);
   U124 : AOI22_X1 port map( A1 => A_ns(39), A2 => n397, B1 => A_s(39), B2 => 
                           n398, ZN => n485);
   U125 : INV_X1 port map( A => A_s(38), ZN => n484);
   U126 : INV_X1 port map( A => A_ns(38), ZN => n483);
   U127 : OAI221_X1 port map( B1 => n393, B2 => n486, C1 => n392, C2 => n487, A
                           => n488, ZN => O_3_port);
   U128 : AOI22_X1 port map( A1 => A_ns(2), A2 => n397, B1 => A_s(2), B2 => 
                           n398, ZN => n488);
   U129 : INV_X1 port map( A => A_s(1), ZN => n487);
   U130 : INV_X1 port map( A => A_ns(1), ZN => n486);
   U131 : OAI221_X1 port map( B1 => n393, B2 => n489, C1 => n392, C2 => n490, A
                           => n491, ZN => O_39_port);
   U132 : AOI22_X1 port map( A1 => A_ns(38), A2 => n397, B1 => A_s(38), B2 => 
                           n398, ZN => n491);
   U133 : INV_X1 port map( A => A_s(37), ZN => n490);
   U134 : INV_X1 port map( A => A_ns(37), ZN => n489);
   U135 : OAI221_X1 port map( B1 => n393, B2 => n492, C1 => n392, C2 => n493, A
                           => n494, ZN => O_38_port);
   U136 : AOI22_X1 port map( A1 => A_ns(37), A2 => n397, B1 => A_s(37), B2 => 
                           n398, ZN => n494);
   U137 : INV_X1 port map( A => A_s(36), ZN => n493);
   U138 : INV_X1 port map( A => A_ns(36), ZN => n492);
   U139 : OAI221_X1 port map( B1 => n393, B2 => n495, C1 => n392, C2 => n496, A
                           => n497, ZN => O_37_port);
   U140 : AOI22_X1 port map( A1 => A_ns(36), A2 => n397, B1 => A_s(36), B2 => 
                           n398, ZN => n497);
   U141 : INV_X1 port map( A => A_s(35), ZN => n496);
   U142 : INV_X1 port map( A => A_ns(35), ZN => n495);
   U143 : OAI221_X1 port map( B1 => n393, B2 => n498, C1 => n392, C2 => n499, A
                           => n500, ZN => O_36_port);
   U144 : AOI22_X1 port map( A1 => A_ns(35), A2 => n397, B1 => A_s(35), B2 => 
                           n398, ZN => n500);
   U145 : INV_X1 port map( A => A_s(34), ZN => n499);
   U146 : INV_X1 port map( A => A_ns(34), ZN => n498);
   U147 : OAI221_X1 port map( B1 => n393, B2 => n501, C1 => n392, C2 => n502, A
                           => n503, ZN => O_35_port);
   U148 : AOI22_X1 port map( A1 => A_ns(34), A2 => n397, B1 => A_s(34), B2 => 
                           n398, ZN => n503);
   U149 : INV_X1 port map( A => A_s(33), ZN => n502);
   U150 : INV_X1 port map( A => A_ns(33), ZN => n501);
   U151 : OAI221_X1 port map( B1 => n393, B2 => n504, C1 => n392, C2 => n505, A
                           => n506, ZN => O_34_port);
   U152 : AOI22_X1 port map( A1 => A_ns(33), A2 => n397, B1 => A_s(33), B2 => 
                           n398, ZN => n506);
   U153 : INV_X1 port map( A => A_s(32), ZN => n505);
   U154 : INV_X1 port map( A => A_ns(32), ZN => n504);
   U155 : OAI221_X1 port map( B1 => n393, B2 => n507, C1 => n392, C2 => n508, A
                           => n509, ZN => O_33_port);
   U156 : AOI22_X1 port map( A1 => A_ns(32), A2 => n397, B1 => A_s(32), B2 => 
                           n398, ZN => n509);
   U157 : INV_X1 port map( A => A_s(31), ZN => n508);
   U158 : INV_X1 port map( A => A_ns(31), ZN => n507);
   U159 : OAI221_X1 port map( B1 => n393, B2 => n510, C1 => n392, C2 => n511, A
                           => n512, ZN => O_32_port);
   U160 : AOI22_X1 port map( A1 => A_ns(31), A2 => n397, B1 => A_s(31), B2 => 
                           n398, ZN => n512);
   U161 : INV_X1 port map( A => A_s(30), ZN => n511);
   U162 : INV_X1 port map( A => A_ns(30), ZN => n510);
   U163 : OAI221_X1 port map( B1 => n393, B2 => n513, C1 => n392, C2 => n514, A
                           => n515, ZN => O_31_port);
   U164 : AOI22_X1 port map( A1 => A_ns(30), A2 => n397, B1 => A_s(30), B2 => 
                           n398, ZN => n515);
   U165 : INV_X1 port map( A => A_s(29), ZN => n514);
   U166 : INV_X1 port map( A => A_ns(29), ZN => n513);
   U167 : OAI221_X1 port map( B1 => n393, B2 => n516, C1 => n392, C2 => n517, A
                           => n518, ZN => O_30_port);
   U168 : AOI22_X1 port map( A1 => A_ns(29), A2 => n397, B1 => A_s(29), B2 => 
                           n398, ZN => n518);
   U169 : INV_X1 port map( A => A_s(28), ZN => n517);
   U170 : INV_X1 port map( A => A_ns(28), ZN => n516);
   U171 : OAI221_X1 port map( B1 => n393, B2 => n519, C1 => n392, C2 => n520, A
                           => n521, ZN => O_2_port);
   U172 : AOI22_X1 port map( A1 => A_ns(1), A2 => n397, B1 => A_s(1), B2 => 
                           n398, ZN => n521);
   U173 : OAI221_X1 port map( B1 => n393, B2 => n522, C1 => n392, C2 => n523, A
                           => n524, ZN => O_29_port);
   U174 : AOI22_X1 port map( A1 => A_ns(28), A2 => n397, B1 => A_s(28), B2 => 
                           n398, ZN => n524);
   U175 : INV_X1 port map( A => A_s(27), ZN => n523);
   U176 : INV_X1 port map( A => A_ns(27), ZN => n522);
   U177 : OAI221_X1 port map( B1 => n393, B2 => n525, C1 => n392, C2 => n526, A
                           => n527, ZN => O_28_port);
   U178 : AOI22_X1 port map( A1 => A_ns(27), A2 => n397, B1 => A_s(27), B2 => 
                           n398, ZN => n527);
   U179 : INV_X1 port map( A => A_s(26), ZN => n526);
   U180 : INV_X1 port map( A => A_ns(26), ZN => n525);
   U181 : OAI221_X1 port map( B1 => n393, B2 => n528, C1 => n392, C2 => n529, A
                           => n530, ZN => O_27_port);
   U182 : AOI22_X1 port map( A1 => A_ns(26), A2 => n397, B1 => A_s(26), B2 => 
                           n398, ZN => n530);
   U183 : INV_X1 port map( A => A_s(25), ZN => n529);
   U184 : INV_X1 port map( A => A_ns(25), ZN => n528);
   U185 : OAI221_X1 port map( B1 => n393, B2 => n531, C1 => n392, C2 => n532, A
                           => n533, ZN => O_26_port);
   U186 : AOI22_X1 port map( A1 => A_ns(25), A2 => n397, B1 => A_s(25), B2 => 
                           n398, ZN => n533);
   U187 : INV_X1 port map( A => A_s(24), ZN => n532);
   U188 : INV_X1 port map( A => A_ns(24), ZN => n531);
   U189 : OAI221_X1 port map( B1 => n393, B2 => n534, C1 => n392, C2 => n535, A
                           => n536, ZN => O_25_port);
   U190 : AOI22_X1 port map( A1 => A_ns(24), A2 => n397, B1 => A_s(24), B2 => 
                           n398, ZN => n536);
   U191 : INV_X1 port map( A => A_s(23), ZN => n535);
   U192 : INV_X1 port map( A => A_ns(23), ZN => n534);
   U193 : OAI221_X1 port map( B1 => n393, B2 => n537, C1 => n392, C2 => n538, A
                           => n539, ZN => O_24_port);
   U194 : AOI22_X1 port map( A1 => A_ns(23), A2 => n397, B1 => A_s(23), B2 => 
                           n398, ZN => n539);
   U195 : INV_X1 port map( A => A_s(22), ZN => n538);
   U196 : INV_X1 port map( A => A_ns(22), ZN => n537);
   U197 : OAI221_X1 port map( B1 => n393, B2 => n540, C1 => n392, C2 => n541, A
                           => n542, ZN => O_23_port);
   U198 : AOI22_X1 port map( A1 => A_ns(22), A2 => n397, B1 => A_s(22), B2 => 
                           n398, ZN => n542);
   U199 : INV_X1 port map( A => A_s(21), ZN => n541);
   U200 : INV_X1 port map( A => A_ns(21), ZN => n540);
   U201 : OAI221_X1 port map( B1 => n393, B2 => n543, C1 => n392, C2 => n544, A
                           => n545, ZN => O_22_port);
   U202 : AOI22_X1 port map( A1 => A_ns(21), A2 => n397, B1 => A_s(21), B2 => 
                           n398, ZN => n545);
   U203 : INV_X1 port map( A => A_s(20), ZN => n544);
   U204 : INV_X1 port map( A => A_ns(20), ZN => n543);
   U205 : OAI221_X1 port map( B1 => n393, B2 => n546, C1 => n392, C2 => n547, A
                           => n548, ZN => O_21_port);
   U206 : AOI22_X1 port map( A1 => A_ns(20), A2 => n397, B1 => A_s(20), B2 => 
                           n398, ZN => n548);
   U207 : INV_X1 port map( A => A_s(19), ZN => n547);
   U208 : INV_X1 port map( A => A_ns(19), ZN => n546);
   U209 : OAI221_X1 port map( B1 => n393, B2 => n549, C1 => n392, C2 => n550, A
                           => n551, ZN => O_20_port);
   U210 : AOI22_X1 port map( A1 => A_ns(19), A2 => n397, B1 => A_s(19), B2 => 
                           n398, ZN => n551);
   U211 : INV_X1 port map( A => A_s(18), ZN => n550);
   U212 : INV_X1 port map( A => A_ns(18), ZN => n549);
   U213 : OAI22_X1 port map( A1 => n552, A2 => n520, B1 => n553, B2 => n519, ZN
                           => O_1_port);
   U214 : INV_X1 port map( A => A_ns(0), ZN => n519);
   U215 : INV_X1 port map( A => A_s(0), ZN => n520);
   U216 : OAI221_X1 port map( B1 => n393, B2 => n554, C1 => n392, C2 => n555, A
                           => n556, ZN => O_19_port);
   U217 : AOI22_X1 port map( A1 => A_ns(18), A2 => n397, B1 => A_s(18), B2 => 
                           n398, ZN => n556);
   U218 : INV_X1 port map( A => A_s(17), ZN => n555);
   U219 : INV_X1 port map( A => A_ns(17), ZN => n554);
   U220 : OAI221_X1 port map( B1 => n393, B2 => n557, C1 => n392, C2 => n558, A
                           => n559, ZN => O_18_port);
   U221 : AOI22_X1 port map( A1 => A_ns(17), A2 => n397, B1 => A_s(17), B2 => 
                           n398, ZN => n559);
   U222 : INV_X1 port map( A => A_s(16), ZN => n558);
   U223 : INV_X1 port map( A => A_ns(16), ZN => n557);
   U224 : OAI221_X1 port map( B1 => n393, B2 => n560, C1 => n392, C2 => n561, A
                           => n562, ZN => O_17_port);
   U225 : AOI22_X1 port map( A1 => A_ns(16), A2 => n397, B1 => A_s(16), B2 => 
                           n398, ZN => n562);
   U226 : INV_X1 port map( A => A_s(15), ZN => n561);
   U227 : INV_X1 port map( A => A_ns(15), ZN => n560);
   U228 : OAI221_X1 port map( B1 => n393, B2 => n563, C1 => n392, C2 => n564, A
                           => n565, ZN => O_16_port);
   U229 : AOI22_X1 port map( A1 => A_ns(15), A2 => n397, B1 => A_s(15), B2 => 
                           n398, ZN => n565);
   U230 : INV_X1 port map( A => A_s(14), ZN => n564);
   U231 : INV_X1 port map( A => A_ns(14), ZN => n563);
   U232 : OAI221_X1 port map( B1 => n393, B2 => n566, C1 => n392, C2 => n567, A
                           => n568, ZN => O_15_port);
   U233 : AOI22_X1 port map( A1 => A_ns(14), A2 => n397, B1 => A_s(14), B2 => 
                           n398, ZN => n568);
   U234 : INV_X1 port map( A => A_s(13), ZN => n567);
   U235 : INV_X1 port map( A => A_ns(13), ZN => n566);
   U236 : OAI221_X1 port map( B1 => n393, B2 => n569, C1 => n392, C2 => n570, A
                           => n571, ZN => O_14_port);
   U237 : AOI22_X1 port map( A1 => A_ns(13), A2 => n397, B1 => A_s(13), B2 => 
                           n398, ZN => n571);
   U238 : INV_X1 port map( A => A_s(12), ZN => n570);
   U239 : INV_X1 port map( A => A_ns(12), ZN => n569);
   U240 : OAI221_X1 port map( B1 => n393, B2 => n572, C1 => n392, C2 => n573, A
                           => n574, ZN => O_13_port);
   U241 : AOI22_X1 port map( A1 => A_ns(12), A2 => n397, B1 => A_s(12), B2 => 
                           n398, ZN => n574);
   U242 : INV_X1 port map( A => A_s(11), ZN => n573);
   U243 : INV_X1 port map( A => A_ns(11), ZN => n572);
   U244 : OAI221_X1 port map( B1 => n393, B2 => n575, C1 => n392, C2 => n576, A
                           => n577, ZN => O_12_port);
   U245 : AOI22_X1 port map( A1 => A_ns(11), A2 => n397, B1 => A_s(11), B2 => 
                           n398, ZN => n577);
   U246 : INV_X1 port map( A => A_s(10), ZN => n576);
   U247 : INV_X1 port map( A => A_ns(10), ZN => n575);
   U248 : OAI221_X1 port map( B1 => n393, B2 => n578, C1 => n392, C2 => n579, A
                           => n580, ZN => O_11_port);
   U249 : AOI22_X1 port map( A1 => A_ns(10), A2 => n397, B1 => A_s(10), B2 => 
                           n398, ZN => n580);
   U250 : INV_X1 port map( A => A_s(9), ZN => n579);
   U251 : INV_X1 port map( A => A_ns(9), ZN => n578);
   U252 : OAI221_X1 port map( B1 => n581, B2 => n393, C1 => n582, C2 => n392, A
                           => n583, ZN => O_10_port);
   U253 : AOI22_X1 port map( A1 => A_ns(9), A2 => n397, B1 => A_s(9), B2 => 
                           n398, ZN => n583);
   U254 : NAND2_X1 port map( A1 => n584, A2 => n552, ZN => n553);
   U255 : NAND2_X1 port map( A1 => n584, A2 => n585, ZN => n552);
   U256 : XOR2_X1 port map( A => B(19), B => B(20), Z => n584);
   U257 : INV_X1 port map( A => A_s(8), ZN => n582);
   U258 : INV_X1 port map( A => B(21), ZN => n585);
   U259 : INV_X1 port map( A => A_ns(8), ZN => n581);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity BOOTHENC_NBIT64_i18 is

   port( A, A_n, A_ns, A_s, B : in std_logic_vector (63 downto 0);  O, A_so, 
         A_nso : out std_logic_vector (63 downto 0));

end BOOTHENC_NBIT64_i18;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT64_i18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, O_63_port, O_62_port, O_61_port, O_60_port, O_59_port,
      O_58_port, O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, 
      O_52_port, O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, 
      O_46_port, O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, 
      O_40_port, O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, 
      O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, 
      O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, 
      O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, 
      O_16_port, O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, 
      O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, 
      O_3_port, O_2_port, O_1_port, n391, n392, n393, n394, n395, n396, n397, 
      n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, 
      n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, 
      n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, 
      n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, 
      n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, 
      n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, 
      n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, 
      n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, 
      n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, 
      n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, 
      n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, 
      n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, 
      n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, 
      n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, 
      n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, 
      n578, n579, n580, n581, n582, n583, n584, n585 : std_logic;

begin
   O <= ( O_63_port, O_62_port, O_61_port, O_60_port, O_59_port, O_58_port, 
      O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, O_52_port, 
      O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, O_46_port, 
      O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, O_40_port, 
      O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, 
      O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, 
      O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, 
      O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, O_16_port, 
      O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, O_10_port, 
      O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, O_3_port, 
      O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(61), A_s(60), A_s(59), A_s(58), A_s(57), A_s(56), A_s(55), 
      A_s(54), A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), 
      A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), 
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   A_nso <= ( A_s(61), A_s(60), A_s(59), A_s(58), A_s(57), A_s(56), A_s(55), 
      A_s(54), A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), 
      A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), 
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : AND3_X1 port map( A1 => B(18), A2 => n585, A3 => B(17), ZN => n391);
   U3 : INV_X4 port map( A => n391, ZN => n392);
   U4 : INV_X4 port map( A => n552, ZN => n398);
   U5 : OR3_X4 port map( A1 => B(17), A2 => B(18), A3 => n585, ZN => n393);
   U6 : INV_X4 port map( A => n553, ZN => n397);
   U7 : OAI221_X1 port map( B1 => n393, B2 => n394, C1 => n392, C2 => n395, A 
                           => n396, ZN => O_9_port);
   U8 : AOI22_X1 port map( A1 => A_ns(8), A2 => n397, B1 => A_s(8), B2 => n398,
                           ZN => n396);
   U9 : INV_X1 port map( A => A_s(7), ZN => n395);
   U10 : INV_X1 port map( A => A_ns(7), ZN => n394);
   U11 : OAI221_X1 port map( B1 => n393, B2 => n399, C1 => n392, C2 => n400, A 
                           => n401, ZN => O_8_port);
   U12 : AOI22_X1 port map( A1 => A_ns(7), A2 => n397, B1 => A_s(7), B2 => n398
                           , ZN => n401);
   U13 : INV_X1 port map( A => A_s(6), ZN => n400);
   U14 : INV_X1 port map( A => A_ns(6), ZN => n399);
   U15 : OAI221_X1 port map( B1 => n393, B2 => n402, C1 => n392, C2 => n403, A 
                           => n404, ZN => O_7_port);
   U16 : AOI22_X1 port map( A1 => A_ns(6), A2 => n397, B1 => A_s(6), B2 => n398
                           , ZN => n404);
   U17 : INV_X1 port map( A => A_s(5), ZN => n403);
   U18 : INV_X1 port map( A => A_ns(5), ZN => n402);
   U19 : OAI221_X1 port map( B1 => n393, B2 => n405, C1 => n392, C2 => n406, A 
                           => n407, ZN => O_6_port);
   U20 : AOI22_X1 port map( A1 => A_ns(5), A2 => n397, B1 => A_s(5), B2 => n398
                           , ZN => n407);
   U21 : INV_X1 port map( A => A_s(4), ZN => n406);
   U22 : INV_X1 port map( A => A_ns(4), ZN => n405);
   U23 : OAI221_X1 port map( B1 => n393, B2 => n408, C1 => n392, C2 => n409, A 
                           => n410, ZN => O_63_port);
   U24 : AOI22_X1 port map( A1 => A_ns(62), A2 => n397, B1 => A_s(62), B2 => 
                           n398, ZN => n410);
   U25 : INV_X1 port map( A => A_s(61), ZN => n409);
   U26 : INV_X1 port map( A => A_ns(61), ZN => n408);
   U27 : OAI221_X1 port map( B1 => n393, B2 => n411, C1 => n392, C2 => n412, A 
                           => n413, ZN => O_62_port);
   U28 : AOI22_X1 port map( A1 => A_ns(61), A2 => n397, B1 => A_s(61), B2 => 
                           n398, ZN => n413);
   U29 : INV_X1 port map( A => A_s(60), ZN => n412);
   U30 : INV_X1 port map( A => A_ns(60), ZN => n411);
   U31 : OAI221_X1 port map( B1 => n393, B2 => n414, C1 => n392, C2 => n415, A 
                           => n416, ZN => O_61_port);
   U32 : AOI22_X1 port map( A1 => A_ns(60), A2 => n397, B1 => A_s(60), B2 => 
                           n398, ZN => n416);
   U33 : INV_X1 port map( A => A_s(59), ZN => n415);
   U34 : INV_X1 port map( A => A_ns(59), ZN => n414);
   U35 : OAI221_X1 port map( B1 => n393, B2 => n417, C1 => n392, C2 => n418, A 
                           => n419, ZN => O_60_port);
   U36 : AOI22_X1 port map( A1 => A_ns(59), A2 => n397, B1 => A_s(59), B2 => 
                           n398, ZN => n419);
   U37 : INV_X1 port map( A => A_s(58), ZN => n418);
   U38 : INV_X1 port map( A => A_ns(58), ZN => n417);
   U39 : OAI221_X1 port map( B1 => n393, B2 => n420, C1 => n392, C2 => n421, A 
                           => n422, ZN => O_5_port);
   U40 : AOI22_X1 port map( A1 => A_ns(4), A2 => n397, B1 => A_s(4), B2 => n398
                           , ZN => n422);
   U41 : INV_X1 port map( A => A_s(3), ZN => n421);
   U42 : INV_X1 port map( A => A_ns(3), ZN => n420);
   U43 : OAI221_X1 port map( B1 => n393, B2 => n423, C1 => n392, C2 => n424, A 
                           => n425, ZN => O_59_port);
   U44 : AOI22_X1 port map( A1 => A_ns(58), A2 => n397, B1 => A_s(58), B2 => 
                           n398, ZN => n425);
   U45 : INV_X1 port map( A => A_s(57), ZN => n424);
   U46 : INV_X1 port map( A => A_ns(57), ZN => n423);
   U47 : OAI221_X1 port map( B1 => n393, B2 => n426, C1 => n392, C2 => n427, A 
                           => n428, ZN => O_58_port);
   U48 : AOI22_X1 port map( A1 => A_ns(57), A2 => n397, B1 => A_s(57), B2 => 
                           n398, ZN => n428);
   U49 : INV_X1 port map( A => A_s(56), ZN => n427);
   U50 : INV_X1 port map( A => A_ns(56), ZN => n426);
   U51 : OAI221_X1 port map( B1 => n393, B2 => n429, C1 => n392, C2 => n430, A 
                           => n431, ZN => O_57_port);
   U52 : AOI22_X1 port map( A1 => A_ns(56), A2 => n397, B1 => A_s(56), B2 => 
                           n398, ZN => n431);
   U53 : INV_X1 port map( A => A_s(55), ZN => n430);
   U54 : INV_X1 port map( A => A_ns(55), ZN => n429);
   U55 : OAI221_X1 port map( B1 => n393, B2 => n432, C1 => n392, C2 => n433, A 
                           => n434, ZN => O_56_port);
   U56 : AOI22_X1 port map( A1 => A_ns(55), A2 => n397, B1 => A_s(55), B2 => 
                           n398, ZN => n434);
   U57 : INV_X1 port map( A => A_s(54), ZN => n433);
   U58 : INV_X1 port map( A => A_ns(54), ZN => n432);
   U59 : OAI221_X1 port map( B1 => n393, B2 => n435, C1 => n392, C2 => n436, A 
                           => n437, ZN => O_55_port);
   U60 : AOI22_X1 port map( A1 => A_ns(54), A2 => n397, B1 => A_s(54), B2 => 
                           n398, ZN => n437);
   U61 : INV_X1 port map( A => A_s(53), ZN => n436);
   U62 : INV_X1 port map( A => A_ns(53), ZN => n435);
   U63 : OAI221_X1 port map( B1 => n393, B2 => n438, C1 => n392, C2 => n439, A 
                           => n440, ZN => O_54_port);
   U64 : AOI22_X1 port map( A1 => A_ns(53), A2 => n397, B1 => A_s(53), B2 => 
                           n398, ZN => n440);
   U65 : INV_X1 port map( A => A_s(52), ZN => n439);
   U66 : INV_X1 port map( A => A_ns(52), ZN => n438);
   U67 : OAI221_X1 port map( B1 => n393, B2 => n441, C1 => n392, C2 => n442, A 
                           => n443, ZN => O_53_port);
   U68 : AOI22_X1 port map( A1 => A_ns(52), A2 => n397, B1 => A_s(52), B2 => 
                           n398, ZN => n443);
   U69 : INV_X1 port map( A => A_s(51), ZN => n442);
   U70 : INV_X1 port map( A => A_ns(51), ZN => n441);
   U71 : OAI221_X1 port map( B1 => n393, B2 => n444, C1 => n392, C2 => n445, A 
                           => n446, ZN => O_52_port);
   U72 : AOI22_X1 port map( A1 => A_ns(51), A2 => n397, B1 => A_s(51), B2 => 
                           n398, ZN => n446);
   U73 : INV_X1 port map( A => A_s(50), ZN => n445);
   U74 : INV_X1 port map( A => A_ns(50), ZN => n444);
   U75 : OAI221_X1 port map( B1 => n393, B2 => n447, C1 => n392, C2 => n448, A 
                           => n449, ZN => O_51_port);
   U76 : AOI22_X1 port map( A1 => A_ns(50), A2 => n397, B1 => A_s(50), B2 => 
                           n398, ZN => n449);
   U77 : INV_X1 port map( A => A_s(49), ZN => n448);
   U78 : INV_X1 port map( A => A_ns(49), ZN => n447);
   U79 : OAI221_X1 port map( B1 => n393, B2 => n450, C1 => n392, C2 => n451, A 
                           => n452, ZN => O_50_port);
   U80 : AOI22_X1 port map( A1 => A_ns(49), A2 => n397, B1 => A_s(49), B2 => 
                           n398, ZN => n452);
   U81 : INV_X1 port map( A => A_s(48), ZN => n451);
   U82 : INV_X1 port map( A => A_ns(48), ZN => n450);
   U83 : OAI221_X1 port map( B1 => n393, B2 => n453, C1 => n392, C2 => n454, A 
                           => n455, ZN => O_4_port);
   U84 : AOI22_X1 port map( A1 => A_ns(3), A2 => n397, B1 => A_s(3), B2 => n398
                           , ZN => n455);
   U85 : INV_X1 port map( A => A_s(2), ZN => n454);
   U86 : INV_X1 port map( A => A_ns(2), ZN => n453);
   U87 : OAI221_X1 port map( B1 => n393, B2 => n456, C1 => n392, C2 => n457, A 
                           => n458, ZN => O_49_port);
   U88 : AOI22_X1 port map( A1 => A_ns(48), A2 => n397, B1 => A_s(48), B2 => 
                           n398, ZN => n458);
   U89 : INV_X1 port map( A => A_s(47), ZN => n457);
   U90 : INV_X1 port map( A => A_ns(47), ZN => n456);
   U91 : OAI221_X1 port map( B1 => n393, B2 => n459, C1 => n392, C2 => n460, A 
                           => n461, ZN => O_48_port);
   U92 : AOI22_X1 port map( A1 => A_ns(47), A2 => n397, B1 => A_s(47), B2 => 
                           n398, ZN => n461);
   U93 : INV_X1 port map( A => A_s(46), ZN => n460);
   U94 : INV_X1 port map( A => A_ns(46), ZN => n459);
   U95 : OAI221_X1 port map( B1 => n393, B2 => n462, C1 => n392, C2 => n463, A 
                           => n464, ZN => O_47_port);
   U96 : AOI22_X1 port map( A1 => A_ns(46), A2 => n397, B1 => A_s(46), B2 => 
                           n398, ZN => n464);
   U97 : INV_X1 port map( A => A_s(45), ZN => n463);
   U98 : INV_X1 port map( A => A_ns(45), ZN => n462);
   U99 : OAI221_X1 port map( B1 => n393, B2 => n465, C1 => n392, C2 => n466, A 
                           => n467, ZN => O_46_port);
   U100 : AOI22_X1 port map( A1 => A_ns(45), A2 => n397, B1 => A_s(45), B2 => 
                           n398, ZN => n467);
   U101 : INV_X1 port map( A => A_s(44), ZN => n466);
   U102 : INV_X1 port map( A => A_ns(44), ZN => n465);
   U103 : OAI221_X1 port map( B1 => n393, B2 => n468, C1 => n392, C2 => n469, A
                           => n470, ZN => O_45_port);
   U104 : AOI22_X1 port map( A1 => A_ns(44), A2 => n397, B1 => A_s(44), B2 => 
                           n398, ZN => n470);
   U105 : INV_X1 port map( A => A_s(43), ZN => n469);
   U106 : INV_X1 port map( A => A_ns(43), ZN => n468);
   U107 : OAI221_X1 port map( B1 => n393, B2 => n471, C1 => n392, C2 => n472, A
                           => n473, ZN => O_44_port);
   U108 : AOI22_X1 port map( A1 => A_ns(43), A2 => n397, B1 => A_s(43), B2 => 
                           n398, ZN => n473);
   U109 : INV_X1 port map( A => A_s(42), ZN => n472);
   U110 : INV_X1 port map( A => A_ns(42), ZN => n471);
   U111 : OAI221_X1 port map( B1 => n393, B2 => n474, C1 => n392, C2 => n475, A
                           => n476, ZN => O_43_port);
   U112 : AOI22_X1 port map( A1 => A_ns(42), A2 => n397, B1 => A_s(42), B2 => 
                           n398, ZN => n476);
   U113 : INV_X1 port map( A => A_s(41), ZN => n475);
   U114 : INV_X1 port map( A => A_ns(41), ZN => n474);
   U115 : OAI221_X1 port map( B1 => n393, B2 => n477, C1 => n392, C2 => n478, A
                           => n479, ZN => O_42_port);
   U116 : AOI22_X1 port map( A1 => A_ns(41), A2 => n397, B1 => A_s(41), B2 => 
                           n398, ZN => n479);
   U117 : INV_X1 port map( A => A_s(40), ZN => n478);
   U118 : INV_X1 port map( A => A_ns(40), ZN => n477);
   U119 : OAI221_X1 port map( B1 => n393, B2 => n480, C1 => n392, C2 => n481, A
                           => n482, ZN => O_41_port);
   U120 : AOI22_X1 port map( A1 => A_ns(40), A2 => n397, B1 => A_s(40), B2 => 
                           n398, ZN => n482);
   U121 : INV_X1 port map( A => A_s(39), ZN => n481);
   U122 : INV_X1 port map( A => A_ns(39), ZN => n480);
   U123 : OAI221_X1 port map( B1 => n393, B2 => n483, C1 => n392, C2 => n484, A
                           => n485, ZN => O_40_port);
   U124 : AOI22_X1 port map( A1 => A_ns(39), A2 => n397, B1 => A_s(39), B2 => 
                           n398, ZN => n485);
   U125 : INV_X1 port map( A => A_s(38), ZN => n484);
   U126 : INV_X1 port map( A => A_ns(38), ZN => n483);
   U127 : OAI221_X1 port map( B1 => n393, B2 => n486, C1 => n392, C2 => n487, A
                           => n488, ZN => O_3_port);
   U128 : AOI22_X1 port map( A1 => A_ns(2), A2 => n397, B1 => A_s(2), B2 => 
                           n398, ZN => n488);
   U129 : INV_X1 port map( A => A_s(1), ZN => n487);
   U130 : INV_X1 port map( A => A_ns(1), ZN => n486);
   U131 : OAI221_X1 port map( B1 => n393, B2 => n489, C1 => n392, C2 => n490, A
                           => n491, ZN => O_39_port);
   U132 : AOI22_X1 port map( A1 => A_ns(38), A2 => n397, B1 => A_s(38), B2 => 
                           n398, ZN => n491);
   U133 : INV_X1 port map( A => A_s(37), ZN => n490);
   U134 : INV_X1 port map( A => A_ns(37), ZN => n489);
   U135 : OAI221_X1 port map( B1 => n393, B2 => n492, C1 => n392, C2 => n493, A
                           => n494, ZN => O_38_port);
   U136 : AOI22_X1 port map( A1 => A_ns(37), A2 => n397, B1 => A_s(37), B2 => 
                           n398, ZN => n494);
   U137 : INV_X1 port map( A => A_s(36), ZN => n493);
   U138 : INV_X1 port map( A => A_ns(36), ZN => n492);
   U139 : OAI221_X1 port map( B1 => n393, B2 => n495, C1 => n392, C2 => n496, A
                           => n497, ZN => O_37_port);
   U140 : AOI22_X1 port map( A1 => A_ns(36), A2 => n397, B1 => A_s(36), B2 => 
                           n398, ZN => n497);
   U141 : INV_X1 port map( A => A_s(35), ZN => n496);
   U142 : INV_X1 port map( A => A_ns(35), ZN => n495);
   U143 : OAI221_X1 port map( B1 => n393, B2 => n498, C1 => n392, C2 => n499, A
                           => n500, ZN => O_36_port);
   U144 : AOI22_X1 port map( A1 => A_ns(35), A2 => n397, B1 => A_s(35), B2 => 
                           n398, ZN => n500);
   U145 : INV_X1 port map( A => A_s(34), ZN => n499);
   U146 : INV_X1 port map( A => A_ns(34), ZN => n498);
   U147 : OAI221_X1 port map( B1 => n393, B2 => n501, C1 => n392, C2 => n502, A
                           => n503, ZN => O_35_port);
   U148 : AOI22_X1 port map( A1 => A_ns(34), A2 => n397, B1 => A_s(34), B2 => 
                           n398, ZN => n503);
   U149 : INV_X1 port map( A => A_s(33), ZN => n502);
   U150 : INV_X1 port map( A => A_ns(33), ZN => n501);
   U151 : OAI221_X1 port map( B1 => n393, B2 => n504, C1 => n392, C2 => n505, A
                           => n506, ZN => O_34_port);
   U152 : AOI22_X1 port map( A1 => A_ns(33), A2 => n397, B1 => A_s(33), B2 => 
                           n398, ZN => n506);
   U153 : INV_X1 port map( A => A_s(32), ZN => n505);
   U154 : INV_X1 port map( A => A_ns(32), ZN => n504);
   U155 : OAI221_X1 port map( B1 => n393, B2 => n507, C1 => n392, C2 => n508, A
                           => n509, ZN => O_33_port);
   U156 : AOI22_X1 port map( A1 => A_ns(32), A2 => n397, B1 => A_s(32), B2 => 
                           n398, ZN => n509);
   U157 : INV_X1 port map( A => A_s(31), ZN => n508);
   U158 : INV_X1 port map( A => A_ns(31), ZN => n507);
   U159 : OAI221_X1 port map( B1 => n393, B2 => n510, C1 => n392, C2 => n511, A
                           => n512, ZN => O_32_port);
   U160 : AOI22_X1 port map( A1 => A_ns(31), A2 => n397, B1 => A_s(31), B2 => 
                           n398, ZN => n512);
   U161 : INV_X1 port map( A => A_s(30), ZN => n511);
   U162 : INV_X1 port map( A => A_ns(30), ZN => n510);
   U163 : OAI221_X1 port map( B1 => n393, B2 => n513, C1 => n392, C2 => n514, A
                           => n515, ZN => O_31_port);
   U164 : AOI22_X1 port map( A1 => A_ns(30), A2 => n397, B1 => A_s(30), B2 => 
                           n398, ZN => n515);
   U165 : INV_X1 port map( A => A_s(29), ZN => n514);
   U166 : INV_X1 port map( A => A_ns(29), ZN => n513);
   U167 : OAI221_X1 port map( B1 => n393, B2 => n516, C1 => n392, C2 => n517, A
                           => n518, ZN => O_30_port);
   U168 : AOI22_X1 port map( A1 => A_ns(29), A2 => n397, B1 => A_s(29), B2 => 
                           n398, ZN => n518);
   U169 : INV_X1 port map( A => A_s(28), ZN => n517);
   U170 : INV_X1 port map( A => A_ns(28), ZN => n516);
   U171 : OAI221_X1 port map( B1 => n393, B2 => n519, C1 => n392, C2 => n520, A
                           => n521, ZN => O_2_port);
   U172 : AOI22_X1 port map( A1 => A_ns(1), A2 => n397, B1 => A_s(1), B2 => 
                           n398, ZN => n521);
   U173 : OAI221_X1 port map( B1 => n393, B2 => n522, C1 => n392, C2 => n523, A
                           => n524, ZN => O_29_port);
   U174 : AOI22_X1 port map( A1 => A_ns(28), A2 => n397, B1 => A_s(28), B2 => 
                           n398, ZN => n524);
   U175 : INV_X1 port map( A => A_s(27), ZN => n523);
   U176 : INV_X1 port map( A => A_ns(27), ZN => n522);
   U177 : OAI221_X1 port map( B1 => n393, B2 => n525, C1 => n392, C2 => n526, A
                           => n527, ZN => O_28_port);
   U178 : AOI22_X1 port map( A1 => A_ns(27), A2 => n397, B1 => A_s(27), B2 => 
                           n398, ZN => n527);
   U179 : INV_X1 port map( A => A_s(26), ZN => n526);
   U180 : INV_X1 port map( A => A_ns(26), ZN => n525);
   U181 : OAI221_X1 port map( B1 => n393, B2 => n528, C1 => n392, C2 => n529, A
                           => n530, ZN => O_27_port);
   U182 : AOI22_X1 port map( A1 => A_ns(26), A2 => n397, B1 => A_s(26), B2 => 
                           n398, ZN => n530);
   U183 : INV_X1 port map( A => A_s(25), ZN => n529);
   U184 : INV_X1 port map( A => A_ns(25), ZN => n528);
   U185 : OAI221_X1 port map( B1 => n393, B2 => n531, C1 => n392, C2 => n532, A
                           => n533, ZN => O_26_port);
   U186 : AOI22_X1 port map( A1 => A_ns(25), A2 => n397, B1 => A_s(25), B2 => 
                           n398, ZN => n533);
   U187 : INV_X1 port map( A => A_s(24), ZN => n532);
   U188 : INV_X1 port map( A => A_ns(24), ZN => n531);
   U189 : OAI221_X1 port map( B1 => n393, B2 => n534, C1 => n392, C2 => n535, A
                           => n536, ZN => O_25_port);
   U190 : AOI22_X1 port map( A1 => A_ns(24), A2 => n397, B1 => A_s(24), B2 => 
                           n398, ZN => n536);
   U191 : INV_X1 port map( A => A_s(23), ZN => n535);
   U192 : INV_X1 port map( A => A_ns(23), ZN => n534);
   U193 : OAI221_X1 port map( B1 => n393, B2 => n537, C1 => n392, C2 => n538, A
                           => n539, ZN => O_24_port);
   U194 : AOI22_X1 port map( A1 => A_ns(23), A2 => n397, B1 => A_s(23), B2 => 
                           n398, ZN => n539);
   U195 : INV_X1 port map( A => A_s(22), ZN => n538);
   U196 : INV_X1 port map( A => A_ns(22), ZN => n537);
   U197 : OAI221_X1 port map( B1 => n393, B2 => n540, C1 => n392, C2 => n541, A
                           => n542, ZN => O_23_port);
   U198 : AOI22_X1 port map( A1 => A_ns(22), A2 => n397, B1 => A_s(22), B2 => 
                           n398, ZN => n542);
   U199 : INV_X1 port map( A => A_s(21), ZN => n541);
   U200 : INV_X1 port map( A => A_ns(21), ZN => n540);
   U201 : OAI221_X1 port map( B1 => n393, B2 => n543, C1 => n392, C2 => n544, A
                           => n545, ZN => O_22_port);
   U202 : AOI22_X1 port map( A1 => A_ns(21), A2 => n397, B1 => A_s(21), B2 => 
                           n398, ZN => n545);
   U203 : INV_X1 port map( A => A_s(20), ZN => n544);
   U204 : INV_X1 port map( A => A_ns(20), ZN => n543);
   U205 : OAI221_X1 port map( B1 => n393, B2 => n546, C1 => n392, C2 => n547, A
                           => n548, ZN => O_21_port);
   U206 : AOI22_X1 port map( A1 => A_ns(20), A2 => n397, B1 => A_s(20), B2 => 
                           n398, ZN => n548);
   U207 : INV_X1 port map( A => A_s(19), ZN => n547);
   U208 : INV_X1 port map( A => A_ns(19), ZN => n546);
   U209 : OAI221_X1 port map( B1 => n393, B2 => n549, C1 => n392, C2 => n550, A
                           => n551, ZN => O_20_port);
   U210 : AOI22_X1 port map( A1 => A_ns(19), A2 => n397, B1 => A_s(19), B2 => 
                           n398, ZN => n551);
   U211 : INV_X1 port map( A => A_s(18), ZN => n550);
   U212 : INV_X1 port map( A => A_ns(18), ZN => n549);
   U213 : OAI22_X1 port map( A1 => n552, A2 => n520, B1 => n553, B2 => n519, ZN
                           => O_1_port);
   U214 : INV_X1 port map( A => A_ns(0), ZN => n519);
   U215 : INV_X1 port map( A => A_s(0), ZN => n520);
   U216 : OAI221_X1 port map( B1 => n393, B2 => n554, C1 => n392, C2 => n555, A
                           => n556, ZN => O_19_port);
   U217 : AOI22_X1 port map( A1 => A_ns(18), A2 => n397, B1 => A_s(18), B2 => 
                           n398, ZN => n556);
   U218 : INV_X1 port map( A => A_s(17), ZN => n555);
   U219 : INV_X1 port map( A => A_ns(17), ZN => n554);
   U220 : OAI221_X1 port map( B1 => n393, B2 => n557, C1 => n392, C2 => n558, A
                           => n559, ZN => O_18_port);
   U221 : AOI22_X1 port map( A1 => A_ns(17), A2 => n397, B1 => A_s(17), B2 => 
                           n398, ZN => n559);
   U222 : INV_X1 port map( A => A_s(16), ZN => n558);
   U223 : INV_X1 port map( A => A_ns(16), ZN => n557);
   U224 : OAI221_X1 port map( B1 => n393, B2 => n560, C1 => n392, C2 => n561, A
                           => n562, ZN => O_17_port);
   U225 : AOI22_X1 port map( A1 => A_ns(16), A2 => n397, B1 => A_s(16), B2 => 
                           n398, ZN => n562);
   U226 : INV_X1 port map( A => A_s(15), ZN => n561);
   U227 : INV_X1 port map( A => A_ns(15), ZN => n560);
   U228 : OAI221_X1 port map( B1 => n393, B2 => n563, C1 => n392, C2 => n564, A
                           => n565, ZN => O_16_port);
   U229 : AOI22_X1 port map( A1 => A_ns(15), A2 => n397, B1 => A_s(15), B2 => 
                           n398, ZN => n565);
   U230 : INV_X1 port map( A => A_s(14), ZN => n564);
   U231 : INV_X1 port map( A => A_ns(14), ZN => n563);
   U232 : OAI221_X1 port map( B1 => n393, B2 => n566, C1 => n392, C2 => n567, A
                           => n568, ZN => O_15_port);
   U233 : AOI22_X1 port map( A1 => A_ns(14), A2 => n397, B1 => A_s(14), B2 => 
                           n398, ZN => n568);
   U234 : INV_X1 port map( A => A_s(13), ZN => n567);
   U235 : INV_X1 port map( A => A_ns(13), ZN => n566);
   U236 : OAI221_X1 port map( B1 => n393, B2 => n569, C1 => n392, C2 => n570, A
                           => n571, ZN => O_14_port);
   U237 : AOI22_X1 port map( A1 => A_ns(13), A2 => n397, B1 => A_s(13), B2 => 
                           n398, ZN => n571);
   U238 : INV_X1 port map( A => A_s(12), ZN => n570);
   U239 : INV_X1 port map( A => A_ns(12), ZN => n569);
   U240 : OAI221_X1 port map( B1 => n393, B2 => n572, C1 => n392, C2 => n573, A
                           => n574, ZN => O_13_port);
   U241 : AOI22_X1 port map( A1 => A_ns(12), A2 => n397, B1 => A_s(12), B2 => 
                           n398, ZN => n574);
   U242 : INV_X1 port map( A => A_s(11), ZN => n573);
   U243 : INV_X1 port map( A => A_ns(11), ZN => n572);
   U244 : OAI221_X1 port map( B1 => n393, B2 => n575, C1 => n392, C2 => n576, A
                           => n577, ZN => O_12_port);
   U245 : AOI22_X1 port map( A1 => A_ns(11), A2 => n397, B1 => A_s(11), B2 => 
                           n398, ZN => n577);
   U246 : INV_X1 port map( A => A_s(10), ZN => n576);
   U247 : INV_X1 port map( A => A_ns(10), ZN => n575);
   U248 : OAI221_X1 port map( B1 => n393, B2 => n578, C1 => n392, C2 => n579, A
                           => n580, ZN => O_11_port);
   U249 : AOI22_X1 port map( A1 => A_ns(10), A2 => n397, B1 => A_s(10), B2 => 
                           n398, ZN => n580);
   U250 : INV_X1 port map( A => A_s(9), ZN => n579);
   U251 : INV_X1 port map( A => A_ns(9), ZN => n578);
   U252 : OAI221_X1 port map( B1 => n581, B2 => n393, C1 => n582, C2 => n392, A
                           => n583, ZN => O_10_port);
   U253 : AOI22_X1 port map( A1 => A_ns(9), A2 => n397, B1 => A_s(9), B2 => 
                           n398, ZN => n583);
   U254 : NAND2_X1 port map( A1 => n584, A2 => n552, ZN => n553);
   U255 : NAND2_X1 port map( A1 => n584, A2 => n585, ZN => n552);
   U256 : XOR2_X1 port map( A => B(17), B => B(18), Z => n584);
   U257 : INV_X1 port map( A => A_s(8), ZN => n582);
   U258 : INV_X1 port map( A => B(19), ZN => n585);
   U259 : INV_X1 port map( A => A_ns(8), ZN => n581);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity BOOTHENC_NBIT64_i16 is

   port( A, A_n, A_ns, A_s, B : in std_logic_vector (63 downto 0);  O, A_so, 
         A_nso : out std_logic_vector (63 downto 0));

end BOOTHENC_NBIT64_i16;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT64_i16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, O_63_port, O_62_port, O_61_port, O_60_port, O_59_port,
      O_58_port, O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, 
      O_52_port, O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, 
      O_46_port, O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, 
      O_40_port, O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, 
      O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, 
      O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, 
      O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, 
      O_16_port, O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, 
      O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, 
      O_3_port, O_2_port, O_1_port, n391, n392, n393, n394, n395, n396, n397, 
      n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, 
      n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, 
      n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, 
      n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, 
      n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, 
      n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, 
      n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, 
      n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, 
      n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, 
      n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, 
      n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, 
      n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, 
      n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, 
      n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, 
      n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, 
      n578, n579, n580, n581, n582, n583, n584, n585 : std_logic;

begin
   O <= ( O_63_port, O_62_port, O_61_port, O_60_port, O_59_port, O_58_port, 
      O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, O_52_port, 
      O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, O_46_port, 
      O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, O_40_port, 
      O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, 
      O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, 
      O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, 
      O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, O_16_port, 
      O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, O_10_port, 
      O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, O_3_port, 
      O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(61), A_s(60), A_s(59), A_s(58), A_s(57), A_s(56), A_s(55), 
      A_s(54), A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), 
      A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), 
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   A_nso <= ( A_s(61), A_s(60), A_s(59), A_s(58), A_s(57), A_s(56), A_s(55), 
      A_s(54), A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), 
      A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), 
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : AND3_X1 port map( A1 => B(16), A2 => n585, A3 => B(15), ZN => n391);
   U3 : INV_X4 port map( A => n391, ZN => n392);
   U4 : INV_X4 port map( A => n552, ZN => n398);
   U5 : OR3_X4 port map( A1 => B(15), A2 => B(16), A3 => n585, ZN => n393);
   U6 : INV_X4 port map( A => n553, ZN => n397);
   U7 : OAI221_X1 port map( B1 => n393, B2 => n394, C1 => n392, C2 => n395, A 
                           => n396, ZN => O_9_port);
   U8 : AOI22_X1 port map( A1 => A_ns(8), A2 => n397, B1 => A_s(8), B2 => n398,
                           ZN => n396);
   U9 : INV_X1 port map( A => A_s(7), ZN => n395);
   U10 : INV_X1 port map( A => A_ns(7), ZN => n394);
   U11 : OAI221_X1 port map( B1 => n393, B2 => n399, C1 => n392, C2 => n400, A 
                           => n401, ZN => O_8_port);
   U12 : AOI22_X1 port map( A1 => A_ns(7), A2 => n397, B1 => A_s(7), B2 => n398
                           , ZN => n401);
   U13 : INV_X1 port map( A => A_s(6), ZN => n400);
   U14 : INV_X1 port map( A => A_ns(6), ZN => n399);
   U15 : OAI221_X1 port map( B1 => n393, B2 => n402, C1 => n392, C2 => n403, A 
                           => n404, ZN => O_7_port);
   U16 : AOI22_X1 port map( A1 => A_ns(6), A2 => n397, B1 => A_s(6), B2 => n398
                           , ZN => n404);
   U17 : INV_X1 port map( A => A_s(5), ZN => n403);
   U18 : INV_X1 port map( A => A_ns(5), ZN => n402);
   U19 : OAI221_X1 port map( B1 => n393, B2 => n405, C1 => n392, C2 => n406, A 
                           => n407, ZN => O_6_port);
   U20 : AOI22_X1 port map( A1 => A_ns(5), A2 => n397, B1 => A_s(5), B2 => n398
                           , ZN => n407);
   U21 : INV_X1 port map( A => A_s(4), ZN => n406);
   U22 : INV_X1 port map( A => A_ns(4), ZN => n405);
   U23 : OAI221_X1 port map( B1 => n393, B2 => n408, C1 => n392, C2 => n409, A 
                           => n410, ZN => O_63_port);
   U24 : AOI22_X1 port map( A1 => A_ns(62), A2 => n397, B1 => A_s(62), B2 => 
                           n398, ZN => n410);
   U25 : INV_X1 port map( A => A_s(61), ZN => n409);
   U26 : INV_X1 port map( A => A_ns(61), ZN => n408);
   U27 : OAI221_X1 port map( B1 => n393, B2 => n411, C1 => n392, C2 => n412, A 
                           => n413, ZN => O_62_port);
   U28 : AOI22_X1 port map( A1 => A_ns(61), A2 => n397, B1 => A_s(61), B2 => 
                           n398, ZN => n413);
   U29 : INV_X1 port map( A => A_s(60), ZN => n412);
   U30 : INV_X1 port map( A => A_ns(60), ZN => n411);
   U31 : OAI221_X1 port map( B1 => n393, B2 => n414, C1 => n392, C2 => n415, A 
                           => n416, ZN => O_61_port);
   U32 : AOI22_X1 port map( A1 => A_ns(60), A2 => n397, B1 => A_s(60), B2 => 
                           n398, ZN => n416);
   U33 : INV_X1 port map( A => A_s(59), ZN => n415);
   U34 : INV_X1 port map( A => A_ns(59), ZN => n414);
   U35 : OAI221_X1 port map( B1 => n393, B2 => n417, C1 => n392, C2 => n418, A 
                           => n419, ZN => O_60_port);
   U36 : AOI22_X1 port map( A1 => A_ns(59), A2 => n397, B1 => A_s(59), B2 => 
                           n398, ZN => n419);
   U37 : INV_X1 port map( A => A_s(58), ZN => n418);
   U38 : INV_X1 port map( A => A_ns(58), ZN => n417);
   U39 : OAI221_X1 port map( B1 => n393, B2 => n420, C1 => n392, C2 => n421, A 
                           => n422, ZN => O_5_port);
   U40 : AOI22_X1 port map( A1 => A_ns(4), A2 => n397, B1 => A_s(4), B2 => n398
                           , ZN => n422);
   U41 : INV_X1 port map( A => A_s(3), ZN => n421);
   U42 : INV_X1 port map( A => A_ns(3), ZN => n420);
   U43 : OAI221_X1 port map( B1 => n393, B2 => n423, C1 => n392, C2 => n424, A 
                           => n425, ZN => O_59_port);
   U44 : AOI22_X1 port map( A1 => A_ns(58), A2 => n397, B1 => A_s(58), B2 => 
                           n398, ZN => n425);
   U45 : INV_X1 port map( A => A_s(57), ZN => n424);
   U46 : INV_X1 port map( A => A_ns(57), ZN => n423);
   U47 : OAI221_X1 port map( B1 => n393, B2 => n426, C1 => n392, C2 => n427, A 
                           => n428, ZN => O_58_port);
   U48 : AOI22_X1 port map( A1 => A_ns(57), A2 => n397, B1 => A_s(57), B2 => 
                           n398, ZN => n428);
   U49 : INV_X1 port map( A => A_s(56), ZN => n427);
   U50 : INV_X1 port map( A => A_ns(56), ZN => n426);
   U51 : OAI221_X1 port map( B1 => n393, B2 => n429, C1 => n392, C2 => n430, A 
                           => n431, ZN => O_57_port);
   U52 : AOI22_X1 port map( A1 => A_ns(56), A2 => n397, B1 => A_s(56), B2 => 
                           n398, ZN => n431);
   U53 : INV_X1 port map( A => A_s(55), ZN => n430);
   U54 : INV_X1 port map( A => A_ns(55), ZN => n429);
   U55 : OAI221_X1 port map( B1 => n393, B2 => n432, C1 => n392, C2 => n433, A 
                           => n434, ZN => O_56_port);
   U56 : AOI22_X1 port map( A1 => A_ns(55), A2 => n397, B1 => A_s(55), B2 => 
                           n398, ZN => n434);
   U57 : INV_X1 port map( A => A_s(54), ZN => n433);
   U58 : INV_X1 port map( A => A_ns(54), ZN => n432);
   U59 : OAI221_X1 port map( B1 => n393, B2 => n435, C1 => n392, C2 => n436, A 
                           => n437, ZN => O_55_port);
   U60 : AOI22_X1 port map( A1 => A_ns(54), A2 => n397, B1 => A_s(54), B2 => 
                           n398, ZN => n437);
   U61 : INV_X1 port map( A => A_s(53), ZN => n436);
   U62 : INV_X1 port map( A => A_ns(53), ZN => n435);
   U63 : OAI221_X1 port map( B1 => n393, B2 => n438, C1 => n392, C2 => n439, A 
                           => n440, ZN => O_54_port);
   U64 : AOI22_X1 port map( A1 => A_ns(53), A2 => n397, B1 => A_s(53), B2 => 
                           n398, ZN => n440);
   U65 : INV_X1 port map( A => A_s(52), ZN => n439);
   U66 : INV_X1 port map( A => A_ns(52), ZN => n438);
   U67 : OAI221_X1 port map( B1 => n393, B2 => n441, C1 => n392, C2 => n442, A 
                           => n443, ZN => O_53_port);
   U68 : AOI22_X1 port map( A1 => A_ns(52), A2 => n397, B1 => A_s(52), B2 => 
                           n398, ZN => n443);
   U69 : INV_X1 port map( A => A_s(51), ZN => n442);
   U70 : INV_X1 port map( A => A_ns(51), ZN => n441);
   U71 : OAI221_X1 port map( B1 => n393, B2 => n444, C1 => n392, C2 => n445, A 
                           => n446, ZN => O_52_port);
   U72 : AOI22_X1 port map( A1 => A_ns(51), A2 => n397, B1 => A_s(51), B2 => 
                           n398, ZN => n446);
   U73 : INV_X1 port map( A => A_s(50), ZN => n445);
   U74 : INV_X1 port map( A => A_ns(50), ZN => n444);
   U75 : OAI221_X1 port map( B1 => n393, B2 => n447, C1 => n392, C2 => n448, A 
                           => n449, ZN => O_51_port);
   U76 : AOI22_X1 port map( A1 => A_ns(50), A2 => n397, B1 => A_s(50), B2 => 
                           n398, ZN => n449);
   U77 : INV_X1 port map( A => A_s(49), ZN => n448);
   U78 : INV_X1 port map( A => A_ns(49), ZN => n447);
   U79 : OAI221_X1 port map( B1 => n393, B2 => n450, C1 => n392, C2 => n451, A 
                           => n452, ZN => O_50_port);
   U80 : AOI22_X1 port map( A1 => A_ns(49), A2 => n397, B1 => A_s(49), B2 => 
                           n398, ZN => n452);
   U81 : INV_X1 port map( A => A_s(48), ZN => n451);
   U82 : INV_X1 port map( A => A_ns(48), ZN => n450);
   U83 : OAI221_X1 port map( B1 => n393, B2 => n453, C1 => n392, C2 => n454, A 
                           => n455, ZN => O_4_port);
   U84 : AOI22_X1 port map( A1 => A_ns(3), A2 => n397, B1 => A_s(3), B2 => n398
                           , ZN => n455);
   U85 : INV_X1 port map( A => A_s(2), ZN => n454);
   U86 : INV_X1 port map( A => A_ns(2), ZN => n453);
   U87 : OAI221_X1 port map( B1 => n393, B2 => n456, C1 => n392, C2 => n457, A 
                           => n458, ZN => O_49_port);
   U88 : AOI22_X1 port map( A1 => A_ns(48), A2 => n397, B1 => A_s(48), B2 => 
                           n398, ZN => n458);
   U89 : INV_X1 port map( A => A_s(47), ZN => n457);
   U90 : INV_X1 port map( A => A_ns(47), ZN => n456);
   U91 : OAI221_X1 port map( B1 => n393, B2 => n459, C1 => n392, C2 => n460, A 
                           => n461, ZN => O_48_port);
   U92 : AOI22_X1 port map( A1 => A_ns(47), A2 => n397, B1 => A_s(47), B2 => 
                           n398, ZN => n461);
   U93 : INV_X1 port map( A => A_s(46), ZN => n460);
   U94 : INV_X1 port map( A => A_ns(46), ZN => n459);
   U95 : OAI221_X1 port map( B1 => n393, B2 => n462, C1 => n392, C2 => n463, A 
                           => n464, ZN => O_47_port);
   U96 : AOI22_X1 port map( A1 => A_ns(46), A2 => n397, B1 => A_s(46), B2 => 
                           n398, ZN => n464);
   U97 : INV_X1 port map( A => A_s(45), ZN => n463);
   U98 : INV_X1 port map( A => A_ns(45), ZN => n462);
   U99 : OAI221_X1 port map( B1 => n393, B2 => n465, C1 => n392, C2 => n466, A 
                           => n467, ZN => O_46_port);
   U100 : AOI22_X1 port map( A1 => A_ns(45), A2 => n397, B1 => A_s(45), B2 => 
                           n398, ZN => n467);
   U101 : INV_X1 port map( A => A_s(44), ZN => n466);
   U102 : INV_X1 port map( A => A_ns(44), ZN => n465);
   U103 : OAI221_X1 port map( B1 => n393, B2 => n468, C1 => n392, C2 => n469, A
                           => n470, ZN => O_45_port);
   U104 : AOI22_X1 port map( A1 => A_ns(44), A2 => n397, B1 => A_s(44), B2 => 
                           n398, ZN => n470);
   U105 : INV_X1 port map( A => A_s(43), ZN => n469);
   U106 : INV_X1 port map( A => A_ns(43), ZN => n468);
   U107 : OAI221_X1 port map( B1 => n393, B2 => n471, C1 => n392, C2 => n472, A
                           => n473, ZN => O_44_port);
   U108 : AOI22_X1 port map( A1 => A_ns(43), A2 => n397, B1 => A_s(43), B2 => 
                           n398, ZN => n473);
   U109 : INV_X1 port map( A => A_s(42), ZN => n472);
   U110 : INV_X1 port map( A => A_ns(42), ZN => n471);
   U111 : OAI221_X1 port map( B1 => n393, B2 => n474, C1 => n392, C2 => n475, A
                           => n476, ZN => O_43_port);
   U112 : AOI22_X1 port map( A1 => A_ns(42), A2 => n397, B1 => A_s(42), B2 => 
                           n398, ZN => n476);
   U113 : INV_X1 port map( A => A_s(41), ZN => n475);
   U114 : INV_X1 port map( A => A_ns(41), ZN => n474);
   U115 : OAI221_X1 port map( B1 => n393, B2 => n477, C1 => n392, C2 => n478, A
                           => n479, ZN => O_42_port);
   U116 : AOI22_X1 port map( A1 => A_ns(41), A2 => n397, B1 => A_s(41), B2 => 
                           n398, ZN => n479);
   U117 : INV_X1 port map( A => A_s(40), ZN => n478);
   U118 : INV_X1 port map( A => A_ns(40), ZN => n477);
   U119 : OAI221_X1 port map( B1 => n393, B2 => n480, C1 => n392, C2 => n481, A
                           => n482, ZN => O_41_port);
   U120 : AOI22_X1 port map( A1 => A_ns(40), A2 => n397, B1 => A_s(40), B2 => 
                           n398, ZN => n482);
   U121 : INV_X1 port map( A => A_s(39), ZN => n481);
   U122 : INV_X1 port map( A => A_ns(39), ZN => n480);
   U123 : OAI221_X1 port map( B1 => n393, B2 => n483, C1 => n392, C2 => n484, A
                           => n485, ZN => O_40_port);
   U124 : AOI22_X1 port map( A1 => A_ns(39), A2 => n397, B1 => A_s(39), B2 => 
                           n398, ZN => n485);
   U125 : INV_X1 port map( A => A_s(38), ZN => n484);
   U126 : INV_X1 port map( A => A_ns(38), ZN => n483);
   U127 : OAI221_X1 port map( B1 => n393, B2 => n486, C1 => n392, C2 => n487, A
                           => n488, ZN => O_3_port);
   U128 : AOI22_X1 port map( A1 => A_ns(2), A2 => n397, B1 => A_s(2), B2 => 
                           n398, ZN => n488);
   U129 : INV_X1 port map( A => A_s(1), ZN => n487);
   U130 : INV_X1 port map( A => A_ns(1), ZN => n486);
   U131 : OAI221_X1 port map( B1 => n393, B2 => n489, C1 => n392, C2 => n490, A
                           => n491, ZN => O_39_port);
   U132 : AOI22_X1 port map( A1 => A_ns(38), A2 => n397, B1 => A_s(38), B2 => 
                           n398, ZN => n491);
   U133 : INV_X1 port map( A => A_s(37), ZN => n490);
   U134 : INV_X1 port map( A => A_ns(37), ZN => n489);
   U135 : OAI221_X1 port map( B1 => n393, B2 => n492, C1 => n392, C2 => n493, A
                           => n494, ZN => O_38_port);
   U136 : AOI22_X1 port map( A1 => A_ns(37), A2 => n397, B1 => A_s(37), B2 => 
                           n398, ZN => n494);
   U137 : INV_X1 port map( A => A_s(36), ZN => n493);
   U138 : INV_X1 port map( A => A_ns(36), ZN => n492);
   U139 : OAI221_X1 port map( B1 => n393, B2 => n495, C1 => n392, C2 => n496, A
                           => n497, ZN => O_37_port);
   U140 : AOI22_X1 port map( A1 => A_ns(36), A2 => n397, B1 => A_s(36), B2 => 
                           n398, ZN => n497);
   U141 : INV_X1 port map( A => A_s(35), ZN => n496);
   U142 : INV_X1 port map( A => A_ns(35), ZN => n495);
   U143 : OAI221_X1 port map( B1 => n393, B2 => n498, C1 => n392, C2 => n499, A
                           => n500, ZN => O_36_port);
   U144 : AOI22_X1 port map( A1 => A_ns(35), A2 => n397, B1 => A_s(35), B2 => 
                           n398, ZN => n500);
   U145 : INV_X1 port map( A => A_s(34), ZN => n499);
   U146 : INV_X1 port map( A => A_ns(34), ZN => n498);
   U147 : OAI221_X1 port map( B1 => n393, B2 => n501, C1 => n392, C2 => n502, A
                           => n503, ZN => O_35_port);
   U148 : AOI22_X1 port map( A1 => A_ns(34), A2 => n397, B1 => A_s(34), B2 => 
                           n398, ZN => n503);
   U149 : INV_X1 port map( A => A_s(33), ZN => n502);
   U150 : INV_X1 port map( A => A_ns(33), ZN => n501);
   U151 : OAI221_X1 port map( B1 => n393, B2 => n504, C1 => n392, C2 => n505, A
                           => n506, ZN => O_34_port);
   U152 : AOI22_X1 port map( A1 => A_ns(33), A2 => n397, B1 => A_s(33), B2 => 
                           n398, ZN => n506);
   U153 : INV_X1 port map( A => A_s(32), ZN => n505);
   U154 : INV_X1 port map( A => A_ns(32), ZN => n504);
   U155 : OAI221_X1 port map( B1 => n393, B2 => n507, C1 => n392, C2 => n508, A
                           => n509, ZN => O_33_port);
   U156 : AOI22_X1 port map( A1 => A_ns(32), A2 => n397, B1 => A_s(32), B2 => 
                           n398, ZN => n509);
   U157 : INV_X1 port map( A => A_s(31), ZN => n508);
   U158 : INV_X1 port map( A => A_ns(31), ZN => n507);
   U159 : OAI221_X1 port map( B1 => n393, B2 => n510, C1 => n392, C2 => n511, A
                           => n512, ZN => O_32_port);
   U160 : AOI22_X1 port map( A1 => A_ns(31), A2 => n397, B1 => A_s(31), B2 => 
                           n398, ZN => n512);
   U161 : INV_X1 port map( A => A_s(30), ZN => n511);
   U162 : INV_X1 port map( A => A_ns(30), ZN => n510);
   U163 : OAI221_X1 port map( B1 => n393, B2 => n513, C1 => n392, C2 => n514, A
                           => n515, ZN => O_31_port);
   U164 : AOI22_X1 port map( A1 => A_ns(30), A2 => n397, B1 => A_s(30), B2 => 
                           n398, ZN => n515);
   U165 : INV_X1 port map( A => A_s(29), ZN => n514);
   U166 : INV_X1 port map( A => A_ns(29), ZN => n513);
   U167 : OAI221_X1 port map( B1 => n393, B2 => n516, C1 => n392, C2 => n517, A
                           => n518, ZN => O_30_port);
   U168 : AOI22_X1 port map( A1 => A_ns(29), A2 => n397, B1 => A_s(29), B2 => 
                           n398, ZN => n518);
   U169 : INV_X1 port map( A => A_s(28), ZN => n517);
   U170 : INV_X1 port map( A => A_ns(28), ZN => n516);
   U171 : OAI221_X1 port map( B1 => n393, B2 => n519, C1 => n392, C2 => n520, A
                           => n521, ZN => O_2_port);
   U172 : AOI22_X1 port map( A1 => A_ns(1), A2 => n397, B1 => A_s(1), B2 => 
                           n398, ZN => n521);
   U173 : OAI221_X1 port map( B1 => n393, B2 => n522, C1 => n392, C2 => n523, A
                           => n524, ZN => O_29_port);
   U174 : AOI22_X1 port map( A1 => A_ns(28), A2 => n397, B1 => A_s(28), B2 => 
                           n398, ZN => n524);
   U175 : INV_X1 port map( A => A_s(27), ZN => n523);
   U176 : INV_X1 port map( A => A_ns(27), ZN => n522);
   U177 : OAI221_X1 port map( B1 => n393, B2 => n525, C1 => n392, C2 => n526, A
                           => n527, ZN => O_28_port);
   U178 : AOI22_X1 port map( A1 => A_ns(27), A2 => n397, B1 => A_s(27), B2 => 
                           n398, ZN => n527);
   U179 : INV_X1 port map( A => A_s(26), ZN => n526);
   U180 : INV_X1 port map( A => A_ns(26), ZN => n525);
   U181 : OAI221_X1 port map( B1 => n393, B2 => n528, C1 => n392, C2 => n529, A
                           => n530, ZN => O_27_port);
   U182 : AOI22_X1 port map( A1 => A_ns(26), A2 => n397, B1 => A_s(26), B2 => 
                           n398, ZN => n530);
   U183 : INV_X1 port map( A => A_s(25), ZN => n529);
   U184 : INV_X1 port map( A => A_ns(25), ZN => n528);
   U185 : OAI221_X1 port map( B1 => n393, B2 => n531, C1 => n392, C2 => n532, A
                           => n533, ZN => O_26_port);
   U186 : AOI22_X1 port map( A1 => A_ns(25), A2 => n397, B1 => A_s(25), B2 => 
                           n398, ZN => n533);
   U187 : INV_X1 port map( A => A_s(24), ZN => n532);
   U188 : INV_X1 port map( A => A_ns(24), ZN => n531);
   U189 : OAI221_X1 port map( B1 => n393, B2 => n534, C1 => n392, C2 => n535, A
                           => n536, ZN => O_25_port);
   U190 : AOI22_X1 port map( A1 => A_ns(24), A2 => n397, B1 => A_s(24), B2 => 
                           n398, ZN => n536);
   U191 : INV_X1 port map( A => A_s(23), ZN => n535);
   U192 : INV_X1 port map( A => A_ns(23), ZN => n534);
   U193 : OAI221_X1 port map( B1 => n393, B2 => n537, C1 => n392, C2 => n538, A
                           => n539, ZN => O_24_port);
   U194 : AOI22_X1 port map( A1 => A_ns(23), A2 => n397, B1 => A_s(23), B2 => 
                           n398, ZN => n539);
   U195 : INV_X1 port map( A => A_s(22), ZN => n538);
   U196 : INV_X1 port map( A => A_ns(22), ZN => n537);
   U197 : OAI221_X1 port map( B1 => n393, B2 => n540, C1 => n392, C2 => n541, A
                           => n542, ZN => O_23_port);
   U198 : AOI22_X1 port map( A1 => A_ns(22), A2 => n397, B1 => A_s(22), B2 => 
                           n398, ZN => n542);
   U199 : INV_X1 port map( A => A_s(21), ZN => n541);
   U200 : INV_X1 port map( A => A_ns(21), ZN => n540);
   U201 : OAI221_X1 port map( B1 => n393, B2 => n543, C1 => n392, C2 => n544, A
                           => n545, ZN => O_22_port);
   U202 : AOI22_X1 port map( A1 => A_ns(21), A2 => n397, B1 => A_s(21), B2 => 
                           n398, ZN => n545);
   U203 : INV_X1 port map( A => A_s(20), ZN => n544);
   U204 : INV_X1 port map( A => A_ns(20), ZN => n543);
   U205 : OAI221_X1 port map( B1 => n393, B2 => n546, C1 => n392, C2 => n547, A
                           => n548, ZN => O_21_port);
   U206 : AOI22_X1 port map( A1 => A_ns(20), A2 => n397, B1 => A_s(20), B2 => 
                           n398, ZN => n548);
   U207 : INV_X1 port map( A => A_s(19), ZN => n547);
   U208 : INV_X1 port map( A => A_ns(19), ZN => n546);
   U209 : OAI221_X1 port map( B1 => n393, B2 => n549, C1 => n392, C2 => n550, A
                           => n551, ZN => O_20_port);
   U210 : AOI22_X1 port map( A1 => A_ns(19), A2 => n397, B1 => A_s(19), B2 => 
                           n398, ZN => n551);
   U211 : INV_X1 port map( A => A_s(18), ZN => n550);
   U212 : INV_X1 port map( A => A_ns(18), ZN => n549);
   U213 : OAI22_X1 port map( A1 => n552, A2 => n520, B1 => n553, B2 => n519, ZN
                           => O_1_port);
   U214 : INV_X1 port map( A => A_ns(0), ZN => n519);
   U215 : INV_X1 port map( A => A_s(0), ZN => n520);
   U216 : OAI221_X1 port map( B1 => n393, B2 => n554, C1 => n392, C2 => n555, A
                           => n556, ZN => O_19_port);
   U217 : AOI22_X1 port map( A1 => A_ns(18), A2 => n397, B1 => A_s(18), B2 => 
                           n398, ZN => n556);
   U218 : INV_X1 port map( A => A_s(17), ZN => n555);
   U219 : INV_X1 port map( A => A_ns(17), ZN => n554);
   U220 : OAI221_X1 port map( B1 => n393, B2 => n557, C1 => n392, C2 => n558, A
                           => n559, ZN => O_18_port);
   U221 : AOI22_X1 port map( A1 => A_ns(17), A2 => n397, B1 => A_s(17), B2 => 
                           n398, ZN => n559);
   U222 : INV_X1 port map( A => A_s(16), ZN => n558);
   U223 : INV_X1 port map( A => A_ns(16), ZN => n557);
   U224 : OAI221_X1 port map( B1 => n393, B2 => n560, C1 => n392, C2 => n561, A
                           => n562, ZN => O_17_port);
   U225 : AOI22_X1 port map( A1 => A_ns(16), A2 => n397, B1 => A_s(16), B2 => 
                           n398, ZN => n562);
   U226 : INV_X1 port map( A => A_s(15), ZN => n561);
   U227 : INV_X1 port map( A => A_ns(15), ZN => n560);
   U228 : OAI221_X1 port map( B1 => n393, B2 => n563, C1 => n392, C2 => n564, A
                           => n565, ZN => O_16_port);
   U229 : AOI22_X1 port map( A1 => A_ns(15), A2 => n397, B1 => A_s(15), B2 => 
                           n398, ZN => n565);
   U230 : INV_X1 port map( A => A_s(14), ZN => n564);
   U231 : INV_X1 port map( A => A_ns(14), ZN => n563);
   U232 : OAI221_X1 port map( B1 => n393, B2 => n566, C1 => n392, C2 => n567, A
                           => n568, ZN => O_15_port);
   U233 : AOI22_X1 port map( A1 => A_ns(14), A2 => n397, B1 => A_s(14), B2 => 
                           n398, ZN => n568);
   U234 : INV_X1 port map( A => A_s(13), ZN => n567);
   U235 : INV_X1 port map( A => A_ns(13), ZN => n566);
   U236 : OAI221_X1 port map( B1 => n393, B2 => n569, C1 => n392, C2 => n570, A
                           => n571, ZN => O_14_port);
   U237 : AOI22_X1 port map( A1 => A_ns(13), A2 => n397, B1 => A_s(13), B2 => 
                           n398, ZN => n571);
   U238 : INV_X1 port map( A => A_s(12), ZN => n570);
   U239 : INV_X1 port map( A => A_ns(12), ZN => n569);
   U240 : OAI221_X1 port map( B1 => n393, B2 => n572, C1 => n392, C2 => n573, A
                           => n574, ZN => O_13_port);
   U241 : AOI22_X1 port map( A1 => A_ns(12), A2 => n397, B1 => A_s(12), B2 => 
                           n398, ZN => n574);
   U242 : INV_X1 port map( A => A_s(11), ZN => n573);
   U243 : INV_X1 port map( A => A_ns(11), ZN => n572);
   U244 : OAI221_X1 port map( B1 => n393, B2 => n575, C1 => n392, C2 => n576, A
                           => n577, ZN => O_12_port);
   U245 : AOI22_X1 port map( A1 => A_ns(11), A2 => n397, B1 => A_s(11), B2 => 
                           n398, ZN => n577);
   U246 : INV_X1 port map( A => A_s(10), ZN => n576);
   U247 : INV_X1 port map( A => A_ns(10), ZN => n575);
   U248 : OAI221_X1 port map( B1 => n393, B2 => n578, C1 => n392, C2 => n579, A
                           => n580, ZN => O_11_port);
   U249 : AOI22_X1 port map( A1 => A_ns(10), A2 => n397, B1 => A_s(10), B2 => 
                           n398, ZN => n580);
   U250 : INV_X1 port map( A => A_s(9), ZN => n579);
   U251 : INV_X1 port map( A => A_ns(9), ZN => n578);
   U252 : OAI221_X1 port map( B1 => n581, B2 => n393, C1 => n582, C2 => n392, A
                           => n583, ZN => O_10_port);
   U253 : AOI22_X1 port map( A1 => A_ns(9), A2 => n397, B1 => A_s(9), B2 => 
                           n398, ZN => n583);
   U254 : NAND2_X1 port map( A1 => n584, A2 => n552, ZN => n553);
   U255 : NAND2_X1 port map( A1 => n584, A2 => n585, ZN => n552);
   U256 : XOR2_X1 port map( A => B(15), B => B(16), Z => n584);
   U257 : INV_X1 port map( A => A_s(8), ZN => n582);
   U258 : INV_X1 port map( A => B(17), ZN => n585);
   U259 : INV_X1 port map( A => A_ns(8), ZN => n581);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity BOOTHENC_NBIT64_i14 is

   port( A, A_n, A_ns, A_s, B : in std_logic_vector (63 downto 0);  O, A_so, 
         A_nso : out std_logic_vector (63 downto 0));

end BOOTHENC_NBIT64_i14;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT64_i14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, O_63_port, O_62_port, O_61_port, O_60_port, O_59_port,
      O_58_port, O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, 
      O_52_port, O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, 
      O_46_port, O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, 
      O_40_port, O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, 
      O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, 
      O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, 
      O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, 
      O_16_port, O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, 
      O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, 
      O_3_port, O_2_port, O_1_port, n391, n392, n393, n394, n395, n396, n397, 
      n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, 
      n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, 
      n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, 
      n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, 
      n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, 
      n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, 
      n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, 
      n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, 
      n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, 
      n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, 
      n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, 
      n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, 
      n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, 
      n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, 
      n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, 
      n578, n579, n580, n581, n582, n583, n584, n585 : std_logic;

begin
   O <= ( O_63_port, O_62_port, O_61_port, O_60_port, O_59_port, O_58_port, 
      O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, O_52_port, 
      O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, O_46_port, 
      O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, O_40_port, 
      O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, 
      O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, 
      O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, 
      O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, O_16_port, 
      O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, O_10_port, 
      O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, O_3_port, 
      O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(61), A_s(60), A_s(59), A_s(58), A_s(57), A_s(56), A_s(55), 
      A_s(54), A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), 
      A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), 
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   A_nso <= ( A_s(61), A_s(60), A_s(59), A_s(58), A_s(57), A_s(56), A_s(55), 
      A_s(54), A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), 
      A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), 
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : AND3_X1 port map( A1 => B(14), A2 => n585, A3 => B(13), ZN => n391);
   U3 : INV_X4 port map( A => n391, ZN => n392);
   U4 : INV_X4 port map( A => n552, ZN => n398);
   U5 : OR3_X4 port map( A1 => B(13), A2 => B(14), A3 => n585, ZN => n393);
   U6 : INV_X4 port map( A => n553, ZN => n397);
   U7 : OAI221_X1 port map( B1 => n393, B2 => n394, C1 => n392, C2 => n395, A 
                           => n396, ZN => O_9_port);
   U8 : AOI22_X1 port map( A1 => A_ns(8), A2 => n397, B1 => A_s(8), B2 => n398,
                           ZN => n396);
   U9 : INV_X1 port map( A => A_s(7), ZN => n395);
   U10 : INV_X1 port map( A => A_ns(7), ZN => n394);
   U11 : OAI221_X1 port map( B1 => n393, B2 => n399, C1 => n392, C2 => n400, A 
                           => n401, ZN => O_8_port);
   U12 : AOI22_X1 port map( A1 => A_ns(7), A2 => n397, B1 => A_s(7), B2 => n398
                           , ZN => n401);
   U13 : INV_X1 port map( A => A_s(6), ZN => n400);
   U14 : INV_X1 port map( A => A_ns(6), ZN => n399);
   U15 : OAI221_X1 port map( B1 => n393, B2 => n402, C1 => n392, C2 => n403, A 
                           => n404, ZN => O_7_port);
   U16 : AOI22_X1 port map( A1 => A_ns(6), A2 => n397, B1 => A_s(6), B2 => n398
                           , ZN => n404);
   U17 : INV_X1 port map( A => A_s(5), ZN => n403);
   U18 : INV_X1 port map( A => A_ns(5), ZN => n402);
   U19 : OAI221_X1 port map( B1 => n393, B2 => n405, C1 => n392, C2 => n406, A 
                           => n407, ZN => O_6_port);
   U20 : AOI22_X1 port map( A1 => A_ns(5), A2 => n397, B1 => A_s(5), B2 => n398
                           , ZN => n407);
   U21 : INV_X1 port map( A => A_s(4), ZN => n406);
   U22 : INV_X1 port map( A => A_ns(4), ZN => n405);
   U23 : OAI221_X1 port map( B1 => n393, B2 => n408, C1 => n392, C2 => n409, A 
                           => n410, ZN => O_63_port);
   U24 : AOI22_X1 port map( A1 => A_ns(62), A2 => n397, B1 => A_s(62), B2 => 
                           n398, ZN => n410);
   U25 : INV_X1 port map( A => A_s(61), ZN => n409);
   U26 : INV_X1 port map( A => A_ns(61), ZN => n408);
   U27 : OAI221_X1 port map( B1 => n393, B2 => n411, C1 => n392, C2 => n412, A 
                           => n413, ZN => O_62_port);
   U28 : AOI22_X1 port map( A1 => A_ns(61), A2 => n397, B1 => A_s(61), B2 => 
                           n398, ZN => n413);
   U29 : INV_X1 port map( A => A_s(60), ZN => n412);
   U30 : INV_X1 port map( A => A_ns(60), ZN => n411);
   U31 : OAI221_X1 port map( B1 => n393, B2 => n414, C1 => n392, C2 => n415, A 
                           => n416, ZN => O_61_port);
   U32 : AOI22_X1 port map( A1 => A_ns(60), A2 => n397, B1 => A_s(60), B2 => 
                           n398, ZN => n416);
   U33 : INV_X1 port map( A => A_s(59), ZN => n415);
   U34 : INV_X1 port map( A => A_ns(59), ZN => n414);
   U35 : OAI221_X1 port map( B1 => n393, B2 => n417, C1 => n392, C2 => n418, A 
                           => n419, ZN => O_60_port);
   U36 : AOI22_X1 port map( A1 => A_ns(59), A2 => n397, B1 => A_s(59), B2 => 
                           n398, ZN => n419);
   U37 : INV_X1 port map( A => A_s(58), ZN => n418);
   U38 : INV_X1 port map( A => A_ns(58), ZN => n417);
   U39 : OAI221_X1 port map( B1 => n393, B2 => n420, C1 => n392, C2 => n421, A 
                           => n422, ZN => O_5_port);
   U40 : AOI22_X1 port map( A1 => A_ns(4), A2 => n397, B1 => A_s(4), B2 => n398
                           , ZN => n422);
   U41 : INV_X1 port map( A => A_s(3), ZN => n421);
   U42 : INV_X1 port map( A => A_ns(3), ZN => n420);
   U43 : OAI221_X1 port map( B1 => n393, B2 => n423, C1 => n392, C2 => n424, A 
                           => n425, ZN => O_59_port);
   U44 : AOI22_X1 port map( A1 => A_ns(58), A2 => n397, B1 => A_s(58), B2 => 
                           n398, ZN => n425);
   U45 : INV_X1 port map( A => A_s(57), ZN => n424);
   U46 : INV_X1 port map( A => A_ns(57), ZN => n423);
   U47 : OAI221_X1 port map( B1 => n393, B2 => n426, C1 => n392, C2 => n427, A 
                           => n428, ZN => O_58_port);
   U48 : AOI22_X1 port map( A1 => A_ns(57), A2 => n397, B1 => A_s(57), B2 => 
                           n398, ZN => n428);
   U49 : INV_X1 port map( A => A_s(56), ZN => n427);
   U50 : INV_X1 port map( A => A_ns(56), ZN => n426);
   U51 : OAI221_X1 port map( B1 => n393, B2 => n429, C1 => n392, C2 => n430, A 
                           => n431, ZN => O_57_port);
   U52 : AOI22_X1 port map( A1 => A_ns(56), A2 => n397, B1 => A_s(56), B2 => 
                           n398, ZN => n431);
   U53 : INV_X1 port map( A => A_s(55), ZN => n430);
   U54 : INV_X1 port map( A => A_ns(55), ZN => n429);
   U55 : OAI221_X1 port map( B1 => n393, B2 => n432, C1 => n392, C2 => n433, A 
                           => n434, ZN => O_56_port);
   U56 : AOI22_X1 port map( A1 => A_ns(55), A2 => n397, B1 => A_s(55), B2 => 
                           n398, ZN => n434);
   U57 : INV_X1 port map( A => A_s(54), ZN => n433);
   U58 : INV_X1 port map( A => A_ns(54), ZN => n432);
   U59 : OAI221_X1 port map( B1 => n393, B2 => n435, C1 => n392, C2 => n436, A 
                           => n437, ZN => O_55_port);
   U60 : AOI22_X1 port map( A1 => A_ns(54), A2 => n397, B1 => A_s(54), B2 => 
                           n398, ZN => n437);
   U61 : INV_X1 port map( A => A_s(53), ZN => n436);
   U62 : INV_X1 port map( A => A_ns(53), ZN => n435);
   U63 : OAI221_X1 port map( B1 => n393, B2 => n438, C1 => n392, C2 => n439, A 
                           => n440, ZN => O_54_port);
   U64 : AOI22_X1 port map( A1 => A_ns(53), A2 => n397, B1 => A_s(53), B2 => 
                           n398, ZN => n440);
   U65 : INV_X1 port map( A => A_s(52), ZN => n439);
   U66 : INV_X1 port map( A => A_ns(52), ZN => n438);
   U67 : OAI221_X1 port map( B1 => n393, B2 => n441, C1 => n392, C2 => n442, A 
                           => n443, ZN => O_53_port);
   U68 : AOI22_X1 port map( A1 => A_ns(52), A2 => n397, B1 => A_s(52), B2 => 
                           n398, ZN => n443);
   U69 : INV_X1 port map( A => A_s(51), ZN => n442);
   U70 : INV_X1 port map( A => A_ns(51), ZN => n441);
   U71 : OAI221_X1 port map( B1 => n393, B2 => n444, C1 => n392, C2 => n445, A 
                           => n446, ZN => O_52_port);
   U72 : AOI22_X1 port map( A1 => A_ns(51), A2 => n397, B1 => A_s(51), B2 => 
                           n398, ZN => n446);
   U73 : INV_X1 port map( A => A_s(50), ZN => n445);
   U74 : INV_X1 port map( A => A_ns(50), ZN => n444);
   U75 : OAI221_X1 port map( B1 => n393, B2 => n447, C1 => n392, C2 => n448, A 
                           => n449, ZN => O_51_port);
   U76 : AOI22_X1 port map( A1 => A_ns(50), A2 => n397, B1 => A_s(50), B2 => 
                           n398, ZN => n449);
   U77 : INV_X1 port map( A => A_s(49), ZN => n448);
   U78 : INV_X1 port map( A => A_ns(49), ZN => n447);
   U79 : OAI221_X1 port map( B1 => n393, B2 => n450, C1 => n392, C2 => n451, A 
                           => n452, ZN => O_50_port);
   U80 : AOI22_X1 port map( A1 => A_ns(49), A2 => n397, B1 => A_s(49), B2 => 
                           n398, ZN => n452);
   U81 : INV_X1 port map( A => A_s(48), ZN => n451);
   U82 : INV_X1 port map( A => A_ns(48), ZN => n450);
   U83 : OAI221_X1 port map( B1 => n393, B2 => n453, C1 => n392, C2 => n454, A 
                           => n455, ZN => O_4_port);
   U84 : AOI22_X1 port map( A1 => A_ns(3), A2 => n397, B1 => A_s(3), B2 => n398
                           , ZN => n455);
   U85 : INV_X1 port map( A => A_s(2), ZN => n454);
   U86 : INV_X1 port map( A => A_ns(2), ZN => n453);
   U87 : OAI221_X1 port map( B1 => n393, B2 => n456, C1 => n392, C2 => n457, A 
                           => n458, ZN => O_49_port);
   U88 : AOI22_X1 port map( A1 => A_ns(48), A2 => n397, B1 => A_s(48), B2 => 
                           n398, ZN => n458);
   U89 : INV_X1 port map( A => A_s(47), ZN => n457);
   U90 : INV_X1 port map( A => A_ns(47), ZN => n456);
   U91 : OAI221_X1 port map( B1 => n393, B2 => n459, C1 => n392, C2 => n460, A 
                           => n461, ZN => O_48_port);
   U92 : AOI22_X1 port map( A1 => A_ns(47), A2 => n397, B1 => A_s(47), B2 => 
                           n398, ZN => n461);
   U93 : INV_X1 port map( A => A_s(46), ZN => n460);
   U94 : INV_X1 port map( A => A_ns(46), ZN => n459);
   U95 : OAI221_X1 port map( B1 => n393, B2 => n462, C1 => n392, C2 => n463, A 
                           => n464, ZN => O_47_port);
   U96 : AOI22_X1 port map( A1 => A_ns(46), A2 => n397, B1 => A_s(46), B2 => 
                           n398, ZN => n464);
   U97 : INV_X1 port map( A => A_s(45), ZN => n463);
   U98 : INV_X1 port map( A => A_ns(45), ZN => n462);
   U99 : OAI221_X1 port map( B1 => n393, B2 => n465, C1 => n392, C2 => n466, A 
                           => n467, ZN => O_46_port);
   U100 : AOI22_X1 port map( A1 => A_ns(45), A2 => n397, B1 => A_s(45), B2 => 
                           n398, ZN => n467);
   U101 : INV_X1 port map( A => A_s(44), ZN => n466);
   U102 : INV_X1 port map( A => A_ns(44), ZN => n465);
   U103 : OAI221_X1 port map( B1 => n393, B2 => n468, C1 => n392, C2 => n469, A
                           => n470, ZN => O_45_port);
   U104 : AOI22_X1 port map( A1 => A_ns(44), A2 => n397, B1 => A_s(44), B2 => 
                           n398, ZN => n470);
   U105 : INV_X1 port map( A => A_s(43), ZN => n469);
   U106 : INV_X1 port map( A => A_ns(43), ZN => n468);
   U107 : OAI221_X1 port map( B1 => n393, B2 => n471, C1 => n392, C2 => n472, A
                           => n473, ZN => O_44_port);
   U108 : AOI22_X1 port map( A1 => A_ns(43), A2 => n397, B1 => A_s(43), B2 => 
                           n398, ZN => n473);
   U109 : INV_X1 port map( A => A_s(42), ZN => n472);
   U110 : INV_X1 port map( A => A_ns(42), ZN => n471);
   U111 : OAI221_X1 port map( B1 => n393, B2 => n474, C1 => n392, C2 => n475, A
                           => n476, ZN => O_43_port);
   U112 : AOI22_X1 port map( A1 => A_ns(42), A2 => n397, B1 => A_s(42), B2 => 
                           n398, ZN => n476);
   U113 : INV_X1 port map( A => A_s(41), ZN => n475);
   U114 : INV_X1 port map( A => A_ns(41), ZN => n474);
   U115 : OAI221_X1 port map( B1 => n393, B2 => n477, C1 => n392, C2 => n478, A
                           => n479, ZN => O_42_port);
   U116 : AOI22_X1 port map( A1 => A_ns(41), A2 => n397, B1 => A_s(41), B2 => 
                           n398, ZN => n479);
   U117 : INV_X1 port map( A => A_s(40), ZN => n478);
   U118 : INV_X1 port map( A => A_ns(40), ZN => n477);
   U119 : OAI221_X1 port map( B1 => n393, B2 => n480, C1 => n392, C2 => n481, A
                           => n482, ZN => O_41_port);
   U120 : AOI22_X1 port map( A1 => A_ns(40), A2 => n397, B1 => A_s(40), B2 => 
                           n398, ZN => n482);
   U121 : INV_X1 port map( A => A_s(39), ZN => n481);
   U122 : INV_X1 port map( A => A_ns(39), ZN => n480);
   U123 : OAI221_X1 port map( B1 => n393, B2 => n483, C1 => n392, C2 => n484, A
                           => n485, ZN => O_40_port);
   U124 : AOI22_X1 port map( A1 => A_ns(39), A2 => n397, B1 => A_s(39), B2 => 
                           n398, ZN => n485);
   U125 : INV_X1 port map( A => A_s(38), ZN => n484);
   U126 : INV_X1 port map( A => A_ns(38), ZN => n483);
   U127 : OAI221_X1 port map( B1 => n393, B2 => n486, C1 => n392, C2 => n487, A
                           => n488, ZN => O_3_port);
   U128 : AOI22_X1 port map( A1 => A_ns(2), A2 => n397, B1 => A_s(2), B2 => 
                           n398, ZN => n488);
   U129 : INV_X1 port map( A => A_s(1), ZN => n487);
   U130 : INV_X1 port map( A => A_ns(1), ZN => n486);
   U131 : OAI221_X1 port map( B1 => n393, B2 => n489, C1 => n392, C2 => n490, A
                           => n491, ZN => O_39_port);
   U132 : AOI22_X1 port map( A1 => A_ns(38), A2 => n397, B1 => A_s(38), B2 => 
                           n398, ZN => n491);
   U133 : INV_X1 port map( A => A_s(37), ZN => n490);
   U134 : INV_X1 port map( A => A_ns(37), ZN => n489);
   U135 : OAI221_X1 port map( B1 => n393, B2 => n492, C1 => n392, C2 => n493, A
                           => n494, ZN => O_38_port);
   U136 : AOI22_X1 port map( A1 => A_ns(37), A2 => n397, B1 => A_s(37), B2 => 
                           n398, ZN => n494);
   U137 : INV_X1 port map( A => A_s(36), ZN => n493);
   U138 : INV_X1 port map( A => A_ns(36), ZN => n492);
   U139 : OAI221_X1 port map( B1 => n393, B2 => n495, C1 => n392, C2 => n496, A
                           => n497, ZN => O_37_port);
   U140 : AOI22_X1 port map( A1 => A_ns(36), A2 => n397, B1 => A_s(36), B2 => 
                           n398, ZN => n497);
   U141 : INV_X1 port map( A => A_s(35), ZN => n496);
   U142 : INV_X1 port map( A => A_ns(35), ZN => n495);
   U143 : OAI221_X1 port map( B1 => n393, B2 => n498, C1 => n392, C2 => n499, A
                           => n500, ZN => O_36_port);
   U144 : AOI22_X1 port map( A1 => A_ns(35), A2 => n397, B1 => A_s(35), B2 => 
                           n398, ZN => n500);
   U145 : INV_X1 port map( A => A_s(34), ZN => n499);
   U146 : INV_X1 port map( A => A_ns(34), ZN => n498);
   U147 : OAI221_X1 port map( B1 => n393, B2 => n501, C1 => n392, C2 => n502, A
                           => n503, ZN => O_35_port);
   U148 : AOI22_X1 port map( A1 => A_ns(34), A2 => n397, B1 => A_s(34), B2 => 
                           n398, ZN => n503);
   U149 : INV_X1 port map( A => A_s(33), ZN => n502);
   U150 : INV_X1 port map( A => A_ns(33), ZN => n501);
   U151 : OAI221_X1 port map( B1 => n393, B2 => n504, C1 => n392, C2 => n505, A
                           => n506, ZN => O_34_port);
   U152 : AOI22_X1 port map( A1 => A_ns(33), A2 => n397, B1 => A_s(33), B2 => 
                           n398, ZN => n506);
   U153 : INV_X1 port map( A => A_s(32), ZN => n505);
   U154 : INV_X1 port map( A => A_ns(32), ZN => n504);
   U155 : OAI221_X1 port map( B1 => n393, B2 => n507, C1 => n392, C2 => n508, A
                           => n509, ZN => O_33_port);
   U156 : AOI22_X1 port map( A1 => A_ns(32), A2 => n397, B1 => A_s(32), B2 => 
                           n398, ZN => n509);
   U157 : INV_X1 port map( A => A_s(31), ZN => n508);
   U158 : INV_X1 port map( A => A_ns(31), ZN => n507);
   U159 : OAI221_X1 port map( B1 => n393, B2 => n510, C1 => n392, C2 => n511, A
                           => n512, ZN => O_32_port);
   U160 : AOI22_X1 port map( A1 => A_ns(31), A2 => n397, B1 => A_s(31), B2 => 
                           n398, ZN => n512);
   U161 : INV_X1 port map( A => A_s(30), ZN => n511);
   U162 : INV_X1 port map( A => A_ns(30), ZN => n510);
   U163 : OAI221_X1 port map( B1 => n393, B2 => n513, C1 => n392, C2 => n514, A
                           => n515, ZN => O_31_port);
   U164 : AOI22_X1 port map( A1 => A_ns(30), A2 => n397, B1 => A_s(30), B2 => 
                           n398, ZN => n515);
   U165 : INV_X1 port map( A => A_s(29), ZN => n514);
   U166 : INV_X1 port map( A => A_ns(29), ZN => n513);
   U167 : OAI221_X1 port map( B1 => n393, B2 => n516, C1 => n392, C2 => n517, A
                           => n518, ZN => O_30_port);
   U168 : AOI22_X1 port map( A1 => A_ns(29), A2 => n397, B1 => A_s(29), B2 => 
                           n398, ZN => n518);
   U169 : INV_X1 port map( A => A_s(28), ZN => n517);
   U170 : INV_X1 port map( A => A_ns(28), ZN => n516);
   U171 : OAI221_X1 port map( B1 => n393, B2 => n519, C1 => n392, C2 => n520, A
                           => n521, ZN => O_2_port);
   U172 : AOI22_X1 port map( A1 => A_ns(1), A2 => n397, B1 => A_s(1), B2 => 
                           n398, ZN => n521);
   U173 : OAI221_X1 port map( B1 => n393, B2 => n522, C1 => n392, C2 => n523, A
                           => n524, ZN => O_29_port);
   U174 : AOI22_X1 port map( A1 => A_ns(28), A2 => n397, B1 => A_s(28), B2 => 
                           n398, ZN => n524);
   U175 : INV_X1 port map( A => A_s(27), ZN => n523);
   U176 : INV_X1 port map( A => A_ns(27), ZN => n522);
   U177 : OAI221_X1 port map( B1 => n393, B2 => n525, C1 => n392, C2 => n526, A
                           => n527, ZN => O_28_port);
   U178 : AOI22_X1 port map( A1 => A_ns(27), A2 => n397, B1 => A_s(27), B2 => 
                           n398, ZN => n527);
   U179 : INV_X1 port map( A => A_s(26), ZN => n526);
   U180 : INV_X1 port map( A => A_ns(26), ZN => n525);
   U181 : OAI221_X1 port map( B1 => n393, B2 => n528, C1 => n392, C2 => n529, A
                           => n530, ZN => O_27_port);
   U182 : AOI22_X1 port map( A1 => A_ns(26), A2 => n397, B1 => A_s(26), B2 => 
                           n398, ZN => n530);
   U183 : INV_X1 port map( A => A_s(25), ZN => n529);
   U184 : INV_X1 port map( A => A_ns(25), ZN => n528);
   U185 : OAI221_X1 port map( B1 => n393, B2 => n531, C1 => n392, C2 => n532, A
                           => n533, ZN => O_26_port);
   U186 : AOI22_X1 port map( A1 => A_ns(25), A2 => n397, B1 => A_s(25), B2 => 
                           n398, ZN => n533);
   U187 : INV_X1 port map( A => A_s(24), ZN => n532);
   U188 : INV_X1 port map( A => A_ns(24), ZN => n531);
   U189 : OAI221_X1 port map( B1 => n393, B2 => n534, C1 => n392, C2 => n535, A
                           => n536, ZN => O_25_port);
   U190 : AOI22_X1 port map( A1 => A_ns(24), A2 => n397, B1 => A_s(24), B2 => 
                           n398, ZN => n536);
   U191 : INV_X1 port map( A => A_s(23), ZN => n535);
   U192 : INV_X1 port map( A => A_ns(23), ZN => n534);
   U193 : OAI221_X1 port map( B1 => n393, B2 => n537, C1 => n392, C2 => n538, A
                           => n539, ZN => O_24_port);
   U194 : AOI22_X1 port map( A1 => A_ns(23), A2 => n397, B1 => A_s(23), B2 => 
                           n398, ZN => n539);
   U195 : INV_X1 port map( A => A_s(22), ZN => n538);
   U196 : INV_X1 port map( A => A_ns(22), ZN => n537);
   U197 : OAI221_X1 port map( B1 => n393, B2 => n540, C1 => n392, C2 => n541, A
                           => n542, ZN => O_23_port);
   U198 : AOI22_X1 port map( A1 => A_ns(22), A2 => n397, B1 => A_s(22), B2 => 
                           n398, ZN => n542);
   U199 : INV_X1 port map( A => A_s(21), ZN => n541);
   U200 : INV_X1 port map( A => A_ns(21), ZN => n540);
   U201 : OAI221_X1 port map( B1 => n393, B2 => n543, C1 => n392, C2 => n544, A
                           => n545, ZN => O_22_port);
   U202 : AOI22_X1 port map( A1 => A_ns(21), A2 => n397, B1 => A_s(21), B2 => 
                           n398, ZN => n545);
   U203 : INV_X1 port map( A => A_s(20), ZN => n544);
   U204 : INV_X1 port map( A => A_ns(20), ZN => n543);
   U205 : OAI221_X1 port map( B1 => n393, B2 => n546, C1 => n392, C2 => n547, A
                           => n548, ZN => O_21_port);
   U206 : AOI22_X1 port map( A1 => A_ns(20), A2 => n397, B1 => A_s(20), B2 => 
                           n398, ZN => n548);
   U207 : INV_X1 port map( A => A_s(19), ZN => n547);
   U208 : INV_X1 port map( A => A_ns(19), ZN => n546);
   U209 : OAI221_X1 port map( B1 => n393, B2 => n549, C1 => n392, C2 => n550, A
                           => n551, ZN => O_20_port);
   U210 : AOI22_X1 port map( A1 => A_ns(19), A2 => n397, B1 => A_s(19), B2 => 
                           n398, ZN => n551);
   U211 : INV_X1 port map( A => A_s(18), ZN => n550);
   U212 : INV_X1 port map( A => A_ns(18), ZN => n549);
   U213 : OAI22_X1 port map( A1 => n552, A2 => n520, B1 => n553, B2 => n519, ZN
                           => O_1_port);
   U214 : INV_X1 port map( A => A_ns(0), ZN => n519);
   U215 : INV_X1 port map( A => A_s(0), ZN => n520);
   U216 : OAI221_X1 port map( B1 => n393, B2 => n554, C1 => n392, C2 => n555, A
                           => n556, ZN => O_19_port);
   U217 : AOI22_X1 port map( A1 => A_ns(18), A2 => n397, B1 => A_s(18), B2 => 
                           n398, ZN => n556);
   U218 : INV_X1 port map( A => A_s(17), ZN => n555);
   U219 : INV_X1 port map( A => A_ns(17), ZN => n554);
   U220 : OAI221_X1 port map( B1 => n393, B2 => n557, C1 => n392, C2 => n558, A
                           => n559, ZN => O_18_port);
   U221 : AOI22_X1 port map( A1 => A_ns(17), A2 => n397, B1 => A_s(17), B2 => 
                           n398, ZN => n559);
   U222 : INV_X1 port map( A => A_s(16), ZN => n558);
   U223 : INV_X1 port map( A => A_ns(16), ZN => n557);
   U224 : OAI221_X1 port map( B1 => n393, B2 => n560, C1 => n392, C2 => n561, A
                           => n562, ZN => O_17_port);
   U225 : AOI22_X1 port map( A1 => A_ns(16), A2 => n397, B1 => A_s(16), B2 => 
                           n398, ZN => n562);
   U226 : INV_X1 port map( A => A_s(15), ZN => n561);
   U227 : INV_X1 port map( A => A_ns(15), ZN => n560);
   U228 : OAI221_X1 port map( B1 => n393, B2 => n563, C1 => n392, C2 => n564, A
                           => n565, ZN => O_16_port);
   U229 : AOI22_X1 port map( A1 => A_ns(15), A2 => n397, B1 => A_s(15), B2 => 
                           n398, ZN => n565);
   U230 : INV_X1 port map( A => A_s(14), ZN => n564);
   U231 : INV_X1 port map( A => A_ns(14), ZN => n563);
   U232 : OAI221_X1 port map( B1 => n393, B2 => n566, C1 => n392, C2 => n567, A
                           => n568, ZN => O_15_port);
   U233 : AOI22_X1 port map( A1 => A_ns(14), A2 => n397, B1 => A_s(14), B2 => 
                           n398, ZN => n568);
   U234 : INV_X1 port map( A => A_s(13), ZN => n567);
   U235 : INV_X1 port map( A => A_ns(13), ZN => n566);
   U236 : OAI221_X1 port map( B1 => n393, B2 => n569, C1 => n392, C2 => n570, A
                           => n571, ZN => O_14_port);
   U237 : AOI22_X1 port map( A1 => A_ns(13), A2 => n397, B1 => A_s(13), B2 => 
                           n398, ZN => n571);
   U238 : INV_X1 port map( A => A_s(12), ZN => n570);
   U239 : INV_X1 port map( A => A_ns(12), ZN => n569);
   U240 : OAI221_X1 port map( B1 => n393, B2 => n572, C1 => n392, C2 => n573, A
                           => n574, ZN => O_13_port);
   U241 : AOI22_X1 port map( A1 => A_ns(12), A2 => n397, B1 => A_s(12), B2 => 
                           n398, ZN => n574);
   U242 : INV_X1 port map( A => A_s(11), ZN => n573);
   U243 : INV_X1 port map( A => A_ns(11), ZN => n572);
   U244 : OAI221_X1 port map( B1 => n393, B2 => n575, C1 => n392, C2 => n576, A
                           => n577, ZN => O_12_port);
   U245 : AOI22_X1 port map( A1 => A_ns(11), A2 => n397, B1 => A_s(11), B2 => 
                           n398, ZN => n577);
   U246 : INV_X1 port map( A => A_s(10), ZN => n576);
   U247 : INV_X1 port map( A => A_ns(10), ZN => n575);
   U248 : OAI221_X1 port map( B1 => n393, B2 => n578, C1 => n392, C2 => n579, A
                           => n580, ZN => O_11_port);
   U249 : AOI22_X1 port map( A1 => A_ns(10), A2 => n397, B1 => A_s(10), B2 => 
                           n398, ZN => n580);
   U250 : INV_X1 port map( A => A_s(9), ZN => n579);
   U251 : INV_X1 port map( A => A_ns(9), ZN => n578);
   U252 : OAI221_X1 port map( B1 => n581, B2 => n393, C1 => n582, C2 => n392, A
                           => n583, ZN => O_10_port);
   U253 : AOI22_X1 port map( A1 => A_ns(9), A2 => n397, B1 => A_s(9), B2 => 
                           n398, ZN => n583);
   U254 : NAND2_X1 port map( A1 => n584, A2 => n552, ZN => n553);
   U255 : NAND2_X1 port map( A1 => n584, A2 => n585, ZN => n552);
   U256 : XOR2_X1 port map( A => B(13), B => B(14), Z => n584);
   U257 : INV_X1 port map( A => A_s(8), ZN => n582);
   U258 : INV_X1 port map( A => B(15), ZN => n585);
   U259 : INV_X1 port map( A => A_ns(8), ZN => n581);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity BOOTHENC_NBIT64_i12 is

   port( A, A_n, A_ns, A_s, B : in std_logic_vector (63 downto 0);  O, A_so, 
         A_nso : out std_logic_vector (63 downto 0));

end BOOTHENC_NBIT64_i12;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT64_i12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, O_63_port, O_62_port, O_61_port, O_60_port, O_59_port,
      O_58_port, O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, 
      O_52_port, O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, 
      O_46_port, O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, 
      O_40_port, O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, 
      O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, 
      O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, 
      O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, 
      O_16_port, O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, 
      O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, 
      O_3_port, O_2_port, O_1_port, n391, n392, n393, n394, n395, n396, n397, 
      n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, 
      n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, 
      n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, 
      n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, 
      n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, 
      n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, 
      n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, 
      n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, 
      n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, 
      n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, 
      n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, 
      n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, 
      n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, 
      n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, 
      n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, 
      n578, n579, n580, n581, n582, n583, n584, n585 : std_logic;

begin
   O <= ( O_63_port, O_62_port, O_61_port, O_60_port, O_59_port, O_58_port, 
      O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, O_52_port, 
      O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, O_46_port, 
      O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, O_40_port, 
      O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, 
      O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, 
      O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, 
      O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, O_16_port, 
      O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, O_10_port, 
      O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, O_3_port, 
      O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(61), A_s(60), A_s(59), A_s(58), A_s(57), A_s(56), A_s(55), 
      A_s(54), A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), 
      A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), 
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   A_nso <= ( A_s(61), A_s(60), A_s(59), A_s(58), A_s(57), A_s(56), A_s(55), 
      A_s(54), A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), 
      A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), 
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : AND3_X1 port map( A1 => B(12), A2 => n585, A3 => B(11), ZN => n391);
   U3 : INV_X4 port map( A => n391, ZN => n392);
   U4 : INV_X4 port map( A => n552, ZN => n398);
   U5 : OR3_X4 port map( A1 => B(11), A2 => B(12), A3 => n585, ZN => n393);
   U6 : INV_X4 port map( A => n553, ZN => n397);
   U7 : OAI221_X1 port map( B1 => n393, B2 => n394, C1 => n392, C2 => n395, A 
                           => n396, ZN => O_9_port);
   U8 : AOI22_X1 port map( A1 => A_ns(8), A2 => n397, B1 => A_s(8), B2 => n398,
                           ZN => n396);
   U9 : INV_X1 port map( A => A_s(7), ZN => n395);
   U10 : INV_X1 port map( A => A_ns(7), ZN => n394);
   U11 : OAI221_X1 port map( B1 => n393, B2 => n399, C1 => n392, C2 => n400, A 
                           => n401, ZN => O_8_port);
   U12 : AOI22_X1 port map( A1 => A_ns(7), A2 => n397, B1 => A_s(7), B2 => n398
                           , ZN => n401);
   U13 : INV_X1 port map( A => A_s(6), ZN => n400);
   U14 : INV_X1 port map( A => A_ns(6), ZN => n399);
   U15 : OAI221_X1 port map( B1 => n393, B2 => n402, C1 => n392, C2 => n403, A 
                           => n404, ZN => O_7_port);
   U16 : AOI22_X1 port map( A1 => A_ns(6), A2 => n397, B1 => A_s(6), B2 => n398
                           , ZN => n404);
   U17 : INV_X1 port map( A => A_s(5), ZN => n403);
   U18 : INV_X1 port map( A => A_ns(5), ZN => n402);
   U19 : OAI221_X1 port map( B1 => n393, B2 => n405, C1 => n392, C2 => n406, A 
                           => n407, ZN => O_6_port);
   U20 : AOI22_X1 port map( A1 => A_ns(5), A2 => n397, B1 => A_s(5), B2 => n398
                           , ZN => n407);
   U21 : INV_X1 port map( A => A_s(4), ZN => n406);
   U22 : INV_X1 port map( A => A_ns(4), ZN => n405);
   U23 : OAI221_X1 port map( B1 => n393, B2 => n408, C1 => n392, C2 => n409, A 
                           => n410, ZN => O_63_port);
   U24 : AOI22_X1 port map( A1 => A_ns(62), A2 => n397, B1 => A_s(62), B2 => 
                           n398, ZN => n410);
   U25 : INV_X1 port map( A => A_s(61), ZN => n409);
   U26 : INV_X1 port map( A => A_ns(61), ZN => n408);
   U27 : OAI221_X1 port map( B1 => n393, B2 => n411, C1 => n392, C2 => n412, A 
                           => n413, ZN => O_62_port);
   U28 : AOI22_X1 port map( A1 => A_ns(61), A2 => n397, B1 => A_s(61), B2 => 
                           n398, ZN => n413);
   U29 : INV_X1 port map( A => A_s(60), ZN => n412);
   U30 : INV_X1 port map( A => A_ns(60), ZN => n411);
   U31 : OAI221_X1 port map( B1 => n393, B2 => n414, C1 => n392, C2 => n415, A 
                           => n416, ZN => O_61_port);
   U32 : AOI22_X1 port map( A1 => A_ns(60), A2 => n397, B1 => A_s(60), B2 => 
                           n398, ZN => n416);
   U33 : INV_X1 port map( A => A_s(59), ZN => n415);
   U34 : INV_X1 port map( A => A_ns(59), ZN => n414);
   U35 : OAI221_X1 port map( B1 => n393, B2 => n417, C1 => n392, C2 => n418, A 
                           => n419, ZN => O_60_port);
   U36 : AOI22_X1 port map( A1 => A_ns(59), A2 => n397, B1 => A_s(59), B2 => 
                           n398, ZN => n419);
   U37 : INV_X1 port map( A => A_s(58), ZN => n418);
   U38 : INV_X1 port map( A => A_ns(58), ZN => n417);
   U39 : OAI221_X1 port map( B1 => n393, B2 => n420, C1 => n392, C2 => n421, A 
                           => n422, ZN => O_5_port);
   U40 : AOI22_X1 port map( A1 => A_ns(4), A2 => n397, B1 => A_s(4), B2 => n398
                           , ZN => n422);
   U41 : INV_X1 port map( A => A_s(3), ZN => n421);
   U42 : INV_X1 port map( A => A_ns(3), ZN => n420);
   U43 : OAI221_X1 port map( B1 => n393, B2 => n423, C1 => n392, C2 => n424, A 
                           => n425, ZN => O_59_port);
   U44 : AOI22_X1 port map( A1 => A_ns(58), A2 => n397, B1 => A_s(58), B2 => 
                           n398, ZN => n425);
   U45 : INV_X1 port map( A => A_s(57), ZN => n424);
   U46 : INV_X1 port map( A => A_ns(57), ZN => n423);
   U47 : OAI221_X1 port map( B1 => n393, B2 => n426, C1 => n392, C2 => n427, A 
                           => n428, ZN => O_58_port);
   U48 : AOI22_X1 port map( A1 => A_ns(57), A2 => n397, B1 => A_s(57), B2 => 
                           n398, ZN => n428);
   U49 : INV_X1 port map( A => A_s(56), ZN => n427);
   U50 : INV_X1 port map( A => A_ns(56), ZN => n426);
   U51 : OAI221_X1 port map( B1 => n393, B2 => n429, C1 => n392, C2 => n430, A 
                           => n431, ZN => O_57_port);
   U52 : AOI22_X1 port map( A1 => A_ns(56), A2 => n397, B1 => A_s(56), B2 => 
                           n398, ZN => n431);
   U53 : INV_X1 port map( A => A_s(55), ZN => n430);
   U54 : INV_X1 port map( A => A_ns(55), ZN => n429);
   U55 : OAI221_X1 port map( B1 => n393, B2 => n432, C1 => n392, C2 => n433, A 
                           => n434, ZN => O_56_port);
   U56 : AOI22_X1 port map( A1 => A_ns(55), A2 => n397, B1 => A_s(55), B2 => 
                           n398, ZN => n434);
   U57 : INV_X1 port map( A => A_s(54), ZN => n433);
   U58 : INV_X1 port map( A => A_ns(54), ZN => n432);
   U59 : OAI221_X1 port map( B1 => n393, B2 => n435, C1 => n392, C2 => n436, A 
                           => n437, ZN => O_55_port);
   U60 : AOI22_X1 port map( A1 => A_ns(54), A2 => n397, B1 => A_s(54), B2 => 
                           n398, ZN => n437);
   U61 : INV_X1 port map( A => A_s(53), ZN => n436);
   U62 : INV_X1 port map( A => A_ns(53), ZN => n435);
   U63 : OAI221_X1 port map( B1 => n393, B2 => n438, C1 => n392, C2 => n439, A 
                           => n440, ZN => O_54_port);
   U64 : AOI22_X1 port map( A1 => A_ns(53), A2 => n397, B1 => A_s(53), B2 => 
                           n398, ZN => n440);
   U65 : INV_X1 port map( A => A_s(52), ZN => n439);
   U66 : INV_X1 port map( A => A_ns(52), ZN => n438);
   U67 : OAI221_X1 port map( B1 => n393, B2 => n441, C1 => n392, C2 => n442, A 
                           => n443, ZN => O_53_port);
   U68 : AOI22_X1 port map( A1 => A_ns(52), A2 => n397, B1 => A_s(52), B2 => 
                           n398, ZN => n443);
   U69 : INV_X1 port map( A => A_s(51), ZN => n442);
   U70 : INV_X1 port map( A => A_ns(51), ZN => n441);
   U71 : OAI221_X1 port map( B1 => n393, B2 => n444, C1 => n392, C2 => n445, A 
                           => n446, ZN => O_52_port);
   U72 : AOI22_X1 port map( A1 => A_ns(51), A2 => n397, B1 => A_s(51), B2 => 
                           n398, ZN => n446);
   U73 : INV_X1 port map( A => A_s(50), ZN => n445);
   U74 : INV_X1 port map( A => A_ns(50), ZN => n444);
   U75 : OAI221_X1 port map( B1 => n393, B2 => n447, C1 => n392, C2 => n448, A 
                           => n449, ZN => O_51_port);
   U76 : AOI22_X1 port map( A1 => A_ns(50), A2 => n397, B1 => A_s(50), B2 => 
                           n398, ZN => n449);
   U77 : INV_X1 port map( A => A_s(49), ZN => n448);
   U78 : INV_X1 port map( A => A_ns(49), ZN => n447);
   U79 : OAI221_X1 port map( B1 => n393, B2 => n450, C1 => n392, C2 => n451, A 
                           => n452, ZN => O_50_port);
   U80 : AOI22_X1 port map( A1 => A_ns(49), A2 => n397, B1 => A_s(49), B2 => 
                           n398, ZN => n452);
   U81 : INV_X1 port map( A => A_s(48), ZN => n451);
   U82 : INV_X1 port map( A => A_ns(48), ZN => n450);
   U83 : OAI221_X1 port map( B1 => n393, B2 => n453, C1 => n392, C2 => n454, A 
                           => n455, ZN => O_4_port);
   U84 : AOI22_X1 port map( A1 => A_ns(3), A2 => n397, B1 => A_s(3), B2 => n398
                           , ZN => n455);
   U85 : INV_X1 port map( A => A_s(2), ZN => n454);
   U86 : INV_X1 port map( A => A_ns(2), ZN => n453);
   U87 : OAI221_X1 port map( B1 => n393, B2 => n456, C1 => n392, C2 => n457, A 
                           => n458, ZN => O_49_port);
   U88 : AOI22_X1 port map( A1 => A_ns(48), A2 => n397, B1 => A_s(48), B2 => 
                           n398, ZN => n458);
   U89 : INV_X1 port map( A => A_s(47), ZN => n457);
   U90 : INV_X1 port map( A => A_ns(47), ZN => n456);
   U91 : OAI221_X1 port map( B1 => n393, B2 => n459, C1 => n392, C2 => n460, A 
                           => n461, ZN => O_48_port);
   U92 : AOI22_X1 port map( A1 => A_ns(47), A2 => n397, B1 => A_s(47), B2 => 
                           n398, ZN => n461);
   U93 : INV_X1 port map( A => A_s(46), ZN => n460);
   U94 : INV_X1 port map( A => A_ns(46), ZN => n459);
   U95 : OAI221_X1 port map( B1 => n393, B2 => n462, C1 => n392, C2 => n463, A 
                           => n464, ZN => O_47_port);
   U96 : AOI22_X1 port map( A1 => A_ns(46), A2 => n397, B1 => A_s(46), B2 => 
                           n398, ZN => n464);
   U97 : INV_X1 port map( A => A_s(45), ZN => n463);
   U98 : INV_X1 port map( A => A_ns(45), ZN => n462);
   U99 : OAI221_X1 port map( B1 => n393, B2 => n465, C1 => n392, C2 => n466, A 
                           => n467, ZN => O_46_port);
   U100 : AOI22_X1 port map( A1 => A_ns(45), A2 => n397, B1 => A_s(45), B2 => 
                           n398, ZN => n467);
   U101 : INV_X1 port map( A => A_s(44), ZN => n466);
   U102 : INV_X1 port map( A => A_ns(44), ZN => n465);
   U103 : OAI221_X1 port map( B1 => n393, B2 => n468, C1 => n392, C2 => n469, A
                           => n470, ZN => O_45_port);
   U104 : AOI22_X1 port map( A1 => A_ns(44), A2 => n397, B1 => A_s(44), B2 => 
                           n398, ZN => n470);
   U105 : INV_X1 port map( A => A_s(43), ZN => n469);
   U106 : INV_X1 port map( A => A_ns(43), ZN => n468);
   U107 : OAI221_X1 port map( B1 => n393, B2 => n471, C1 => n392, C2 => n472, A
                           => n473, ZN => O_44_port);
   U108 : AOI22_X1 port map( A1 => A_ns(43), A2 => n397, B1 => A_s(43), B2 => 
                           n398, ZN => n473);
   U109 : INV_X1 port map( A => A_s(42), ZN => n472);
   U110 : INV_X1 port map( A => A_ns(42), ZN => n471);
   U111 : OAI221_X1 port map( B1 => n393, B2 => n474, C1 => n392, C2 => n475, A
                           => n476, ZN => O_43_port);
   U112 : AOI22_X1 port map( A1 => A_ns(42), A2 => n397, B1 => A_s(42), B2 => 
                           n398, ZN => n476);
   U113 : INV_X1 port map( A => A_s(41), ZN => n475);
   U114 : INV_X1 port map( A => A_ns(41), ZN => n474);
   U115 : OAI221_X1 port map( B1 => n393, B2 => n477, C1 => n392, C2 => n478, A
                           => n479, ZN => O_42_port);
   U116 : AOI22_X1 port map( A1 => A_ns(41), A2 => n397, B1 => A_s(41), B2 => 
                           n398, ZN => n479);
   U117 : INV_X1 port map( A => A_s(40), ZN => n478);
   U118 : INV_X1 port map( A => A_ns(40), ZN => n477);
   U119 : OAI221_X1 port map( B1 => n393, B2 => n480, C1 => n392, C2 => n481, A
                           => n482, ZN => O_41_port);
   U120 : AOI22_X1 port map( A1 => A_ns(40), A2 => n397, B1 => A_s(40), B2 => 
                           n398, ZN => n482);
   U121 : INV_X1 port map( A => A_s(39), ZN => n481);
   U122 : INV_X1 port map( A => A_ns(39), ZN => n480);
   U123 : OAI221_X1 port map( B1 => n393, B2 => n483, C1 => n392, C2 => n484, A
                           => n485, ZN => O_40_port);
   U124 : AOI22_X1 port map( A1 => A_ns(39), A2 => n397, B1 => A_s(39), B2 => 
                           n398, ZN => n485);
   U125 : INV_X1 port map( A => A_s(38), ZN => n484);
   U126 : INV_X1 port map( A => A_ns(38), ZN => n483);
   U127 : OAI221_X1 port map( B1 => n393, B2 => n486, C1 => n392, C2 => n487, A
                           => n488, ZN => O_3_port);
   U128 : AOI22_X1 port map( A1 => A_ns(2), A2 => n397, B1 => A_s(2), B2 => 
                           n398, ZN => n488);
   U129 : INV_X1 port map( A => A_s(1), ZN => n487);
   U130 : INV_X1 port map( A => A_ns(1), ZN => n486);
   U131 : OAI221_X1 port map( B1 => n393, B2 => n489, C1 => n392, C2 => n490, A
                           => n491, ZN => O_39_port);
   U132 : AOI22_X1 port map( A1 => A_ns(38), A2 => n397, B1 => A_s(38), B2 => 
                           n398, ZN => n491);
   U133 : INV_X1 port map( A => A_s(37), ZN => n490);
   U134 : INV_X1 port map( A => A_ns(37), ZN => n489);
   U135 : OAI221_X1 port map( B1 => n393, B2 => n492, C1 => n392, C2 => n493, A
                           => n494, ZN => O_38_port);
   U136 : AOI22_X1 port map( A1 => A_ns(37), A2 => n397, B1 => A_s(37), B2 => 
                           n398, ZN => n494);
   U137 : INV_X1 port map( A => A_s(36), ZN => n493);
   U138 : INV_X1 port map( A => A_ns(36), ZN => n492);
   U139 : OAI221_X1 port map( B1 => n393, B2 => n495, C1 => n392, C2 => n496, A
                           => n497, ZN => O_37_port);
   U140 : AOI22_X1 port map( A1 => A_ns(36), A2 => n397, B1 => A_s(36), B2 => 
                           n398, ZN => n497);
   U141 : INV_X1 port map( A => A_s(35), ZN => n496);
   U142 : INV_X1 port map( A => A_ns(35), ZN => n495);
   U143 : OAI221_X1 port map( B1 => n393, B2 => n498, C1 => n392, C2 => n499, A
                           => n500, ZN => O_36_port);
   U144 : AOI22_X1 port map( A1 => A_ns(35), A2 => n397, B1 => A_s(35), B2 => 
                           n398, ZN => n500);
   U145 : INV_X1 port map( A => A_s(34), ZN => n499);
   U146 : INV_X1 port map( A => A_ns(34), ZN => n498);
   U147 : OAI221_X1 port map( B1 => n393, B2 => n501, C1 => n392, C2 => n502, A
                           => n503, ZN => O_35_port);
   U148 : AOI22_X1 port map( A1 => A_ns(34), A2 => n397, B1 => A_s(34), B2 => 
                           n398, ZN => n503);
   U149 : INV_X1 port map( A => A_s(33), ZN => n502);
   U150 : INV_X1 port map( A => A_ns(33), ZN => n501);
   U151 : OAI221_X1 port map( B1 => n393, B2 => n504, C1 => n392, C2 => n505, A
                           => n506, ZN => O_34_port);
   U152 : AOI22_X1 port map( A1 => A_ns(33), A2 => n397, B1 => A_s(33), B2 => 
                           n398, ZN => n506);
   U153 : INV_X1 port map( A => A_s(32), ZN => n505);
   U154 : INV_X1 port map( A => A_ns(32), ZN => n504);
   U155 : OAI221_X1 port map( B1 => n393, B2 => n507, C1 => n392, C2 => n508, A
                           => n509, ZN => O_33_port);
   U156 : AOI22_X1 port map( A1 => A_ns(32), A2 => n397, B1 => A_s(32), B2 => 
                           n398, ZN => n509);
   U157 : INV_X1 port map( A => A_s(31), ZN => n508);
   U158 : INV_X1 port map( A => A_ns(31), ZN => n507);
   U159 : OAI221_X1 port map( B1 => n393, B2 => n510, C1 => n392, C2 => n511, A
                           => n512, ZN => O_32_port);
   U160 : AOI22_X1 port map( A1 => A_ns(31), A2 => n397, B1 => A_s(31), B2 => 
                           n398, ZN => n512);
   U161 : INV_X1 port map( A => A_s(30), ZN => n511);
   U162 : INV_X1 port map( A => A_ns(30), ZN => n510);
   U163 : OAI221_X1 port map( B1 => n393, B2 => n513, C1 => n392, C2 => n514, A
                           => n515, ZN => O_31_port);
   U164 : AOI22_X1 port map( A1 => A_ns(30), A2 => n397, B1 => A_s(30), B2 => 
                           n398, ZN => n515);
   U165 : INV_X1 port map( A => A_s(29), ZN => n514);
   U166 : INV_X1 port map( A => A_ns(29), ZN => n513);
   U167 : OAI221_X1 port map( B1 => n393, B2 => n516, C1 => n392, C2 => n517, A
                           => n518, ZN => O_30_port);
   U168 : AOI22_X1 port map( A1 => A_ns(29), A2 => n397, B1 => A_s(29), B2 => 
                           n398, ZN => n518);
   U169 : INV_X1 port map( A => A_s(28), ZN => n517);
   U170 : INV_X1 port map( A => A_ns(28), ZN => n516);
   U171 : OAI221_X1 port map( B1 => n393, B2 => n519, C1 => n392, C2 => n520, A
                           => n521, ZN => O_2_port);
   U172 : AOI22_X1 port map( A1 => A_ns(1), A2 => n397, B1 => A_s(1), B2 => 
                           n398, ZN => n521);
   U173 : OAI221_X1 port map( B1 => n393, B2 => n522, C1 => n392, C2 => n523, A
                           => n524, ZN => O_29_port);
   U174 : AOI22_X1 port map( A1 => A_ns(28), A2 => n397, B1 => A_s(28), B2 => 
                           n398, ZN => n524);
   U175 : INV_X1 port map( A => A_s(27), ZN => n523);
   U176 : INV_X1 port map( A => A_ns(27), ZN => n522);
   U177 : OAI221_X1 port map( B1 => n393, B2 => n525, C1 => n392, C2 => n526, A
                           => n527, ZN => O_28_port);
   U178 : AOI22_X1 port map( A1 => A_ns(27), A2 => n397, B1 => A_s(27), B2 => 
                           n398, ZN => n527);
   U179 : INV_X1 port map( A => A_s(26), ZN => n526);
   U180 : INV_X1 port map( A => A_ns(26), ZN => n525);
   U181 : OAI221_X1 port map( B1 => n393, B2 => n528, C1 => n392, C2 => n529, A
                           => n530, ZN => O_27_port);
   U182 : AOI22_X1 port map( A1 => A_ns(26), A2 => n397, B1 => A_s(26), B2 => 
                           n398, ZN => n530);
   U183 : INV_X1 port map( A => A_s(25), ZN => n529);
   U184 : INV_X1 port map( A => A_ns(25), ZN => n528);
   U185 : OAI221_X1 port map( B1 => n393, B2 => n531, C1 => n392, C2 => n532, A
                           => n533, ZN => O_26_port);
   U186 : AOI22_X1 port map( A1 => A_ns(25), A2 => n397, B1 => A_s(25), B2 => 
                           n398, ZN => n533);
   U187 : INV_X1 port map( A => A_s(24), ZN => n532);
   U188 : INV_X1 port map( A => A_ns(24), ZN => n531);
   U189 : OAI221_X1 port map( B1 => n393, B2 => n534, C1 => n392, C2 => n535, A
                           => n536, ZN => O_25_port);
   U190 : AOI22_X1 port map( A1 => A_ns(24), A2 => n397, B1 => A_s(24), B2 => 
                           n398, ZN => n536);
   U191 : INV_X1 port map( A => A_s(23), ZN => n535);
   U192 : INV_X1 port map( A => A_ns(23), ZN => n534);
   U193 : OAI221_X1 port map( B1 => n393, B2 => n537, C1 => n392, C2 => n538, A
                           => n539, ZN => O_24_port);
   U194 : AOI22_X1 port map( A1 => A_ns(23), A2 => n397, B1 => A_s(23), B2 => 
                           n398, ZN => n539);
   U195 : INV_X1 port map( A => A_s(22), ZN => n538);
   U196 : INV_X1 port map( A => A_ns(22), ZN => n537);
   U197 : OAI221_X1 port map( B1 => n393, B2 => n540, C1 => n392, C2 => n541, A
                           => n542, ZN => O_23_port);
   U198 : AOI22_X1 port map( A1 => A_ns(22), A2 => n397, B1 => A_s(22), B2 => 
                           n398, ZN => n542);
   U199 : INV_X1 port map( A => A_s(21), ZN => n541);
   U200 : INV_X1 port map( A => A_ns(21), ZN => n540);
   U201 : OAI221_X1 port map( B1 => n393, B2 => n543, C1 => n392, C2 => n544, A
                           => n545, ZN => O_22_port);
   U202 : AOI22_X1 port map( A1 => A_ns(21), A2 => n397, B1 => A_s(21), B2 => 
                           n398, ZN => n545);
   U203 : INV_X1 port map( A => A_s(20), ZN => n544);
   U204 : INV_X1 port map( A => A_ns(20), ZN => n543);
   U205 : OAI221_X1 port map( B1 => n393, B2 => n546, C1 => n392, C2 => n547, A
                           => n548, ZN => O_21_port);
   U206 : AOI22_X1 port map( A1 => A_ns(20), A2 => n397, B1 => A_s(20), B2 => 
                           n398, ZN => n548);
   U207 : INV_X1 port map( A => A_s(19), ZN => n547);
   U208 : INV_X1 port map( A => A_ns(19), ZN => n546);
   U209 : OAI221_X1 port map( B1 => n393, B2 => n549, C1 => n392, C2 => n550, A
                           => n551, ZN => O_20_port);
   U210 : AOI22_X1 port map( A1 => A_ns(19), A2 => n397, B1 => A_s(19), B2 => 
                           n398, ZN => n551);
   U211 : INV_X1 port map( A => A_s(18), ZN => n550);
   U212 : INV_X1 port map( A => A_ns(18), ZN => n549);
   U213 : OAI22_X1 port map( A1 => n552, A2 => n520, B1 => n553, B2 => n519, ZN
                           => O_1_port);
   U214 : INV_X1 port map( A => A_ns(0), ZN => n519);
   U215 : INV_X1 port map( A => A_s(0), ZN => n520);
   U216 : OAI221_X1 port map( B1 => n393, B2 => n554, C1 => n392, C2 => n555, A
                           => n556, ZN => O_19_port);
   U217 : AOI22_X1 port map( A1 => A_ns(18), A2 => n397, B1 => A_s(18), B2 => 
                           n398, ZN => n556);
   U218 : INV_X1 port map( A => A_s(17), ZN => n555);
   U219 : INV_X1 port map( A => A_ns(17), ZN => n554);
   U220 : OAI221_X1 port map( B1 => n393, B2 => n557, C1 => n392, C2 => n558, A
                           => n559, ZN => O_18_port);
   U221 : AOI22_X1 port map( A1 => A_ns(17), A2 => n397, B1 => A_s(17), B2 => 
                           n398, ZN => n559);
   U222 : INV_X1 port map( A => A_s(16), ZN => n558);
   U223 : INV_X1 port map( A => A_ns(16), ZN => n557);
   U224 : OAI221_X1 port map( B1 => n393, B2 => n560, C1 => n392, C2 => n561, A
                           => n562, ZN => O_17_port);
   U225 : AOI22_X1 port map( A1 => A_ns(16), A2 => n397, B1 => A_s(16), B2 => 
                           n398, ZN => n562);
   U226 : INV_X1 port map( A => A_s(15), ZN => n561);
   U227 : INV_X1 port map( A => A_ns(15), ZN => n560);
   U228 : OAI221_X1 port map( B1 => n393, B2 => n563, C1 => n392, C2 => n564, A
                           => n565, ZN => O_16_port);
   U229 : AOI22_X1 port map( A1 => A_ns(15), A2 => n397, B1 => A_s(15), B2 => 
                           n398, ZN => n565);
   U230 : INV_X1 port map( A => A_s(14), ZN => n564);
   U231 : INV_X1 port map( A => A_ns(14), ZN => n563);
   U232 : OAI221_X1 port map( B1 => n393, B2 => n566, C1 => n392, C2 => n567, A
                           => n568, ZN => O_15_port);
   U233 : AOI22_X1 port map( A1 => A_ns(14), A2 => n397, B1 => A_s(14), B2 => 
                           n398, ZN => n568);
   U234 : INV_X1 port map( A => A_s(13), ZN => n567);
   U235 : INV_X1 port map( A => A_ns(13), ZN => n566);
   U236 : OAI221_X1 port map( B1 => n393, B2 => n569, C1 => n392, C2 => n570, A
                           => n571, ZN => O_14_port);
   U237 : AOI22_X1 port map( A1 => A_ns(13), A2 => n397, B1 => A_s(13), B2 => 
                           n398, ZN => n571);
   U238 : INV_X1 port map( A => A_s(12), ZN => n570);
   U239 : INV_X1 port map( A => A_ns(12), ZN => n569);
   U240 : OAI221_X1 port map( B1 => n393, B2 => n572, C1 => n392, C2 => n573, A
                           => n574, ZN => O_13_port);
   U241 : AOI22_X1 port map( A1 => A_ns(12), A2 => n397, B1 => A_s(12), B2 => 
                           n398, ZN => n574);
   U242 : INV_X1 port map( A => A_s(11), ZN => n573);
   U243 : INV_X1 port map( A => A_ns(11), ZN => n572);
   U244 : OAI221_X1 port map( B1 => n393, B2 => n575, C1 => n392, C2 => n576, A
                           => n577, ZN => O_12_port);
   U245 : AOI22_X1 port map( A1 => A_ns(11), A2 => n397, B1 => A_s(11), B2 => 
                           n398, ZN => n577);
   U246 : INV_X1 port map( A => A_s(10), ZN => n576);
   U247 : INV_X1 port map( A => A_ns(10), ZN => n575);
   U248 : OAI221_X1 port map( B1 => n393, B2 => n578, C1 => n392, C2 => n579, A
                           => n580, ZN => O_11_port);
   U249 : AOI22_X1 port map( A1 => A_ns(10), A2 => n397, B1 => A_s(10), B2 => 
                           n398, ZN => n580);
   U250 : INV_X1 port map( A => A_s(9), ZN => n579);
   U251 : INV_X1 port map( A => A_ns(9), ZN => n578);
   U252 : OAI221_X1 port map( B1 => n581, B2 => n393, C1 => n582, C2 => n392, A
                           => n583, ZN => O_10_port);
   U253 : AOI22_X1 port map( A1 => A_ns(9), A2 => n397, B1 => A_s(9), B2 => 
                           n398, ZN => n583);
   U254 : NAND2_X1 port map( A1 => n584, A2 => n552, ZN => n553);
   U255 : NAND2_X1 port map( A1 => n584, A2 => n585, ZN => n552);
   U256 : XOR2_X1 port map( A => B(11), B => B(12), Z => n584);
   U257 : INV_X1 port map( A => A_s(8), ZN => n582);
   U258 : INV_X1 port map( A => B(13), ZN => n585);
   U259 : INV_X1 port map( A => A_ns(8), ZN => n581);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity BOOTHENC_NBIT64_i10 is

   port( A, A_n, A_ns, A_s, B : in std_logic_vector (63 downto 0);  O, A_so, 
         A_nso : out std_logic_vector (63 downto 0));

end BOOTHENC_NBIT64_i10;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT64_i10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, O_63_port, O_62_port, O_61_port, O_60_port, O_59_port,
      O_58_port, O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, 
      O_52_port, O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, 
      O_46_port, O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, 
      O_40_port, O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, 
      O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, 
      O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, 
      O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, 
      O_16_port, O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, 
      O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, 
      O_3_port, O_2_port, O_1_port, n391, n392, n393, n394, n395, n396, n397, 
      n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, 
      n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, 
      n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, 
      n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, 
      n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, 
      n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, 
      n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, 
      n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, 
      n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, 
      n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, 
      n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, 
      n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, 
      n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, 
      n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, 
      n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, 
      n578, n579, n580, n581, n582, n583, n584, n585 : std_logic;

begin
   O <= ( O_63_port, O_62_port, O_61_port, O_60_port, O_59_port, O_58_port, 
      O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, O_52_port, 
      O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, O_46_port, 
      O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, O_40_port, 
      O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, 
      O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, 
      O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, 
      O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, O_16_port, 
      O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, O_10_port, 
      O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, O_3_port, 
      O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(61), A_s(60), A_s(59), A_s(58), A_s(57), A_s(56), A_s(55), 
      A_s(54), A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), 
      A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), 
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   A_nso <= ( A_s(61), A_s(60), A_s(59), A_s(58), A_s(57), A_s(56), A_s(55), 
      A_s(54), A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), 
      A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), 
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : AND3_X1 port map( A1 => B(9), A2 => n585, A3 => B(10), ZN => n391);
   U3 : INV_X4 port map( A => n391, ZN => n392);
   U4 : INV_X4 port map( A => n552, ZN => n398);
   U5 : OR3_X4 port map( A1 => B(10), A2 => B(9), A3 => n585, ZN => n393);
   U6 : INV_X4 port map( A => n553, ZN => n397);
   U7 : OAI221_X1 port map( B1 => n393, B2 => n394, C1 => n392, C2 => n395, A 
                           => n396, ZN => O_9_port);
   U8 : AOI22_X1 port map( A1 => A_ns(8), A2 => n397, B1 => A_s(8), B2 => n398,
                           ZN => n396);
   U9 : INV_X1 port map( A => A_s(7), ZN => n395);
   U10 : INV_X1 port map( A => A_ns(7), ZN => n394);
   U11 : OAI221_X1 port map( B1 => n393, B2 => n399, C1 => n392, C2 => n400, A 
                           => n401, ZN => O_8_port);
   U12 : AOI22_X1 port map( A1 => A_ns(7), A2 => n397, B1 => A_s(7), B2 => n398
                           , ZN => n401);
   U13 : INV_X1 port map( A => A_s(6), ZN => n400);
   U14 : INV_X1 port map( A => A_ns(6), ZN => n399);
   U15 : OAI221_X1 port map( B1 => n393, B2 => n402, C1 => n392, C2 => n403, A 
                           => n404, ZN => O_7_port);
   U16 : AOI22_X1 port map( A1 => A_ns(6), A2 => n397, B1 => A_s(6), B2 => n398
                           , ZN => n404);
   U17 : INV_X1 port map( A => A_s(5), ZN => n403);
   U18 : INV_X1 port map( A => A_ns(5), ZN => n402);
   U19 : OAI221_X1 port map( B1 => n393, B2 => n405, C1 => n392, C2 => n406, A 
                           => n407, ZN => O_6_port);
   U20 : AOI22_X1 port map( A1 => A_ns(5), A2 => n397, B1 => A_s(5), B2 => n398
                           , ZN => n407);
   U21 : INV_X1 port map( A => A_s(4), ZN => n406);
   U22 : INV_X1 port map( A => A_ns(4), ZN => n405);
   U23 : OAI221_X1 port map( B1 => n393, B2 => n408, C1 => n392, C2 => n409, A 
                           => n410, ZN => O_63_port);
   U24 : AOI22_X1 port map( A1 => A_ns(62), A2 => n397, B1 => A_s(62), B2 => 
                           n398, ZN => n410);
   U25 : INV_X1 port map( A => A_s(61), ZN => n409);
   U26 : INV_X1 port map( A => A_ns(61), ZN => n408);
   U27 : OAI221_X1 port map( B1 => n393, B2 => n411, C1 => n392, C2 => n412, A 
                           => n413, ZN => O_62_port);
   U28 : AOI22_X1 port map( A1 => A_ns(61), A2 => n397, B1 => A_s(61), B2 => 
                           n398, ZN => n413);
   U29 : INV_X1 port map( A => A_s(60), ZN => n412);
   U30 : INV_X1 port map( A => A_ns(60), ZN => n411);
   U31 : OAI221_X1 port map( B1 => n393, B2 => n414, C1 => n392, C2 => n415, A 
                           => n416, ZN => O_61_port);
   U32 : AOI22_X1 port map( A1 => A_ns(60), A2 => n397, B1 => A_s(60), B2 => 
                           n398, ZN => n416);
   U33 : INV_X1 port map( A => A_s(59), ZN => n415);
   U34 : INV_X1 port map( A => A_ns(59), ZN => n414);
   U35 : OAI221_X1 port map( B1 => n393, B2 => n417, C1 => n392, C2 => n418, A 
                           => n419, ZN => O_60_port);
   U36 : AOI22_X1 port map( A1 => A_ns(59), A2 => n397, B1 => A_s(59), B2 => 
                           n398, ZN => n419);
   U37 : INV_X1 port map( A => A_s(58), ZN => n418);
   U38 : INV_X1 port map( A => A_ns(58), ZN => n417);
   U39 : OAI221_X1 port map( B1 => n393, B2 => n420, C1 => n392, C2 => n421, A 
                           => n422, ZN => O_5_port);
   U40 : AOI22_X1 port map( A1 => A_ns(4), A2 => n397, B1 => A_s(4), B2 => n398
                           , ZN => n422);
   U41 : INV_X1 port map( A => A_s(3), ZN => n421);
   U42 : INV_X1 port map( A => A_ns(3), ZN => n420);
   U43 : OAI221_X1 port map( B1 => n393, B2 => n423, C1 => n392, C2 => n424, A 
                           => n425, ZN => O_59_port);
   U44 : AOI22_X1 port map( A1 => A_ns(58), A2 => n397, B1 => A_s(58), B2 => 
                           n398, ZN => n425);
   U45 : INV_X1 port map( A => A_s(57), ZN => n424);
   U46 : INV_X1 port map( A => A_ns(57), ZN => n423);
   U47 : OAI221_X1 port map( B1 => n393, B2 => n426, C1 => n392, C2 => n427, A 
                           => n428, ZN => O_58_port);
   U48 : AOI22_X1 port map( A1 => A_ns(57), A2 => n397, B1 => A_s(57), B2 => 
                           n398, ZN => n428);
   U49 : INV_X1 port map( A => A_s(56), ZN => n427);
   U50 : INV_X1 port map( A => A_ns(56), ZN => n426);
   U51 : OAI221_X1 port map( B1 => n393, B2 => n429, C1 => n392, C2 => n430, A 
                           => n431, ZN => O_57_port);
   U52 : AOI22_X1 port map( A1 => A_ns(56), A2 => n397, B1 => A_s(56), B2 => 
                           n398, ZN => n431);
   U53 : INV_X1 port map( A => A_s(55), ZN => n430);
   U54 : INV_X1 port map( A => A_ns(55), ZN => n429);
   U55 : OAI221_X1 port map( B1 => n393, B2 => n432, C1 => n392, C2 => n433, A 
                           => n434, ZN => O_56_port);
   U56 : AOI22_X1 port map( A1 => A_ns(55), A2 => n397, B1 => A_s(55), B2 => 
                           n398, ZN => n434);
   U57 : INV_X1 port map( A => A_s(54), ZN => n433);
   U58 : INV_X1 port map( A => A_ns(54), ZN => n432);
   U59 : OAI221_X1 port map( B1 => n393, B2 => n435, C1 => n392, C2 => n436, A 
                           => n437, ZN => O_55_port);
   U60 : AOI22_X1 port map( A1 => A_ns(54), A2 => n397, B1 => A_s(54), B2 => 
                           n398, ZN => n437);
   U61 : INV_X1 port map( A => A_s(53), ZN => n436);
   U62 : INV_X1 port map( A => A_ns(53), ZN => n435);
   U63 : OAI221_X1 port map( B1 => n393, B2 => n438, C1 => n392, C2 => n439, A 
                           => n440, ZN => O_54_port);
   U64 : AOI22_X1 port map( A1 => A_ns(53), A2 => n397, B1 => A_s(53), B2 => 
                           n398, ZN => n440);
   U65 : INV_X1 port map( A => A_s(52), ZN => n439);
   U66 : INV_X1 port map( A => A_ns(52), ZN => n438);
   U67 : OAI221_X1 port map( B1 => n393, B2 => n441, C1 => n392, C2 => n442, A 
                           => n443, ZN => O_53_port);
   U68 : AOI22_X1 port map( A1 => A_ns(52), A2 => n397, B1 => A_s(52), B2 => 
                           n398, ZN => n443);
   U69 : INV_X1 port map( A => A_s(51), ZN => n442);
   U70 : INV_X1 port map( A => A_ns(51), ZN => n441);
   U71 : OAI221_X1 port map( B1 => n393, B2 => n444, C1 => n392, C2 => n445, A 
                           => n446, ZN => O_52_port);
   U72 : AOI22_X1 port map( A1 => A_ns(51), A2 => n397, B1 => A_s(51), B2 => 
                           n398, ZN => n446);
   U73 : INV_X1 port map( A => A_s(50), ZN => n445);
   U74 : INV_X1 port map( A => A_ns(50), ZN => n444);
   U75 : OAI221_X1 port map( B1 => n393, B2 => n447, C1 => n392, C2 => n448, A 
                           => n449, ZN => O_51_port);
   U76 : AOI22_X1 port map( A1 => A_ns(50), A2 => n397, B1 => A_s(50), B2 => 
                           n398, ZN => n449);
   U77 : INV_X1 port map( A => A_s(49), ZN => n448);
   U78 : INV_X1 port map( A => A_ns(49), ZN => n447);
   U79 : OAI221_X1 port map( B1 => n393, B2 => n450, C1 => n392, C2 => n451, A 
                           => n452, ZN => O_50_port);
   U80 : AOI22_X1 port map( A1 => A_ns(49), A2 => n397, B1 => A_s(49), B2 => 
                           n398, ZN => n452);
   U81 : INV_X1 port map( A => A_s(48), ZN => n451);
   U82 : INV_X1 port map( A => A_ns(48), ZN => n450);
   U83 : OAI221_X1 port map( B1 => n393, B2 => n453, C1 => n392, C2 => n454, A 
                           => n455, ZN => O_4_port);
   U84 : AOI22_X1 port map( A1 => A_ns(3), A2 => n397, B1 => A_s(3), B2 => n398
                           , ZN => n455);
   U85 : INV_X1 port map( A => A_s(2), ZN => n454);
   U86 : INV_X1 port map( A => A_ns(2), ZN => n453);
   U87 : OAI221_X1 port map( B1 => n393, B2 => n456, C1 => n392, C2 => n457, A 
                           => n458, ZN => O_49_port);
   U88 : AOI22_X1 port map( A1 => A_ns(48), A2 => n397, B1 => A_s(48), B2 => 
                           n398, ZN => n458);
   U89 : INV_X1 port map( A => A_s(47), ZN => n457);
   U90 : INV_X1 port map( A => A_ns(47), ZN => n456);
   U91 : OAI221_X1 port map( B1 => n393, B2 => n459, C1 => n392, C2 => n460, A 
                           => n461, ZN => O_48_port);
   U92 : AOI22_X1 port map( A1 => A_ns(47), A2 => n397, B1 => A_s(47), B2 => 
                           n398, ZN => n461);
   U93 : INV_X1 port map( A => A_s(46), ZN => n460);
   U94 : INV_X1 port map( A => A_ns(46), ZN => n459);
   U95 : OAI221_X1 port map( B1 => n393, B2 => n462, C1 => n392, C2 => n463, A 
                           => n464, ZN => O_47_port);
   U96 : AOI22_X1 port map( A1 => A_ns(46), A2 => n397, B1 => A_s(46), B2 => 
                           n398, ZN => n464);
   U97 : INV_X1 port map( A => A_s(45), ZN => n463);
   U98 : INV_X1 port map( A => A_ns(45), ZN => n462);
   U99 : OAI221_X1 port map( B1 => n393, B2 => n465, C1 => n392, C2 => n466, A 
                           => n467, ZN => O_46_port);
   U100 : AOI22_X1 port map( A1 => A_ns(45), A2 => n397, B1 => A_s(45), B2 => 
                           n398, ZN => n467);
   U101 : INV_X1 port map( A => A_s(44), ZN => n466);
   U102 : INV_X1 port map( A => A_ns(44), ZN => n465);
   U103 : OAI221_X1 port map( B1 => n393, B2 => n468, C1 => n392, C2 => n469, A
                           => n470, ZN => O_45_port);
   U104 : AOI22_X1 port map( A1 => A_ns(44), A2 => n397, B1 => A_s(44), B2 => 
                           n398, ZN => n470);
   U105 : INV_X1 port map( A => A_s(43), ZN => n469);
   U106 : INV_X1 port map( A => A_ns(43), ZN => n468);
   U107 : OAI221_X1 port map( B1 => n393, B2 => n471, C1 => n392, C2 => n472, A
                           => n473, ZN => O_44_port);
   U108 : AOI22_X1 port map( A1 => A_ns(43), A2 => n397, B1 => A_s(43), B2 => 
                           n398, ZN => n473);
   U109 : INV_X1 port map( A => A_s(42), ZN => n472);
   U110 : INV_X1 port map( A => A_ns(42), ZN => n471);
   U111 : OAI221_X1 port map( B1 => n393, B2 => n474, C1 => n392, C2 => n475, A
                           => n476, ZN => O_43_port);
   U112 : AOI22_X1 port map( A1 => A_ns(42), A2 => n397, B1 => A_s(42), B2 => 
                           n398, ZN => n476);
   U113 : INV_X1 port map( A => A_s(41), ZN => n475);
   U114 : INV_X1 port map( A => A_ns(41), ZN => n474);
   U115 : OAI221_X1 port map( B1 => n393, B2 => n477, C1 => n392, C2 => n478, A
                           => n479, ZN => O_42_port);
   U116 : AOI22_X1 port map( A1 => A_ns(41), A2 => n397, B1 => A_s(41), B2 => 
                           n398, ZN => n479);
   U117 : INV_X1 port map( A => A_s(40), ZN => n478);
   U118 : INV_X1 port map( A => A_ns(40), ZN => n477);
   U119 : OAI221_X1 port map( B1 => n393, B2 => n480, C1 => n392, C2 => n481, A
                           => n482, ZN => O_41_port);
   U120 : AOI22_X1 port map( A1 => A_ns(40), A2 => n397, B1 => A_s(40), B2 => 
                           n398, ZN => n482);
   U121 : INV_X1 port map( A => A_s(39), ZN => n481);
   U122 : INV_X1 port map( A => A_ns(39), ZN => n480);
   U123 : OAI221_X1 port map( B1 => n393, B2 => n483, C1 => n392, C2 => n484, A
                           => n485, ZN => O_40_port);
   U124 : AOI22_X1 port map( A1 => A_ns(39), A2 => n397, B1 => A_s(39), B2 => 
                           n398, ZN => n485);
   U125 : INV_X1 port map( A => A_s(38), ZN => n484);
   U126 : INV_X1 port map( A => A_ns(38), ZN => n483);
   U127 : OAI221_X1 port map( B1 => n393, B2 => n486, C1 => n392, C2 => n487, A
                           => n488, ZN => O_3_port);
   U128 : AOI22_X1 port map( A1 => A_ns(2), A2 => n397, B1 => A_s(2), B2 => 
                           n398, ZN => n488);
   U129 : INV_X1 port map( A => A_s(1), ZN => n487);
   U130 : INV_X1 port map( A => A_ns(1), ZN => n486);
   U131 : OAI221_X1 port map( B1 => n393, B2 => n489, C1 => n392, C2 => n490, A
                           => n491, ZN => O_39_port);
   U132 : AOI22_X1 port map( A1 => A_ns(38), A2 => n397, B1 => A_s(38), B2 => 
                           n398, ZN => n491);
   U133 : INV_X1 port map( A => A_s(37), ZN => n490);
   U134 : INV_X1 port map( A => A_ns(37), ZN => n489);
   U135 : OAI221_X1 port map( B1 => n393, B2 => n492, C1 => n392, C2 => n493, A
                           => n494, ZN => O_38_port);
   U136 : AOI22_X1 port map( A1 => A_ns(37), A2 => n397, B1 => A_s(37), B2 => 
                           n398, ZN => n494);
   U137 : INV_X1 port map( A => A_s(36), ZN => n493);
   U138 : INV_X1 port map( A => A_ns(36), ZN => n492);
   U139 : OAI221_X1 port map( B1 => n393, B2 => n495, C1 => n392, C2 => n496, A
                           => n497, ZN => O_37_port);
   U140 : AOI22_X1 port map( A1 => A_ns(36), A2 => n397, B1 => A_s(36), B2 => 
                           n398, ZN => n497);
   U141 : INV_X1 port map( A => A_s(35), ZN => n496);
   U142 : INV_X1 port map( A => A_ns(35), ZN => n495);
   U143 : OAI221_X1 port map( B1 => n393, B2 => n498, C1 => n392, C2 => n499, A
                           => n500, ZN => O_36_port);
   U144 : AOI22_X1 port map( A1 => A_ns(35), A2 => n397, B1 => A_s(35), B2 => 
                           n398, ZN => n500);
   U145 : INV_X1 port map( A => A_s(34), ZN => n499);
   U146 : INV_X1 port map( A => A_ns(34), ZN => n498);
   U147 : OAI221_X1 port map( B1 => n393, B2 => n501, C1 => n392, C2 => n502, A
                           => n503, ZN => O_35_port);
   U148 : AOI22_X1 port map( A1 => A_ns(34), A2 => n397, B1 => A_s(34), B2 => 
                           n398, ZN => n503);
   U149 : INV_X1 port map( A => A_s(33), ZN => n502);
   U150 : INV_X1 port map( A => A_ns(33), ZN => n501);
   U151 : OAI221_X1 port map( B1 => n393, B2 => n504, C1 => n392, C2 => n505, A
                           => n506, ZN => O_34_port);
   U152 : AOI22_X1 port map( A1 => A_ns(33), A2 => n397, B1 => A_s(33), B2 => 
                           n398, ZN => n506);
   U153 : INV_X1 port map( A => A_s(32), ZN => n505);
   U154 : INV_X1 port map( A => A_ns(32), ZN => n504);
   U155 : OAI221_X1 port map( B1 => n393, B2 => n507, C1 => n392, C2 => n508, A
                           => n509, ZN => O_33_port);
   U156 : AOI22_X1 port map( A1 => A_ns(32), A2 => n397, B1 => A_s(32), B2 => 
                           n398, ZN => n509);
   U157 : INV_X1 port map( A => A_s(31), ZN => n508);
   U158 : INV_X1 port map( A => A_ns(31), ZN => n507);
   U159 : OAI221_X1 port map( B1 => n393, B2 => n510, C1 => n392, C2 => n511, A
                           => n512, ZN => O_32_port);
   U160 : AOI22_X1 port map( A1 => A_ns(31), A2 => n397, B1 => A_s(31), B2 => 
                           n398, ZN => n512);
   U161 : INV_X1 port map( A => A_s(30), ZN => n511);
   U162 : INV_X1 port map( A => A_ns(30), ZN => n510);
   U163 : OAI221_X1 port map( B1 => n393, B2 => n513, C1 => n392, C2 => n514, A
                           => n515, ZN => O_31_port);
   U164 : AOI22_X1 port map( A1 => A_ns(30), A2 => n397, B1 => A_s(30), B2 => 
                           n398, ZN => n515);
   U165 : INV_X1 port map( A => A_s(29), ZN => n514);
   U166 : INV_X1 port map( A => A_ns(29), ZN => n513);
   U167 : OAI221_X1 port map( B1 => n393, B2 => n516, C1 => n392, C2 => n517, A
                           => n518, ZN => O_30_port);
   U168 : AOI22_X1 port map( A1 => A_ns(29), A2 => n397, B1 => A_s(29), B2 => 
                           n398, ZN => n518);
   U169 : INV_X1 port map( A => A_s(28), ZN => n517);
   U170 : INV_X1 port map( A => A_ns(28), ZN => n516);
   U171 : OAI221_X1 port map( B1 => n393, B2 => n519, C1 => n392, C2 => n520, A
                           => n521, ZN => O_2_port);
   U172 : AOI22_X1 port map( A1 => A_ns(1), A2 => n397, B1 => A_s(1), B2 => 
                           n398, ZN => n521);
   U173 : OAI221_X1 port map( B1 => n393, B2 => n522, C1 => n392, C2 => n523, A
                           => n524, ZN => O_29_port);
   U174 : AOI22_X1 port map( A1 => A_ns(28), A2 => n397, B1 => A_s(28), B2 => 
                           n398, ZN => n524);
   U175 : INV_X1 port map( A => A_s(27), ZN => n523);
   U176 : INV_X1 port map( A => A_ns(27), ZN => n522);
   U177 : OAI221_X1 port map( B1 => n393, B2 => n525, C1 => n392, C2 => n526, A
                           => n527, ZN => O_28_port);
   U178 : AOI22_X1 port map( A1 => A_ns(27), A2 => n397, B1 => A_s(27), B2 => 
                           n398, ZN => n527);
   U179 : INV_X1 port map( A => A_s(26), ZN => n526);
   U180 : INV_X1 port map( A => A_ns(26), ZN => n525);
   U181 : OAI221_X1 port map( B1 => n393, B2 => n528, C1 => n392, C2 => n529, A
                           => n530, ZN => O_27_port);
   U182 : AOI22_X1 port map( A1 => A_ns(26), A2 => n397, B1 => A_s(26), B2 => 
                           n398, ZN => n530);
   U183 : INV_X1 port map( A => A_s(25), ZN => n529);
   U184 : INV_X1 port map( A => A_ns(25), ZN => n528);
   U185 : OAI221_X1 port map( B1 => n393, B2 => n531, C1 => n392, C2 => n532, A
                           => n533, ZN => O_26_port);
   U186 : AOI22_X1 port map( A1 => A_ns(25), A2 => n397, B1 => A_s(25), B2 => 
                           n398, ZN => n533);
   U187 : INV_X1 port map( A => A_s(24), ZN => n532);
   U188 : INV_X1 port map( A => A_ns(24), ZN => n531);
   U189 : OAI221_X1 port map( B1 => n393, B2 => n534, C1 => n392, C2 => n535, A
                           => n536, ZN => O_25_port);
   U190 : AOI22_X1 port map( A1 => A_ns(24), A2 => n397, B1 => A_s(24), B2 => 
                           n398, ZN => n536);
   U191 : INV_X1 port map( A => A_s(23), ZN => n535);
   U192 : INV_X1 port map( A => A_ns(23), ZN => n534);
   U193 : OAI221_X1 port map( B1 => n393, B2 => n537, C1 => n392, C2 => n538, A
                           => n539, ZN => O_24_port);
   U194 : AOI22_X1 port map( A1 => A_ns(23), A2 => n397, B1 => A_s(23), B2 => 
                           n398, ZN => n539);
   U195 : INV_X1 port map( A => A_s(22), ZN => n538);
   U196 : INV_X1 port map( A => A_ns(22), ZN => n537);
   U197 : OAI221_X1 port map( B1 => n393, B2 => n540, C1 => n392, C2 => n541, A
                           => n542, ZN => O_23_port);
   U198 : AOI22_X1 port map( A1 => A_ns(22), A2 => n397, B1 => A_s(22), B2 => 
                           n398, ZN => n542);
   U199 : INV_X1 port map( A => A_s(21), ZN => n541);
   U200 : INV_X1 port map( A => A_ns(21), ZN => n540);
   U201 : OAI221_X1 port map( B1 => n393, B2 => n543, C1 => n392, C2 => n544, A
                           => n545, ZN => O_22_port);
   U202 : AOI22_X1 port map( A1 => A_ns(21), A2 => n397, B1 => A_s(21), B2 => 
                           n398, ZN => n545);
   U203 : INV_X1 port map( A => A_s(20), ZN => n544);
   U204 : INV_X1 port map( A => A_ns(20), ZN => n543);
   U205 : OAI221_X1 port map( B1 => n393, B2 => n546, C1 => n392, C2 => n547, A
                           => n548, ZN => O_21_port);
   U206 : AOI22_X1 port map( A1 => A_ns(20), A2 => n397, B1 => A_s(20), B2 => 
                           n398, ZN => n548);
   U207 : INV_X1 port map( A => A_s(19), ZN => n547);
   U208 : INV_X1 port map( A => A_ns(19), ZN => n546);
   U209 : OAI221_X1 port map( B1 => n393, B2 => n549, C1 => n392, C2 => n550, A
                           => n551, ZN => O_20_port);
   U210 : AOI22_X1 port map( A1 => A_ns(19), A2 => n397, B1 => A_s(19), B2 => 
                           n398, ZN => n551);
   U211 : INV_X1 port map( A => A_s(18), ZN => n550);
   U212 : INV_X1 port map( A => A_ns(18), ZN => n549);
   U213 : OAI22_X1 port map( A1 => n552, A2 => n520, B1 => n553, B2 => n519, ZN
                           => O_1_port);
   U214 : INV_X1 port map( A => A_ns(0), ZN => n519);
   U215 : INV_X1 port map( A => A_s(0), ZN => n520);
   U216 : OAI221_X1 port map( B1 => n393, B2 => n554, C1 => n392, C2 => n555, A
                           => n556, ZN => O_19_port);
   U217 : AOI22_X1 port map( A1 => A_ns(18), A2 => n397, B1 => A_s(18), B2 => 
                           n398, ZN => n556);
   U218 : INV_X1 port map( A => A_s(17), ZN => n555);
   U219 : INV_X1 port map( A => A_ns(17), ZN => n554);
   U220 : OAI221_X1 port map( B1 => n393, B2 => n557, C1 => n392, C2 => n558, A
                           => n559, ZN => O_18_port);
   U221 : AOI22_X1 port map( A1 => A_ns(17), A2 => n397, B1 => A_s(17), B2 => 
                           n398, ZN => n559);
   U222 : INV_X1 port map( A => A_s(16), ZN => n558);
   U223 : INV_X1 port map( A => A_ns(16), ZN => n557);
   U224 : OAI221_X1 port map( B1 => n393, B2 => n560, C1 => n392, C2 => n561, A
                           => n562, ZN => O_17_port);
   U225 : AOI22_X1 port map( A1 => A_ns(16), A2 => n397, B1 => A_s(16), B2 => 
                           n398, ZN => n562);
   U226 : INV_X1 port map( A => A_s(15), ZN => n561);
   U227 : INV_X1 port map( A => A_ns(15), ZN => n560);
   U228 : OAI221_X1 port map( B1 => n393, B2 => n563, C1 => n392, C2 => n564, A
                           => n565, ZN => O_16_port);
   U229 : AOI22_X1 port map( A1 => A_ns(15), A2 => n397, B1 => A_s(15), B2 => 
                           n398, ZN => n565);
   U230 : INV_X1 port map( A => A_s(14), ZN => n564);
   U231 : INV_X1 port map( A => A_ns(14), ZN => n563);
   U232 : OAI221_X1 port map( B1 => n393, B2 => n566, C1 => n392, C2 => n567, A
                           => n568, ZN => O_15_port);
   U233 : AOI22_X1 port map( A1 => A_ns(14), A2 => n397, B1 => A_s(14), B2 => 
                           n398, ZN => n568);
   U234 : INV_X1 port map( A => A_s(13), ZN => n567);
   U235 : INV_X1 port map( A => A_ns(13), ZN => n566);
   U236 : OAI221_X1 port map( B1 => n393, B2 => n569, C1 => n392, C2 => n570, A
                           => n571, ZN => O_14_port);
   U237 : AOI22_X1 port map( A1 => A_ns(13), A2 => n397, B1 => A_s(13), B2 => 
                           n398, ZN => n571);
   U238 : INV_X1 port map( A => A_s(12), ZN => n570);
   U239 : INV_X1 port map( A => A_ns(12), ZN => n569);
   U240 : OAI221_X1 port map( B1 => n393, B2 => n572, C1 => n392, C2 => n573, A
                           => n574, ZN => O_13_port);
   U241 : AOI22_X1 port map( A1 => A_ns(12), A2 => n397, B1 => A_s(12), B2 => 
                           n398, ZN => n574);
   U242 : INV_X1 port map( A => A_s(11), ZN => n573);
   U243 : INV_X1 port map( A => A_ns(11), ZN => n572);
   U244 : OAI221_X1 port map( B1 => n393, B2 => n575, C1 => n392, C2 => n576, A
                           => n577, ZN => O_12_port);
   U245 : AOI22_X1 port map( A1 => A_ns(11), A2 => n397, B1 => A_s(11), B2 => 
                           n398, ZN => n577);
   U246 : INV_X1 port map( A => A_s(10), ZN => n576);
   U247 : INV_X1 port map( A => A_ns(10), ZN => n575);
   U248 : OAI221_X1 port map( B1 => n393, B2 => n578, C1 => n392, C2 => n579, A
                           => n580, ZN => O_11_port);
   U249 : AOI22_X1 port map( A1 => A_ns(10), A2 => n397, B1 => A_s(10), B2 => 
                           n398, ZN => n580);
   U250 : INV_X1 port map( A => A_s(9), ZN => n579);
   U251 : INV_X1 port map( A => A_ns(9), ZN => n578);
   U252 : OAI221_X1 port map( B1 => n581, B2 => n393, C1 => n582, C2 => n392, A
                           => n583, ZN => O_10_port);
   U253 : AOI22_X1 port map( A1 => A_ns(9), A2 => n397, B1 => A_s(9), B2 => 
                           n398, ZN => n583);
   U254 : NAND2_X1 port map( A1 => n584, A2 => n552, ZN => n553);
   U255 : NAND2_X1 port map( A1 => n584, A2 => n585, ZN => n552);
   U256 : XOR2_X1 port map( A => B(10), B => B(9), Z => n584);
   U257 : INV_X1 port map( A => A_s(8), ZN => n582);
   U258 : INV_X1 port map( A => B(11), ZN => n585);
   U259 : INV_X1 port map( A => A_ns(8), ZN => n581);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity BOOTHENC_NBIT64_i8 is

   port( A, A_n, A_ns, A_s, B : in std_logic_vector (63 downto 0);  O, A_so, 
         A_nso : out std_logic_vector (63 downto 0));

end BOOTHENC_NBIT64_i8;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT64_i8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, O_63_port, O_62_port, O_61_port, O_60_port, O_59_port,
      O_58_port, O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, 
      O_52_port, O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, 
      O_46_port, O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, 
      O_40_port, O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, 
      O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, 
      O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, 
      O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, 
      O_16_port, O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, 
      O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, 
      O_3_port, O_2_port, O_1_port, n391, n392, n393, n394, n395, n396, n397, 
      n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, 
      n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, 
      n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, 
      n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, 
      n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, 
      n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, 
      n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, 
      n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, 
      n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, 
      n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, 
      n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, 
      n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, 
      n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, 
      n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, 
      n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, 
      n578, n579, n580, n581, n582, n583, n584, n585 : std_logic;

begin
   O <= ( O_63_port, O_62_port, O_61_port, O_60_port, O_59_port, O_58_port, 
      O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, O_52_port, 
      O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, O_46_port, 
      O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, O_40_port, 
      O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, 
      O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, 
      O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, 
      O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, O_16_port, 
      O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, O_10_port, 
      O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, O_3_port, 
      O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(61), A_s(60), A_s(59), A_s(58), A_s(57), A_s(56), A_s(55), 
      A_s(54), A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), 
      A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), 
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   A_nso <= ( A_s(61), A_s(60), A_s(59), A_s(58), A_s(57), A_s(56), A_s(55), 
      A_s(54), A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), 
      A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), 
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : AND3_X1 port map( A1 => B(8), A2 => n585, A3 => B(7), ZN => n391);
   U3 : INV_X4 port map( A => n391, ZN => n392);
   U4 : INV_X4 port map( A => n552, ZN => n398);
   U5 : OR3_X4 port map( A1 => B(7), A2 => B(8), A3 => n585, ZN => n393);
   U6 : INV_X4 port map( A => n553, ZN => n397);
   U7 : OAI221_X1 port map( B1 => n393, B2 => n394, C1 => n392, C2 => n395, A 
                           => n396, ZN => O_9_port);
   U8 : AOI22_X1 port map( A1 => A_ns(8), A2 => n397, B1 => A_s(8), B2 => n398,
                           ZN => n396);
   U9 : INV_X1 port map( A => A_s(7), ZN => n395);
   U10 : INV_X1 port map( A => A_ns(7), ZN => n394);
   U11 : OAI221_X1 port map( B1 => n393, B2 => n399, C1 => n392, C2 => n400, A 
                           => n401, ZN => O_8_port);
   U12 : AOI22_X1 port map( A1 => A_ns(7), A2 => n397, B1 => A_s(7), B2 => n398
                           , ZN => n401);
   U13 : INV_X1 port map( A => A_s(6), ZN => n400);
   U14 : INV_X1 port map( A => A_ns(6), ZN => n399);
   U15 : OAI221_X1 port map( B1 => n393, B2 => n402, C1 => n392, C2 => n403, A 
                           => n404, ZN => O_7_port);
   U16 : AOI22_X1 port map( A1 => A_ns(6), A2 => n397, B1 => A_s(6), B2 => n398
                           , ZN => n404);
   U17 : INV_X1 port map( A => A_s(5), ZN => n403);
   U18 : INV_X1 port map( A => A_ns(5), ZN => n402);
   U19 : OAI221_X1 port map( B1 => n393, B2 => n405, C1 => n392, C2 => n406, A 
                           => n407, ZN => O_6_port);
   U20 : AOI22_X1 port map( A1 => A_ns(5), A2 => n397, B1 => A_s(5), B2 => n398
                           , ZN => n407);
   U21 : INV_X1 port map( A => A_s(4), ZN => n406);
   U22 : INV_X1 port map( A => A_ns(4), ZN => n405);
   U23 : OAI221_X1 port map( B1 => n393, B2 => n408, C1 => n392, C2 => n409, A 
                           => n410, ZN => O_63_port);
   U24 : AOI22_X1 port map( A1 => A_ns(62), A2 => n397, B1 => A_s(62), B2 => 
                           n398, ZN => n410);
   U25 : INV_X1 port map( A => A_s(61), ZN => n409);
   U26 : INV_X1 port map( A => A_ns(61), ZN => n408);
   U27 : OAI221_X1 port map( B1 => n393, B2 => n411, C1 => n392, C2 => n412, A 
                           => n413, ZN => O_62_port);
   U28 : AOI22_X1 port map( A1 => A_ns(61), A2 => n397, B1 => A_s(61), B2 => 
                           n398, ZN => n413);
   U29 : INV_X1 port map( A => A_s(60), ZN => n412);
   U30 : INV_X1 port map( A => A_ns(60), ZN => n411);
   U31 : OAI221_X1 port map( B1 => n393, B2 => n414, C1 => n392, C2 => n415, A 
                           => n416, ZN => O_61_port);
   U32 : AOI22_X1 port map( A1 => A_ns(60), A2 => n397, B1 => A_s(60), B2 => 
                           n398, ZN => n416);
   U33 : INV_X1 port map( A => A_s(59), ZN => n415);
   U34 : INV_X1 port map( A => A_ns(59), ZN => n414);
   U35 : OAI221_X1 port map( B1 => n393, B2 => n417, C1 => n392, C2 => n418, A 
                           => n419, ZN => O_60_port);
   U36 : AOI22_X1 port map( A1 => A_ns(59), A2 => n397, B1 => A_s(59), B2 => 
                           n398, ZN => n419);
   U37 : INV_X1 port map( A => A_s(58), ZN => n418);
   U38 : INV_X1 port map( A => A_ns(58), ZN => n417);
   U39 : OAI221_X1 port map( B1 => n393, B2 => n420, C1 => n392, C2 => n421, A 
                           => n422, ZN => O_5_port);
   U40 : AOI22_X1 port map( A1 => A_ns(4), A2 => n397, B1 => A_s(4), B2 => n398
                           , ZN => n422);
   U41 : INV_X1 port map( A => A_s(3), ZN => n421);
   U42 : INV_X1 port map( A => A_ns(3), ZN => n420);
   U43 : OAI221_X1 port map( B1 => n393, B2 => n423, C1 => n392, C2 => n424, A 
                           => n425, ZN => O_59_port);
   U44 : AOI22_X1 port map( A1 => A_ns(58), A2 => n397, B1 => A_s(58), B2 => 
                           n398, ZN => n425);
   U45 : INV_X1 port map( A => A_s(57), ZN => n424);
   U46 : INV_X1 port map( A => A_ns(57), ZN => n423);
   U47 : OAI221_X1 port map( B1 => n393, B2 => n426, C1 => n392, C2 => n427, A 
                           => n428, ZN => O_58_port);
   U48 : AOI22_X1 port map( A1 => A_ns(57), A2 => n397, B1 => A_s(57), B2 => 
                           n398, ZN => n428);
   U49 : INV_X1 port map( A => A_s(56), ZN => n427);
   U50 : INV_X1 port map( A => A_ns(56), ZN => n426);
   U51 : OAI221_X1 port map( B1 => n393, B2 => n429, C1 => n392, C2 => n430, A 
                           => n431, ZN => O_57_port);
   U52 : AOI22_X1 port map( A1 => A_ns(56), A2 => n397, B1 => A_s(56), B2 => 
                           n398, ZN => n431);
   U53 : INV_X1 port map( A => A_s(55), ZN => n430);
   U54 : INV_X1 port map( A => A_ns(55), ZN => n429);
   U55 : OAI221_X1 port map( B1 => n393, B2 => n432, C1 => n392, C2 => n433, A 
                           => n434, ZN => O_56_port);
   U56 : AOI22_X1 port map( A1 => A_ns(55), A2 => n397, B1 => A_s(55), B2 => 
                           n398, ZN => n434);
   U57 : INV_X1 port map( A => A_s(54), ZN => n433);
   U58 : INV_X1 port map( A => A_ns(54), ZN => n432);
   U59 : OAI221_X1 port map( B1 => n393, B2 => n435, C1 => n392, C2 => n436, A 
                           => n437, ZN => O_55_port);
   U60 : AOI22_X1 port map( A1 => A_ns(54), A2 => n397, B1 => A_s(54), B2 => 
                           n398, ZN => n437);
   U61 : INV_X1 port map( A => A_s(53), ZN => n436);
   U62 : INV_X1 port map( A => A_ns(53), ZN => n435);
   U63 : OAI221_X1 port map( B1 => n393, B2 => n438, C1 => n392, C2 => n439, A 
                           => n440, ZN => O_54_port);
   U64 : AOI22_X1 port map( A1 => A_ns(53), A2 => n397, B1 => A_s(53), B2 => 
                           n398, ZN => n440);
   U65 : INV_X1 port map( A => A_s(52), ZN => n439);
   U66 : INV_X1 port map( A => A_ns(52), ZN => n438);
   U67 : OAI221_X1 port map( B1 => n393, B2 => n441, C1 => n392, C2 => n442, A 
                           => n443, ZN => O_53_port);
   U68 : AOI22_X1 port map( A1 => A_ns(52), A2 => n397, B1 => A_s(52), B2 => 
                           n398, ZN => n443);
   U69 : INV_X1 port map( A => A_s(51), ZN => n442);
   U70 : INV_X1 port map( A => A_ns(51), ZN => n441);
   U71 : OAI221_X1 port map( B1 => n393, B2 => n444, C1 => n392, C2 => n445, A 
                           => n446, ZN => O_52_port);
   U72 : AOI22_X1 port map( A1 => A_ns(51), A2 => n397, B1 => A_s(51), B2 => 
                           n398, ZN => n446);
   U73 : INV_X1 port map( A => A_s(50), ZN => n445);
   U74 : INV_X1 port map( A => A_ns(50), ZN => n444);
   U75 : OAI221_X1 port map( B1 => n393, B2 => n447, C1 => n392, C2 => n448, A 
                           => n449, ZN => O_51_port);
   U76 : AOI22_X1 port map( A1 => A_ns(50), A2 => n397, B1 => A_s(50), B2 => 
                           n398, ZN => n449);
   U77 : INV_X1 port map( A => A_s(49), ZN => n448);
   U78 : INV_X1 port map( A => A_ns(49), ZN => n447);
   U79 : OAI221_X1 port map( B1 => n393, B2 => n450, C1 => n392, C2 => n451, A 
                           => n452, ZN => O_50_port);
   U80 : AOI22_X1 port map( A1 => A_ns(49), A2 => n397, B1 => A_s(49), B2 => 
                           n398, ZN => n452);
   U81 : INV_X1 port map( A => A_s(48), ZN => n451);
   U82 : INV_X1 port map( A => A_ns(48), ZN => n450);
   U83 : OAI221_X1 port map( B1 => n393, B2 => n453, C1 => n392, C2 => n454, A 
                           => n455, ZN => O_4_port);
   U84 : AOI22_X1 port map( A1 => A_ns(3), A2 => n397, B1 => A_s(3), B2 => n398
                           , ZN => n455);
   U85 : INV_X1 port map( A => A_s(2), ZN => n454);
   U86 : INV_X1 port map( A => A_ns(2), ZN => n453);
   U87 : OAI221_X1 port map( B1 => n393, B2 => n456, C1 => n392, C2 => n457, A 
                           => n458, ZN => O_49_port);
   U88 : AOI22_X1 port map( A1 => A_ns(48), A2 => n397, B1 => A_s(48), B2 => 
                           n398, ZN => n458);
   U89 : INV_X1 port map( A => A_s(47), ZN => n457);
   U90 : INV_X1 port map( A => A_ns(47), ZN => n456);
   U91 : OAI221_X1 port map( B1 => n393, B2 => n459, C1 => n392, C2 => n460, A 
                           => n461, ZN => O_48_port);
   U92 : AOI22_X1 port map( A1 => A_ns(47), A2 => n397, B1 => A_s(47), B2 => 
                           n398, ZN => n461);
   U93 : INV_X1 port map( A => A_s(46), ZN => n460);
   U94 : INV_X1 port map( A => A_ns(46), ZN => n459);
   U95 : OAI221_X1 port map( B1 => n393, B2 => n462, C1 => n392, C2 => n463, A 
                           => n464, ZN => O_47_port);
   U96 : AOI22_X1 port map( A1 => A_ns(46), A2 => n397, B1 => A_s(46), B2 => 
                           n398, ZN => n464);
   U97 : INV_X1 port map( A => A_s(45), ZN => n463);
   U98 : INV_X1 port map( A => A_ns(45), ZN => n462);
   U99 : OAI221_X1 port map( B1 => n393, B2 => n465, C1 => n392, C2 => n466, A 
                           => n467, ZN => O_46_port);
   U100 : AOI22_X1 port map( A1 => A_ns(45), A2 => n397, B1 => A_s(45), B2 => 
                           n398, ZN => n467);
   U101 : INV_X1 port map( A => A_s(44), ZN => n466);
   U102 : INV_X1 port map( A => A_ns(44), ZN => n465);
   U103 : OAI221_X1 port map( B1 => n393, B2 => n468, C1 => n392, C2 => n469, A
                           => n470, ZN => O_45_port);
   U104 : AOI22_X1 port map( A1 => A_ns(44), A2 => n397, B1 => A_s(44), B2 => 
                           n398, ZN => n470);
   U105 : INV_X1 port map( A => A_s(43), ZN => n469);
   U106 : INV_X1 port map( A => A_ns(43), ZN => n468);
   U107 : OAI221_X1 port map( B1 => n393, B2 => n471, C1 => n392, C2 => n472, A
                           => n473, ZN => O_44_port);
   U108 : AOI22_X1 port map( A1 => A_ns(43), A2 => n397, B1 => A_s(43), B2 => 
                           n398, ZN => n473);
   U109 : INV_X1 port map( A => A_s(42), ZN => n472);
   U110 : INV_X1 port map( A => A_ns(42), ZN => n471);
   U111 : OAI221_X1 port map( B1 => n393, B2 => n474, C1 => n392, C2 => n475, A
                           => n476, ZN => O_43_port);
   U112 : AOI22_X1 port map( A1 => A_ns(42), A2 => n397, B1 => A_s(42), B2 => 
                           n398, ZN => n476);
   U113 : INV_X1 port map( A => A_s(41), ZN => n475);
   U114 : INV_X1 port map( A => A_ns(41), ZN => n474);
   U115 : OAI221_X1 port map( B1 => n393, B2 => n477, C1 => n392, C2 => n478, A
                           => n479, ZN => O_42_port);
   U116 : AOI22_X1 port map( A1 => A_ns(41), A2 => n397, B1 => A_s(41), B2 => 
                           n398, ZN => n479);
   U117 : INV_X1 port map( A => A_s(40), ZN => n478);
   U118 : INV_X1 port map( A => A_ns(40), ZN => n477);
   U119 : OAI221_X1 port map( B1 => n393, B2 => n480, C1 => n392, C2 => n481, A
                           => n482, ZN => O_41_port);
   U120 : AOI22_X1 port map( A1 => A_ns(40), A2 => n397, B1 => A_s(40), B2 => 
                           n398, ZN => n482);
   U121 : INV_X1 port map( A => A_s(39), ZN => n481);
   U122 : INV_X1 port map( A => A_ns(39), ZN => n480);
   U123 : OAI221_X1 port map( B1 => n393, B2 => n483, C1 => n392, C2 => n484, A
                           => n485, ZN => O_40_port);
   U124 : AOI22_X1 port map( A1 => A_ns(39), A2 => n397, B1 => A_s(39), B2 => 
                           n398, ZN => n485);
   U125 : INV_X1 port map( A => A_s(38), ZN => n484);
   U126 : INV_X1 port map( A => A_ns(38), ZN => n483);
   U127 : OAI221_X1 port map( B1 => n393, B2 => n486, C1 => n392, C2 => n487, A
                           => n488, ZN => O_3_port);
   U128 : AOI22_X1 port map( A1 => A_ns(2), A2 => n397, B1 => A_s(2), B2 => 
                           n398, ZN => n488);
   U129 : INV_X1 port map( A => A_s(1), ZN => n487);
   U130 : INV_X1 port map( A => A_ns(1), ZN => n486);
   U131 : OAI221_X1 port map( B1 => n393, B2 => n489, C1 => n392, C2 => n490, A
                           => n491, ZN => O_39_port);
   U132 : AOI22_X1 port map( A1 => A_ns(38), A2 => n397, B1 => A_s(38), B2 => 
                           n398, ZN => n491);
   U133 : INV_X1 port map( A => A_s(37), ZN => n490);
   U134 : INV_X1 port map( A => A_ns(37), ZN => n489);
   U135 : OAI221_X1 port map( B1 => n393, B2 => n492, C1 => n392, C2 => n493, A
                           => n494, ZN => O_38_port);
   U136 : AOI22_X1 port map( A1 => A_ns(37), A2 => n397, B1 => A_s(37), B2 => 
                           n398, ZN => n494);
   U137 : INV_X1 port map( A => A_s(36), ZN => n493);
   U138 : INV_X1 port map( A => A_ns(36), ZN => n492);
   U139 : OAI221_X1 port map( B1 => n393, B2 => n495, C1 => n392, C2 => n496, A
                           => n497, ZN => O_37_port);
   U140 : AOI22_X1 port map( A1 => A_ns(36), A2 => n397, B1 => A_s(36), B2 => 
                           n398, ZN => n497);
   U141 : INV_X1 port map( A => A_s(35), ZN => n496);
   U142 : INV_X1 port map( A => A_ns(35), ZN => n495);
   U143 : OAI221_X1 port map( B1 => n393, B2 => n498, C1 => n392, C2 => n499, A
                           => n500, ZN => O_36_port);
   U144 : AOI22_X1 port map( A1 => A_ns(35), A2 => n397, B1 => A_s(35), B2 => 
                           n398, ZN => n500);
   U145 : INV_X1 port map( A => A_s(34), ZN => n499);
   U146 : INV_X1 port map( A => A_ns(34), ZN => n498);
   U147 : OAI221_X1 port map( B1 => n393, B2 => n501, C1 => n392, C2 => n502, A
                           => n503, ZN => O_35_port);
   U148 : AOI22_X1 port map( A1 => A_ns(34), A2 => n397, B1 => A_s(34), B2 => 
                           n398, ZN => n503);
   U149 : INV_X1 port map( A => A_s(33), ZN => n502);
   U150 : INV_X1 port map( A => A_ns(33), ZN => n501);
   U151 : OAI221_X1 port map( B1 => n393, B2 => n504, C1 => n392, C2 => n505, A
                           => n506, ZN => O_34_port);
   U152 : AOI22_X1 port map( A1 => A_ns(33), A2 => n397, B1 => A_s(33), B2 => 
                           n398, ZN => n506);
   U153 : INV_X1 port map( A => A_s(32), ZN => n505);
   U154 : INV_X1 port map( A => A_ns(32), ZN => n504);
   U155 : OAI221_X1 port map( B1 => n393, B2 => n507, C1 => n392, C2 => n508, A
                           => n509, ZN => O_33_port);
   U156 : AOI22_X1 port map( A1 => A_ns(32), A2 => n397, B1 => A_s(32), B2 => 
                           n398, ZN => n509);
   U157 : INV_X1 port map( A => A_s(31), ZN => n508);
   U158 : INV_X1 port map( A => A_ns(31), ZN => n507);
   U159 : OAI221_X1 port map( B1 => n393, B2 => n510, C1 => n392, C2 => n511, A
                           => n512, ZN => O_32_port);
   U160 : AOI22_X1 port map( A1 => A_ns(31), A2 => n397, B1 => A_s(31), B2 => 
                           n398, ZN => n512);
   U161 : INV_X1 port map( A => A_s(30), ZN => n511);
   U162 : INV_X1 port map( A => A_ns(30), ZN => n510);
   U163 : OAI221_X1 port map( B1 => n393, B2 => n513, C1 => n392, C2 => n514, A
                           => n515, ZN => O_31_port);
   U164 : AOI22_X1 port map( A1 => A_ns(30), A2 => n397, B1 => A_s(30), B2 => 
                           n398, ZN => n515);
   U165 : INV_X1 port map( A => A_s(29), ZN => n514);
   U166 : INV_X1 port map( A => A_ns(29), ZN => n513);
   U167 : OAI221_X1 port map( B1 => n393, B2 => n516, C1 => n392, C2 => n517, A
                           => n518, ZN => O_30_port);
   U168 : AOI22_X1 port map( A1 => A_ns(29), A2 => n397, B1 => A_s(29), B2 => 
                           n398, ZN => n518);
   U169 : INV_X1 port map( A => A_s(28), ZN => n517);
   U170 : INV_X1 port map( A => A_ns(28), ZN => n516);
   U171 : OAI221_X1 port map( B1 => n393, B2 => n519, C1 => n392, C2 => n520, A
                           => n521, ZN => O_2_port);
   U172 : AOI22_X1 port map( A1 => A_ns(1), A2 => n397, B1 => A_s(1), B2 => 
                           n398, ZN => n521);
   U173 : OAI221_X1 port map( B1 => n393, B2 => n522, C1 => n392, C2 => n523, A
                           => n524, ZN => O_29_port);
   U174 : AOI22_X1 port map( A1 => A_ns(28), A2 => n397, B1 => A_s(28), B2 => 
                           n398, ZN => n524);
   U175 : INV_X1 port map( A => A_s(27), ZN => n523);
   U176 : INV_X1 port map( A => A_ns(27), ZN => n522);
   U177 : OAI221_X1 port map( B1 => n393, B2 => n525, C1 => n392, C2 => n526, A
                           => n527, ZN => O_28_port);
   U178 : AOI22_X1 port map( A1 => A_ns(27), A2 => n397, B1 => A_s(27), B2 => 
                           n398, ZN => n527);
   U179 : INV_X1 port map( A => A_s(26), ZN => n526);
   U180 : INV_X1 port map( A => A_ns(26), ZN => n525);
   U181 : OAI221_X1 port map( B1 => n393, B2 => n528, C1 => n392, C2 => n529, A
                           => n530, ZN => O_27_port);
   U182 : AOI22_X1 port map( A1 => A_ns(26), A2 => n397, B1 => A_s(26), B2 => 
                           n398, ZN => n530);
   U183 : INV_X1 port map( A => A_s(25), ZN => n529);
   U184 : INV_X1 port map( A => A_ns(25), ZN => n528);
   U185 : OAI221_X1 port map( B1 => n393, B2 => n531, C1 => n392, C2 => n532, A
                           => n533, ZN => O_26_port);
   U186 : AOI22_X1 port map( A1 => A_ns(25), A2 => n397, B1 => A_s(25), B2 => 
                           n398, ZN => n533);
   U187 : INV_X1 port map( A => A_s(24), ZN => n532);
   U188 : INV_X1 port map( A => A_ns(24), ZN => n531);
   U189 : OAI221_X1 port map( B1 => n393, B2 => n534, C1 => n392, C2 => n535, A
                           => n536, ZN => O_25_port);
   U190 : AOI22_X1 port map( A1 => A_ns(24), A2 => n397, B1 => A_s(24), B2 => 
                           n398, ZN => n536);
   U191 : INV_X1 port map( A => A_s(23), ZN => n535);
   U192 : INV_X1 port map( A => A_ns(23), ZN => n534);
   U193 : OAI221_X1 port map( B1 => n393, B2 => n537, C1 => n392, C2 => n538, A
                           => n539, ZN => O_24_port);
   U194 : AOI22_X1 port map( A1 => A_ns(23), A2 => n397, B1 => A_s(23), B2 => 
                           n398, ZN => n539);
   U195 : INV_X1 port map( A => A_s(22), ZN => n538);
   U196 : INV_X1 port map( A => A_ns(22), ZN => n537);
   U197 : OAI221_X1 port map( B1 => n393, B2 => n540, C1 => n392, C2 => n541, A
                           => n542, ZN => O_23_port);
   U198 : AOI22_X1 port map( A1 => A_ns(22), A2 => n397, B1 => A_s(22), B2 => 
                           n398, ZN => n542);
   U199 : INV_X1 port map( A => A_s(21), ZN => n541);
   U200 : INV_X1 port map( A => A_ns(21), ZN => n540);
   U201 : OAI221_X1 port map( B1 => n393, B2 => n543, C1 => n392, C2 => n544, A
                           => n545, ZN => O_22_port);
   U202 : AOI22_X1 port map( A1 => A_ns(21), A2 => n397, B1 => A_s(21), B2 => 
                           n398, ZN => n545);
   U203 : INV_X1 port map( A => A_s(20), ZN => n544);
   U204 : INV_X1 port map( A => A_ns(20), ZN => n543);
   U205 : OAI221_X1 port map( B1 => n393, B2 => n546, C1 => n392, C2 => n547, A
                           => n548, ZN => O_21_port);
   U206 : AOI22_X1 port map( A1 => A_ns(20), A2 => n397, B1 => A_s(20), B2 => 
                           n398, ZN => n548);
   U207 : INV_X1 port map( A => A_s(19), ZN => n547);
   U208 : INV_X1 port map( A => A_ns(19), ZN => n546);
   U209 : OAI221_X1 port map( B1 => n393, B2 => n549, C1 => n392, C2 => n550, A
                           => n551, ZN => O_20_port);
   U210 : AOI22_X1 port map( A1 => A_ns(19), A2 => n397, B1 => A_s(19), B2 => 
                           n398, ZN => n551);
   U211 : INV_X1 port map( A => A_s(18), ZN => n550);
   U212 : INV_X1 port map( A => A_ns(18), ZN => n549);
   U213 : OAI22_X1 port map( A1 => n552, A2 => n520, B1 => n553, B2 => n519, ZN
                           => O_1_port);
   U214 : INV_X1 port map( A => A_ns(0), ZN => n519);
   U215 : INV_X1 port map( A => A_s(0), ZN => n520);
   U216 : OAI221_X1 port map( B1 => n393, B2 => n554, C1 => n392, C2 => n555, A
                           => n556, ZN => O_19_port);
   U217 : AOI22_X1 port map( A1 => A_ns(18), A2 => n397, B1 => A_s(18), B2 => 
                           n398, ZN => n556);
   U218 : INV_X1 port map( A => A_s(17), ZN => n555);
   U219 : INV_X1 port map( A => A_ns(17), ZN => n554);
   U220 : OAI221_X1 port map( B1 => n393, B2 => n557, C1 => n392, C2 => n558, A
                           => n559, ZN => O_18_port);
   U221 : AOI22_X1 port map( A1 => A_ns(17), A2 => n397, B1 => A_s(17), B2 => 
                           n398, ZN => n559);
   U222 : INV_X1 port map( A => A_s(16), ZN => n558);
   U223 : INV_X1 port map( A => A_ns(16), ZN => n557);
   U224 : OAI221_X1 port map( B1 => n393, B2 => n560, C1 => n392, C2 => n561, A
                           => n562, ZN => O_17_port);
   U225 : AOI22_X1 port map( A1 => A_ns(16), A2 => n397, B1 => A_s(16), B2 => 
                           n398, ZN => n562);
   U226 : INV_X1 port map( A => A_s(15), ZN => n561);
   U227 : INV_X1 port map( A => A_ns(15), ZN => n560);
   U228 : OAI221_X1 port map( B1 => n393, B2 => n563, C1 => n392, C2 => n564, A
                           => n565, ZN => O_16_port);
   U229 : AOI22_X1 port map( A1 => A_ns(15), A2 => n397, B1 => A_s(15), B2 => 
                           n398, ZN => n565);
   U230 : INV_X1 port map( A => A_s(14), ZN => n564);
   U231 : INV_X1 port map( A => A_ns(14), ZN => n563);
   U232 : OAI221_X1 port map( B1 => n393, B2 => n566, C1 => n392, C2 => n567, A
                           => n568, ZN => O_15_port);
   U233 : AOI22_X1 port map( A1 => A_ns(14), A2 => n397, B1 => A_s(14), B2 => 
                           n398, ZN => n568);
   U234 : INV_X1 port map( A => A_s(13), ZN => n567);
   U235 : INV_X1 port map( A => A_ns(13), ZN => n566);
   U236 : OAI221_X1 port map( B1 => n393, B2 => n569, C1 => n392, C2 => n570, A
                           => n571, ZN => O_14_port);
   U237 : AOI22_X1 port map( A1 => A_ns(13), A2 => n397, B1 => A_s(13), B2 => 
                           n398, ZN => n571);
   U238 : INV_X1 port map( A => A_s(12), ZN => n570);
   U239 : INV_X1 port map( A => A_ns(12), ZN => n569);
   U240 : OAI221_X1 port map( B1 => n393, B2 => n572, C1 => n392, C2 => n573, A
                           => n574, ZN => O_13_port);
   U241 : AOI22_X1 port map( A1 => A_ns(12), A2 => n397, B1 => A_s(12), B2 => 
                           n398, ZN => n574);
   U242 : INV_X1 port map( A => A_s(11), ZN => n573);
   U243 : INV_X1 port map( A => A_ns(11), ZN => n572);
   U244 : OAI221_X1 port map( B1 => n393, B2 => n575, C1 => n392, C2 => n576, A
                           => n577, ZN => O_12_port);
   U245 : AOI22_X1 port map( A1 => A_ns(11), A2 => n397, B1 => A_s(11), B2 => 
                           n398, ZN => n577);
   U246 : INV_X1 port map( A => A_s(10), ZN => n576);
   U247 : INV_X1 port map( A => A_ns(10), ZN => n575);
   U248 : OAI221_X1 port map( B1 => n393, B2 => n578, C1 => n392, C2 => n579, A
                           => n580, ZN => O_11_port);
   U249 : AOI22_X1 port map( A1 => A_ns(10), A2 => n397, B1 => A_s(10), B2 => 
                           n398, ZN => n580);
   U250 : INV_X1 port map( A => A_s(9), ZN => n579);
   U251 : INV_X1 port map( A => A_ns(9), ZN => n578);
   U252 : OAI221_X1 port map( B1 => n581, B2 => n393, C1 => n582, C2 => n392, A
                           => n583, ZN => O_10_port);
   U253 : AOI22_X1 port map( A1 => A_ns(9), A2 => n397, B1 => A_s(9), B2 => 
                           n398, ZN => n583);
   U254 : NAND2_X1 port map( A1 => n584, A2 => n552, ZN => n553);
   U255 : NAND2_X1 port map( A1 => n584, A2 => n585, ZN => n552);
   U256 : XOR2_X1 port map( A => B(7), B => B(8), Z => n584);
   U257 : INV_X1 port map( A => A_s(8), ZN => n582);
   U258 : INV_X1 port map( A => B(9), ZN => n585);
   U259 : INV_X1 port map( A => A_ns(8), ZN => n581);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity BOOTHENC_NBIT64_i6 is

   port( A, A_n, A_ns, A_s, B : in std_logic_vector (63 downto 0);  O, A_so, 
         A_nso : out std_logic_vector (63 downto 0));

end BOOTHENC_NBIT64_i6;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT64_i6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, O_63_port, O_62_port, O_61_port, O_60_port, O_59_port,
      O_58_port, O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, 
      O_52_port, O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, 
      O_46_port, O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, 
      O_40_port, O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, 
      O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, 
      O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, 
      O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, 
      O_16_port, O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, 
      O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, 
      O_3_port, O_2_port, O_1_port, n391, n392, n393, n394, n395, n396, n397, 
      n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, 
      n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, 
      n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, 
      n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, 
      n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, 
      n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, 
      n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, 
      n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, 
      n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, 
      n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, 
      n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, 
      n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, 
      n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, 
      n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, 
      n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, 
      n578, n579, n580, n581, n582, n583, n584, n585 : std_logic;

begin
   O <= ( O_63_port, O_62_port, O_61_port, O_60_port, O_59_port, O_58_port, 
      O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, O_52_port, 
      O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, O_46_port, 
      O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, O_40_port, 
      O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, 
      O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, 
      O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, 
      O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, O_16_port, 
      O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, O_10_port, 
      O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, O_3_port, 
      O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(61), A_s(60), A_s(59), A_s(58), A_s(57), A_s(56), A_s(55), 
      A_s(54), A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), 
      A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), 
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   A_nso <= ( A_s(61), A_s(60), A_s(59), A_s(58), A_s(57), A_s(56), A_s(55), 
      A_s(54), A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), 
      A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), 
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : AND3_X1 port map( A1 => B(6), A2 => n585, A3 => B(5), ZN => n391);
   U3 : INV_X4 port map( A => n391, ZN => n392);
   U4 : INV_X4 port map( A => n552, ZN => n398);
   U5 : OR3_X4 port map( A1 => B(5), A2 => B(6), A3 => n585, ZN => n393);
   U6 : INV_X4 port map( A => n553, ZN => n397);
   U7 : OAI221_X1 port map( B1 => n393, B2 => n394, C1 => n392, C2 => n395, A 
                           => n396, ZN => O_9_port);
   U8 : AOI22_X1 port map( A1 => A_ns(8), A2 => n397, B1 => A_s(8), B2 => n398,
                           ZN => n396);
   U9 : INV_X1 port map( A => A_s(7), ZN => n395);
   U10 : INV_X1 port map( A => A_ns(7), ZN => n394);
   U11 : OAI221_X1 port map( B1 => n393, B2 => n399, C1 => n392, C2 => n400, A 
                           => n401, ZN => O_8_port);
   U12 : AOI22_X1 port map( A1 => A_ns(7), A2 => n397, B1 => A_s(7), B2 => n398
                           , ZN => n401);
   U13 : INV_X1 port map( A => A_s(6), ZN => n400);
   U14 : INV_X1 port map( A => A_ns(6), ZN => n399);
   U15 : OAI221_X1 port map( B1 => n393, B2 => n402, C1 => n392, C2 => n403, A 
                           => n404, ZN => O_7_port);
   U16 : AOI22_X1 port map( A1 => A_ns(6), A2 => n397, B1 => A_s(6), B2 => n398
                           , ZN => n404);
   U17 : INV_X1 port map( A => A_s(5), ZN => n403);
   U18 : INV_X1 port map( A => A_ns(5), ZN => n402);
   U19 : OAI221_X1 port map( B1 => n393, B2 => n405, C1 => n392, C2 => n406, A 
                           => n407, ZN => O_6_port);
   U20 : AOI22_X1 port map( A1 => A_ns(5), A2 => n397, B1 => A_s(5), B2 => n398
                           , ZN => n407);
   U21 : INV_X1 port map( A => A_s(4), ZN => n406);
   U22 : INV_X1 port map( A => A_ns(4), ZN => n405);
   U23 : OAI221_X1 port map( B1 => n393, B2 => n408, C1 => n392, C2 => n409, A 
                           => n410, ZN => O_63_port);
   U24 : AOI22_X1 port map( A1 => A_ns(62), A2 => n397, B1 => A_s(62), B2 => 
                           n398, ZN => n410);
   U25 : INV_X1 port map( A => A_s(61), ZN => n409);
   U26 : INV_X1 port map( A => A_ns(61), ZN => n408);
   U27 : OAI221_X1 port map( B1 => n393, B2 => n411, C1 => n392, C2 => n412, A 
                           => n413, ZN => O_62_port);
   U28 : AOI22_X1 port map( A1 => A_ns(61), A2 => n397, B1 => A_s(61), B2 => 
                           n398, ZN => n413);
   U29 : INV_X1 port map( A => A_s(60), ZN => n412);
   U30 : INV_X1 port map( A => A_ns(60), ZN => n411);
   U31 : OAI221_X1 port map( B1 => n393, B2 => n414, C1 => n392, C2 => n415, A 
                           => n416, ZN => O_61_port);
   U32 : AOI22_X1 port map( A1 => A_ns(60), A2 => n397, B1 => A_s(60), B2 => 
                           n398, ZN => n416);
   U33 : INV_X1 port map( A => A_s(59), ZN => n415);
   U34 : INV_X1 port map( A => A_ns(59), ZN => n414);
   U35 : OAI221_X1 port map( B1 => n393, B2 => n417, C1 => n392, C2 => n418, A 
                           => n419, ZN => O_60_port);
   U36 : AOI22_X1 port map( A1 => A_ns(59), A2 => n397, B1 => A_s(59), B2 => 
                           n398, ZN => n419);
   U37 : INV_X1 port map( A => A_s(58), ZN => n418);
   U38 : INV_X1 port map( A => A_ns(58), ZN => n417);
   U39 : OAI221_X1 port map( B1 => n393, B2 => n420, C1 => n392, C2 => n421, A 
                           => n422, ZN => O_5_port);
   U40 : AOI22_X1 port map( A1 => A_ns(4), A2 => n397, B1 => A_s(4), B2 => n398
                           , ZN => n422);
   U41 : INV_X1 port map( A => A_s(3), ZN => n421);
   U42 : INV_X1 port map( A => A_ns(3), ZN => n420);
   U43 : OAI221_X1 port map( B1 => n393, B2 => n423, C1 => n392, C2 => n424, A 
                           => n425, ZN => O_59_port);
   U44 : AOI22_X1 port map( A1 => A_ns(58), A2 => n397, B1 => A_s(58), B2 => 
                           n398, ZN => n425);
   U45 : INV_X1 port map( A => A_s(57), ZN => n424);
   U46 : INV_X1 port map( A => A_ns(57), ZN => n423);
   U47 : OAI221_X1 port map( B1 => n393, B2 => n426, C1 => n392, C2 => n427, A 
                           => n428, ZN => O_58_port);
   U48 : AOI22_X1 port map( A1 => A_ns(57), A2 => n397, B1 => A_s(57), B2 => 
                           n398, ZN => n428);
   U49 : INV_X1 port map( A => A_s(56), ZN => n427);
   U50 : INV_X1 port map( A => A_ns(56), ZN => n426);
   U51 : OAI221_X1 port map( B1 => n393, B2 => n429, C1 => n392, C2 => n430, A 
                           => n431, ZN => O_57_port);
   U52 : AOI22_X1 port map( A1 => A_ns(56), A2 => n397, B1 => A_s(56), B2 => 
                           n398, ZN => n431);
   U53 : INV_X1 port map( A => A_s(55), ZN => n430);
   U54 : INV_X1 port map( A => A_ns(55), ZN => n429);
   U55 : OAI221_X1 port map( B1 => n393, B2 => n432, C1 => n392, C2 => n433, A 
                           => n434, ZN => O_56_port);
   U56 : AOI22_X1 port map( A1 => A_ns(55), A2 => n397, B1 => A_s(55), B2 => 
                           n398, ZN => n434);
   U57 : INV_X1 port map( A => A_s(54), ZN => n433);
   U58 : INV_X1 port map( A => A_ns(54), ZN => n432);
   U59 : OAI221_X1 port map( B1 => n393, B2 => n435, C1 => n392, C2 => n436, A 
                           => n437, ZN => O_55_port);
   U60 : AOI22_X1 port map( A1 => A_ns(54), A2 => n397, B1 => A_s(54), B2 => 
                           n398, ZN => n437);
   U61 : INV_X1 port map( A => A_s(53), ZN => n436);
   U62 : INV_X1 port map( A => A_ns(53), ZN => n435);
   U63 : OAI221_X1 port map( B1 => n393, B2 => n438, C1 => n392, C2 => n439, A 
                           => n440, ZN => O_54_port);
   U64 : AOI22_X1 port map( A1 => A_ns(53), A2 => n397, B1 => A_s(53), B2 => 
                           n398, ZN => n440);
   U65 : INV_X1 port map( A => A_s(52), ZN => n439);
   U66 : INV_X1 port map( A => A_ns(52), ZN => n438);
   U67 : OAI221_X1 port map( B1 => n393, B2 => n441, C1 => n392, C2 => n442, A 
                           => n443, ZN => O_53_port);
   U68 : AOI22_X1 port map( A1 => A_ns(52), A2 => n397, B1 => A_s(52), B2 => 
                           n398, ZN => n443);
   U69 : INV_X1 port map( A => A_s(51), ZN => n442);
   U70 : INV_X1 port map( A => A_ns(51), ZN => n441);
   U71 : OAI221_X1 port map( B1 => n393, B2 => n444, C1 => n392, C2 => n445, A 
                           => n446, ZN => O_52_port);
   U72 : AOI22_X1 port map( A1 => A_ns(51), A2 => n397, B1 => A_s(51), B2 => 
                           n398, ZN => n446);
   U73 : INV_X1 port map( A => A_s(50), ZN => n445);
   U74 : INV_X1 port map( A => A_ns(50), ZN => n444);
   U75 : OAI221_X1 port map( B1 => n393, B2 => n447, C1 => n392, C2 => n448, A 
                           => n449, ZN => O_51_port);
   U76 : AOI22_X1 port map( A1 => A_ns(50), A2 => n397, B1 => A_s(50), B2 => 
                           n398, ZN => n449);
   U77 : INV_X1 port map( A => A_s(49), ZN => n448);
   U78 : INV_X1 port map( A => A_ns(49), ZN => n447);
   U79 : OAI221_X1 port map( B1 => n393, B2 => n450, C1 => n392, C2 => n451, A 
                           => n452, ZN => O_50_port);
   U80 : AOI22_X1 port map( A1 => A_ns(49), A2 => n397, B1 => A_s(49), B2 => 
                           n398, ZN => n452);
   U81 : INV_X1 port map( A => A_s(48), ZN => n451);
   U82 : INV_X1 port map( A => A_ns(48), ZN => n450);
   U83 : OAI221_X1 port map( B1 => n393, B2 => n453, C1 => n392, C2 => n454, A 
                           => n455, ZN => O_4_port);
   U84 : AOI22_X1 port map( A1 => A_ns(3), A2 => n397, B1 => A_s(3), B2 => n398
                           , ZN => n455);
   U85 : INV_X1 port map( A => A_s(2), ZN => n454);
   U86 : INV_X1 port map( A => A_ns(2), ZN => n453);
   U87 : OAI221_X1 port map( B1 => n393, B2 => n456, C1 => n392, C2 => n457, A 
                           => n458, ZN => O_49_port);
   U88 : AOI22_X1 port map( A1 => A_ns(48), A2 => n397, B1 => A_s(48), B2 => 
                           n398, ZN => n458);
   U89 : INV_X1 port map( A => A_s(47), ZN => n457);
   U90 : INV_X1 port map( A => A_ns(47), ZN => n456);
   U91 : OAI221_X1 port map( B1 => n393, B2 => n459, C1 => n392, C2 => n460, A 
                           => n461, ZN => O_48_port);
   U92 : AOI22_X1 port map( A1 => A_ns(47), A2 => n397, B1 => A_s(47), B2 => 
                           n398, ZN => n461);
   U93 : INV_X1 port map( A => A_s(46), ZN => n460);
   U94 : INV_X1 port map( A => A_ns(46), ZN => n459);
   U95 : OAI221_X1 port map( B1 => n393, B2 => n462, C1 => n392, C2 => n463, A 
                           => n464, ZN => O_47_port);
   U96 : AOI22_X1 port map( A1 => A_ns(46), A2 => n397, B1 => A_s(46), B2 => 
                           n398, ZN => n464);
   U97 : INV_X1 port map( A => A_s(45), ZN => n463);
   U98 : INV_X1 port map( A => A_ns(45), ZN => n462);
   U99 : OAI221_X1 port map( B1 => n393, B2 => n465, C1 => n392, C2 => n466, A 
                           => n467, ZN => O_46_port);
   U100 : AOI22_X1 port map( A1 => A_ns(45), A2 => n397, B1 => A_s(45), B2 => 
                           n398, ZN => n467);
   U101 : INV_X1 port map( A => A_s(44), ZN => n466);
   U102 : INV_X1 port map( A => A_ns(44), ZN => n465);
   U103 : OAI221_X1 port map( B1 => n393, B2 => n468, C1 => n392, C2 => n469, A
                           => n470, ZN => O_45_port);
   U104 : AOI22_X1 port map( A1 => A_ns(44), A2 => n397, B1 => A_s(44), B2 => 
                           n398, ZN => n470);
   U105 : INV_X1 port map( A => A_s(43), ZN => n469);
   U106 : INV_X1 port map( A => A_ns(43), ZN => n468);
   U107 : OAI221_X1 port map( B1 => n393, B2 => n471, C1 => n392, C2 => n472, A
                           => n473, ZN => O_44_port);
   U108 : AOI22_X1 port map( A1 => A_ns(43), A2 => n397, B1 => A_s(43), B2 => 
                           n398, ZN => n473);
   U109 : INV_X1 port map( A => A_s(42), ZN => n472);
   U110 : INV_X1 port map( A => A_ns(42), ZN => n471);
   U111 : OAI221_X1 port map( B1 => n393, B2 => n474, C1 => n392, C2 => n475, A
                           => n476, ZN => O_43_port);
   U112 : AOI22_X1 port map( A1 => A_ns(42), A2 => n397, B1 => A_s(42), B2 => 
                           n398, ZN => n476);
   U113 : INV_X1 port map( A => A_s(41), ZN => n475);
   U114 : INV_X1 port map( A => A_ns(41), ZN => n474);
   U115 : OAI221_X1 port map( B1 => n393, B2 => n477, C1 => n392, C2 => n478, A
                           => n479, ZN => O_42_port);
   U116 : AOI22_X1 port map( A1 => A_ns(41), A2 => n397, B1 => A_s(41), B2 => 
                           n398, ZN => n479);
   U117 : INV_X1 port map( A => A_s(40), ZN => n478);
   U118 : INV_X1 port map( A => A_ns(40), ZN => n477);
   U119 : OAI221_X1 port map( B1 => n393, B2 => n480, C1 => n392, C2 => n481, A
                           => n482, ZN => O_41_port);
   U120 : AOI22_X1 port map( A1 => A_ns(40), A2 => n397, B1 => A_s(40), B2 => 
                           n398, ZN => n482);
   U121 : INV_X1 port map( A => A_s(39), ZN => n481);
   U122 : INV_X1 port map( A => A_ns(39), ZN => n480);
   U123 : OAI221_X1 port map( B1 => n393, B2 => n483, C1 => n392, C2 => n484, A
                           => n485, ZN => O_40_port);
   U124 : AOI22_X1 port map( A1 => A_ns(39), A2 => n397, B1 => A_s(39), B2 => 
                           n398, ZN => n485);
   U125 : INV_X1 port map( A => A_s(38), ZN => n484);
   U126 : INV_X1 port map( A => A_ns(38), ZN => n483);
   U127 : OAI221_X1 port map( B1 => n393, B2 => n486, C1 => n392, C2 => n487, A
                           => n488, ZN => O_3_port);
   U128 : AOI22_X1 port map( A1 => A_ns(2), A2 => n397, B1 => A_s(2), B2 => 
                           n398, ZN => n488);
   U129 : INV_X1 port map( A => A_s(1), ZN => n487);
   U130 : INV_X1 port map( A => A_ns(1), ZN => n486);
   U131 : OAI221_X1 port map( B1 => n393, B2 => n489, C1 => n392, C2 => n490, A
                           => n491, ZN => O_39_port);
   U132 : AOI22_X1 port map( A1 => A_ns(38), A2 => n397, B1 => A_s(38), B2 => 
                           n398, ZN => n491);
   U133 : INV_X1 port map( A => A_s(37), ZN => n490);
   U134 : INV_X1 port map( A => A_ns(37), ZN => n489);
   U135 : OAI221_X1 port map( B1 => n393, B2 => n492, C1 => n392, C2 => n493, A
                           => n494, ZN => O_38_port);
   U136 : AOI22_X1 port map( A1 => A_ns(37), A2 => n397, B1 => A_s(37), B2 => 
                           n398, ZN => n494);
   U137 : INV_X1 port map( A => A_s(36), ZN => n493);
   U138 : INV_X1 port map( A => A_ns(36), ZN => n492);
   U139 : OAI221_X1 port map( B1 => n393, B2 => n495, C1 => n392, C2 => n496, A
                           => n497, ZN => O_37_port);
   U140 : AOI22_X1 port map( A1 => A_ns(36), A2 => n397, B1 => A_s(36), B2 => 
                           n398, ZN => n497);
   U141 : INV_X1 port map( A => A_s(35), ZN => n496);
   U142 : INV_X1 port map( A => A_ns(35), ZN => n495);
   U143 : OAI221_X1 port map( B1 => n393, B2 => n498, C1 => n392, C2 => n499, A
                           => n500, ZN => O_36_port);
   U144 : AOI22_X1 port map( A1 => A_ns(35), A2 => n397, B1 => A_s(35), B2 => 
                           n398, ZN => n500);
   U145 : INV_X1 port map( A => A_s(34), ZN => n499);
   U146 : INV_X1 port map( A => A_ns(34), ZN => n498);
   U147 : OAI221_X1 port map( B1 => n393, B2 => n501, C1 => n392, C2 => n502, A
                           => n503, ZN => O_35_port);
   U148 : AOI22_X1 port map( A1 => A_ns(34), A2 => n397, B1 => A_s(34), B2 => 
                           n398, ZN => n503);
   U149 : INV_X1 port map( A => A_s(33), ZN => n502);
   U150 : INV_X1 port map( A => A_ns(33), ZN => n501);
   U151 : OAI221_X1 port map( B1 => n393, B2 => n504, C1 => n392, C2 => n505, A
                           => n506, ZN => O_34_port);
   U152 : AOI22_X1 port map( A1 => A_ns(33), A2 => n397, B1 => A_s(33), B2 => 
                           n398, ZN => n506);
   U153 : INV_X1 port map( A => A_s(32), ZN => n505);
   U154 : INV_X1 port map( A => A_ns(32), ZN => n504);
   U155 : OAI221_X1 port map( B1 => n393, B2 => n507, C1 => n392, C2 => n508, A
                           => n509, ZN => O_33_port);
   U156 : AOI22_X1 port map( A1 => A_ns(32), A2 => n397, B1 => A_s(32), B2 => 
                           n398, ZN => n509);
   U157 : INV_X1 port map( A => A_s(31), ZN => n508);
   U158 : INV_X1 port map( A => A_ns(31), ZN => n507);
   U159 : OAI221_X1 port map( B1 => n393, B2 => n510, C1 => n392, C2 => n511, A
                           => n512, ZN => O_32_port);
   U160 : AOI22_X1 port map( A1 => A_ns(31), A2 => n397, B1 => A_s(31), B2 => 
                           n398, ZN => n512);
   U161 : INV_X1 port map( A => A_s(30), ZN => n511);
   U162 : INV_X1 port map( A => A_ns(30), ZN => n510);
   U163 : OAI221_X1 port map( B1 => n393, B2 => n513, C1 => n392, C2 => n514, A
                           => n515, ZN => O_31_port);
   U164 : AOI22_X1 port map( A1 => A_ns(30), A2 => n397, B1 => A_s(30), B2 => 
                           n398, ZN => n515);
   U165 : INV_X1 port map( A => A_s(29), ZN => n514);
   U166 : INV_X1 port map( A => A_ns(29), ZN => n513);
   U167 : OAI221_X1 port map( B1 => n393, B2 => n516, C1 => n392, C2 => n517, A
                           => n518, ZN => O_30_port);
   U168 : AOI22_X1 port map( A1 => A_ns(29), A2 => n397, B1 => A_s(29), B2 => 
                           n398, ZN => n518);
   U169 : INV_X1 port map( A => A_s(28), ZN => n517);
   U170 : INV_X1 port map( A => A_ns(28), ZN => n516);
   U171 : OAI221_X1 port map( B1 => n393, B2 => n519, C1 => n392, C2 => n520, A
                           => n521, ZN => O_2_port);
   U172 : AOI22_X1 port map( A1 => A_ns(1), A2 => n397, B1 => A_s(1), B2 => 
                           n398, ZN => n521);
   U173 : OAI221_X1 port map( B1 => n393, B2 => n522, C1 => n392, C2 => n523, A
                           => n524, ZN => O_29_port);
   U174 : AOI22_X1 port map( A1 => A_ns(28), A2 => n397, B1 => A_s(28), B2 => 
                           n398, ZN => n524);
   U175 : INV_X1 port map( A => A_s(27), ZN => n523);
   U176 : INV_X1 port map( A => A_ns(27), ZN => n522);
   U177 : OAI221_X1 port map( B1 => n393, B2 => n525, C1 => n392, C2 => n526, A
                           => n527, ZN => O_28_port);
   U178 : AOI22_X1 port map( A1 => A_ns(27), A2 => n397, B1 => A_s(27), B2 => 
                           n398, ZN => n527);
   U179 : INV_X1 port map( A => A_s(26), ZN => n526);
   U180 : INV_X1 port map( A => A_ns(26), ZN => n525);
   U181 : OAI221_X1 port map( B1 => n393, B2 => n528, C1 => n392, C2 => n529, A
                           => n530, ZN => O_27_port);
   U182 : AOI22_X1 port map( A1 => A_ns(26), A2 => n397, B1 => A_s(26), B2 => 
                           n398, ZN => n530);
   U183 : INV_X1 port map( A => A_s(25), ZN => n529);
   U184 : INV_X1 port map( A => A_ns(25), ZN => n528);
   U185 : OAI221_X1 port map( B1 => n393, B2 => n531, C1 => n392, C2 => n532, A
                           => n533, ZN => O_26_port);
   U186 : AOI22_X1 port map( A1 => A_ns(25), A2 => n397, B1 => A_s(25), B2 => 
                           n398, ZN => n533);
   U187 : INV_X1 port map( A => A_s(24), ZN => n532);
   U188 : INV_X1 port map( A => A_ns(24), ZN => n531);
   U189 : OAI221_X1 port map( B1 => n393, B2 => n534, C1 => n392, C2 => n535, A
                           => n536, ZN => O_25_port);
   U190 : AOI22_X1 port map( A1 => A_ns(24), A2 => n397, B1 => A_s(24), B2 => 
                           n398, ZN => n536);
   U191 : INV_X1 port map( A => A_s(23), ZN => n535);
   U192 : INV_X1 port map( A => A_ns(23), ZN => n534);
   U193 : OAI221_X1 port map( B1 => n393, B2 => n537, C1 => n392, C2 => n538, A
                           => n539, ZN => O_24_port);
   U194 : AOI22_X1 port map( A1 => A_ns(23), A2 => n397, B1 => A_s(23), B2 => 
                           n398, ZN => n539);
   U195 : INV_X1 port map( A => A_s(22), ZN => n538);
   U196 : INV_X1 port map( A => A_ns(22), ZN => n537);
   U197 : OAI221_X1 port map( B1 => n393, B2 => n540, C1 => n392, C2 => n541, A
                           => n542, ZN => O_23_port);
   U198 : AOI22_X1 port map( A1 => A_ns(22), A2 => n397, B1 => A_s(22), B2 => 
                           n398, ZN => n542);
   U199 : INV_X1 port map( A => A_s(21), ZN => n541);
   U200 : INV_X1 port map( A => A_ns(21), ZN => n540);
   U201 : OAI221_X1 port map( B1 => n393, B2 => n543, C1 => n392, C2 => n544, A
                           => n545, ZN => O_22_port);
   U202 : AOI22_X1 port map( A1 => A_ns(21), A2 => n397, B1 => A_s(21), B2 => 
                           n398, ZN => n545);
   U203 : INV_X1 port map( A => A_s(20), ZN => n544);
   U204 : INV_X1 port map( A => A_ns(20), ZN => n543);
   U205 : OAI221_X1 port map( B1 => n393, B2 => n546, C1 => n392, C2 => n547, A
                           => n548, ZN => O_21_port);
   U206 : AOI22_X1 port map( A1 => A_ns(20), A2 => n397, B1 => A_s(20), B2 => 
                           n398, ZN => n548);
   U207 : INV_X1 port map( A => A_s(19), ZN => n547);
   U208 : INV_X1 port map( A => A_ns(19), ZN => n546);
   U209 : OAI221_X1 port map( B1 => n393, B2 => n549, C1 => n392, C2 => n550, A
                           => n551, ZN => O_20_port);
   U210 : AOI22_X1 port map( A1 => A_ns(19), A2 => n397, B1 => A_s(19), B2 => 
                           n398, ZN => n551);
   U211 : INV_X1 port map( A => A_s(18), ZN => n550);
   U212 : INV_X1 port map( A => A_ns(18), ZN => n549);
   U213 : OAI22_X1 port map( A1 => n552, A2 => n520, B1 => n553, B2 => n519, ZN
                           => O_1_port);
   U214 : INV_X1 port map( A => A_ns(0), ZN => n519);
   U215 : INV_X1 port map( A => A_s(0), ZN => n520);
   U216 : OAI221_X1 port map( B1 => n393, B2 => n554, C1 => n392, C2 => n555, A
                           => n556, ZN => O_19_port);
   U217 : AOI22_X1 port map( A1 => A_ns(18), A2 => n397, B1 => A_s(18), B2 => 
                           n398, ZN => n556);
   U218 : INV_X1 port map( A => A_s(17), ZN => n555);
   U219 : INV_X1 port map( A => A_ns(17), ZN => n554);
   U220 : OAI221_X1 port map( B1 => n393, B2 => n557, C1 => n392, C2 => n558, A
                           => n559, ZN => O_18_port);
   U221 : AOI22_X1 port map( A1 => A_ns(17), A2 => n397, B1 => A_s(17), B2 => 
                           n398, ZN => n559);
   U222 : INV_X1 port map( A => A_s(16), ZN => n558);
   U223 : INV_X1 port map( A => A_ns(16), ZN => n557);
   U224 : OAI221_X1 port map( B1 => n393, B2 => n560, C1 => n392, C2 => n561, A
                           => n562, ZN => O_17_port);
   U225 : AOI22_X1 port map( A1 => A_ns(16), A2 => n397, B1 => A_s(16), B2 => 
                           n398, ZN => n562);
   U226 : INV_X1 port map( A => A_s(15), ZN => n561);
   U227 : INV_X1 port map( A => A_ns(15), ZN => n560);
   U228 : OAI221_X1 port map( B1 => n393, B2 => n563, C1 => n392, C2 => n564, A
                           => n565, ZN => O_16_port);
   U229 : AOI22_X1 port map( A1 => A_ns(15), A2 => n397, B1 => A_s(15), B2 => 
                           n398, ZN => n565);
   U230 : INV_X1 port map( A => A_s(14), ZN => n564);
   U231 : INV_X1 port map( A => A_ns(14), ZN => n563);
   U232 : OAI221_X1 port map( B1 => n393, B2 => n566, C1 => n392, C2 => n567, A
                           => n568, ZN => O_15_port);
   U233 : AOI22_X1 port map( A1 => A_ns(14), A2 => n397, B1 => A_s(14), B2 => 
                           n398, ZN => n568);
   U234 : INV_X1 port map( A => A_s(13), ZN => n567);
   U235 : INV_X1 port map( A => A_ns(13), ZN => n566);
   U236 : OAI221_X1 port map( B1 => n393, B2 => n569, C1 => n392, C2 => n570, A
                           => n571, ZN => O_14_port);
   U237 : AOI22_X1 port map( A1 => A_ns(13), A2 => n397, B1 => A_s(13), B2 => 
                           n398, ZN => n571);
   U238 : INV_X1 port map( A => A_s(12), ZN => n570);
   U239 : INV_X1 port map( A => A_ns(12), ZN => n569);
   U240 : OAI221_X1 port map( B1 => n393, B2 => n572, C1 => n392, C2 => n573, A
                           => n574, ZN => O_13_port);
   U241 : AOI22_X1 port map( A1 => A_ns(12), A2 => n397, B1 => A_s(12), B2 => 
                           n398, ZN => n574);
   U242 : INV_X1 port map( A => A_s(11), ZN => n573);
   U243 : INV_X1 port map( A => A_ns(11), ZN => n572);
   U244 : OAI221_X1 port map( B1 => n393, B2 => n575, C1 => n392, C2 => n576, A
                           => n577, ZN => O_12_port);
   U245 : AOI22_X1 port map( A1 => A_ns(11), A2 => n397, B1 => A_s(11), B2 => 
                           n398, ZN => n577);
   U246 : INV_X1 port map( A => A_s(10), ZN => n576);
   U247 : INV_X1 port map( A => A_ns(10), ZN => n575);
   U248 : OAI221_X1 port map( B1 => n393, B2 => n578, C1 => n392, C2 => n579, A
                           => n580, ZN => O_11_port);
   U249 : AOI22_X1 port map( A1 => A_ns(10), A2 => n397, B1 => A_s(10), B2 => 
                           n398, ZN => n580);
   U250 : INV_X1 port map( A => A_s(9), ZN => n579);
   U251 : INV_X1 port map( A => A_ns(9), ZN => n578);
   U252 : OAI221_X1 port map( B1 => n581, B2 => n393, C1 => n582, C2 => n392, A
                           => n583, ZN => O_10_port);
   U253 : AOI22_X1 port map( A1 => A_ns(9), A2 => n397, B1 => A_s(9), B2 => 
                           n398, ZN => n583);
   U254 : NAND2_X1 port map( A1 => n584, A2 => n552, ZN => n553);
   U255 : NAND2_X1 port map( A1 => n584, A2 => n585, ZN => n552);
   U256 : XOR2_X1 port map( A => B(5), B => B(6), Z => n584);
   U257 : INV_X1 port map( A => A_s(8), ZN => n582);
   U258 : INV_X1 port map( A => B(7), ZN => n585);
   U259 : INV_X1 port map( A => A_ns(8), ZN => n581);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity BOOTHENC_NBIT64_i4 is

   port( A, A_n, A_ns, A_s, B : in std_logic_vector (63 downto 0);  O, A_so, 
         A_nso : out std_logic_vector (63 downto 0));

end BOOTHENC_NBIT64_i4;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT64_i4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, O_63_port, O_62_port, O_61_port, O_60_port, O_59_port,
      O_58_port, O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, 
      O_52_port, O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, 
      O_46_port, O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, 
      O_40_port, O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, 
      O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, 
      O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, 
      O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, 
      O_16_port, O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, 
      O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, 
      O_3_port, O_2_port, O_1_port, n391, n392, n393, n394, n395, n396, n397, 
      n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, 
      n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, 
      n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, 
      n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, 
      n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, 
      n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, 
      n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, 
      n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, 
      n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, 
      n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, 
      n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, 
      n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, 
      n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, 
      n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, 
      n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, 
      n578, n579, n580, n581, n582, n583, n584, n585 : std_logic;

begin
   O <= ( O_63_port, O_62_port, O_61_port, O_60_port, O_59_port, O_58_port, 
      O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, O_52_port, 
      O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, O_46_port, 
      O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, O_40_port, 
      O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, 
      O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, 
      O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, 
      O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, O_16_port, 
      O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, O_10_port, 
      O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, O_3_port, 
      O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(61), A_s(60), A_s(59), A_s(58), A_s(57), A_s(56), A_s(55), 
      A_s(54), A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), 
      A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), 
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   A_nso <= ( A_s(61), A_s(60), A_s(59), A_s(58), A_s(57), A_s(56), A_s(55), 
      A_s(54), A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), 
      A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), 
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : AND3_X1 port map( A1 => B(4), A2 => n585, A3 => B(3), ZN => n391);
   U3 : INV_X4 port map( A => n391, ZN => n392);
   U4 : INV_X4 port map( A => n552, ZN => n398);
   U5 : OR3_X4 port map( A1 => B(3), A2 => B(4), A3 => n585, ZN => n393);
   U6 : INV_X4 port map( A => n553, ZN => n397);
   U7 : OAI221_X1 port map( B1 => n393, B2 => n394, C1 => n392, C2 => n395, A 
                           => n396, ZN => O_9_port);
   U8 : AOI22_X1 port map( A1 => A_ns(8), A2 => n397, B1 => A_s(8), B2 => n398,
                           ZN => n396);
   U9 : INV_X1 port map( A => A_s(7), ZN => n395);
   U10 : INV_X1 port map( A => A_ns(7), ZN => n394);
   U11 : OAI221_X1 port map( B1 => n393, B2 => n399, C1 => n392, C2 => n400, A 
                           => n401, ZN => O_8_port);
   U12 : AOI22_X1 port map( A1 => A_ns(7), A2 => n397, B1 => A_s(7), B2 => n398
                           , ZN => n401);
   U13 : INV_X1 port map( A => A_s(6), ZN => n400);
   U14 : INV_X1 port map( A => A_ns(6), ZN => n399);
   U15 : OAI221_X1 port map( B1 => n393, B2 => n402, C1 => n392, C2 => n403, A 
                           => n404, ZN => O_7_port);
   U16 : AOI22_X1 port map( A1 => A_ns(6), A2 => n397, B1 => A_s(6), B2 => n398
                           , ZN => n404);
   U17 : INV_X1 port map( A => A_s(5), ZN => n403);
   U18 : INV_X1 port map( A => A_ns(5), ZN => n402);
   U19 : OAI221_X1 port map( B1 => n393, B2 => n405, C1 => n392, C2 => n406, A 
                           => n407, ZN => O_6_port);
   U20 : AOI22_X1 port map( A1 => A_ns(5), A2 => n397, B1 => A_s(5), B2 => n398
                           , ZN => n407);
   U21 : INV_X1 port map( A => A_s(4), ZN => n406);
   U22 : INV_X1 port map( A => A_ns(4), ZN => n405);
   U23 : OAI221_X1 port map( B1 => n393, B2 => n408, C1 => n392, C2 => n409, A 
                           => n410, ZN => O_63_port);
   U24 : AOI22_X1 port map( A1 => A_ns(62), A2 => n397, B1 => A_s(62), B2 => 
                           n398, ZN => n410);
   U25 : INV_X1 port map( A => A_s(61), ZN => n409);
   U26 : INV_X1 port map( A => A_ns(61), ZN => n408);
   U27 : OAI221_X1 port map( B1 => n393, B2 => n411, C1 => n392, C2 => n412, A 
                           => n413, ZN => O_62_port);
   U28 : AOI22_X1 port map( A1 => A_ns(61), A2 => n397, B1 => A_s(61), B2 => 
                           n398, ZN => n413);
   U29 : INV_X1 port map( A => A_s(60), ZN => n412);
   U30 : INV_X1 port map( A => A_ns(60), ZN => n411);
   U31 : OAI221_X1 port map( B1 => n393, B2 => n414, C1 => n392, C2 => n415, A 
                           => n416, ZN => O_61_port);
   U32 : AOI22_X1 port map( A1 => A_ns(60), A2 => n397, B1 => A_s(60), B2 => 
                           n398, ZN => n416);
   U33 : INV_X1 port map( A => A_s(59), ZN => n415);
   U34 : INV_X1 port map( A => A_ns(59), ZN => n414);
   U35 : OAI221_X1 port map( B1 => n393, B2 => n417, C1 => n392, C2 => n418, A 
                           => n419, ZN => O_60_port);
   U36 : AOI22_X1 port map( A1 => A_ns(59), A2 => n397, B1 => A_s(59), B2 => 
                           n398, ZN => n419);
   U37 : INV_X1 port map( A => A_s(58), ZN => n418);
   U38 : INV_X1 port map( A => A_ns(58), ZN => n417);
   U39 : OAI221_X1 port map( B1 => n393, B2 => n420, C1 => n392, C2 => n421, A 
                           => n422, ZN => O_5_port);
   U40 : AOI22_X1 port map( A1 => A_ns(4), A2 => n397, B1 => A_s(4), B2 => n398
                           , ZN => n422);
   U41 : INV_X1 port map( A => A_s(3), ZN => n421);
   U42 : INV_X1 port map( A => A_ns(3), ZN => n420);
   U43 : OAI221_X1 port map( B1 => n393, B2 => n423, C1 => n392, C2 => n424, A 
                           => n425, ZN => O_59_port);
   U44 : AOI22_X1 port map( A1 => A_ns(58), A2 => n397, B1 => A_s(58), B2 => 
                           n398, ZN => n425);
   U45 : INV_X1 port map( A => A_s(57), ZN => n424);
   U46 : INV_X1 port map( A => A_ns(57), ZN => n423);
   U47 : OAI221_X1 port map( B1 => n393, B2 => n426, C1 => n392, C2 => n427, A 
                           => n428, ZN => O_58_port);
   U48 : AOI22_X1 port map( A1 => A_ns(57), A2 => n397, B1 => A_s(57), B2 => 
                           n398, ZN => n428);
   U49 : INV_X1 port map( A => A_s(56), ZN => n427);
   U50 : INV_X1 port map( A => A_ns(56), ZN => n426);
   U51 : OAI221_X1 port map( B1 => n393, B2 => n429, C1 => n392, C2 => n430, A 
                           => n431, ZN => O_57_port);
   U52 : AOI22_X1 port map( A1 => A_ns(56), A2 => n397, B1 => A_s(56), B2 => 
                           n398, ZN => n431);
   U53 : INV_X1 port map( A => A_s(55), ZN => n430);
   U54 : INV_X1 port map( A => A_ns(55), ZN => n429);
   U55 : OAI221_X1 port map( B1 => n393, B2 => n432, C1 => n392, C2 => n433, A 
                           => n434, ZN => O_56_port);
   U56 : AOI22_X1 port map( A1 => A_ns(55), A2 => n397, B1 => A_s(55), B2 => 
                           n398, ZN => n434);
   U57 : INV_X1 port map( A => A_s(54), ZN => n433);
   U58 : INV_X1 port map( A => A_ns(54), ZN => n432);
   U59 : OAI221_X1 port map( B1 => n393, B2 => n435, C1 => n392, C2 => n436, A 
                           => n437, ZN => O_55_port);
   U60 : AOI22_X1 port map( A1 => A_ns(54), A2 => n397, B1 => A_s(54), B2 => 
                           n398, ZN => n437);
   U61 : INV_X1 port map( A => A_s(53), ZN => n436);
   U62 : INV_X1 port map( A => A_ns(53), ZN => n435);
   U63 : OAI221_X1 port map( B1 => n393, B2 => n438, C1 => n392, C2 => n439, A 
                           => n440, ZN => O_54_port);
   U64 : AOI22_X1 port map( A1 => A_ns(53), A2 => n397, B1 => A_s(53), B2 => 
                           n398, ZN => n440);
   U65 : INV_X1 port map( A => A_s(52), ZN => n439);
   U66 : INV_X1 port map( A => A_ns(52), ZN => n438);
   U67 : OAI221_X1 port map( B1 => n393, B2 => n441, C1 => n392, C2 => n442, A 
                           => n443, ZN => O_53_port);
   U68 : AOI22_X1 port map( A1 => A_ns(52), A2 => n397, B1 => A_s(52), B2 => 
                           n398, ZN => n443);
   U69 : INV_X1 port map( A => A_s(51), ZN => n442);
   U70 : INV_X1 port map( A => A_ns(51), ZN => n441);
   U71 : OAI221_X1 port map( B1 => n393, B2 => n444, C1 => n392, C2 => n445, A 
                           => n446, ZN => O_52_port);
   U72 : AOI22_X1 port map( A1 => A_ns(51), A2 => n397, B1 => A_s(51), B2 => 
                           n398, ZN => n446);
   U73 : INV_X1 port map( A => A_s(50), ZN => n445);
   U74 : INV_X1 port map( A => A_ns(50), ZN => n444);
   U75 : OAI221_X1 port map( B1 => n393, B2 => n447, C1 => n392, C2 => n448, A 
                           => n449, ZN => O_51_port);
   U76 : AOI22_X1 port map( A1 => A_ns(50), A2 => n397, B1 => A_s(50), B2 => 
                           n398, ZN => n449);
   U77 : INV_X1 port map( A => A_s(49), ZN => n448);
   U78 : INV_X1 port map( A => A_ns(49), ZN => n447);
   U79 : OAI221_X1 port map( B1 => n393, B2 => n450, C1 => n392, C2 => n451, A 
                           => n452, ZN => O_50_port);
   U80 : AOI22_X1 port map( A1 => A_ns(49), A2 => n397, B1 => A_s(49), B2 => 
                           n398, ZN => n452);
   U81 : INV_X1 port map( A => A_s(48), ZN => n451);
   U82 : INV_X1 port map( A => A_ns(48), ZN => n450);
   U83 : OAI221_X1 port map( B1 => n393, B2 => n453, C1 => n392, C2 => n454, A 
                           => n455, ZN => O_4_port);
   U84 : AOI22_X1 port map( A1 => A_ns(3), A2 => n397, B1 => A_s(3), B2 => n398
                           , ZN => n455);
   U85 : INV_X1 port map( A => A_s(2), ZN => n454);
   U86 : INV_X1 port map( A => A_ns(2), ZN => n453);
   U87 : OAI221_X1 port map( B1 => n393, B2 => n456, C1 => n392, C2 => n457, A 
                           => n458, ZN => O_49_port);
   U88 : AOI22_X1 port map( A1 => A_ns(48), A2 => n397, B1 => A_s(48), B2 => 
                           n398, ZN => n458);
   U89 : INV_X1 port map( A => A_s(47), ZN => n457);
   U90 : INV_X1 port map( A => A_ns(47), ZN => n456);
   U91 : OAI221_X1 port map( B1 => n393, B2 => n459, C1 => n392, C2 => n460, A 
                           => n461, ZN => O_48_port);
   U92 : AOI22_X1 port map( A1 => A_ns(47), A2 => n397, B1 => A_s(47), B2 => 
                           n398, ZN => n461);
   U93 : INV_X1 port map( A => A_s(46), ZN => n460);
   U94 : INV_X1 port map( A => A_ns(46), ZN => n459);
   U95 : OAI221_X1 port map( B1 => n393, B2 => n462, C1 => n392, C2 => n463, A 
                           => n464, ZN => O_47_port);
   U96 : AOI22_X1 port map( A1 => A_ns(46), A2 => n397, B1 => A_s(46), B2 => 
                           n398, ZN => n464);
   U97 : INV_X1 port map( A => A_s(45), ZN => n463);
   U98 : INV_X1 port map( A => A_ns(45), ZN => n462);
   U99 : OAI221_X1 port map( B1 => n393, B2 => n465, C1 => n392, C2 => n466, A 
                           => n467, ZN => O_46_port);
   U100 : AOI22_X1 port map( A1 => A_ns(45), A2 => n397, B1 => A_s(45), B2 => 
                           n398, ZN => n467);
   U101 : INV_X1 port map( A => A_s(44), ZN => n466);
   U102 : INV_X1 port map( A => A_ns(44), ZN => n465);
   U103 : OAI221_X1 port map( B1 => n393, B2 => n468, C1 => n392, C2 => n469, A
                           => n470, ZN => O_45_port);
   U104 : AOI22_X1 port map( A1 => A_ns(44), A2 => n397, B1 => A_s(44), B2 => 
                           n398, ZN => n470);
   U105 : INV_X1 port map( A => A_s(43), ZN => n469);
   U106 : INV_X1 port map( A => A_ns(43), ZN => n468);
   U107 : OAI221_X1 port map( B1 => n393, B2 => n471, C1 => n392, C2 => n472, A
                           => n473, ZN => O_44_port);
   U108 : AOI22_X1 port map( A1 => A_ns(43), A2 => n397, B1 => A_s(43), B2 => 
                           n398, ZN => n473);
   U109 : INV_X1 port map( A => A_s(42), ZN => n472);
   U110 : INV_X1 port map( A => A_ns(42), ZN => n471);
   U111 : OAI221_X1 port map( B1 => n393, B2 => n474, C1 => n392, C2 => n475, A
                           => n476, ZN => O_43_port);
   U112 : AOI22_X1 port map( A1 => A_ns(42), A2 => n397, B1 => A_s(42), B2 => 
                           n398, ZN => n476);
   U113 : INV_X1 port map( A => A_s(41), ZN => n475);
   U114 : INV_X1 port map( A => A_ns(41), ZN => n474);
   U115 : OAI221_X1 port map( B1 => n393, B2 => n477, C1 => n392, C2 => n478, A
                           => n479, ZN => O_42_port);
   U116 : AOI22_X1 port map( A1 => A_ns(41), A2 => n397, B1 => A_s(41), B2 => 
                           n398, ZN => n479);
   U117 : INV_X1 port map( A => A_s(40), ZN => n478);
   U118 : INV_X1 port map( A => A_ns(40), ZN => n477);
   U119 : OAI221_X1 port map( B1 => n393, B2 => n480, C1 => n392, C2 => n481, A
                           => n482, ZN => O_41_port);
   U120 : AOI22_X1 port map( A1 => A_ns(40), A2 => n397, B1 => A_s(40), B2 => 
                           n398, ZN => n482);
   U121 : INV_X1 port map( A => A_s(39), ZN => n481);
   U122 : INV_X1 port map( A => A_ns(39), ZN => n480);
   U123 : OAI221_X1 port map( B1 => n393, B2 => n483, C1 => n392, C2 => n484, A
                           => n485, ZN => O_40_port);
   U124 : AOI22_X1 port map( A1 => A_ns(39), A2 => n397, B1 => A_s(39), B2 => 
                           n398, ZN => n485);
   U125 : INV_X1 port map( A => A_s(38), ZN => n484);
   U126 : INV_X1 port map( A => A_ns(38), ZN => n483);
   U127 : OAI221_X1 port map( B1 => n393, B2 => n486, C1 => n392, C2 => n487, A
                           => n488, ZN => O_3_port);
   U128 : AOI22_X1 port map( A1 => A_ns(2), A2 => n397, B1 => A_s(2), B2 => 
                           n398, ZN => n488);
   U129 : INV_X1 port map( A => A_s(1), ZN => n487);
   U130 : INV_X1 port map( A => A_ns(1), ZN => n486);
   U131 : OAI221_X1 port map( B1 => n393, B2 => n489, C1 => n392, C2 => n490, A
                           => n491, ZN => O_39_port);
   U132 : AOI22_X1 port map( A1 => A_ns(38), A2 => n397, B1 => A_s(38), B2 => 
                           n398, ZN => n491);
   U133 : INV_X1 port map( A => A_s(37), ZN => n490);
   U134 : INV_X1 port map( A => A_ns(37), ZN => n489);
   U135 : OAI221_X1 port map( B1 => n393, B2 => n492, C1 => n392, C2 => n493, A
                           => n494, ZN => O_38_port);
   U136 : AOI22_X1 port map( A1 => A_ns(37), A2 => n397, B1 => A_s(37), B2 => 
                           n398, ZN => n494);
   U137 : INV_X1 port map( A => A_s(36), ZN => n493);
   U138 : INV_X1 port map( A => A_ns(36), ZN => n492);
   U139 : OAI221_X1 port map( B1 => n393, B2 => n495, C1 => n392, C2 => n496, A
                           => n497, ZN => O_37_port);
   U140 : AOI22_X1 port map( A1 => A_ns(36), A2 => n397, B1 => A_s(36), B2 => 
                           n398, ZN => n497);
   U141 : INV_X1 port map( A => A_s(35), ZN => n496);
   U142 : INV_X1 port map( A => A_ns(35), ZN => n495);
   U143 : OAI221_X1 port map( B1 => n393, B2 => n498, C1 => n392, C2 => n499, A
                           => n500, ZN => O_36_port);
   U144 : AOI22_X1 port map( A1 => A_ns(35), A2 => n397, B1 => A_s(35), B2 => 
                           n398, ZN => n500);
   U145 : INV_X1 port map( A => A_s(34), ZN => n499);
   U146 : INV_X1 port map( A => A_ns(34), ZN => n498);
   U147 : OAI221_X1 port map( B1 => n393, B2 => n501, C1 => n392, C2 => n502, A
                           => n503, ZN => O_35_port);
   U148 : AOI22_X1 port map( A1 => A_ns(34), A2 => n397, B1 => A_s(34), B2 => 
                           n398, ZN => n503);
   U149 : INV_X1 port map( A => A_s(33), ZN => n502);
   U150 : INV_X1 port map( A => A_ns(33), ZN => n501);
   U151 : OAI221_X1 port map( B1 => n393, B2 => n504, C1 => n392, C2 => n505, A
                           => n506, ZN => O_34_port);
   U152 : AOI22_X1 port map( A1 => A_ns(33), A2 => n397, B1 => A_s(33), B2 => 
                           n398, ZN => n506);
   U153 : INV_X1 port map( A => A_s(32), ZN => n505);
   U154 : INV_X1 port map( A => A_ns(32), ZN => n504);
   U155 : OAI221_X1 port map( B1 => n393, B2 => n507, C1 => n392, C2 => n508, A
                           => n509, ZN => O_33_port);
   U156 : AOI22_X1 port map( A1 => A_ns(32), A2 => n397, B1 => A_s(32), B2 => 
                           n398, ZN => n509);
   U157 : INV_X1 port map( A => A_s(31), ZN => n508);
   U158 : INV_X1 port map( A => A_ns(31), ZN => n507);
   U159 : OAI221_X1 port map( B1 => n393, B2 => n510, C1 => n392, C2 => n511, A
                           => n512, ZN => O_32_port);
   U160 : AOI22_X1 port map( A1 => A_ns(31), A2 => n397, B1 => A_s(31), B2 => 
                           n398, ZN => n512);
   U161 : INV_X1 port map( A => A_s(30), ZN => n511);
   U162 : INV_X1 port map( A => A_ns(30), ZN => n510);
   U163 : OAI221_X1 port map( B1 => n393, B2 => n513, C1 => n392, C2 => n514, A
                           => n515, ZN => O_31_port);
   U164 : AOI22_X1 port map( A1 => A_ns(30), A2 => n397, B1 => A_s(30), B2 => 
                           n398, ZN => n515);
   U165 : INV_X1 port map( A => A_s(29), ZN => n514);
   U166 : INV_X1 port map( A => A_ns(29), ZN => n513);
   U167 : OAI221_X1 port map( B1 => n393, B2 => n516, C1 => n392, C2 => n517, A
                           => n518, ZN => O_30_port);
   U168 : AOI22_X1 port map( A1 => A_ns(29), A2 => n397, B1 => A_s(29), B2 => 
                           n398, ZN => n518);
   U169 : INV_X1 port map( A => A_s(28), ZN => n517);
   U170 : INV_X1 port map( A => A_ns(28), ZN => n516);
   U171 : OAI221_X1 port map( B1 => n393, B2 => n519, C1 => n392, C2 => n520, A
                           => n521, ZN => O_2_port);
   U172 : AOI22_X1 port map( A1 => A_ns(1), A2 => n397, B1 => A_s(1), B2 => 
                           n398, ZN => n521);
   U173 : OAI221_X1 port map( B1 => n393, B2 => n522, C1 => n392, C2 => n523, A
                           => n524, ZN => O_29_port);
   U174 : AOI22_X1 port map( A1 => A_ns(28), A2 => n397, B1 => A_s(28), B2 => 
                           n398, ZN => n524);
   U175 : INV_X1 port map( A => A_s(27), ZN => n523);
   U176 : INV_X1 port map( A => A_ns(27), ZN => n522);
   U177 : OAI221_X1 port map( B1 => n393, B2 => n525, C1 => n392, C2 => n526, A
                           => n527, ZN => O_28_port);
   U178 : AOI22_X1 port map( A1 => A_ns(27), A2 => n397, B1 => A_s(27), B2 => 
                           n398, ZN => n527);
   U179 : INV_X1 port map( A => A_s(26), ZN => n526);
   U180 : INV_X1 port map( A => A_ns(26), ZN => n525);
   U181 : OAI221_X1 port map( B1 => n393, B2 => n528, C1 => n392, C2 => n529, A
                           => n530, ZN => O_27_port);
   U182 : AOI22_X1 port map( A1 => A_ns(26), A2 => n397, B1 => A_s(26), B2 => 
                           n398, ZN => n530);
   U183 : INV_X1 port map( A => A_s(25), ZN => n529);
   U184 : INV_X1 port map( A => A_ns(25), ZN => n528);
   U185 : OAI221_X1 port map( B1 => n393, B2 => n531, C1 => n392, C2 => n532, A
                           => n533, ZN => O_26_port);
   U186 : AOI22_X1 port map( A1 => A_ns(25), A2 => n397, B1 => A_s(25), B2 => 
                           n398, ZN => n533);
   U187 : INV_X1 port map( A => A_s(24), ZN => n532);
   U188 : INV_X1 port map( A => A_ns(24), ZN => n531);
   U189 : OAI221_X1 port map( B1 => n393, B2 => n534, C1 => n392, C2 => n535, A
                           => n536, ZN => O_25_port);
   U190 : AOI22_X1 port map( A1 => A_ns(24), A2 => n397, B1 => A_s(24), B2 => 
                           n398, ZN => n536);
   U191 : INV_X1 port map( A => A_s(23), ZN => n535);
   U192 : INV_X1 port map( A => A_ns(23), ZN => n534);
   U193 : OAI221_X1 port map( B1 => n393, B2 => n537, C1 => n392, C2 => n538, A
                           => n539, ZN => O_24_port);
   U194 : AOI22_X1 port map( A1 => A_ns(23), A2 => n397, B1 => A_s(23), B2 => 
                           n398, ZN => n539);
   U195 : INV_X1 port map( A => A_s(22), ZN => n538);
   U196 : INV_X1 port map( A => A_ns(22), ZN => n537);
   U197 : OAI221_X1 port map( B1 => n393, B2 => n540, C1 => n392, C2 => n541, A
                           => n542, ZN => O_23_port);
   U198 : AOI22_X1 port map( A1 => A_ns(22), A2 => n397, B1 => A_s(22), B2 => 
                           n398, ZN => n542);
   U199 : INV_X1 port map( A => A_s(21), ZN => n541);
   U200 : INV_X1 port map( A => A_ns(21), ZN => n540);
   U201 : OAI221_X1 port map( B1 => n393, B2 => n543, C1 => n392, C2 => n544, A
                           => n545, ZN => O_22_port);
   U202 : AOI22_X1 port map( A1 => A_ns(21), A2 => n397, B1 => A_s(21), B2 => 
                           n398, ZN => n545);
   U203 : INV_X1 port map( A => A_s(20), ZN => n544);
   U204 : INV_X1 port map( A => A_ns(20), ZN => n543);
   U205 : OAI221_X1 port map( B1 => n393, B2 => n546, C1 => n392, C2 => n547, A
                           => n548, ZN => O_21_port);
   U206 : AOI22_X1 port map( A1 => A_ns(20), A2 => n397, B1 => A_s(20), B2 => 
                           n398, ZN => n548);
   U207 : INV_X1 port map( A => A_s(19), ZN => n547);
   U208 : INV_X1 port map( A => A_ns(19), ZN => n546);
   U209 : OAI221_X1 port map( B1 => n393, B2 => n549, C1 => n392, C2 => n550, A
                           => n551, ZN => O_20_port);
   U210 : AOI22_X1 port map( A1 => A_ns(19), A2 => n397, B1 => A_s(19), B2 => 
                           n398, ZN => n551);
   U211 : INV_X1 port map( A => A_s(18), ZN => n550);
   U212 : INV_X1 port map( A => A_ns(18), ZN => n549);
   U213 : OAI22_X1 port map( A1 => n552, A2 => n520, B1 => n553, B2 => n519, ZN
                           => O_1_port);
   U214 : INV_X1 port map( A => A_ns(0), ZN => n519);
   U215 : INV_X1 port map( A => A_s(0), ZN => n520);
   U216 : OAI221_X1 port map( B1 => n393, B2 => n554, C1 => n392, C2 => n555, A
                           => n556, ZN => O_19_port);
   U217 : AOI22_X1 port map( A1 => A_ns(18), A2 => n397, B1 => A_s(18), B2 => 
                           n398, ZN => n556);
   U218 : INV_X1 port map( A => A_s(17), ZN => n555);
   U219 : INV_X1 port map( A => A_ns(17), ZN => n554);
   U220 : OAI221_X1 port map( B1 => n393, B2 => n557, C1 => n392, C2 => n558, A
                           => n559, ZN => O_18_port);
   U221 : AOI22_X1 port map( A1 => A_ns(17), A2 => n397, B1 => A_s(17), B2 => 
                           n398, ZN => n559);
   U222 : INV_X1 port map( A => A_s(16), ZN => n558);
   U223 : INV_X1 port map( A => A_ns(16), ZN => n557);
   U224 : OAI221_X1 port map( B1 => n393, B2 => n560, C1 => n392, C2 => n561, A
                           => n562, ZN => O_17_port);
   U225 : AOI22_X1 port map( A1 => A_ns(16), A2 => n397, B1 => A_s(16), B2 => 
                           n398, ZN => n562);
   U226 : INV_X1 port map( A => A_s(15), ZN => n561);
   U227 : INV_X1 port map( A => A_ns(15), ZN => n560);
   U228 : OAI221_X1 port map( B1 => n393, B2 => n563, C1 => n392, C2 => n564, A
                           => n565, ZN => O_16_port);
   U229 : AOI22_X1 port map( A1 => A_ns(15), A2 => n397, B1 => A_s(15), B2 => 
                           n398, ZN => n565);
   U230 : INV_X1 port map( A => A_s(14), ZN => n564);
   U231 : INV_X1 port map( A => A_ns(14), ZN => n563);
   U232 : OAI221_X1 port map( B1 => n393, B2 => n566, C1 => n392, C2 => n567, A
                           => n568, ZN => O_15_port);
   U233 : AOI22_X1 port map( A1 => A_ns(14), A2 => n397, B1 => A_s(14), B2 => 
                           n398, ZN => n568);
   U234 : INV_X1 port map( A => A_s(13), ZN => n567);
   U235 : INV_X1 port map( A => A_ns(13), ZN => n566);
   U236 : OAI221_X1 port map( B1 => n393, B2 => n569, C1 => n392, C2 => n570, A
                           => n571, ZN => O_14_port);
   U237 : AOI22_X1 port map( A1 => A_ns(13), A2 => n397, B1 => A_s(13), B2 => 
                           n398, ZN => n571);
   U238 : INV_X1 port map( A => A_s(12), ZN => n570);
   U239 : INV_X1 port map( A => A_ns(12), ZN => n569);
   U240 : OAI221_X1 port map( B1 => n393, B2 => n572, C1 => n392, C2 => n573, A
                           => n574, ZN => O_13_port);
   U241 : AOI22_X1 port map( A1 => A_ns(12), A2 => n397, B1 => A_s(12), B2 => 
                           n398, ZN => n574);
   U242 : INV_X1 port map( A => A_s(11), ZN => n573);
   U243 : INV_X1 port map( A => A_ns(11), ZN => n572);
   U244 : OAI221_X1 port map( B1 => n393, B2 => n575, C1 => n392, C2 => n576, A
                           => n577, ZN => O_12_port);
   U245 : AOI22_X1 port map( A1 => A_ns(11), A2 => n397, B1 => A_s(11), B2 => 
                           n398, ZN => n577);
   U246 : INV_X1 port map( A => A_s(10), ZN => n576);
   U247 : INV_X1 port map( A => A_ns(10), ZN => n575);
   U248 : OAI221_X1 port map( B1 => n393, B2 => n578, C1 => n392, C2 => n579, A
                           => n580, ZN => O_11_port);
   U249 : AOI22_X1 port map( A1 => A_ns(10), A2 => n397, B1 => A_s(10), B2 => 
                           n398, ZN => n580);
   U250 : INV_X1 port map( A => A_s(9), ZN => n579);
   U251 : INV_X1 port map( A => A_ns(9), ZN => n578);
   U252 : OAI221_X1 port map( B1 => n581, B2 => n393, C1 => n582, C2 => n392, A
                           => n583, ZN => O_10_port);
   U253 : AOI22_X1 port map( A1 => A_ns(9), A2 => n397, B1 => A_s(9), B2 => 
                           n398, ZN => n583);
   U254 : NAND2_X1 port map( A1 => n584, A2 => n552, ZN => n553);
   U255 : NAND2_X1 port map( A1 => n584, A2 => n585, ZN => n552);
   U256 : XOR2_X1 port map( A => B(3), B => B(4), Z => n584);
   U257 : INV_X1 port map( A => A_s(8), ZN => n582);
   U258 : INV_X1 port map( A => B(5), ZN => n585);
   U259 : INV_X1 port map( A => A_ns(8), ZN => n581);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity BOOTHENC_NBIT64_i2 is

   port( A, A_n, A_ns, A_s, B : in std_logic_vector (63 downto 0);  O, A_so, 
         A_nso : out std_logic_vector (63 downto 0));

end BOOTHENC_NBIT64_i2;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT64_i2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, O_63_port, O_62_port, O_61_port, O_60_port, O_59_port,
      O_58_port, O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, 
      O_52_port, O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, 
      O_46_port, O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, 
      O_40_port, O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, 
      O_34_port, O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, 
      O_28_port, O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, 
      O_22_port, O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, 
      O_16_port, O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, 
      O_10_port, O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, 
      O_3_port, O_2_port, O_1_port, n391, n392, n393, n394, n395, n396, n397, 
      n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, 
      n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, 
      n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, 
      n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, 
      n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, 
      n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, 
      n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, 
      n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, 
      n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, 
      n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, 
      n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, 
      n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, 
      n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, 
      n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, 
      n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, 
      n578, n579, n580, n581, n582, n583, n584, n585 : std_logic;

begin
   O <= ( O_63_port, O_62_port, O_61_port, O_60_port, O_59_port, O_58_port, 
      O_57_port, O_56_port, O_55_port, O_54_port, O_53_port, O_52_port, 
      O_51_port, O_50_port, O_49_port, O_48_port, O_47_port, O_46_port, 
      O_45_port, O_44_port, O_43_port, O_42_port, O_41_port, O_40_port, 
      O_39_port, O_38_port, O_37_port, O_36_port, O_35_port, O_34_port, 
      O_33_port, O_32_port, O_31_port, O_30_port, O_29_port, O_28_port, 
      O_27_port, O_26_port, O_25_port, O_24_port, O_23_port, O_22_port, 
      O_21_port, O_20_port, O_19_port, O_18_port, O_17_port, O_16_port, 
      O_15_port, O_14_port, O_13_port, O_12_port, O_11_port, O_10_port, 
      O_9_port, O_8_port, O_7_port, O_6_port, O_5_port, O_4_port, O_3_port, 
      O_2_port, O_1_port, X_Logic0_port );
   A_so <= ( A_s(61), A_s(60), A_s(59), A_s(58), A_s(57), A_s(56), A_s(55), 
      A_s(54), A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), 
      A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), 
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   A_nso <= ( A_s(61), A_s(60), A_s(59), A_s(58), A_s(57), A_s(56), A_s(55), 
      A_s(54), A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), A_s(47), 
      A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), A_s(39), 
      A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), A_s(31), 
      A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), A_s(23), 
      A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), A_s(15), 
      A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), A_s(7), 
      A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), X_Logic0_port, 
      X_Logic0_port );
   
   X_Logic0_port <= '0';
   U2 : AND3_X1 port map( A1 => B(2), A2 => n585, A3 => B(1), ZN => n391);
   U3 : INV_X4 port map( A => n391, ZN => n392);
   U4 : INV_X4 port map( A => n552, ZN => n398);
   U5 : OR3_X4 port map( A1 => B(1), A2 => B(2), A3 => n585, ZN => n393);
   U6 : INV_X4 port map( A => n553, ZN => n397);
   U7 : OAI221_X1 port map( B1 => n393, B2 => n394, C1 => n392, C2 => n395, A 
                           => n396, ZN => O_9_port);
   U8 : AOI22_X1 port map( A1 => A_ns(8), A2 => n397, B1 => A_s(8), B2 => n398,
                           ZN => n396);
   U9 : INV_X1 port map( A => A_s(7), ZN => n395);
   U10 : INV_X1 port map( A => A_ns(7), ZN => n394);
   U11 : OAI221_X1 port map( B1 => n393, B2 => n399, C1 => n392, C2 => n400, A 
                           => n401, ZN => O_8_port);
   U12 : AOI22_X1 port map( A1 => A_ns(7), A2 => n397, B1 => A_s(7), B2 => n398
                           , ZN => n401);
   U13 : INV_X1 port map( A => A_s(6), ZN => n400);
   U14 : INV_X1 port map( A => A_ns(6), ZN => n399);
   U15 : OAI221_X1 port map( B1 => n393, B2 => n402, C1 => n392, C2 => n403, A 
                           => n404, ZN => O_7_port);
   U16 : AOI22_X1 port map( A1 => A_ns(6), A2 => n397, B1 => A_s(6), B2 => n398
                           , ZN => n404);
   U17 : INV_X1 port map( A => A_s(5), ZN => n403);
   U18 : INV_X1 port map( A => A_ns(5), ZN => n402);
   U19 : OAI221_X1 port map( B1 => n393, B2 => n405, C1 => n392, C2 => n406, A 
                           => n407, ZN => O_6_port);
   U20 : AOI22_X1 port map( A1 => A_ns(5), A2 => n397, B1 => A_s(5), B2 => n398
                           , ZN => n407);
   U21 : INV_X1 port map( A => A_s(4), ZN => n406);
   U22 : INV_X1 port map( A => A_ns(4), ZN => n405);
   U23 : OAI221_X1 port map( B1 => n393, B2 => n408, C1 => n392, C2 => n409, A 
                           => n410, ZN => O_63_port);
   U24 : AOI22_X1 port map( A1 => A_ns(62), A2 => n397, B1 => A_s(62), B2 => 
                           n398, ZN => n410);
   U25 : INV_X1 port map( A => A_s(61), ZN => n409);
   U26 : INV_X1 port map( A => A_ns(61), ZN => n408);
   U27 : OAI221_X1 port map( B1 => n393, B2 => n411, C1 => n392, C2 => n412, A 
                           => n413, ZN => O_62_port);
   U28 : AOI22_X1 port map( A1 => A_ns(61), A2 => n397, B1 => A_s(61), B2 => 
                           n398, ZN => n413);
   U29 : INV_X1 port map( A => A_s(60), ZN => n412);
   U30 : INV_X1 port map( A => A_ns(60), ZN => n411);
   U31 : OAI221_X1 port map( B1 => n393, B2 => n414, C1 => n392, C2 => n415, A 
                           => n416, ZN => O_61_port);
   U32 : AOI22_X1 port map( A1 => A_ns(60), A2 => n397, B1 => A_s(60), B2 => 
                           n398, ZN => n416);
   U33 : INV_X1 port map( A => A_s(59), ZN => n415);
   U34 : INV_X1 port map( A => A_ns(59), ZN => n414);
   U35 : OAI221_X1 port map( B1 => n393, B2 => n417, C1 => n392, C2 => n418, A 
                           => n419, ZN => O_60_port);
   U36 : AOI22_X1 port map( A1 => A_ns(59), A2 => n397, B1 => A_s(59), B2 => 
                           n398, ZN => n419);
   U37 : INV_X1 port map( A => A_s(58), ZN => n418);
   U38 : INV_X1 port map( A => A_ns(58), ZN => n417);
   U39 : OAI221_X1 port map( B1 => n393, B2 => n420, C1 => n392, C2 => n421, A 
                           => n422, ZN => O_5_port);
   U40 : AOI22_X1 port map( A1 => A_ns(4), A2 => n397, B1 => A_s(4), B2 => n398
                           , ZN => n422);
   U41 : INV_X1 port map( A => A_s(3), ZN => n421);
   U42 : INV_X1 port map( A => A_ns(3), ZN => n420);
   U43 : OAI221_X1 port map( B1 => n393, B2 => n423, C1 => n392, C2 => n424, A 
                           => n425, ZN => O_59_port);
   U44 : AOI22_X1 port map( A1 => A_ns(58), A2 => n397, B1 => A_s(58), B2 => 
                           n398, ZN => n425);
   U45 : INV_X1 port map( A => A_s(57), ZN => n424);
   U46 : INV_X1 port map( A => A_ns(57), ZN => n423);
   U47 : OAI221_X1 port map( B1 => n393, B2 => n426, C1 => n392, C2 => n427, A 
                           => n428, ZN => O_58_port);
   U48 : AOI22_X1 port map( A1 => A_ns(57), A2 => n397, B1 => A_s(57), B2 => 
                           n398, ZN => n428);
   U49 : INV_X1 port map( A => A_s(56), ZN => n427);
   U50 : INV_X1 port map( A => A_ns(56), ZN => n426);
   U51 : OAI221_X1 port map( B1 => n393, B2 => n429, C1 => n392, C2 => n430, A 
                           => n431, ZN => O_57_port);
   U52 : AOI22_X1 port map( A1 => A_ns(56), A2 => n397, B1 => A_s(56), B2 => 
                           n398, ZN => n431);
   U53 : INV_X1 port map( A => A_s(55), ZN => n430);
   U54 : INV_X1 port map( A => A_ns(55), ZN => n429);
   U55 : OAI221_X1 port map( B1 => n393, B2 => n432, C1 => n392, C2 => n433, A 
                           => n434, ZN => O_56_port);
   U56 : AOI22_X1 port map( A1 => A_ns(55), A2 => n397, B1 => A_s(55), B2 => 
                           n398, ZN => n434);
   U57 : INV_X1 port map( A => A_s(54), ZN => n433);
   U58 : INV_X1 port map( A => A_ns(54), ZN => n432);
   U59 : OAI221_X1 port map( B1 => n393, B2 => n435, C1 => n392, C2 => n436, A 
                           => n437, ZN => O_55_port);
   U60 : AOI22_X1 port map( A1 => A_ns(54), A2 => n397, B1 => A_s(54), B2 => 
                           n398, ZN => n437);
   U61 : INV_X1 port map( A => A_s(53), ZN => n436);
   U62 : INV_X1 port map( A => A_ns(53), ZN => n435);
   U63 : OAI221_X1 port map( B1 => n393, B2 => n438, C1 => n392, C2 => n439, A 
                           => n440, ZN => O_54_port);
   U64 : AOI22_X1 port map( A1 => A_ns(53), A2 => n397, B1 => A_s(53), B2 => 
                           n398, ZN => n440);
   U65 : INV_X1 port map( A => A_s(52), ZN => n439);
   U66 : INV_X1 port map( A => A_ns(52), ZN => n438);
   U67 : OAI221_X1 port map( B1 => n393, B2 => n441, C1 => n392, C2 => n442, A 
                           => n443, ZN => O_53_port);
   U68 : AOI22_X1 port map( A1 => A_ns(52), A2 => n397, B1 => A_s(52), B2 => 
                           n398, ZN => n443);
   U69 : INV_X1 port map( A => A_s(51), ZN => n442);
   U70 : INV_X1 port map( A => A_ns(51), ZN => n441);
   U71 : OAI221_X1 port map( B1 => n393, B2 => n444, C1 => n392, C2 => n445, A 
                           => n446, ZN => O_52_port);
   U72 : AOI22_X1 port map( A1 => A_ns(51), A2 => n397, B1 => A_s(51), B2 => 
                           n398, ZN => n446);
   U73 : INV_X1 port map( A => A_s(50), ZN => n445);
   U74 : INV_X1 port map( A => A_ns(50), ZN => n444);
   U75 : OAI221_X1 port map( B1 => n393, B2 => n447, C1 => n392, C2 => n448, A 
                           => n449, ZN => O_51_port);
   U76 : AOI22_X1 port map( A1 => A_ns(50), A2 => n397, B1 => A_s(50), B2 => 
                           n398, ZN => n449);
   U77 : INV_X1 port map( A => A_s(49), ZN => n448);
   U78 : INV_X1 port map( A => A_ns(49), ZN => n447);
   U79 : OAI221_X1 port map( B1 => n393, B2 => n450, C1 => n392, C2 => n451, A 
                           => n452, ZN => O_50_port);
   U80 : AOI22_X1 port map( A1 => A_ns(49), A2 => n397, B1 => A_s(49), B2 => 
                           n398, ZN => n452);
   U81 : INV_X1 port map( A => A_s(48), ZN => n451);
   U82 : INV_X1 port map( A => A_ns(48), ZN => n450);
   U83 : OAI221_X1 port map( B1 => n393, B2 => n453, C1 => n392, C2 => n454, A 
                           => n455, ZN => O_4_port);
   U84 : AOI22_X1 port map( A1 => A_ns(3), A2 => n397, B1 => A_s(3), B2 => n398
                           , ZN => n455);
   U85 : INV_X1 port map( A => A_s(2), ZN => n454);
   U86 : INV_X1 port map( A => A_ns(2), ZN => n453);
   U87 : OAI221_X1 port map( B1 => n393, B2 => n456, C1 => n392, C2 => n457, A 
                           => n458, ZN => O_49_port);
   U88 : AOI22_X1 port map( A1 => A_ns(48), A2 => n397, B1 => A_s(48), B2 => 
                           n398, ZN => n458);
   U89 : INV_X1 port map( A => A_s(47), ZN => n457);
   U90 : INV_X1 port map( A => A_ns(47), ZN => n456);
   U91 : OAI221_X1 port map( B1 => n393, B2 => n459, C1 => n392, C2 => n460, A 
                           => n461, ZN => O_48_port);
   U92 : AOI22_X1 port map( A1 => A_ns(47), A2 => n397, B1 => A_s(47), B2 => 
                           n398, ZN => n461);
   U93 : INV_X1 port map( A => A_s(46), ZN => n460);
   U94 : INV_X1 port map( A => A_ns(46), ZN => n459);
   U95 : OAI221_X1 port map( B1 => n393, B2 => n462, C1 => n392, C2 => n463, A 
                           => n464, ZN => O_47_port);
   U96 : AOI22_X1 port map( A1 => A_ns(46), A2 => n397, B1 => A_s(46), B2 => 
                           n398, ZN => n464);
   U97 : INV_X1 port map( A => A_s(45), ZN => n463);
   U98 : INV_X1 port map( A => A_ns(45), ZN => n462);
   U99 : OAI221_X1 port map( B1 => n393, B2 => n465, C1 => n392, C2 => n466, A 
                           => n467, ZN => O_46_port);
   U100 : AOI22_X1 port map( A1 => A_ns(45), A2 => n397, B1 => A_s(45), B2 => 
                           n398, ZN => n467);
   U101 : INV_X1 port map( A => A_s(44), ZN => n466);
   U102 : INV_X1 port map( A => A_ns(44), ZN => n465);
   U103 : OAI221_X1 port map( B1 => n393, B2 => n468, C1 => n392, C2 => n469, A
                           => n470, ZN => O_45_port);
   U104 : AOI22_X1 port map( A1 => A_ns(44), A2 => n397, B1 => A_s(44), B2 => 
                           n398, ZN => n470);
   U105 : INV_X1 port map( A => A_s(43), ZN => n469);
   U106 : INV_X1 port map( A => A_ns(43), ZN => n468);
   U107 : OAI221_X1 port map( B1 => n393, B2 => n471, C1 => n392, C2 => n472, A
                           => n473, ZN => O_44_port);
   U108 : AOI22_X1 port map( A1 => A_ns(43), A2 => n397, B1 => A_s(43), B2 => 
                           n398, ZN => n473);
   U109 : INV_X1 port map( A => A_s(42), ZN => n472);
   U110 : INV_X1 port map( A => A_ns(42), ZN => n471);
   U111 : OAI221_X1 port map( B1 => n393, B2 => n474, C1 => n392, C2 => n475, A
                           => n476, ZN => O_43_port);
   U112 : AOI22_X1 port map( A1 => A_ns(42), A2 => n397, B1 => A_s(42), B2 => 
                           n398, ZN => n476);
   U113 : INV_X1 port map( A => A_s(41), ZN => n475);
   U114 : INV_X1 port map( A => A_ns(41), ZN => n474);
   U115 : OAI221_X1 port map( B1 => n393, B2 => n477, C1 => n392, C2 => n478, A
                           => n479, ZN => O_42_port);
   U116 : AOI22_X1 port map( A1 => A_ns(41), A2 => n397, B1 => A_s(41), B2 => 
                           n398, ZN => n479);
   U117 : INV_X1 port map( A => A_s(40), ZN => n478);
   U118 : INV_X1 port map( A => A_ns(40), ZN => n477);
   U119 : OAI221_X1 port map( B1 => n393, B2 => n480, C1 => n392, C2 => n481, A
                           => n482, ZN => O_41_port);
   U120 : AOI22_X1 port map( A1 => A_ns(40), A2 => n397, B1 => A_s(40), B2 => 
                           n398, ZN => n482);
   U121 : INV_X1 port map( A => A_s(39), ZN => n481);
   U122 : INV_X1 port map( A => A_ns(39), ZN => n480);
   U123 : OAI221_X1 port map( B1 => n393, B2 => n483, C1 => n392, C2 => n484, A
                           => n485, ZN => O_40_port);
   U124 : AOI22_X1 port map( A1 => A_ns(39), A2 => n397, B1 => A_s(39), B2 => 
                           n398, ZN => n485);
   U125 : INV_X1 port map( A => A_s(38), ZN => n484);
   U126 : INV_X1 port map( A => A_ns(38), ZN => n483);
   U127 : OAI221_X1 port map( B1 => n393, B2 => n486, C1 => n392, C2 => n487, A
                           => n488, ZN => O_3_port);
   U128 : AOI22_X1 port map( A1 => A_ns(2), A2 => n397, B1 => A_s(2), B2 => 
                           n398, ZN => n488);
   U129 : INV_X1 port map( A => A_s(1), ZN => n487);
   U130 : INV_X1 port map( A => A_ns(1), ZN => n486);
   U131 : OAI221_X1 port map( B1 => n393, B2 => n489, C1 => n392, C2 => n490, A
                           => n491, ZN => O_39_port);
   U132 : AOI22_X1 port map( A1 => A_ns(38), A2 => n397, B1 => A_s(38), B2 => 
                           n398, ZN => n491);
   U133 : INV_X1 port map( A => A_s(37), ZN => n490);
   U134 : INV_X1 port map( A => A_ns(37), ZN => n489);
   U135 : OAI221_X1 port map( B1 => n393, B2 => n492, C1 => n392, C2 => n493, A
                           => n494, ZN => O_38_port);
   U136 : AOI22_X1 port map( A1 => A_ns(37), A2 => n397, B1 => A_s(37), B2 => 
                           n398, ZN => n494);
   U137 : INV_X1 port map( A => A_s(36), ZN => n493);
   U138 : INV_X1 port map( A => A_ns(36), ZN => n492);
   U139 : OAI221_X1 port map( B1 => n393, B2 => n495, C1 => n392, C2 => n496, A
                           => n497, ZN => O_37_port);
   U140 : AOI22_X1 port map( A1 => A_ns(36), A2 => n397, B1 => A_s(36), B2 => 
                           n398, ZN => n497);
   U141 : INV_X1 port map( A => A_s(35), ZN => n496);
   U142 : INV_X1 port map( A => A_ns(35), ZN => n495);
   U143 : OAI221_X1 port map( B1 => n393, B2 => n498, C1 => n392, C2 => n499, A
                           => n500, ZN => O_36_port);
   U144 : AOI22_X1 port map( A1 => A_ns(35), A2 => n397, B1 => A_s(35), B2 => 
                           n398, ZN => n500);
   U145 : INV_X1 port map( A => A_s(34), ZN => n499);
   U146 : INV_X1 port map( A => A_ns(34), ZN => n498);
   U147 : OAI221_X1 port map( B1 => n393, B2 => n501, C1 => n392, C2 => n502, A
                           => n503, ZN => O_35_port);
   U148 : AOI22_X1 port map( A1 => A_ns(34), A2 => n397, B1 => A_s(34), B2 => 
                           n398, ZN => n503);
   U149 : INV_X1 port map( A => A_s(33), ZN => n502);
   U150 : INV_X1 port map( A => A_ns(33), ZN => n501);
   U151 : OAI221_X1 port map( B1 => n393, B2 => n504, C1 => n392, C2 => n505, A
                           => n506, ZN => O_34_port);
   U152 : AOI22_X1 port map( A1 => A_ns(33), A2 => n397, B1 => A_s(33), B2 => 
                           n398, ZN => n506);
   U153 : INV_X1 port map( A => A_s(32), ZN => n505);
   U154 : INV_X1 port map( A => A_ns(32), ZN => n504);
   U155 : OAI221_X1 port map( B1 => n393, B2 => n507, C1 => n392, C2 => n508, A
                           => n509, ZN => O_33_port);
   U156 : AOI22_X1 port map( A1 => A_ns(32), A2 => n397, B1 => A_s(32), B2 => 
                           n398, ZN => n509);
   U157 : INV_X1 port map( A => A_s(31), ZN => n508);
   U158 : INV_X1 port map( A => A_ns(31), ZN => n507);
   U159 : OAI221_X1 port map( B1 => n393, B2 => n510, C1 => n392, C2 => n511, A
                           => n512, ZN => O_32_port);
   U160 : AOI22_X1 port map( A1 => A_ns(31), A2 => n397, B1 => A_s(31), B2 => 
                           n398, ZN => n512);
   U161 : INV_X1 port map( A => A_s(30), ZN => n511);
   U162 : INV_X1 port map( A => A_ns(30), ZN => n510);
   U163 : OAI221_X1 port map( B1 => n393, B2 => n513, C1 => n392, C2 => n514, A
                           => n515, ZN => O_31_port);
   U164 : AOI22_X1 port map( A1 => A_ns(30), A2 => n397, B1 => A_s(30), B2 => 
                           n398, ZN => n515);
   U165 : INV_X1 port map( A => A_s(29), ZN => n514);
   U166 : INV_X1 port map( A => A_ns(29), ZN => n513);
   U167 : OAI221_X1 port map( B1 => n393, B2 => n516, C1 => n392, C2 => n517, A
                           => n518, ZN => O_30_port);
   U168 : AOI22_X1 port map( A1 => A_ns(29), A2 => n397, B1 => A_s(29), B2 => 
                           n398, ZN => n518);
   U169 : INV_X1 port map( A => A_s(28), ZN => n517);
   U170 : INV_X1 port map( A => A_ns(28), ZN => n516);
   U171 : OAI221_X1 port map( B1 => n393, B2 => n519, C1 => n392, C2 => n520, A
                           => n521, ZN => O_2_port);
   U172 : AOI22_X1 port map( A1 => A_ns(1), A2 => n397, B1 => A_s(1), B2 => 
                           n398, ZN => n521);
   U173 : OAI221_X1 port map( B1 => n393, B2 => n522, C1 => n392, C2 => n523, A
                           => n524, ZN => O_29_port);
   U174 : AOI22_X1 port map( A1 => A_ns(28), A2 => n397, B1 => A_s(28), B2 => 
                           n398, ZN => n524);
   U175 : INV_X1 port map( A => A_s(27), ZN => n523);
   U176 : INV_X1 port map( A => A_ns(27), ZN => n522);
   U177 : OAI221_X1 port map( B1 => n393, B2 => n525, C1 => n392, C2 => n526, A
                           => n527, ZN => O_28_port);
   U178 : AOI22_X1 port map( A1 => A_ns(27), A2 => n397, B1 => A_s(27), B2 => 
                           n398, ZN => n527);
   U179 : INV_X1 port map( A => A_s(26), ZN => n526);
   U180 : INV_X1 port map( A => A_ns(26), ZN => n525);
   U181 : OAI221_X1 port map( B1 => n393, B2 => n528, C1 => n392, C2 => n529, A
                           => n530, ZN => O_27_port);
   U182 : AOI22_X1 port map( A1 => A_ns(26), A2 => n397, B1 => A_s(26), B2 => 
                           n398, ZN => n530);
   U183 : INV_X1 port map( A => A_s(25), ZN => n529);
   U184 : INV_X1 port map( A => A_ns(25), ZN => n528);
   U185 : OAI221_X1 port map( B1 => n393, B2 => n531, C1 => n392, C2 => n532, A
                           => n533, ZN => O_26_port);
   U186 : AOI22_X1 port map( A1 => A_ns(25), A2 => n397, B1 => A_s(25), B2 => 
                           n398, ZN => n533);
   U187 : INV_X1 port map( A => A_s(24), ZN => n532);
   U188 : INV_X1 port map( A => A_ns(24), ZN => n531);
   U189 : OAI221_X1 port map( B1 => n393, B2 => n534, C1 => n392, C2 => n535, A
                           => n536, ZN => O_25_port);
   U190 : AOI22_X1 port map( A1 => A_ns(24), A2 => n397, B1 => A_s(24), B2 => 
                           n398, ZN => n536);
   U191 : INV_X1 port map( A => A_s(23), ZN => n535);
   U192 : INV_X1 port map( A => A_ns(23), ZN => n534);
   U193 : OAI221_X1 port map( B1 => n393, B2 => n537, C1 => n392, C2 => n538, A
                           => n539, ZN => O_24_port);
   U194 : AOI22_X1 port map( A1 => A_ns(23), A2 => n397, B1 => A_s(23), B2 => 
                           n398, ZN => n539);
   U195 : INV_X1 port map( A => A_s(22), ZN => n538);
   U196 : INV_X1 port map( A => A_ns(22), ZN => n537);
   U197 : OAI221_X1 port map( B1 => n393, B2 => n540, C1 => n392, C2 => n541, A
                           => n542, ZN => O_23_port);
   U198 : AOI22_X1 port map( A1 => A_ns(22), A2 => n397, B1 => A_s(22), B2 => 
                           n398, ZN => n542);
   U199 : INV_X1 port map( A => A_s(21), ZN => n541);
   U200 : INV_X1 port map( A => A_ns(21), ZN => n540);
   U201 : OAI221_X1 port map( B1 => n393, B2 => n543, C1 => n392, C2 => n544, A
                           => n545, ZN => O_22_port);
   U202 : AOI22_X1 port map( A1 => A_ns(21), A2 => n397, B1 => A_s(21), B2 => 
                           n398, ZN => n545);
   U203 : INV_X1 port map( A => A_s(20), ZN => n544);
   U204 : INV_X1 port map( A => A_ns(20), ZN => n543);
   U205 : OAI221_X1 port map( B1 => n393, B2 => n546, C1 => n392, C2 => n547, A
                           => n548, ZN => O_21_port);
   U206 : AOI22_X1 port map( A1 => A_ns(20), A2 => n397, B1 => A_s(20), B2 => 
                           n398, ZN => n548);
   U207 : INV_X1 port map( A => A_s(19), ZN => n547);
   U208 : INV_X1 port map( A => A_ns(19), ZN => n546);
   U209 : OAI221_X1 port map( B1 => n393, B2 => n549, C1 => n392, C2 => n550, A
                           => n551, ZN => O_20_port);
   U210 : AOI22_X1 port map( A1 => A_ns(19), A2 => n397, B1 => A_s(19), B2 => 
                           n398, ZN => n551);
   U211 : INV_X1 port map( A => A_s(18), ZN => n550);
   U212 : INV_X1 port map( A => A_ns(18), ZN => n549);
   U213 : OAI22_X1 port map( A1 => n552, A2 => n520, B1 => n553, B2 => n519, ZN
                           => O_1_port);
   U214 : INV_X1 port map( A => A_ns(0), ZN => n519);
   U215 : INV_X1 port map( A => A_s(0), ZN => n520);
   U216 : OAI221_X1 port map( B1 => n393, B2 => n554, C1 => n392, C2 => n555, A
                           => n556, ZN => O_19_port);
   U217 : AOI22_X1 port map( A1 => A_ns(18), A2 => n397, B1 => A_s(18), B2 => 
                           n398, ZN => n556);
   U218 : INV_X1 port map( A => A_s(17), ZN => n555);
   U219 : INV_X1 port map( A => A_ns(17), ZN => n554);
   U220 : OAI221_X1 port map( B1 => n393, B2 => n557, C1 => n392, C2 => n558, A
                           => n559, ZN => O_18_port);
   U221 : AOI22_X1 port map( A1 => A_ns(17), A2 => n397, B1 => A_s(17), B2 => 
                           n398, ZN => n559);
   U222 : INV_X1 port map( A => A_s(16), ZN => n558);
   U223 : INV_X1 port map( A => A_ns(16), ZN => n557);
   U224 : OAI221_X1 port map( B1 => n393, B2 => n560, C1 => n392, C2 => n561, A
                           => n562, ZN => O_17_port);
   U225 : AOI22_X1 port map( A1 => A_ns(16), A2 => n397, B1 => A_s(16), B2 => 
                           n398, ZN => n562);
   U226 : INV_X1 port map( A => A_s(15), ZN => n561);
   U227 : INV_X1 port map( A => A_ns(15), ZN => n560);
   U228 : OAI221_X1 port map( B1 => n393, B2 => n563, C1 => n392, C2 => n564, A
                           => n565, ZN => O_16_port);
   U229 : AOI22_X1 port map( A1 => A_ns(15), A2 => n397, B1 => A_s(15), B2 => 
                           n398, ZN => n565);
   U230 : INV_X1 port map( A => A_s(14), ZN => n564);
   U231 : INV_X1 port map( A => A_ns(14), ZN => n563);
   U232 : OAI221_X1 port map( B1 => n393, B2 => n566, C1 => n392, C2 => n567, A
                           => n568, ZN => O_15_port);
   U233 : AOI22_X1 port map( A1 => A_ns(14), A2 => n397, B1 => A_s(14), B2 => 
                           n398, ZN => n568);
   U234 : INV_X1 port map( A => A_s(13), ZN => n567);
   U235 : INV_X1 port map( A => A_ns(13), ZN => n566);
   U236 : OAI221_X1 port map( B1 => n393, B2 => n569, C1 => n392, C2 => n570, A
                           => n571, ZN => O_14_port);
   U237 : AOI22_X1 port map( A1 => A_ns(13), A2 => n397, B1 => A_s(13), B2 => 
                           n398, ZN => n571);
   U238 : INV_X1 port map( A => A_s(12), ZN => n570);
   U239 : INV_X1 port map( A => A_ns(12), ZN => n569);
   U240 : OAI221_X1 port map( B1 => n393, B2 => n572, C1 => n392, C2 => n573, A
                           => n574, ZN => O_13_port);
   U241 : AOI22_X1 port map( A1 => A_ns(12), A2 => n397, B1 => A_s(12), B2 => 
                           n398, ZN => n574);
   U242 : INV_X1 port map( A => A_s(11), ZN => n573);
   U243 : INV_X1 port map( A => A_ns(11), ZN => n572);
   U244 : OAI221_X1 port map( B1 => n393, B2 => n575, C1 => n392, C2 => n576, A
                           => n577, ZN => O_12_port);
   U245 : AOI22_X1 port map( A1 => A_ns(11), A2 => n397, B1 => A_s(11), B2 => 
                           n398, ZN => n577);
   U246 : INV_X1 port map( A => A_s(10), ZN => n576);
   U247 : INV_X1 port map( A => A_ns(10), ZN => n575);
   U248 : OAI221_X1 port map( B1 => n393, B2 => n578, C1 => n392, C2 => n579, A
                           => n580, ZN => O_11_port);
   U249 : AOI22_X1 port map( A1 => A_ns(10), A2 => n397, B1 => A_s(10), B2 => 
                           n398, ZN => n580);
   U250 : INV_X1 port map( A => A_s(9), ZN => n579);
   U251 : INV_X1 port map( A => A_ns(9), ZN => n578);
   U252 : OAI221_X1 port map( B1 => n581, B2 => n393, C1 => n582, C2 => n392, A
                           => n583, ZN => O_10_port);
   U253 : AOI22_X1 port map( A1 => A_ns(9), A2 => n397, B1 => A_s(9), B2 => 
                           n398, ZN => n583);
   U254 : NAND2_X1 port map( A1 => n584, A2 => n552, ZN => n553);
   U255 : NAND2_X1 port map( A1 => n584, A2 => n585, ZN => n552);
   U256 : XOR2_X1 port map( A => B(1), B => B(2), Z => n584);
   U257 : INV_X1 port map( A => A_s(8), ZN => n582);
   U258 : INV_X1 port map( A => B(3), ZN => n585);
   U259 : INV_X1 port map( A => A_ns(8), ZN => n581);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity BOOTHENC_NBIT64_i0 is

   port( A, A_n, A_ns, A_s, B : in std_logic_vector (63 downto 0);  O, A_so, 
         A_nso : out std_logic_vector (63 downto 0));

end BOOTHENC_NBIT64_i0;

architecture SYN_BEHAVIOURAL of BOOTHENC_NBIT64_i0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, n267, n268, n269, n270, n271, n272, n273, n274, n275, 
      n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, 
      n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, 
      n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, 
      n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, 
      n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, 
      n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, 
      n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, 
      n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, 
      n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, 
      n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, 
      n396, n397, n398, n399 : std_logic;

begin
   A_so <= ( A_s(62), A_s(61), A_s(60), A_s(59), A_s(58), A_s(57), A_s(56), 
      A_s(55), A_s(54), A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), 
      A_s(47), A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), 
      A_s(39), A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), 
      A_s(31), A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), 
      A_s(23), A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), 
      A_s(15), A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), 
      A_s(7), A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), 
      X_Logic0_port );
   A_nso <= ( A_s(62), A_s(61), A_s(60), A_s(59), A_s(58), A_s(57), A_s(56), 
      A_s(55), A_s(54), A_s(53), A_s(52), A_s(51), A_s(50), A_s(49), A_s(48), 
      A_s(47), A_s(46), A_s(45), A_s(44), A_s(43), A_s(42), A_s(41), A_s(40), 
      A_s(39), A_s(38), A_s(37), A_s(36), A_s(35), A_s(34), A_s(33), A_s(32), 
      A_s(31), A_s(30), A_s(29), A_s(28), A_s(27), A_s(26), A_s(25), A_s(24), 
      A_s(23), A_s(22), A_s(21), A_s(20), A_s(19), A_s(18), A_s(17), A_s(16), 
      A_s(15), A_s(14), A_s(13), A_s(12), A_s(11), A_s(10), A_s(9), A_s(8), 
      A_s(7), A_s(6), A_s(5), A_s(4), A_s(3), A_s(2), A_s(1), A_s(0), 
      X_Logic0_port );
   
   X_Logic0_port <= '0';
   U3 : INV_X4 port map( A => n280, ZN => n272);
   U4 : OR2_X4 port map( A1 => n398, A2 => B(0), ZN => n267);
   U5 : NAND2_X4 port map( A1 => B(0), A2 => n280, ZN => n269);
   U6 : OAI221_X1 port map( B1 => n267, B2 => n268, C1 => n269, C2 => n270, A 
                           => n271, ZN => O(9));
   U7 : NAND2_X1 port map( A1 => A_s(9), A2 => n272, ZN => n271);
   U8 : OAI221_X1 port map( B1 => n267, B2 => n273, C1 => n268, C2 => n269, A 
                           => n274, ZN => O(8));
   U9 : NAND2_X1 port map( A1 => A_s(8), A2 => n272, ZN => n274);
   U10 : INV_X1 port map( A => A_ns(8), ZN => n268);
   U11 : OAI221_X1 port map( B1 => n267, B2 => n275, C1 => n269, C2 => n273, A 
                           => n276, ZN => O(7));
   U12 : NAND2_X1 port map( A1 => A_s(7), A2 => n272, ZN => n276);
   U13 : INV_X1 port map( A => A_ns(7), ZN => n273);
   U14 : OAI221_X1 port map( B1 => n267, B2 => n277, C1 => n269, C2 => n275, A 
                           => n278, ZN => O(6));
   U15 : NAND2_X1 port map( A1 => A_s(6), A2 => n272, ZN => n278);
   U16 : INV_X1 port map( A => A_ns(6), ZN => n275);
   U17 : OAI222_X1 port map( A1 => n279, A2 => n280, B1 => n281, B2 => n267, C1
                           => n282, C2 => n269, ZN => O(63));
   U18 : INV_X1 port map( A => A_ns(63), ZN => n282);
   U19 : INV_X1 port map( A => A_s(63), ZN => n279);
   U20 : OAI221_X1 port map( B1 => n267, B2 => n283, C1 => n269, C2 => n281, A 
                           => n284, ZN => O(62));
   U21 : NAND2_X1 port map( A1 => A_s(62), A2 => n272, ZN => n284);
   U22 : INV_X1 port map( A => A_ns(62), ZN => n281);
   U23 : OAI221_X1 port map( B1 => n267, B2 => n285, C1 => n269, C2 => n283, A 
                           => n286, ZN => O(61));
   U24 : NAND2_X1 port map( A1 => A_s(61), A2 => n272, ZN => n286);
   U25 : INV_X1 port map( A => A_ns(61), ZN => n283);
   U26 : OAI221_X1 port map( B1 => n267, B2 => n287, C1 => n269, C2 => n285, A 
                           => n288, ZN => O(60));
   U27 : NAND2_X1 port map( A1 => A_s(60), A2 => n272, ZN => n288);
   U28 : INV_X1 port map( A => A_ns(60), ZN => n285);
   U29 : OAI221_X1 port map( B1 => n267, B2 => n289, C1 => n269, C2 => n277, A 
                           => n290, ZN => O(5));
   U30 : NAND2_X1 port map( A1 => A_s(5), A2 => n272, ZN => n290);
   U31 : INV_X1 port map( A => A_ns(5), ZN => n277);
   U32 : OAI221_X1 port map( B1 => n267, B2 => n291, C1 => n269, C2 => n287, A 
                           => n292, ZN => O(59));
   U33 : NAND2_X1 port map( A1 => A_s(59), A2 => n272, ZN => n292);
   U34 : INV_X1 port map( A => A_ns(59), ZN => n287);
   U35 : OAI221_X1 port map( B1 => n267, B2 => n293, C1 => n269, C2 => n291, A 
                           => n294, ZN => O(58));
   U36 : NAND2_X1 port map( A1 => A_s(58), A2 => n272, ZN => n294);
   U37 : INV_X1 port map( A => A_ns(58), ZN => n291);
   U38 : OAI221_X1 port map( B1 => n267, B2 => n295, C1 => n269, C2 => n293, A 
                           => n296, ZN => O(57));
   U39 : NAND2_X1 port map( A1 => A_s(57), A2 => n272, ZN => n296);
   U40 : INV_X1 port map( A => A_ns(57), ZN => n293);
   U41 : OAI221_X1 port map( B1 => n267, B2 => n297, C1 => n269, C2 => n295, A 
                           => n298, ZN => O(56));
   U42 : NAND2_X1 port map( A1 => A_s(56), A2 => n272, ZN => n298);
   U43 : INV_X1 port map( A => A_ns(56), ZN => n295);
   U44 : OAI221_X1 port map( B1 => n267, B2 => n299, C1 => n269, C2 => n297, A 
                           => n300, ZN => O(55));
   U45 : NAND2_X1 port map( A1 => A_s(55), A2 => n272, ZN => n300);
   U46 : INV_X1 port map( A => A_ns(55), ZN => n297);
   U47 : OAI221_X1 port map( B1 => n267, B2 => n301, C1 => n269, C2 => n299, A 
                           => n302, ZN => O(54));
   U48 : NAND2_X1 port map( A1 => A_s(54), A2 => n272, ZN => n302);
   U49 : INV_X1 port map( A => A_ns(54), ZN => n299);
   U50 : OAI221_X1 port map( B1 => n267, B2 => n303, C1 => n269, C2 => n301, A 
                           => n304, ZN => O(53));
   U51 : NAND2_X1 port map( A1 => A_s(53), A2 => n272, ZN => n304);
   U52 : INV_X1 port map( A => A_ns(53), ZN => n301);
   U53 : OAI221_X1 port map( B1 => n267, B2 => n305, C1 => n269, C2 => n303, A 
                           => n306, ZN => O(52));
   U54 : NAND2_X1 port map( A1 => A_s(52), A2 => n272, ZN => n306);
   U55 : INV_X1 port map( A => A_ns(52), ZN => n303);
   U56 : OAI221_X1 port map( B1 => n267, B2 => n307, C1 => n269, C2 => n305, A 
                           => n308, ZN => O(51));
   U57 : NAND2_X1 port map( A1 => A_s(51), A2 => n272, ZN => n308);
   U58 : INV_X1 port map( A => A_ns(51), ZN => n305);
   U59 : OAI221_X1 port map( B1 => n267, B2 => n309, C1 => n269, C2 => n307, A 
                           => n310, ZN => O(50));
   U60 : NAND2_X1 port map( A1 => A_s(50), A2 => n272, ZN => n310);
   U61 : INV_X1 port map( A => A_ns(50), ZN => n307);
   U62 : OAI221_X1 port map( B1 => n267, B2 => n311, C1 => n269, C2 => n289, A 
                           => n312, ZN => O(4));
   U63 : NAND2_X1 port map( A1 => A_s(4), A2 => n272, ZN => n312);
   U64 : INV_X1 port map( A => A_ns(4), ZN => n289);
   U65 : OAI221_X1 port map( B1 => n267, B2 => n313, C1 => n269, C2 => n309, A 
                           => n314, ZN => O(49));
   U66 : NAND2_X1 port map( A1 => A_s(49), A2 => n272, ZN => n314);
   U67 : INV_X1 port map( A => A_ns(49), ZN => n309);
   U68 : OAI221_X1 port map( B1 => n267, B2 => n315, C1 => n269, C2 => n313, A 
                           => n316, ZN => O(48));
   U69 : NAND2_X1 port map( A1 => A_s(48), A2 => n272, ZN => n316);
   U70 : INV_X1 port map( A => A_ns(48), ZN => n313);
   U71 : OAI221_X1 port map( B1 => n267, B2 => n317, C1 => n269, C2 => n315, A 
                           => n318, ZN => O(47));
   U72 : NAND2_X1 port map( A1 => A_s(47), A2 => n272, ZN => n318);
   U73 : INV_X1 port map( A => A_ns(47), ZN => n315);
   U74 : OAI221_X1 port map( B1 => n267, B2 => n319, C1 => n269, C2 => n317, A 
                           => n320, ZN => O(46));
   U75 : NAND2_X1 port map( A1 => A_s(46), A2 => n272, ZN => n320);
   U76 : INV_X1 port map( A => A_ns(46), ZN => n317);
   U77 : OAI221_X1 port map( B1 => n267, B2 => n321, C1 => n269, C2 => n319, A 
                           => n322, ZN => O(45));
   U78 : NAND2_X1 port map( A1 => A_s(45), A2 => n272, ZN => n322);
   U79 : INV_X1 port map( A => A_ns(45), ZN => n319);
   U80 : OAI221_X1 port map( B1 => n267, B2 => n323, C1 => n269, C2 => n321, A 
                           => n324, ZN => O(44));
   U81 : NAND2_X1 port map( A1 => A_s(44), A2 => n272, ZN => n324);
   U82 : INV_X1 port map( A => A_ns(44), ZN => n321);
   U83 : OAI221_X1 port map( B1 => n267, B2 => n325, C1 => n269, C2 => n323, A 
                           => n326, ZN => O(43));
   U84 : NAND2_X1 port map( A1 => A_s(43), A2 => n272, ZN => n326);
   U85 : INV_X1 port map( A => A_ns(43), ZN => n323);
   U86 : OAI221_X1 port map( B1 => n267, B2 => n327, C1 => n269, C2 => n325, A 
                           => n328, ZN => O(42));
   U87 : NAND2_X1 port map( A1 => A_s(42), A2 => n272, ZN => n328);
   U88 : INV_X1 port map( A => A_ns(42), ZN => n325);
   U89 : OAI221_X1 port map( B1 => n267, B2 => n329, C1 => n269, C2 => n327, A 
                           => n330, ZN => O(41));
   U90 : NAND2_X1 port map( A1 => A_s(41), A2 => n272, ZN => n330);
   U91 : INV_X1 port map( A => A_ns(41), ZN => n327);
   U92 : OAI221_X1 port map( B1 => n267, B2 => n331, C1 => n269, C2 => n329, A 
                           => n332, ZN => O(40));
   U93 : NAND2_X1 port map( A1 => A_s(40), A2 => n272, ZN => n332);
   U94 : INV_X1 port map( A => A_ns(40), ZN => n329);
   U95 : OAI221_X1 port map( B1 => n267, B2 => n333, C1 => n269, C2 => n311, A 
                           => n334, ZN => O(3));
   U96 : NAND2_X1 port map( A1 => A_s(3), A2 => n272, ZN => n334);
   U97 : INV_X1 port map( A => A_ns(3), ZN => n311);
   U98 : OAI221_X1 port map( B1 => n267, B2 => n335, C1 => n269, C2 => n331, A 
                           => n336, ZN => O(39));
   U99 : NAND2_X1 port map( A1 => A_s(39), A2 => n272, ZN => n336);
   U100 : INV_X1 port map( A => A_ns(39), ZN => n331);
   U101 : OAI221_X1 port map( B1 => n267, B2 => n337, C1 => n269, C2 => n335, A
                           => n338, ZN => O(38));
   U102 : NAND2_X1 port map( A1 => A_s(38), A2 => n272, ZN => n338);
   U103 : INV_X1 port map( A => A_ns(38), ZN => n335);
   U104 : OAI221_X1 port map( B1 => n267, B2 => n339, C1 => n269, C2 => n337, A
                           => n340, ZN => O(37));
   U105 : NAND2_X1 port map( A1 => A_s(37), A2 => n272, ZN => n340);
   U106 : INV_X1 port map( A => A_ns(37), ZN => n337);
   U107 : OAI221_X1 port map( B1 => n267, B2 => n341, C1 => n269, C2 => n339, A
                           => n342, ZN => O(36));
   U108 : NAND2_X1 port map( A1 => A_s(36), A2 => n272, ZN => n342);
   U109 : INV_X1 port map( A => A_ns(36), ZN => n339);
   U110 : OAI221_X1 port map( B1 => n267, B2 => n343, C1 => n269, C2 => n341, A
                           => n344, ZN => O(35));
   U111 : NAND2_X1 port map( A1 => A_s(35), A2 => n272, ZN => n344);
   U112 : INV_X1 port map( A => A_ns(35), ZN => n341);
   U113 : OAI221_X1 port map( B1 => n267, B2 => n345, C1 => n269, C2 => n343, A
                           => n346, ZN => O(34));
   U114 : NAND2_X1 port map( A1 => A_s(34), A2 => n272, ZN => n346);
   U115 : INV_X1 port map( A => A_ns(34), ZN => n343);
   U116 : OAI221_X1 port map( B1 => n267, B2 => n347, C1 => n269, C2 => n345, A
                           => n348, ZN => O(33));
   U117 : NAND2_X1 port map( A1 => A_s(33), A2 => n272, ZN => n348);
   U118 : INV_X1 port map( A => A_ns(33), ZN => n345);
   U119 : OAI221_X1 port map( B1 => n267, B2 => n349, C1 => n269, C2 => n347, A
                           => n350, ZN => O(32));
   U120 : NAND2_X1 port map( A1 => A_s(32), A2 => n272, ZN => n350);
   U121 : INV_X1 port map( A => A_ns(32), ZN => n347);
   U122 : OAI221_X1 port map( B1 => n267, B2 => n351, C1 => n269, C2 => n349, A
                           => n352, ZN => O(31));
   U123 : NAND2_X1 port map( A1 => A_s(31), A2 => n272, ZN => n352);
   U124 : INV_X1 port map( A => A_ns(31), ZN => n349);
   U125 : OAI221_X1 port map( B1 => n267, B2 => n353, C1 => n269, C2 => n351, A
                           => n354, ZN => O(30));
   U126 : NAND2_X1 port map( A1 => A_s(30), A2 => n272, ZN => n354);
   U127 : INV_X1 port map( A => A_ns(30), ZN => n351);
   U128 : OAI221_X1 port map( B1 => n267, B2 => n355, C1 => n269, C2 => n333, A
                           => n356, ZN => O(2));
   U129 : NAND2_X1 port map( A1 => A_s(2), A2 => n272, ZN => n356);
   U130 : INV_X1 port map( A => A_ns(2), ZN => n333);
   U131 : OAI221_X1 port map( B1 => n267, B2 => n357, C1 => n269, C2 => n353, A
                           => n358, ZN => O(29));
   U132 : NAND2_X1 port map( A1 => A_s(29), A2 => n272, ZN => n358);
   U133 : INV_X1 port map( A => A_ns(29), ZN => n353);
   U134 : OAI221_X1 port map( B1 => n267, B2 => n359, C1 => n269, C2 => n357, A
                           => n360, ZN => O(28));
   U135 : NAND2_X1 port map( A1 => A_s(28), A2 => n272, ZN => n360);
   U136 : INV_X1 port map( A => A_ns(28), ZN => n357);
   U137 : OAI221_X1 port map( B1 => n267, B2 => n361, C1 => n269, C2 => n359, A
                           => n362, ZN => O(27));
   U138 : NAND2_X1 port map( A1 => A_s(27), A2 => n272, ZN => n362);
   U139 : INV_X1 port map( A => A_ns(27), ZN => n359);
   U140 : OAI221_X1 port map( B1 => n267, B2 => n363, C1 => n269, C2 => n361, A
                           => n364, ZN => O(26));
   U141 : NAND2_X1 port map( A1 => A_s(26), A2 => n272, ZN => n364);
   U142 : INV_X1 port map( A => A_ns(26), ZN => n361);
   U143 : OAI221_X1 port map( B1 => n267, B2 => n365, C1 => n269, C2 => n363, A
                           => n366, ZN => O(25));
   U144 : NAND2_X1 port map( A1 => A_s(25), A2 => n272, ZN => n366);
   U145 : INV_X1 port map( A => A_ns(25), ZN => n363);
   U146 : OAI221_X1 port map( B1 => n267, B2 => n367, C1 => n269, C2 => n365, A
                           => n368, ZN => O(24));
   U147 : NAND2_X1 port map( A1 => A_s(24), A2 => n272, ZN => n368);
   U148 : INV_X1 port map( A => A_ns(24), ZN => n365);
   U149 : OAI221_X1 port map( B1 => n267, B2 => n369, C1 => n269, C2 => n367, A
                           => n370, ZN => O(23));
   U150 : NAND2_X1 port map( A1 => A_s(23), A2 => n272, ZN => n370);
   U151 : INV_X1 port map( A => A_ns(23), ZN => n367);
   U152 : OAI221_X1 port map( B1 => n267, B2 => n371, C1 => n269, C2 => n369, A
                           => n372, ZN => O(22));
   U153 : NAND2_X1 port map( A1 => A_s(22), A2 => n272, ZN => n372);
   U154 : INV_X1 port map( A => A_ns(22), ZN => n369);
   U155 : OAI221_X1 port map( B1 => n267, B2 => n373, C1 => n269, C2 => n371, A
                           => n374, ZN => O(21));
   U156 : NAND2_X1 port map( A1 => A_s(21), A2 => n272, ZN => n374);
   U157 : INV_X1 port map( A => A_ns(21), ZN => n371);
   U158 : OAI221_X1 port map( B1 => n267, B2 => n375, C1 => n269, C2 => n373, A
                           => n376, ZN => O(20));
   U159 : NAND2_X1 port map( A1 => A_s(20), A2 => n272, ZN => n376);
   U160 : INV_X1 port map( A => A_ns(20), ZN => n373);
   U161 : OAI221_X1 port map( B1 => n267, B2 => n377, C1 => n269, C2 => n355, A
                           => n378, ZN => O(1));
   U162 : NAND2_X1 port map( A1 => A_s(1), A2 => n272, ZN => n378);
   U163 : INV_X1 port map( A => A_ns(1), ZN => n355);
   U164 : OAI221_X1 port map( B1 => n267, B2 => n379, C1 => n269, C2 => n375, A
                           => n380, ZN => O(19));
   U165 : NAND2_X1 port map( A1 => A_s(19), A2 => n272, ZN => n380);
   U166 : INV_X1 port map( A => A_ns(19), ZN => n375);
   U167 : OAI221_X1 port map( B1 => n267, B2 => n381, C1 => n269, C2 => n379, A
                           => n382, ZN => O(18));
   U168 : NAND2_X1 port map( A1 => A_s(18), A2 => n272, ZN => n382);
   U169 : INV_X1 port map( A => A_ns(18), ZN => n379);
   U170 : OAI221_X1 port map( B1 => n267, B2 => n383, C1 => n269, C2 => n381, A
                           => n384, ZN => O(17));
   U171 : NAND2_X1 port map( A1 => A_s(17), A2 => n272, ZN => n384);
   U172 : INV_X1 port map( A => A_ns(17), ZN => n381);
   U173 : OAI221_X1 port map( B1 => n267, B2 => n385, C1 => n269, C2 => n383, A
                           => n386, ZN => O(16));
   U174 : NAND2_X1 port map( A1 => A_s(16), A2 => n272, ZN => n386);
   U175 : INV_X1 port map( A => A_ns(16), ZN => n383);
   U176 : OAI221_X1 port map( B1 => n267, B2 => n387, C1 => n269, C2 => n385, A
                           => n388, ZN => O(15));
   U177 : NAND2_X1 port map( A1 => A_s(15), A2 => n272, ZN => n388);
   U178 : INV_X1 port map( A => A_ns(15), ZN => n385);
   U179 : OAI221_X1 port map( B1 => n267, B2 => n389, C1 => n269, C2 => n387, A
                           => n390, ZN => O(14));
   U180 : NAND2_X1 port map( A1 => A_s(14), A2 => n272, ZN => n390);
   U181 : INV_X1 port map( A => A_ns(14), ZN => n387);
   U182 : OAI221_X1 port map( B1 => n267, B2 => n391, C1 => n269, C2 => n389, A
                           => n392, ZN => O(13));
   U183 : NAND2_X1 port map( A1 => A_s(13), A2 => n272, ZN => n392);
   U184 : INV_X1 port map( A => A_ns(13), ZN => n389);
   U185 : OAI221_X1 port map( B1 => n267, B2 => n393, C1 => n269, C2 => n391, A
                           => n394, ZN => O(12));
   U186 : NAND2_X1 port map( A1 => A_s(12), A2 => n272, ZN => n394);
   U187 : INV_X1 port map( A => A_ns(12), ZN => n391);
   U188 : OAI221_X1 port map( B1 => n267, B2 => n395, C1 => n269, C2 => n393, A
                           => n396, ZN => O(11));
   U189 : NAND2_X1 port map( A1 => A_s(11), A2 => n272, ZN => n396);
   U190 : INV_X1 port map( A => A_ns(11), ZN => n393);
   U191 : OAI221_X1 port map( B1 => n267, B2 => n270, C1 => n269, C2 => n395, A
                           => n397, ZN => O(10));
   U192 : NAND2_X1 port map( A1 => A_s(10), A2 => n272, ZN => n397);
   U193 : INV_X1 port map( A => A_ns(10), ZN => n395);
   U194 : INV_X1 port map( A => A_ns(9), ZN => n270);
   U195 : OAI22_X1 port map( A1 => n280, A2 => n399, B1 => n269, B2 => n377, ZN
                           => O(0));
   U196 : INV_X1 port map( A => A_ns(0), ZN => n377);
   U197 : INV_X1 port map( A => A_s(0), ZN => n399);
   U198 : NAND2_X1 port map( A1 => B(0), A2 => n398, ZN => n280);
   U199 : INV_X1 port map( A => B(1), ZN => n398);

end SYN_BEHAVIOURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_NBIT32_1.all;

entity BOOTHMUL_NBIT32_1 is

   port( A, B : in std_logic_vector (31 downto 0);  S : out std_logic_vector 
         (63 downto 0));

end BOOTHMUL_NBIT32_1;

architecture SYN_BEHAVIOURAL of BOOTHMUL_NBIT32_1 is

   component BOOTHMUL_NBIT32_1_DW01_sub_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component RCA_NBIT64_16
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT64_17
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT64_18
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT64_19
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT64_20
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT64_21
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT64_22
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT64_23
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT64_24
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT64_25
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT64_26
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT64_27
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT64_28
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT64_29
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_NBIT64_15
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component BOOTHENC_NBIT64_i30
      port( A, A_n, A_ns, A_s, B : in std_logic_vector (63 downto 0);  O, A_so,
            A_nso : out std_logic_vector (63 downto 0));
   end component;
   
   component BOOTHENC_NBIT64_i28
      port( A, A_n, A_ns, A_s, B : in std_logic_vector (63 downto 0);  O, A_so,
            A_nso : out std_logic_vector (63 downto 0));
   end component;
   
   component BOOTHENC_NBIT64_i26
      port( A, A_n, A_ns, A_s, B : in std_logic_vector (63 downto 0);  O, A_so,
            A_nso : out std_logic_vector (63 downto 0));
   end component;
   
   component BOOTHENC_NBIT64_i24
      port( A, A_n, A_ns, A_s, B : in std_logic_vector (63 downto 0);  O, A_so,
            A_nso : out std_logic_vector (63 downto 0));
   end component;
   
   component BOOTHENC_NBIT64_i22
      port( A, A_n, A_ns, A_s, B : in std_logic_vector (63 downto 0);  O, A_so,
            A_nso : out std_logic_vector (63 downto 0));
   end component;
   
   component BOOTHENC_NBIT64_i20
      port( A, A_n, A_ns, A_s, B : in std_logic_vector (63 downto 0);  O, A_so,
            A_nso : out std_logic_vector (63 downto 0));
   end component;
   
   component BOOTHENC_NBIT64_i18
      port( A, A_n, A_ns, A_s, B : in std_logic_vector (63 downto 0);  O, A_so,
            A_nso : out std_logic_vector (63 downto 0));
   end component;
   
   component BOOTHENC_NBIT64_i16
      port( A, A_n, A_ns, A_s, B : in std_logic_vector (63 downto 0);  O, A_so,
            A_nso : out std_logic_vector (63 downto 0));
   end component;
   
   component BOOTHENC_NBIT64_i14
      port( A, A_n, A_ns, A_s, B : in std_logic_vector (63 downto 0);  O, A_so,
            A_nso : out std_logic_vector (63 downto 0));
   end component;
   
   component BOOTHENC_NBIT64_i12
      port( A, A_n, A_ns, A_s, B : in std_logic_vector (63 downto 0);  O, A_so,
            A_nso : out std_logic_vector (63 downto 0));
   end component;
   
   component BOOTHENC_NBIT64_i10
      port( A, A_n, A_ns, A_s, B : in std_logic_vector (63 downto 0);  O, A_so,
            A_nso : out std_logic_vector (63 downto 0));
   end component;
   
   component BOOTHENC_NBIT64_i8
      port( A, A_n, A_ns, A_s, B : in std_logic_vector (63 downto 0);  O, A_so,
            A_nso : out std_logic_vector (63 downto 0));
   end component;
   
   component BOOTHENC_NBIT64_i6
      port( A, A_n, A_ns, A_s, B : in std_logic_vector (63 downto 0);  O, A_so,
            A_nso : out std_logic_vector (63 downto 0));
   end component;
   
   component BOOTHENC_NBIT64_i4
      port( A, A_n, A_ns, A_s, B : in std_logic_vector (63 downto 0);  O, A_so,
            A_nso : out std_logic_vector (63 downto 0));
   end component;
   
   component BOOTHENC_NBIT64_i2
      port( A, A_n, A_ns, A_s, B : in std_logic_vector (63 downto 0);  O, A_so,
            A_nso : out std_logic_vector (63 downto 0));
   end component;
   
   component BOOTHENC_NBIT64_i0
      port( A, A_n, A_ns, A_s, B : in std_logic_vector (63 downto 0);  O, A_so,
            A_nso : out std_logic_vector (63 downto 0));
   end component;
   
   signal X_Logic0_port, A_n_63, A_n_30_port, A_n_29_port, A_n_28_port, 
      A_n_27_port, A_n_26_port, A_n_25_port, A_n_24_port, A_n_23_port, 
      A_n_22_port, A_n_21_port, A_n_20_port, A_n_19_port, A_n_18_port, 
      A_n_17_port, A_n_16_port, A_n_15_port, A_n_14_port, A_n_13_port, 
      A_n_12_port, A_n_11_port, A_n_10_port, A_n_9_port, A_n_8_port, A_n_7_port
      , A_n_6_port, A_n_5_port, A_n_4_port, A_n_3_port, A_n_2_port, A_n_1_port,
      A_n_0_port, SHIFT_1023_port, SHIFT_1022_port, SHIFT_1021_port, 
      SHIFT_1020_port, SHIFT_1019_port, SHIFT_1018_port, SHIFT_1017_port, 
      SHIFT_1016_port, SHIFT_1015_port, SHIFT_1014_port, SHIFT_1013_port, 
      SHIFT_1012_port, SHIFT_1011_port, SHIFT_1010_port, SHIFT_1009_port, 
      SHIFT_1008_port, SHIFT_1007_port, SHIFT_1006_port, SHIFT_1005_port, 
      SHIFT_1004_port, SHIFT_1003_port, SHIFT_1002_port, SHIFT_1001_port, 
      SHIFT_1000_port, SHIFT_999_port, SHIFT_998_port, SHIFT_997_port, 
      SHIFT_996_port, SHIFT_995_port, SHIFT_994_port, SHIFT_993_port, 
      SHIFT_992_port, SHIFT_991_port, SHIFT_990_port, SHIFT_989_port, 
      SHIFT_988_port, SHIFT_987_port, SHIFT_986_port, SHIFT_985_port, 
      SHIFT_984_port, SHIFT_983_port, SHIFT_982_port, SHIFT_981_port, 
      SHIFT_980_port, SHIFT_979_port, SHIFT_978_port, SHIFT_977_port, 
      SHIFT_976_port, SHIFT_975_port, SHIFT_974_port, SHIFT_973_port, 
      SHIFT_972_port, SHIFT_971_port, SHIFT_970_port, SHIFT_969_port, 
      SHIFT_968_port, SHIFT_967_port, SHIFT_966_port, SHIFT_965_port, 
      SHIFT_964_port, SHIFT_963_port, SHIFT_962_port, SHIFT_961_port, 
      SHIFT_960_port, SHIFT_959_port, SHIFT_958_port, SHIFT_957_port, 
      SHIFT_956_port, SHIFT_955_port, SHIFT_954_port, SHIFT_953_port, 
      SHIFT_952_port, SHIFT_951_port, SHIFT_950_port, SHIFT_949_port, 
      SHIFT_948_port, SHIFT_947_port, SHIFT_946_port, SHIFT_945_port, 
      SHIFT_944_port, SHIFT_943_port, SHIFT_942_port, SHIFT_941_port, 
      SHIFT_940_port, SHIFT_939_port, SHIFT_938_port, SHIFT_937_port, 
      SHIFT_936_port, SHIFT_935_port, SHIFT_934_port, SHIFT_933_port, 
      SHIFT_932_port, SHIFT_931_port, SHIFT_930_port, SHIFT_929_port, 
      SHIFT_928_port, SHIFT_927_port, SHIFT_926_port, SHIFT_925_port, 
      SHIFT_924_port, SHIFT_923_port, SHIFT_922_port, SHIFT_921_port, 
      SHIFT_920_port, SHIFT_919_port, SHIFT_918_port, SHIFT_917_port, 
      SHIFT_916_port, SHIFT_915_port, SHIFT_914_port, SHIFT_913_port, 
      SHIFT_912_port, SHIFT_911_port, SHIFT_910_port, SHIFT_909_port, 
      SHIFT_908_port, SHIFT_907_port, SHIFT_906_port, SHIFT_905_port, 
      SHIFT_904_port, SHIFT_903_port, SHIFT_902_port, SHIFT_901_port, 
      SHIFT_900_port, SHIFT_899_port, SHIFT_898_port, SHIFT_897_port, 
      SHIFT_896_port, SHIFT_895_port, SHIFT_894_port, SHIFT_893_port, 
      SHIFT_892_port, SHIFT_891_port, SHIFT_890_port, SHIFT_889_port, 
      SHIFT_888_port, SHIFT_887_port, SHIFT_886_port, SHIFT_885_port, 
      SHIFT_884_port, SHIFT_883_port, SHIFT_882_port, SHIFT_881_port, 
      SHIFT_880_port, SHIFT_879_port, SHIFT_878_port, SHIFT_877_port, 
      SHIFT_876_port, SHIFT_875_port, SHIFT_874_port, SHIFT_873_port, 
      SHIFT_872_port, SHIFT_871_port, SHIFT_870_port, SHIFT_869_port, 
      SHIFT_868_port, SHIFT_867_port, SHIFT_866_port, SHIFT_865_port, 
      SHIFT_864_port, SHIFT_863_port, SHIFT_862_port, SHIFT_861_port, 
      SHIFT_860_port, SHIFT_859_port, SHIFT_858_port, SHIFT_857_port, 
      SHIFT_856_port, SHIFT_855_port, SHIFT_854_port, SHIFT_853_port, 
      SHIFT_852_port, SHIFT_851_port, SHIFT_850_port, SHIFT_849_port, 
      SHIFT_848_port, SHIFT_847_port, SHIFT_846_port, SHIFT_845_port, 
      SHIFT_844_port, SHIFT_843_port, SHIFT_842_port, SHIFT_841_port, 
      SHIFT_840_port, SHIFT_839_port, SHIFT_838_port, SHIFT_837_port, 
      SHIFT_836_port, SHIFT_835_port, SHIFT_834_port, SHIFT_833_port, 
      SHIFT_832_port, SHIFT_831_port, SHIFT_830_port, SHIFT_829_port, 
      SHIFT_828_port, SHIFT_827_port, SHIFT_826_port, SHIFT_825_port, 
      SHIFT_824_port, SHIFT_823_port, SHIFT_822_port, SHIFT_821_port, 
      SHIFT_820_port, SHIFT_819_port, SHIFT_818_port, SHIFT_817_port, 
      SHIFT_816_port, SHIFT_815_port, SHIFT_814_port, SHIFT_813_port, 
      SHIFT_812_port, SHIFT_811_port, SHIFT_810_port, SHIFT_809_port, 
      SHIFT_808_port, SHIFT_807_port, SHIFT_806_port, SHIFT_805_port, 
      SHIFT_804_port, SHIFT_803_port, SHIFT_802_port, SHIFT_801_port, 
      SHIFT_800_port, SHIFT_799_port, SHIFT_798_port, SHIFT_797_port, 
      SHIFT_796_port, SHIFT_795_port, SHIFT_794_port, SHIFT_793_port, 
      SHIFT_792_port, SHIFT_791_port, SHIFT_790_port, SHIFT_789_port, 
      SHIFT_788_port, SHIFT_787_port, SHIFT_786_port, SHIFT_785_port, 
      SHIFT_784_port, SHIFT_783_port, SHIFT_782_port, SHIFT_781_port, 
      SHIFT_780_port, SHIFT_779_port, SHIFT_778_port, SHIFT_777_port, 
      SHIFT_776_port, SHIFT_775_port, SHIFT_774_port, SHIFT_773_port, 
      SHIFT_772_port, SHIFT_771_port, SHIFT_770_port, SHIFT_769_port, 
      SHIFT_768_port, SHIFT_767_port, SHIFT_766_port, SHIFT_765_port, 
      SHIFT_764_port, SHIFT_763_port, SHIFT_762_port, SHIFT_761_port, 
      SHIFT_760_port, SHIFT_759_port, SHIFT_758_port, SHIFT_757_port, 
      SHIFT_756_port, SHIFT_755_port, SHIFT_754_port, SHIFT_753_port, 
      SHIFT_752_port, SHIFT_751_port, SHIFT_750_port, SHIFT_749_port, 
      SHIFT_748_port, SHIFT_747_port, SHIFT_746_port, SHIFT_745_port, 
      SHIFT_744_port, SHIFT_743_port, SHIFT_742_port, SHIFT_741_port, 
      SHIFT_740_port, SHIFT_739_port, SHIFT_738_port, SHIFT_737_port, 
      SHIFT_736_port, SHIFT_735_port, SHIFT_734_port, SHIFT_733_port, 
      SHIFT_732_port, SHIFT_731_port, SHIFT_730_port, SHIFT_729_port, 
      SHIFT_728_port, SHIFT_727_port, SHIFT_726_port, SHIFT_725_port, 
      SHIFT_724_port, SHIFT_723_port, SHIFT_722_port, SHIFT_721_port, 
      SHIFT_720_port, SHIFT_719_port, SHIFT_718_port, SHIFT_717_port, 
      SHIFT_716_port, SHIFT_715_port, SHIFT_714_port, SHIFT_713_port, 
      SHIFT_712_port, SHIFT_711_port, SHIFT_710_port, SHIFT_709_port, 
      SHIFT_708_port, SHIFT_707_port, SHIFT_706_port, SHIFT_705_port, 
      SHIFT_704_port, SHIFT_703_port, SHIFT_702_port, SHIFT_701_port, 
      SHIFT_700_port, SHIFT_699_port, SHIFT_698_port, SHIFT_697_port, 
      SHIFT_696_port, SHIFT_695_port, SHIFT_694_port, SHIFT_693_port, 
      SHIFT_692_port, SHIFT_691_port, SHIFT_690_port, SHIFT_689_port, 
      SHIFT_688_port, SHIFT_687_port, SHIFT_686_port, SHIFT_685_port, 
      SHIFT_684_port, SHIFT_683_port, SHIFT_682_port, SHIFT_681_port, 
      SHIFT_680_port, SHIFT_679_port, SHIFT_678_port, SHIFT_677_port, 
      SHIFT_676_port, SHIFT_675_port, SHIFT_674_port, SHIFT_673_port, 
      SHIFT_672_port, SHIFT_671_port, SHIFT_670_port, SHIFT_669_port, 
      SHIFT_668_port, SHIFT_667_port, SHIFT_666_port, SHIFT_665_port, 
      SHIFT_664_port, SHIFT_663_port, SHIFT_662_port, SHIFT_661_port, 
      SHIFT_660_port, SHIFT_659_port, SHIFT_658_port, SHIFT_657_port, 
      SHIFT_656_port, SHIFT_655_port, SHIFT_654_port, SHIFT_653_port, 
      SHIFT_652_port, SHIFT_651_port, SHIFT_650_port, SHIFT_649_port, 
      SHIFT_648_port, SHIFT_647_port, SHIFT_646_port, SHIFT_645_port, 
      SHIFT_644_port, SHIFT_643_port, SHIFT_642_port, SHIFT_641_port, 
      SHIFT_640_port, SHIFT_639_port, SHIFT_638_port, SHIFT_637_port, 
      SHIFT_636_port, SHIFT_635_port, SHIFT_634_port, SHIFT_633_port, 
      SHIFT_632_port, SHIFT_631_port, SHIFT_630_port, SHIFT_629_port, 
      SHIFT_628_port, SHIFT_627_port, SHIFT_626_port, SHIFT_625_port, 
      SHIFT_624_port, SHIFT_623_port, SHIFT_622_port, SHIFT_621_port, 
      SHIFT_620_port, SHIFT_619_port, SHIFT_618_port, SHIFT_617_port, 
      SHIFT_616_port, SHIFT_615_port, SHIFT_614_port, SHIFT_613_port, 
      SHIFT_612_port, SHIFT_611_port, SHIFT_610_port, SHIFT_609_port, 
      SHIFT_608_port, SHIFT_607_port, SHIFT_606_port, SHIFT_605_port, 
      SHIFT_604_port, SHIFT_603_port, SHIFT_602_port, SHIFT_601_port, 
      SHIFT_600_port, SHIFT_599_port, SHIFT_598_port, SHIFT_597_port, 
      SHIFT_596_port, SHIFT_595_port, SHIFT_594_port, SHIFT_593_port, 
      SHIFT_592_port, SHIFT_591_port, SHIFT_590_port, SHIFT_589_port, 
      SHIFT_588_port, SHIFT_587_port, SHIFT_586_port, SHIFT_585_port, 
      SHIFT_584_port, SHIFT_583_port, SHIFT_582_port, SHIFT_581_port, 
      SHIFT_580_port, SHIFT_579_port, SHIFT_578_port, SHIFT_577_port, 
      SHIFT_576_port, SHIFT_575_port, SHIFT_574_port, SHIFT_573_port, 
      SHIFT_572_port, SHIFT_571_port, SHIFT_570_port, SHIFT_569_port, 
      SHIFT_568_port, SHIFT_567_port, SHIFT_566_port, SHIFT_565_port, 
      SHIFT_564_port, SHIFT_563_port, SHIFT_562_port, SHIFT_561_port, 
      SHIFT_560_port, SHIFT_559_port, SHIFT_558_port, SHIFT_557_port, 
      SHIFT_556_port, SHIFT_555_port, SHIFT_554_port, SHIFT_553_port, 
      SHIFT_552_port, SHIFT_551_port, SHIFT_550_port, SHIFT_549_port, 
      SHIFT_548_port, SHIFT_547_port, SHIFT_546_port, SHIFT_545_port, 
      SHIFT_544_port, SHIFT_543_port, SHIFT_542_port, SHIFT_541_port, 
      SHIFT_540_port, SHIFT_539_port, SHIFT_538_port, SHIFT_537_port, 
      SHIFT_536_port, SHIFT_535_port, SHIFT_534_port, SHIFT_533_port, 
      SHIFT_532_port, SHIFT_531_port, SHIFT_530_port, SHIFT_529_port, 
      SHIFT_528_port, SHIFT_527_port, SHIFT_526_port, SHIFT_525_port, 
      SHIFT_524_port, SHIFT_523_port, SHIFT_522_port, SHIFT_521_port, 
      SHIFT_520_port, SHIFT_519_port, SHIFT_518_port, SHIFT_517_port, 
      SHIFT_516_port, SHIFT_515_port, SHIFT_514_port, SHIFT_513_port, 
      SHIFT_512_port, SHIFT_511_port, SHIFT_510_port, SHIFT_509_port, 
      SHIFT_508_port, SHIFT_507_port, SHIFT_506_port, SHIFT_505_port, 
      SHIFT_504_port, SHIFT_503_port, SHIFT_502_port, SHIFT_501_port, 
      SHIFT_500_port, SHIFT_499_port, SHIFT_498_port, SHIFT_497_port, 
      SHIFT_496_port, SHIFT_495_port, SHIFT_494_port, SHIFT_493_port, 
      SHIFT_492_port, SHIFT_491_port, SHIFT_490_port, SHIFT_489_port, 
      SHIFT_488_port, SHIFT_487_port, SHIFT_486_port, SHIFT_485_port, 
      SHIFT_484_port, SHIFT_483_port, SHIFT_482_port, SHIFT_481_port, 
      SHIFT_480_port, SHIFT_479_port, SHIFT_478_port, SHIFT_477_port, 
      SHIFT_476_port, SHIFT_475_port, SHIFT_474_port, SHIFT_473_port, 
      SHIFT_472_port, SHIFT_471_port, SHIFT_470_port, SHIFT_469_port, 
      SHIFT_468_port, SHIFT_467_port, SHIFT_466_port, SHIFT_465_port, 
      SHIFT_464_port, SHIFT_463_port, SHIFT_462_port, SHIFT_461_port, 
      SHIFT_460_port, SHIFT_459_port, SHIFT_458_port, SHIFT_457_port, 
      SHIFT_456_port, SHIFT_455_port, SHIFT_454_port, SHIFT_453_port, 
      SHIFT_452_port, SHIFT_451_port, SHIFT_450_port, SHIFT_449_port, 
      SHIFT_448_port, SHIFT_447_port, SHIFT_446_port, SHIFT_445_port, 
      SHIFT_444_port, SHIFT_443_port, SHIFT_442_port, SHIFT_441_port, 
      SHIFT_440_port, SHIFT_439_port, SHIFT_438_port, SHIFT_437_port, 
      SHIFT_436_port, SHIFT_435_port, SHIFT_434_port, SHIFT_433_port, 
      SHIFT_432_port, SHIFT_431_port, SHIFT_430_port, SHIFT_429_port, 
      SHIFT_428_port, SHIFT_427_port, SHIFT_426_port, SHIFT_425_port, 
      SHIFT_424_port, SHIFT_423_port, SHIFT_422_port, SHIFT_421_port, 
      SHIFT_420_port, SHIFT_419_port, SHIFT_418_port, SHIFT_417_port, 
      SHIFT_416_port, SHIFT_415_port, SHIFT_414_port, SHIFT_413_port, 
      SHIFT_412_port, SHIFT_411_port, SHIFT_410_port, SHIFT_409_port, 
      SHIFT_408_port, SHIFT_407_port, SHIFT_406_port, SHIFT_405_port, 
      SHIFT_404_port, SHIFT_403_port, SHIFT_402_port, SHIFT_401_port, 
      SHIFT_400_port, SHIFT_399_port, SHIFT_398_port, SHIFT_397_port, 
      SHIFT_396_port, SHIFT_395_port, SHIFT_394_port, SHIFT_393_port, 
      SHIFT_392_port, SHIFT_391_port, SHIFT_390_port, SHIFT_389_port, 
      SHIFT_388_port, SHIFT_387_port, SHIFT_386_port, SHIFT_385_port, 
      SHIFT_384_port, SHIFT_383_port, SHIFT_382_port, SHIFT_381_port, 
      SHIFT_380_port, SHIFT_379_port, SHIFT_378_port, SHIFT_377_port, 
      SHIFT_376_port, SHIFT_375_port, SHIFT_374_port, SHIFT_373_port, 
      SHIFT_372_port, SHIFT_371_port, SHIFT_370_port, SHIFT_369_port, 
      SHIFT_368_port, SHIFT_367_port, SHIFT_366_port, SHIFT_365_port, 
      SHIFT_364_port, SHIFT_363_port, SHIFT_362_port, SHIFT_361_port, 
      SHIFT_360_port, SHIFT_359_port, SHIFT_358_port, SHIFT_357_port, 
      SHIFT_356_port, SHIFT_355_port, SHIFT_354_port, SHIFT_353_port, 
      SHIFT_352_port, SHIFT_351_port, SHIFT_350_port, SHIFT_349_port, 
      SHIFT_348_port, SHIFT_347_port, SHIFT_346_port, SHIFT_345_port, 
      SHIFT_344_port, SHIFT_343_port, SHIFT_342_port, SHIFT_341_port, 
      SHIFT_340_port, SHIFT_339_port, SHIFT_338_port, SHIFT_337_port, 
      SHIFT_336_port, SHIFT_335_port, SHIFT_334_port, SHIFT_333_port, 
      SHIFT_332_port, SHIFT_331_port, SHIFT_330_port, SHIFT_329_port, 
      SHIFT_328_port, SHIFT_327_port, SHIFT_326_port, SHIFT_325_port, 
      SHIFT_324_port, SHIFT_323_port, SHIFT_322_port, SHIFT_321_port, 
      SHIFT_320_port, SHIFT_319_port, SHIFT_318_port, SHIFT_317_port, 
      SHIFT_316_port, SHIFT_315_port, SHIFT_314_port, SHIFT_313_port, 
      SHIFT_312_port, SHIFT_311_port, SHIFT_310_port, SHIFT_309_port, 
      SHIFT_308_port, SHIFT_307_port, SHIFT_306_port, SHIFT_305_port, 
      SHIFT_304_port, SHIFT_303_port, SHIFT_302_port, SHIFT_301_port, 
      SHIFT_300_port, SHIFT_299_port, SHIFT_298_port, SHIFT_297_port, 
      SHIFT_296_port, SHIFT_295_port, SHIFT_294_port, SHIFT_293_port, 
      SHIFT_292_port, SHIFT_291_port, SHIFT_290_port, SHIFT_289_port, 
      SHIFT_288_port, SHIFT_287_port, SHIFT_286_port, SHIFT_285_port, 
      SHIFT_284_port, SHIFT_283_port, SHIFT_282_port, SHIFT_281_port, 
      SHIFT_280_port, SHIFT_279_port, SHIFT_278_port, SHIFT_277_port, 
      SHIFT_276_port, SHIFT_275_port, SHIFT_274_port, SHIFT_273_port, 
      SHIFT_272_port, SHIFT_271_port, SHIFT_270_port, SHIFT_269_port, 
      SHIFT_268_port, SHIFT_267_port, SHIFT_266_port, SHIFT_265_port, 
      SHIFT_264_port, SHIFT_263_port, SHIFT_262_port, SHIFT_261_port, 
      SHIFT_260_port, SHIFT_259_port, SHIFT_258_port, SHIFT_257_port, 
      SHIFT_256_port, SHIFT_255_port, SHIFT_254_port, SHIFT_253_port, 
      SHIFT_252_port, SHIFT_251_port, SHIFT_250_port, SHIFT_249_port, 
      SHIFT_248_port, SHIFT_247_port, SHIFT_246_port, SHIFT_245_port, 
      SHIFT_244_port, SHIFT_243_port, SHIFT_242_port, SHIFT_241_port, 
      SHIFT_240_port, SHIFT_239_port, SHIFT_238_port, SHIFT_237_port, 
      SHIFT_236_port, SHIFT_235_port, SHIFT_234_port, SHIFT_233_port, 
      SHIFT_232_port, SHIFT_231_port, SHIFT_230_port, SHIFT_229_port, 
      SHIFT_228_port, SHIFT_227_port, SHIFT_226_port, SHIFT_225_port, 
      SHIFT_224_port, SHIFT_223_port, SHIFT_222_port, SHIFT_221_port, 
      SHIFT_220_port, SHIFT_219_port, SHIFT_218_port, SHIFT_217_port, 
      SHIFT_216_port, SHIFT_215_port, SHIFT_214_port, SHIFT_213_port, 
      SHIFT_212_port, SHIFT_211_port, SHIFT_210_port, SHIFT_209_port, 
      SHIFT_208_port, SHIFT_207_port, SHIFT_206_port, SHIFT_205_port, 
      SHIFT_204_port, SHIFT_203_port, SHIFT_202_port, SHIFT_201_port, 
      SHIFT_200_port, SHIFT_199_port, SHIFT_198_port, SHIFT_197_port, 
      SHIFT_196_port, SHIFT_195_port, SHIFT_194_port, SHIFT_193_port, 
      SHIFT_192_port, SHIFT_191_port, SHIFT_190_port, SHIFT_189_port, 
      SHIFT_188_port, SHIFT_187_port, SHIFT_186_port, SHIFT_185_port, 
      SHIFT_184_port, SHIFT_183_port, SHIFT_182_port, SHIFT_181_port, 
      SHIFT_180_port, SHIFT_179_port, SHIFT_178_port, SHIFT_177_port, 
      SHIFT_176_port, SHIFT_175_port, SHIFT_174_port, SHIFT_173_port, 
      SHIFT_172_port, SHIFT_171_port, SHIFT_170_port, SHIFT_169_port, 
      SHIFT_168_port, SHIFT_167_port, SHIFT_166_port, SHIFT_165_port, 
      SHIFT_164_port, SHIFT_163_port, SHIFT_162_port, SHIFT_161_port, 
      SHIFT_160_port, SHIFT_159_port, SHIFT_158_port, SHIFT_157_port, 
      SHIFT_156_port, SHIFT_155_port, SHIFT_154_port, SHIFT_153_port, 
      SHIFT_152_port, SHIFT_151_port, SHIFT_150_port, SHIFT_149_port, 
      SHIFT_148_port, SHIFT_147_port, SHIFT_146_port, SHIFT_145_port, 
      SHIFT_144_port, SHIFT_143_port, SHIFT_142_port, SHIFT_141_port, 
      SHIFT_140_port, SHIFT_139_port, SHIFT_138_port, SHIFT_137_port, 
      SHIFT_136_port, SHIFT_135_port, SHIFT_134_port, SHIFT_133_port, 
      SHIFT_132_port, SHIFT_131_port, SHIFT_130_port, SHIFT_129_port, 
      SHIFT_128_port, SHIFT_127_port, SHIFT_126_port, SHIFT_125_port, 
      SHIFT_124_port, SHIFT_123_port, SHIFT_122_port, SHIFT_121_port, 
      SHIFT_120_port, SHIFT_119_port, SHIFT_118_port, SHIFT_117_port, 
      SHIFT_116_port, SHIFT_115_port, SHIFT_114_port, SHIFT_113_port, 
      SHIFT_112_port, SHIFT_111_port, SHIFT_110_port, SHIFT_109_port, 
      SHIFT_108_port, SHIFT_107_port, SHIFT_106_port, SHIFT_105_port, 
      SHIFT_104_port, SHIFT_103_port, SHIFT_102_port, SHIFT_101_port, 
      SHIFT_100_port, SHIFT_99_port, SHIFT_98_port, SHIFT_97_port, 
      SHIFT_96_port, SHIFT_95_port, SHIFT_94_port, SHIFT_93_port, SHIFT_92_port
      , SHIFT_91_port, SHIFT_90_port, SHIFT_89_port, SHIFT_88_port, 
      SHIFT_87_port, SHIFT_86_port, SHIFT_85_port, SHIFT_84_port, SHIFT_83_port
      , SHIFT_82_port, SHIFT_81_port, SHIFT_80_port, SHIFT_79_port, 
      SHIFT_78_port, SHIFT_77_port, SHIFT_76_port, SHIFT_75_port, SHIFT_74_port
      , SHIFT_73_port, SHIFT_72_port, SHIFT_71_port, SHIFT_70_port, 
      SHIFT_69_port, SHIFT_68_port, SHIFT_67_port, SHIFT_66_port, SHIFT_65_port
      , SHIFT_64_port, SHIFT_n_1023_port, SHIFT_n_1022_port, SHIFT_n_1021_port,
      SHIFT_n_1020_port, SHIFT_n_1019_port, SHIFT_n_1018_port, 
      SHIFT_n_1017_port, SHIFT_n_1016_port, SHIFT_n_1015_port, 
      SHIFT_n_1014_port, SHIFT_n_1013_port, SHIFT_n_1012_port, 
      SHIFT_n_1011_port, SHIFT_n_1010_port, SHIFT_n_1009_port, 
      SHIFT_n_1008_port, SHIFT_n_1007_port, SHIFT_n_1006_port, 
      SHIFT_n_1005_port, SHIFT_n_1004_port, SHIFT_n_1003_port, 
      SHIFT_n_1002_port, SHIFT_n_1001_port, SHIFT_n_1000_port, SHIFT_n_999_port
      , SHIFT_n_998_port, SHIFT_n_997_port, SHIFT_n_996_port, SHIFT_n_995_port,
      SHIFT_n_994_port, SHIFT_n_993_port, SHIFT_n_992_port, SHIFT_n_991_port, 
      SHIFT_n_990_port, SHIFT_n_989_port, SHIFT_n_988_port, SHIFT_n_987_port, 
      SHIFT_n_986_port, SHIFT_n_985_port, SHIFT_n_984_port, SHIFT_n_983_port, 
      SHIFT_n_982_port, SHIFT_n_981_port, SHIFT_n_980_port, SHIFT_n_979_port, 
      SHIFT_n_978_port, SHIFT_n_977_port, SHIFT_n_976_port, SHIFT_n_975_port, 
      SHIFT_n_974_port, SHIFT_n_973_port, SHIFT_n_972_port, SHIFT_n_971_port, 
      SHIFT_n_970_port, SHIFT_n_969_port, SHIFT_n_968_port, SHIFT_n_967_port, 
      SHIFT_n_966_port, SHIFT_n_965_port, SHIFT_n_964_port, SHIFT_n_963_port, 
      SHIFT_n_962_port, SHIFT_n_961_port, SHIFT_n_960_port, SHIFT_n_959_port, 
      SHIFT_n_958_port, SHIFT_n_957_port, SHIFT_n_956_port, SHIFT_n_955_port, 
      SHIFT_n_954_port, SHIFT_n_953_port, SHIFT_n_952_port, SHIFT_n_951_port, 
      SHIFT_n_950_port, SHIFT_n_949_port, SHIFT_n_948_port, SHIFT_n_947_port, 
      SHIFT_n_946_port, SHIFT_n_945_port, SHIFT_n_944_port, SHIFT_n_943_port, 
      SHIFT_n_942_port, SHIFT_n_941_port, SHIFT_n_940_port, SHIFT_n_939_port, 
      SHIFT_n_938_port, SHIFT_n_937_port, SHIFT_n_936_port, SHIFT_n_935_port, 
      SHIFT_n_934_port, SHIFT_n_933_port, SHIFT_n_932_port, SHIFT_n_931_port, 
      SHIFT_n_930_port, SHIFT_n_929_port, SHIFT_n_928_port, SHIFT_n_927_port, 
      SHIFT_n_926_port, SHIFT_n_925_port, SHIFT_n_924_port, SHIFT_n_923_port, 
      SHIFT_n_922_port, SHIFT_n_921_port, SHIFT_n_920_port, SHIFT_n_919_port, 
      SHIFT_n_918_port, SHIFT_n_917_port, SHIFT_n_916_port, SHIFT_n_915_port, 
      SHIFT_n_914_port, SHIFT_n_913_port, SHIFT_n_912_port, SHIFT_n_911_port, 
      SHIFT_n_910_port, SHIFT_n_909_port, SHIFT_n_908_port, SHIFT_n_907_port, 
      SHIFT_n_906_port, SHIFT_n_905_port, SHIFT_n_904_port, SHIFT_n_903_port, 
      SHIFT_n_902_port, SHIFT_n_901_port, SHIFT_n_900_port, SHIFT_n_899_port, 
      SHIFT_n_898_port, SHIFT_n_897_port, SHIFT_n_896_port, SHIFT_n_895_port, 
      SHIFT_n_894_port, SHIFT_n_893_port, SHIFT_n_892_port, SHIFT_n_891_port, 
      SHIFT_n_890_port, SHIFT_n_889_port, SHIFT_n_888_port, SHIFT_n_887_port, 
      SHIFT_n_886_port, SHIFT_n_885_port, SHIFT_n_884_port, SHIFT_n_883_port, 
      SHIFT_n_882_port, SHIFT_n_881_port, SHIFT_n_880_port, SHIFT_n_879_port, 
      SHIFT_n_878_port, SHIFT_n_877_port, SHIFT_n_876_port, SHIFT_n_875_port, 
      SHIFT_n_874_port, SHIFT_n_873_port, SHIFT_n_872_port, SHIFT_n_871_port, 
      SHIFT_n_870_port, SHIFT_n_869_port, SHIFT_n_868_port, SHIFT_n_867_port, 
      SHIFT_n_866_port, SHIFT_n_865_port, SHIFT_n_864_port, SHIFT_n_863_port, 
      SHIFT_n_862_port, SHIFT_n_861_port, SHIFT_n_860_port, SHIFT_n_859_port, 
      SHIFT_n_858_port, SHIFT_n_857_port, SHIFT_n_856_port, SHIFT_n_855_port, 
      SHIFT_n_854_port, SHIFT_n_853_port, SHIFT_n_852_port, SHIFT_n_851_port, 
      SHIFT_n_850_port, SHIFT_n_849_port, SHIFT_n_848_port, SHIFT_n_847_port, 
      SHIFT_n_846_port, SHIFT_n_845_port, SHIFT_n_844_port, SHIFT_n_843_port, 
      SHIFT_n_842_port, SHIFT_n_841_port, SHIFT_n_840_port, SHIFT_n_839_port, 
      SHIFT_n_838_port, SHIFT_n_837_port, SHIFT_n_836_port, SHIFT_n_835_port, 
      SHIFT_n_834_port, SHIFT_n_833_port, SHIFT_n_832_port, SHIFT_n_831_port, 
      SHIFT_n_830_port, SHIFT_n_829_port, SHIFT_n_828_port, SHIFT_n_827_port, 
      SHIFT_n_826_port, SHIFT_n_825_port, SHIFT_n_824_port, SHIFT_n_823_port, 
      SHIFT_n_822_port, SHIFT_n_821_port, SHIFT_n_820_port, SHIFT_n_819_port, 
      SHIFT_n_818_port, SHIFT_n_817_port, SHIFT_n_816_port, SHIFT_n_815_port, 
      SHIFT_n_814_port, SHIFT_n_813_port, SHIFT_n_812_port, SHIFT_n_811_port, 
      SHIFT_n_810_port, SHIFT_n_809_port, SHIFT_n_808_port, SHIFT_n_807_port, 
      SHIFT_n_806_port, SHIFT_n_805_port, SHIFT_n_804_port, SHIFT_n_803_port, 
      SHIFT_n_802_port, SHIFT_n_801_port, SHIFT_n_800_port, SHIFT_n_799_port, 
      SHIFT_n_798_port, SHIFT_n_797_port, SHIFT_n_796_port, SHIFT_n_795_port, 
      SHIFT_n_794_port, SHIFT_n_793_port, SHIFT_n_792_port, SHIFT_n_791_port, 
      SHIFT_n_790_port, SHIFT_n_789_port, SHIFT_n_788_port, SHIFT_n_787_port, 
      SHIFT_n_786_port, SHIFT_n_785_port, SHIFT_n_784_port, SHIFT_n_783_port, 
      SHIFT_n_782_port, SHIFT_n_781_port, SHIFT_n_780_port, SHIFT_n_779_port, 
      SHIFT_n_778_port, SHIFT_n_777_port, SHIFT_n_776_port, SHIFT_n_775_port, 
      SHIFT_n_774_port, SHIFT_n_773_port, SHIFT_n_772_port, SHIFT_n_771_port, 
      SHIFT_n_770_port, SHIFT_n_769_port, SHIFT_n_768_port, SHIFT_n_767_port, 
      SHIFT_n_766_port, SHIFT_n_765_port, SHIFT_n_764_port, SHIFT_n_763_port, 
      SHIFT_n_762_port, SHIFT_n_761_port, SHIFT_n_760_port, SHIFT_n_759_port, 
      SHIFT_n_758_port, SHIFT_n_757_port, SHIFT_n_756_port, SHIFT_n_755_port, 
      SHIFT_n_754_port, SHIFT_n_753_port, SHIFT_n_752_port, SHIFT_n_751_port, 
      SHIFT_n_750_port, SHIFT_n_749_port, SHIFT_n_748_port, SHIFT_n_747_port, 
      SHIFT_n_746_port, SHIFT_n_745_port, SHIFT_n_744_port, SHIFT_n_743_port, 
      SHIFT_n_742_port, SHIFT_n_741_port, SHIFT_n_740_port, SHIFT_n_739_port, 
      SHIFT_n_738_port, SHIFT_n_737_port, SHIFT_n_736_port, SHIFT_n_735_port, 
      SHIFT_n_734_port, SHIFT_n_733_port, SHIFT_n_732_port, SHIFT_n_731_port, 
      SHIFT_n_730_port, SHIFT_n_729_port, SHIFT_n_728_port, SHIFT_n_727_port, 
      SHIFT_n_726_port, SHIFT_n_725_port, SHIFT_n_724_port, SHIFT_n_723_port, 
      SHIFT_n_722_port, SHIFT_n_721_port, SHIFT_n_720_port, SHIFT_n_719_port, 
      SHIFT_n_718_port, SHIFT_n_717_port, SHIFT_n_716_port, SHIFT_n_715_port, 
      SHIFT_n_714_port, SHIFT_n_713_port, SHIFT_n_712_port, SHIFT_n_711_port, 
      SHIFT_n_710_port, SHIFT_n_709_port, SHIFT_n_708_port, SHIFT_n_707_port, 
      SHIFT_n_706_port, SHIFT_n_705_port, SHIFT_n_704_port, SHIFT_n_703_port, 
      SHIFT_n_702_port, SHIFT_n_701_port, SHIFT_n_700_port, SHIFT_n_699_port, 
      SHIFT_n_698_port, SHIFT_n_697_port, SHIFT_n_696_port, SHIFT_n_695_port, 
      SHIFT_n_694_port, SHIFT_n_693_port, SHIFT_n_692_port, SHIFT_n_691_port, 
      SHIFT_n_690_port, SHIFT_n_689_port, SHIFT_n_688_port, SHIFT_n_687_port, 
      SHIFT_n_686_port, SHIFT_n_685_port, SHIFT_n_684_port, SHIFT_n_683_port, 
      SHIFT_n_682_port, SHIFT_n_681_port, SHIFT_n_680_port, SHIFT_n_679_port, 
      SHIFT_n_678_port, SHIFT_n_677_port, SHIFT_n_676_port, SHIFT_n_675_port, 
      SHIFT_n_674_port, SHIFT_n_673_port, SHIFT_n_672_port, SHIFT_n_671_port, 
      SHIFT_n_670_port, SHIFT_n_669_port, SHIFT_n_668_port, SHIFT_n_667_port, 
      SHIFT_n_666_port, SHIFT_n_665_port, SHIFT_n_664_port, SHIFT_n_663_port, 
      SHIFT_n_662_port, SHIFT_n_661_port, SHIFT_n_660_port, SHIFT_n_659_port, 
      SHIFT_n_658_port, SHIFT_n_657_port, SHIFT_n_656_port, SHIFT_n_655_port, 
      SHIFT_n_654_port, SHIFT_n_653_port, SHIFT_n_652_port, SHIFT_n_651_port, 
      SHIFT_n_650_port, SHIFT_n_649_port, SHIFT_n_648_port, SHIFT_n_647_port, 
      SHIFT_n_646_port, SHIFT_n_645_port, SHIFT_n_644_port, SHIFT_n_643_port, 
      SHIFT_n_642_port, SHIFT_n_641_port, SHIFT_n_640_port, SHIFT_n_639_port, 
      SHIFT_n_638_port, SHIFT_n_637_port, SHIFT_n_636_port, SHIFT_n_635_port, 
      SHIFT_n_634_port, SHIFT_n_633_port, SHIFT_n_632_port, SHIFT_n_631_port, 
      SHIFT_n_630_port, SHIFT_n_629_port, SHIFT_n_628_port, SHIFT_n_627_port, 
      SHIFT_n_626_port, SHIFT_n_625_port, SHIFT_n_624_port, SHIFT_n_623_port, 
      SHIFT_n_622_port, SHIFT_n_621_port, SHIFT_n_620_port, SHIFT_n_619_port, 
      SHIFT_n_618_port, SHIFT_n_617_port, SHIFT_n_616_port, SHIFT_n_615_port, 
      SHIFT_n_614_port, SHIFT_n_613_port, SHIFT_n_612_port, SHIFT_n_611_port, 
      SHIFT_n_610_port, SHIFT_n_609_port, SHIFT_n_608_port, SHIFT_n_607_port, 
      SHIFT_n_606_port, SHIFT_n_605_port, SHIFT_n_604_port, SHIFT_n_603_port, 
      SHIFT_n_602_port, SHIFT_n_601_port, SHIFT_n_600_port, SHIFT_n_599_port, 
      SHIFT_n_598_port, SHIFT_n_597_port, SHIFT_n_596_port, SHIFT_n_595_port, 
      SHIFT_n_594_port, SHIFT_n_593_port, SHIFT_n_592_port, SHIFT_n_591_port, 
      SHIFT_n_590_port, SHIFT_n_589_port, SHIFT_n_588_port, SHIFT_n_587_port, 
      SHIFT_n_586_port, SHIFT_n_585_port, SHIFT_n_584_port, SHIFT_n_583_port, 
      SHIFT_n_582_port, SHIFT_n_581_port, SHIFT_n_580_port, SHIFT_n_579_port, 
      SHIFT_n_578_port, SHIFT_n_577_port, SHIFT_n_576_port, SHIFT_n_575_port, 
      SHIFT_n_574_port, SHIFT_n_573_port, SHIFT_n_572_port, SHIFT_n_571_port, 
      SHIFT_n_570_port, SHIFT_n_569_port, SHIFT_n_568_port, SHIFT_n_567_port, 
      SHIFT_n_566_port, SHIFT_n_565_port, SHIFT_n_564_port, SHIFT_n_563_port, 
      SHIFT_n_562_port, SHIFT_n_561_port, SHIFT_n_560_port, SHIFT_n_559_port, 
      SHIFT_n_558_port, SHIFT_n_557_port, SHIFT_n_556_port, SHIFT_n_555_port, 
      SHIFT_n_554_port, SHIFT_n_553_port, SHIFT_n_552_port, SHIFT_n_551_port, 
      SHIFT_n_550_port, SHIFT_n_549_port, SHIFT_n_548_port, SHIFT_n_547_port, 
      SHIFT_n_546_port, SHIFT_n_545_port, SHIFT_n_544_port, SHIFT_n_543_port, 
      SHIFT_n_542_port, SHIFT_n_541_port, SHIFT_n_540_port, SHIFT_n_539_port, 
      SHIFT_n_538_port, SHIFT_n_537_port, SHIFT_n_536_port, SHIFT_n_535_port, 
      SHIFT_n_534_port, SHIFT_n_533_port, SHIFT_n_532_port, SHIFT_n_531_port, 
      SHIFT_n_530_port, SHIFT_n_529_port, SHIFT_n_528_port, SHIFT_n_527_port, 
      SHIFT_n_526_port, SHIFT_n_525_port, SHIFT_n_524_port, SHIFT_n_523_port, 
      SHIFT_n_522_port, SHIFT_n_521_port, SHIFT_n_520_port, SHIFT_n_519_port, 
      SHIFT_n_518_port, SHIFT_n_517_port, SHIFT_n_516_port, SHIFT_n_515_port, 
      SHIFT_n_514_port, SHIFT_n_513_port, SHIFT_n_512_port, SHIFT_n_511_port, 
      SHIFT_n_510_port, SHIFT_n_509_port, SHIFT_n_508_port, SHIFT_n_507_port, 
      SHIFT_n_506_port, SHIFT_n_505_port, SHIFT_n_504_port, SHIFT_n_503_port, 
      SHIFT_n_502_port, SHIFT_n_501_port, SHIFT_n_500_port, SHIFT_n_499_port, 
      SHIFT_n_498_port, SHIFT_n_497_port, SHIFT_n_496_port, SHIFT_n_495_port, 
      SHIFT_n_494_port, SHIFT_n_493_port, SHIFT_n_492_port, SHIFT_n_491_port, 
      SHIFT_n_490_port, SHIFT_n_489_port, SHIFT_n_488_port, SHIFT_n_487_port, 
      SHIFT_n_486_port, SHIFT_n_485_port, SHIFT_n_484_port, SHIFT_n_483_port, 
      SHIFT_n_482_port, SHIFT_n_481_port, SHIFT_n_480_port, SHIFT_n_479_port, 
      SHIFT_n_478_port, SHIFT_n_477_port, SHIFT_n_476_port, SHIFT_n_475_port, 
      SHIFT_n_474_port, SHIFT_n_473_port, SHIFT_n_472_port, SHIFT_n_471_port, 
      SHIFT_n_470_port, SHIFT_n_469_port, SHIFT_n_468_port, SHIFT_n_467_port, 
      SHIFT_n_466_port, SHIFT_n_465_port, SHIFT_n_464_port, SHIFT_n_463_port, 
      SHIFT_n_462_port, SHIFT_n_461_port, SHIFT_n_460_port, SHIFT_n_459_port, 
      SHIFT_n_458_port, SHIFT_n_457_port, SHIFT_n_456_port, SHIFT_n_455_port, 
      SHIFT_n_454_port, SHIFT_n_453_port, SHIFT_n_452_port, SHIFT_n_451_port, 
      SHIFT_n_450_port, SHIFT_n_449_port, SHIFT_n_448_port, SHIFT_n_447_port, 
      SHIFT_n_446_port, SHIFT_n_445_port, SHIFT_n_444_port, SHIFT_n_443_port, 
      SHIFT_n_442_port, SHIFT_n_441_port, SHIFT_n_440_port, SHIFT_n_439_port, 
      SHIFT_n_438_port, SHIFT_n_437_port, SHIFT_n_436_port, SHIFT_n_435_port, 
      SHIFT_n_434_port, SHIFT_n_433_port, SHIFT_n_432_port, SHIFT_n_431_port, 
      SHIFT_n_430_port, SHIFT_n_429_port, SHIFT_n_428_port, SHIFT_n_427_port, 
      SHIFT_n_426_port, SHIFT_n_425_port, SHIFT_n_424_port, SHIFT_n_423_port, 
      SHIFT_n_422_port, SHIFT_n_421_port, SHIFT_n_420_port, SHIFT_n_419_port, 
      SHIFT_n_418_port, SHIFT_n_417_port, SHIFT_n_416_port, SHIFT_n_415_port, 
      SHIFT_n_414_port, SHIFT_n_413_port, SHIFT_n_412_port, SHIFT_n_411_port, 
      SHIFT_n_410_port, SHIFT_n_409_port, SHIFT_n_408_port, SHIFT_n_407_port, 
      SHIFT_n_406_port, SHIFT_n_405_port, SHIFT_n_404_port, SHIFT_n_403_port, 
      SHIFT_n_402_port, SHIFT_n_401_port, SHIFT_n_400_port, SHIFT_n_399_port, 
      SHIFT_n_398_port, SHIFT_n_397_port, SHIFT_n_396_port, SHIFT_n_395_port, 
      SHIFT_n_394_port, SHIFT_n_393_port, SHIFT_n_392_port, SHIFT_n_391_port, 
      SHIFT_n_390_port, SHIFT_n_389_port, SHIFT_n_388_port, SHIFT_n_387_port, 
      SHIFT_n_386_port, SHIFT_n_385_port, SHIFT_n_384_port, SHIFT_n_383_port, 
      SHIFT_n_382_port, SHIFT_n_381_port, SHIFT_n_380_port, SHIFT_n_379_port, 
      SHIFT_n_378_port, SHIFT_n_377_port, SHIFT_n_376_port, SHIFT_n_375_port, 
      SHIFT_n_374_port, SHIFT_n_373_port, SHIFT_n_372_port, SHIFT_n_371_port, 
      SHIFT_n_370_port, SHIFT_n_369_port, SHIFT_n_368_port, SHIFT_n_367_port, 
      SHIFT_n_366_port, SHIFT_n_365_port, SHIFT_n_364_port, SHIFT_n_363_port, 
      SHIFT_n_362_port, SHIFT_n_361_port, SHIFT_n_360_port, SHIFT_n_359_port, 
      SHIFT_n_358_port, SHIFT_n_357_port, SHIFT_n_356_port, SHIFT_n_355_port, 
      SHIFT_n_354_port, SHIFT_n_353_port, SHIFT_n_352_port, SHIFT_n_351_port, 
      SHIFT_n_350_port, SHIFT_n_349_port, SHIFT_n_348_port, SHIFT_n_347_port, 
      SHIFT_n_346_port, SHIFT_n_345_port, SHIFT_n_344_port, SHIFT_n_343_port, 
      SHIFT_n_342_port, SHIFT_n_341_port, SHIFT_n_340_port, SHIFT_n_339_port, 
      SHIFT_n_338_port, SHIFT_n_337_port, SHIFT_n_336_port, SHIFT_n_335_port, 
      SHIFT_n_334_port, SHIFT_n_333_port, SHIFT_n_332_port, SHIFT_n_331_port, 
      SHIFT_n_330_port, SHIFT_n_329_port, SHIFT_n_328_port, SHIFT_n_327_port, 
      SHIFT_n_326_port, SHIFT_n_325_port, SHIFT_n_324_port, SHIFT_n_323_port, 
      SHIFT_n_322_port, SHIFT_n_321_port, SHIFT_n_320_port, SHIFT_n_319_port, 
      SHIFT_n_318_port, SHIFT_n_317_port, SHIFT_n_316_port, SHIFT_n_315_port, 
      SHIFT_n_314_port, SHIFT_n_313_port, SHIFT_n_312_port, SHIFT_n_311_port, 
      SHIFT_n_310_port, SHIFT_n_309_port, SHIFT_n_308_port, SHIFT_n_307_port, 
      SHIFT_n_306_port, SHIFT_n_305_port, SHIFT_n_304_port, SHIFT_n_303_port, 
      SHIFT_n_302_port, SHIFT_n_301_port, SHIFT_n_300_port, SHIFT_n_299_port, 
      SHIFT_n_298_port, SHIFT_n_297_port, SHIFT_n_296_port, SHIFT_n_295_port, 
      SHIFT_n_294_port, SHIFT_n_293_port, SHIFT_n_292_port, SHIFT_n_291_port, 
      SHIFT_n_290_port, SHIFT_n_289_port, SHIFT_n_288_port, SHIFT_n_287_port, 
      SHIFT_n_286_port, SHIFT_n_285_port, SHIFT_n_284_port, SHIFT_n_283_port, 
      SHIFT_n_282_port, SHIFT_n_281_port, SHIFT_n_280_port, SHIFT_n_279_port, 
      SHIFT_n_278_port, SHIFT_n_277_port, SHIFT_n_276_port, SHIFT_n_275_port, 
      SHIFT_n_274_port, SHIFT_n_273_port, SHIFT_n_272_port, SHIFT_n_271_port, 
      SHIFT_n_270_port, SHIFT_n_269_port, SHIFT_n_268_port, SHIFT_n_267_port, 
      SHIFT_n_266_port, SHIFT_n_265_port, SHIFT_n_264_port, SHIFT_n_263_port, 
      SHIFT_n_262_port, SHIFT_n_261_port, SHIFT_n_260_port, SHIFT_n_259_port, 
      SHIFT_n_258_port, SHIFT_n_257_port, SHIFT_n_256_port, SHIFT_n_255_port, 
      SHIFT_n_254_port, SHIFT_n_253_port, SHIFT_n_252_port, SHIFT_n_251_port, 
      SHIFT_n_250_port, SHIFT_n_249_port, SHIFT_n_248_port, SHIFT_n_247_port, 
      SHIFT_n_246_port, SHIFT_n_245_port, SHIFT_n_244_port, SHIFT_n_243_port, 
      SHIFT_n_242_port, SHIFT_n_241_port, SHIFT_n_240_port, SHIFT_n_239_port, 
      SHIFT_n_238_port, SHIFT_n_237_port, SHIFT_n_236_port, SHIFT_n_235_port, 
      SHIFT_n_234_port, SHIFT_n_233_port, SHIFT_n_232_port, SHIFT_n_231_port, 
      SHIFT_n_230_port, SHIFT_n_229_port, SHIFT_n_228_port, SHIFT_n_227_port, 
      SHIFT_n_226_port, SHIFT_n_225_port, SHIFT_n_224_port, SHIFT_n_223_port, 
      SHIFT_n_222_port, SHIFT_n_221_port, SHIFT_n_220_port, SHIFT_n_219_port, 
      SHIFT_n_218_port, SHIFT_n_217_port, SHIFT_n_216_port, SHIFT_n_215_port, 
      SHIFT_n_214_port, SHIFT_n_213_port, SHIFT_n_212_port, SHIFT_n_211_port, 
      SHIFT_n_210_port, SHIFT_n_209_port, SHIFT_n_208_port, SHIFT_n_207_port, 
      SHIFT_n_206_port, SHIFT_n_205_port, SHIFT_n_204_port, SHIFT_n_203_port, 
      SHIFT_n_202_port, SHIFT_n_201_port, SHIFT_n_200_port, SHIFT_n_199_port, 
      SHIFT_n_198_port, SHIFT_n_197_port, SHIFT_n_196_port, SHIFT_n_195_port, 
      SHIFT_n_194_port, SHIFT_n_193_port, SHIFT_n_192_port, SHIFT_n_191_port, 
      SHIFT_n_190_port, SHIFT_n_189_port, SHIFT_n_188_port, SHIFT_n_187_port, 
      SHIFT_n_186_port, SHIFT_n_185_port, SHIFT_n_184_port, SHIFT_n_183_port, 
      SHIFT_n_182_port, SHIFT_n_181_port, SHIFT_n_180_port, SHIFT_n_179_port, 
      SHIFT_n_178_port, SHIFT_n_177_port, SHIFT_n_176_port, SHIFT_n_175_port, 
      SHIFT_n_174_port, SHIFT_n_173_port, SHIFT_n_172_port, SHIFT_n_171_port, 
      SHIFT_n_170_port, SHIFT_n_169_port, SHIFT_n_168_port, SHIFT_n_167_port, 
      SHIFT_n_166_port, SHIFT_n_165_port, SHIFT_n_164_port, SHIFT_n_163_port, 
      SHIFT_n_162_port, SHIFT_n_161_port, SHIFT_n_160_port, SHIFT_n_159_port, 
      SHIFT_n_158_port, SHIFT_n_157_port, SHIFT_n_156_port, SHIFT_n_155_port, 
      SHIFT_n_154_port, SHIFT_n_153_port, SHIFT_n_152_port, SHIFT_n_151_port, 
      SHIFT_n_150_port, SHIFT_n_149_port, SHIFT_n_148_port, SHIFT_n_147_port, 
      SHIFT_n_146_port, SHIFT_n_145_port, SHIFT_n_144_port, SHIFT_n_143_port, 
      SHIFT_n_142_port, SHIFT_n_141_port, SHIFT_n_140_port, SHIFT_n_139_port, 
      SHIFT_n_138_port, SHIFT_n_137_port, SHIFT_n_136_port, SHIFT_n_135_port, 
      SHIFT_n_134_port, SHIFT_n_133_port, SHIFT_n_132_port, SHIFT_n_131_port, 
      SHIFT_n_130_port, SHIFT_n_129_port, SHIFT_n_128_port, SHIFT_n_127_port, 
      SHIFT_n_126_port, SHIFT_n_125_port, SHIFT_n_124_port, SHIFT_n_123_port, 
      SHIFT_n_122_port, SHIFT_n_121_port, SHIFT_n_120_port, SHIFT_n_119_port, 
      SHIFT_n_118_port, SHIFT_n_117_port, SHIFT_n_116_port, SHIFT_n_115_port, 
      SHIFT_n_114_port, SHIFT_n_113_port, SHIFT_n_112_port, SHIFT_n_111_port, 
      SHIFT_n_110_port, SHIFT_n_109_port, SHIFT_n_108_port, SHIFT_n_107_port, 
      SHIFT_n_106_port, SHIFT_n_105_port, SHIFT_n_104_port, SHIFT_n_103_port, 
      SHIFT_n_102_port, SHIFT_n_101_port, SHIFT_n_100_port, SHIFT_n_99_port, 
      SHIFT_n_98_port, SHIFT_n_97_port, SHIFT_n_96_port, SHIFT_n_95_port, 
      SHIFT_n_94_port, SHIFT_n_93_port, SHIFT_n_92_port, SHIFT_n_91_port, 
      SHIFT_n_90_port, SHIFT_n_89_port, SHIFT_n_88_port, SHIFT_n_87_port, 
      SHIFT_n_86_port, SHIFT_n_85_port, SHIFT_n_84_port, SHIFT_n_83_port, 
      SHIFT_n_82_port, SHIFT_n_81_port, SHIFT_n_80_port, SHIFT_n_79_port, 
      SHIFT_n_78_port, SHIFT_n_77_port, SHIFT_n_76_port, SHIFT_n_75_port, 
      SHIFT_n_74_port, SHIFT_n_73_port, SHIFT_n_72_port, SHIFT_n_71_port, 
      SHIFT_n_70_port, SHIFT_n_69_port, SHIFT_n_68_port, SHIFT_n_67_port, 
      SHIFT_n_66_port, SHIFT_n_65_port, SHIFT_n_64_port, OTMP_511_port, 
      OTMP_510_port, OTMP_509_port, OTMP_508_port, OTMP_507_port, OTMP_506_port
      , OTMP_505_port, OTMP_504_port, OTMP_503_port, OTMP_502_port, 
      OTMP_501_port, OTMP_500_port, OTMP_499_port, OTMP_498_port, OTMP_497_port
      , OTMP_496_port, OTMP_495_port, OTMP_494_port, OTMP_493_port, 
      OTMP_492_port, OTMP_491_port, OTMP_490_port, OTMP_489_port, OTMP_488_port
      , OTMP_487_port, OTMP_486_port, OTMP_485_port, OTMP_484_port, 
      OTMP_483_port, OTMP_482_port, OTMP_481_port, OTMP_480_port, OTMP_479_port
      , OTMP_478_port, OTMP_477_port, OTMP_476_port, OTMP_475_port, 
      OTMP_474_port, OTMP_473_port, OTMP_472_port, OTMP_471_port, OTMP_470_port
      , OTMP_469_port, OTMP_468_port, OTMP_467_port, OTMP_466_port, 
      OTMP_465_port, OTMP_464_port, OTMP_463_port, OTMP_462_port, OTMP_461_port
      , OTMP_460_port, OTMP_459_port, OTMP_458_port, OTMP_457_port, 
      OTMP_456_port, OTMP_455_port, OTMP_454_port, OTMP_453_port, OTMP_452_port
      , OTMP_451_port, OTMP_450_port, OTMP_449_port, OTMP_448_port, 
      OTMP_447_port, OTMP_446_port, OTMP_445_port, OTMP_444_port, OTMP_443_port
      , OTMP_442_port, OTMP_441_port, OTMP_440_port, OTMP_439_port, 
      OTMP_438_port, OTMP_437_port, OTMP_436_port, OTMP_435_port, OTMP_434_port
      , OTMP_433_port, OTMP_432_port, OTMP_431_port, OTMP_430_port, 
      OTMP_429_port, OTMP_428_port, OTMP_427_port, OTMP_426_port, OTMP_425_port
      , OTMP_424_port, OTMP_423_port, OTMP_422_port, OTMP_421_port, 
      OTMP_420_port, OTMP_419_port, OTMP_418_port, OTMP_417_port, OTMP_416_port
      , OTMP_415_port, OTMP_414_port, OTMP_413_port, OTMP_412_port, 
      OTMP_411_port, OTMP_410_port, OTMP_409_port, OTMP_408_port, OTMP_407_port
      , OTMP_406_port, OTMP_405_port, OTMP_404_port, OTMP_403_port, 
      OTMP_402_port, OTMP_401_port, OTMP_400_port, OTMP_399_port, OTMP_398_port
      , OTMP_397_port, OTMP_396_port, OTMP_395_port, OTMP_394_port, 
      OTMP_393_port, OTMP_392_port, OTMP_391_port, OTMP_390_port, OTMP_389_port
      , OTMP_388_port, OTMP_387_port, OTMP_386_port, OTMP_385_port, 
      OTMP_384_port, OTMP_383_port, OTMP_382_port, OTMP_381_port, OTMP_380_port
      , OTMP_379_port, OTMP_378_port, OTMP_377_port, OTMP_376_port, 
      OTMP_375_port, OTMP_374_port, OTMP_373_port, OTMP_372_port, OTMP_371_port
      , OTMP_370_port, OTMP_369_port, OTMP_368_port, OTMP_367_port, 
      OTMP_366_port, OTMP_365_port, OTMP_364_port, OTMP_363_port, OTMP_362_port
      , OTMP_361_port, OTMP_360_port, OTMP_359_port, OTMP_358_port, 
      OTMP_357_port, OTMP_356_port, OTMP_355_port, OTMP_354_port, OTMP_353_port
      , OTMP_352_port, OTMP_351_port, OTMP_350_port, OTMP_349_port, 
      OTMP_348_port, OTMP_347_port, OTMP_346_port, OTMP_345_port, OTMP_344_port
      , OTMP_343_port, OTMP_342_port, OTMP_341_port, OTMP_340_port, 
      OTMP_339_port, OTMP_338_port, OTMP_337_port, OTMP_336_port, OTMP_335_port
      , OTMP_334_port, OTMP_333_port, OTMP_332_port, OTMP_331_port, 
      OTMP_330_port, OTMP_329_port, OTMP_328_port, OTMP_327_port, OTMP_326_port
      , OTMP_325_port, OTMP_324_port, OTMP_323_port, OTMP_322_port, 
      OTMP_321_port, OTMP_320_port, OTMP_319_port, OTMP_318_port, OTMP_317_port
      , OTMP_316_port, OTMP_315_port, OTMP_314_port, OTMP_313_port, 
      OTMP_312_port, OTMP_311_port, OTMP_310_port, OTMP_309_port, OTMP_308_port
      , OTMP_307_port, OTMP_306_port, OTMP_305_port, OTMP_304_port, 
      OTMP_303_port, OTMP_302_port, OTMP_301_port, OTMP_300_port, OTMP_299_port
      , OTMP_298_port, OTMP_297_port, OTMP_296_port, OTMP_295_port, 
      OTMP_294_port, OTMP_293_port, OTMP_292_port, OTMP_291_port, OTMP_290_port
      , OTMP_289_port, OTMP_288_port, OTMP_287_port, OTMP_286_port, 
      OTMP_285_port, OTMP_284_port, OTMP_283_port, OTMP_282_port, OTMP_281_port
      , OTMP_280_port, OTMP_279_port, OTMP_278_port, OTMP_277_port, 
      OTMP_276_port, OTMP_275_port, OTMP_274_port, OTMP_273_port, OTMP_272_port
      , OTMP_271_port, OTMP_270_port, OTMP_269_port, OTMP_268_port, 
      OTMP_267_port, OTMP_266_port, OTMP_265_port, OTMP_264_port, OTMP_263_port
      , OTMP_262_port, OTMP_261_port, OTMP_260_port, OTMP_259_port, 
      OTMP_258_port, OTMP_257_port, OTMP_256_port, OTMP_255_port, OTMP_254_port
      , OTMP_253_port, OTMP_252_port, OTMP_251_port, OTMP_250_port, 
      OTMP_249_port, OTMP_248_port, OTMP_247_port, OTMP_246_port, OTMP_245_port
      , OTMP_244_port, OTMP_243_port, OTMP_242_port, OTMP_241_port, 
      OTMP_240_port, OTMP_239_port, OTMP_238_port, OTMP_237_port, OTMP_236_port
      , OTMP_235_port, OTMP_234_port, OTMP_233_port, OTMP_232_port, 
      OTMP_231_port, OTMP_230_port, OTMP_229_port, OTMP_228_port, OTMP_227_port
      , OTMP_226_port, OTMP_225_port, OTMP_224_port, OTMP_223_port, 
      OTMP_222_port, OTMP_221_port, OTMP_220_port, OTMP_219_port, OTMP_218_port
      , OTMP_217_port, OTMP_216_port, OTMP_215_port, OTMP_214_port, 
      OTMP_213_port, OTMP_212_port, OTMP_211_port, OTMP_210_port, OTMP_209_port
      , OTMP_208_port, OTMP_207_port, OTMP_206_port, OTMP_205_port, 
      OTMP_204_port, OTMP_203_port, OTMP_202_port, OTMP_201_port, OTMP_200_port
      , OTMP_199_port, OTMP_198_port, OTMP_197_port, OTMP_196_port, 
      OTMP_195_port, OTMP_194_port, OTMP_193_port, OTMP_192_port, OTMP_191_port
      , OTMP_190_port, OTMP_189_port, OTMP_188_port, OTMP_187_port, 
      OTMP_186_port, OTMP_185_port, OTMP_184_port, OTMP_183_port, OTMP_182_port
      , OTMP_181_port, OTMP_180_port, OTMP_179_port, OTMP_178_port, 
      OTMP_177_port, OTMP_176_port, OTMP_175_port, OTMP_174_port, OTMP_173_port
      , OTMP_172_port, OTMP_171_port, OTMP_170_port, OTMP_169_port, 
      OTMP_168_port, OTMP_167_port, OTMP_166_port, OTMP_165_port, OTMP_164_port
      , OTMP_163_port, OTMP_162_port, OTMP_161_port, OTMP_160_port, 
      OTMP_159_port, OTMP_158_port, OTMP_157_port, OTMP_156_port, OTMP_155_port
      , OTMP_154_port, OTMP_153_port, OTMP_152_port, OTMP_151_port, 
      OTMP_150_port, OTMP_149_port, OTMP_148_port, OTMP_147_port, OTMP_146_port
      , OTMP_145_port, OTMP_144_port, OTMP_143_port, OTMP_142_port, 
      OTMP_141_port, OTMP_140_port, OTMP_139_port, OTMP_138_port, OTMP_137_port
      , OTMP_136_port, OTMP_135_port, OTMP_134_port, OTMP_133_port, 
      OTMP_132_port, OTMP_131_port, OTMP_130_port, OTMP_129_port, OTMP_128_port
      , OTMP_127_port, OTMP_126_port, OTMP_125_port, OTMP_124_port, 
      OTMP_123_port, OTMP_122_port, OTMP_121_port, OTMP_120_port, OTMP_119_port
      , OTMP_118_port, OTMP_117_port, OTMP_116_port, OTMP_115_port, 
      OTMP_114_port, OTMP_113_port, OTMP_112_port, OTMP_111_port, OTMP_110_port
      , OTMP_109_port, OTMP_108_port, OTMP_107_port, OTMP_106_port, 
      OTMP_105_port, OTMP_104_port, OTMP_103_port, OTMP_102_port, OTMP_101_port
      , OTMP_100_port, OTMP_99_port, OTMP_98_port, OTMP_97_port, OTMP_96_port, 
      OTMP_95_port, OTMP_94_port, OTMP_93_port, OTMP_92_port, OTMP_91_port, 
      OTMP_90_port, OTMP_89_port, OTMP_88_port, OTMP_87_port, OTMP_86_port, 
      OTMP_85_port, OTMP_84_port, OTMP_83_port, OTMP_82_port, OTMP_81_port, 
      OTMP_80_port, OTMP_79_port, OTMP_78_port, OTMP_77_port, OTMP_76_port, 
      OTMP_75_port, OTMP_74_port, OTMP_73_port, OTMP_72_port, OTMP_71_port, 
      OTMP_70_port, OTMP_69_port, OTMP_68_port, OTMP_67_port, OTMP_66_port, 
      OTMP_65_port, OTMP_64_port, OTMP_63_port, OTMP_62_port, OTMP_61_port, 
      OTMP_60_port, OTMP_59_port, OTMP_58_port, OTMP_57_port, OTMP_56_port, 
      OTMP_55_port, OTMP_54_port, OTMP_53_port, OTMP_52_port, OTMP_51_port, 
      OTMP_50_port, OTMP_49_port, OTMP_48_port, OTMP_47_port, OTMP_46_port, 
      OTMP_45_port, OTMP_44_port, OTMP_43_port, OTMP_42_port, OTMP_41_port, 
      OTMP_40_port, OTMP_39_port, OTMP_38_port, OTMP_37_port, OTMP_36_port, 
      OTMP_35_port, OTMP_34_port, OTMP_33_port, OTMP_32_port, OTMP_31_port, 
      OTMP_30_port, OTMP_29_port, OTMP_28_port, OTMP_27_port, OTMP_26_port, 
      OTMP_25_port, OTMP_24_port, OTMP_23_port, OTMP_22_port, OTMP_21_port, 
      OTMP_20_port, OTMP_19_port, OTMP_18_port, OTMP_17_port, OTMP_16_port, 
      OTMP_15_port, OTMP_14_port, OTMP_13_port, OTMP_12_port, OTMP_11_port, 
      OTMP_10_port, OTMP_9_port, OTMP_8_port, OTMP_7_port, OTMP_6_port, 
      OTMP_5_port, OTMP_4_port, OTMP_3_port, OTMP_2_port, OTMP_1_port, 
      OTMP_0_port, OTMP_1023_port, OTMP_1022_port, OTMP_1021_port, 
      OTMP_1020_port, OTMP_1019_port, OTMP_1018_port, OTMP_1017_port, 
      OTMP_1016_port, OTMP_1015_port, OTMP_1014_port, OTMP_1013_port, 
      OTMP_1012_port, OTMP_1011_port, OTMP_1010_port, OTMP_1009_port, 
      OTMP_1008_port, OTMP_1007_port, OTMP_1006_port, OTMP_1005_port, 
      OTMP_1004_port, OTMP_1003_port, OTMP_1002_port, OTMP_1001_port, 
      OTMP_1000_port, OTMP_999_port, OTMP_998_port, OTMP_997_port, 
      OTMP_996_port, OTMP_995_port, OTMP_994_port, OTMP_993_port, OTMP_992_port
      , OTMP_991_port, OTMP_990_port, OTMP_989_port, OTMP_988_port, 
      OTMP_987_port, OTMP_986_port, OTMP_985_port, OTMP_984_port, OTMP_983_port
      , OTMP_982_port, OTMP_981_port, OTMP_980_port, OTMP_979_port, 
      OTMP_978_port, OTMP_977_port, OTMP_976_port, OTMP_975_port, OTMP_974_port
      , OTMP_973_port, OTMP_972_port, OTMP_971_port, OTMP_970_port, 
      OTMP_969_port, OTMP_968_port, OTMP_967_port, OTMP_966_port, OTMP_965_port
      , OTMP_964_port, OTMP_963_port, OTMP_962_port, OTMP_961_port, 
      OTMP_960_port, OTMP_959_port, OTMP_958_port, OTMP_957_port, OTMP_956_port
      , OTMP_955_port, OTMP_954_port, OTMP_953_port, OTMP_952_port, 
      OTMP_951_port, OTMP_950_port, OTMP_949_port, OTMP_948_port, OTMP_947_port
      , OTMP_946_port, OTMP_945_port, OTMP_944_port, OTMP_943_port, 
      OTMP_942_port, OTMP_941_port, OTMP_940_port, OTMP_939_port, OTMP_938_port
      , OTMP_937_port, OTMP_936_port, OTMP_935_port, OTMP_934_port, 
      OTMP_933_port, OTMP_932_port, OTMP_931_port, OTMP_930_port, OTMP_929_port
      , OTMP_928_port, OTMP_927_port, OTMP_926_port, OTMP_925_port, 
      OTMP_924_port, OTMP_923_port, OTMP_922_port, OTMP_921_port, OTMP_920_port
      , OTMP_919_port, OTMP_918_port, OTMP_917_port, OTMP_916_port, 
      OTMP_915_port, OTMP_914_port, OTMP_913_port, OTMP_912_port, OTMP_911_port
      , OTMP_910_port, OTMP_909_port, OTMP_908_port, OTMP_907_port, 
      OTMP_906_port, OTMP_905_port, OTMP_904_port, OTMP_903_port, OTMP_902_port
      , OTMP_901_port, OTMP_900_port, OTMP_899_port, OTMP_898_port, 
      OTMP_897_port, OTMP_896_port, OTMP_895_port, OTMP_894_port, OTMP_893_port
      , OTMP_892_port, OTMP_891_port, OTMP_890_port, OTMP_889_port, 
      OTMP_888_port, OTMP_887_port, OTMP_886_port, OTMP_885_port, OTMP_884_port
      , OTMP_883_port, OTMP_882_port, OTMP_881_port, OTMP_880_port, 
      OTMP_879_port, OTMP_878_port, OTMP_877_port, OTMP_876_port, OTMP_875_port
      , OTMP_874_port, OTMP_873_port, OTMP_872_port, OTMP_871_port, 
      OTMP_870_port, OTMP_869_port, OTMP_868_port, OTMP_867_port, OTMP_866_port
      , OTMP_865_port, OTMP_864_port, OTMP_863_port, OTMP_862_port, 
      OTMP_861_port, OTMP_860_port, OTMP_859_port, OTMP_858_port, OTMP_857_port
      , OTMP_856_port, OTMP_855_port, OTMP_854_port, OTMP_853_port, 
      OTMP_852_port, OTMP_851_port, OTMP_850_port, OTMP_849_port, OTMP_848_port
      , OTMP_847_port, OTMP_846_port, OTMP_845_port, OTMP_844_port, 
      OTMP_843_port, OTMP_842_port, OTMP_841_port, OTMP_840_port, OTMP_839_port
      , OTMP_838_port, OTMP_837_port, OTMP_836_port, OTMP_835_port, 
      OTMP_834_port, OTMP_833_port, OTMP_832_port, OTMP_831_port, OTMP_830_port
      , OTMP_829_port, OTMP_828_port, OTMP_827_port, OTMP_826_port, 
      OTMP_825_port, OTMP_824_port, OTMP_823_port, OTMP_822_port, OTMP_821_port
      , OTMP_820_port, OTMP_819_port, OTMP_818_port, OTMP_817_port, 
      OTMP_816_port, OTMP_815_port, OTMP_814_port, OTMP_813_port, OTMP_812_port
      , OTMP_811_port, OTMP_810_port, OTMP_809_port, OTMP_808_port, 
      OTMP_807_port, OTMP_806_port, OTMP_805_port, OTMP_804_port, OTMP_803_port
      , OTMP_802_port, OTMP_801_port, OTMP_800_port, OTMP_799_port, 
      OTMP_798_port, OTMP_797_port, OTMP_796_port, OTMP_795_port, OTMP_794_port
      , OTMP_793_port, OTMP_792_port, OTMP_791_port, OTMP_790_port, 
      OTMP_789_port, OTMP_788_port, OTMP_787_port, OTMP_786_port, OTMP_785_port
      , OTMP_784_port, OTMP_783_port, OTMP_782_port, OTMP_781_port, 
      OTMP_780_port, OTMP_779_port, OTMP_778_port, OTMP_777_port, OTMP_776_port
      , OTMP_775_port, OTMP_774_port, OTMP_773_port, OTMP_772_port, 
      OTMP_771_port, OTMP_770_port, OTMP_769_port, OTMP_768_port, OTMP_767_port
      , OTMP_766_port, OTMP_765_port, OTMP_764_port, OTMP_763_port, 
      OTMP_762_port, OTMP_761_port, OTMP_760_port, OTMP_759_port, OTMP_758_port
      , OTMP_757_port, OTMP_756_port, OTMP_755_port, OTMP_754_port, 
      OTMP_753_port, OTMP_752_port, OTMP_751_port, OTMP_750_port, OTMP_749_port
      , OTMP_748_port, OTMP_747_port, OTMP_746_port, OTMP_745_port, 
      OTMP_744_port, OTMP_743_port, OTMP_742_port, OTMP_741_port, OTMP_740_port
      , OTMP_739_port, OTMP_738_port, OTMP_737_port, OTMP_736_port, 
      OTMP_735_port, OTMP_734_port, OTMP_733_port, OTMP_732_port, OTMP_731_port
      , OTMP_730_port, OTMP_729_port, OTMP_728_port, OTMP_727_port, 
      OTMP_726_port, OTMP_725_port, OTMP_724_port, OTMP_723_port, OTMP_722_port
      , OTMP_721_port, OTMP_720_port, OTMP_719_port, OTMP_718_port, 
      OTMP_717_port, OTMP_716_port, OTMP_715_port, OTMP_714_port, OTMP_713_port
      , OTMP_712_port, OTMP_711_port, OTMP_710_port, OTMP_709_port, 
      OTMP_708_port, OTMP_707_port, OTMP_706_port, OTMP_705_port, OTMP_704_port
      , OTMP_703_port, OTMP_702_port, OTMP_701_port, OTMP_700_port, 
      OTMP_699_port, OTMP_698_port, OTMP_697_port, OTMP_696_port, OTMP_695_port
      , OTMP_694_port, OTMP_693_port, OTMP_692_port, OTMP_691_port, 
      OTMP_690_port, OTMP_689_port, OTMP_688_port, OTMP_687_port, OTMP_686_port
      , OTMP_685_port, OTMP_684_port, OTMP_683_port, OTMP_682_port, 
      OTMP_681_port, OTMP_680_port, OTMP_679_port, OTMP_678_port, OTMP_677_port
      , OTMP_676_port, OTMP_675_port, OTMP_674_port, OTMP_673_port, 
      OTMP_672_port, OTMP_671_port, OTMP_670_port, OTMP_669_port, OTMP_668_port
      , OTMP_667_port, OTMP_666_port, OTMP_665_port, OTMP_664_port, 
      OTMP_663_port, OTMP_662_port, OTMP_661_port, OTMP_660_port, OTMP_659_port
      , OTMP_658_port, OTMP_657_port, OTMP_656_port, OTMP_655_port, 
      OTMP_654_port, OTMP_653_port, OTMP_652_port, OTMP_651_port, OTMP_650_port
      , OTMP_649_port, OTMP_648_port, OTMP_647_port, OTMP_646_port, 
      OTMP_645_port, OTMP_644_port, OTMP_643_port, OTMP_642_port, OTMP_641_port
      , OTMP_640_port, OTMP_639_port, OTMP_638_port, OTMP_637_port, 
      OTMP_636_port, OTMP_635_port, OTMP_634_port, OTMP_633_port, OTMP_632_port
      , OTMP_631_port, OTMP_630_port, OTMP_629_port, OTMP_628_port, 
      OTMP_627_port, OTMP_626_port, OTMP_625_port, OTMP_624_port, OTMP_623_port
      , OTMP_622_port, OTMP_621_port, OTMP_620_port, OTMP_619_port, 
      OTMP_618_port, OTMP_617_port, OTMP_616_port, OTMP_615_port, OTMP_614_port
      , OTMP_613_port, OTMP_612_port, OTMP_611_port, OTMP_610_port, 
      OTMP_609_port, OTMP_608_port, OTMP_607_port, OTMP_606_port, OTMP_605_port
      , OTMP_604_port, OTMP_603_port, OTMP_602_port, OTMP_601_port, 
      OTMP_600_port, OTMP_599_port, OTMP_598_port, OTMP_597_port, OTMP_596_port
      , OTMP_595_port, OTMP_594_port, OTMP_593_port, OTMP_592_port, 
      OTMP_591_port, OTMP_590_port, OTMP_589_port, OTMP_588_port, OTMP_587_port
      , OTMP_586_port, OTMP_585_port, OTMP_584_port, OTMP_583_port, 
      OTMP_582_port, OTMP_581_port, OTMP_580_port, OTMP_579_port, OTMP_578_port
      , OTMP_577_port, OTMP_576_port, OTMP_575_port, OTMP_574_port, 
      OTMP_573_port, OTMP_572_port, OTMP_571_port, OTMP_570_port, OTMP_569_port
      , OTMP_568_port, OTMP_567_port, OTMP_566_port, OTMP_565_port, 
      OTMP_564_port, OTMP_563_port, OTMP_562_port, OTMP_561_port, OTMP_560_port
      , OTMP_559_port, OTMP_558_port, OTMP_557_port, OTMP_556_port, 
      OTMP_555_port, OTMP_554_port, OTMP_553_port, OTMP_552_port, OTMP_551_port
      , OTMP_550_port, OTMP_549_port, OTMP_548_port, OTMP_547_port, 
      OTMP_546_port, OTMP_545_port, OTMP_544_port, OTMP_543_port, OTMP_542_port
      , OTMP_541_port, OTMP_540_port, OTMP_539_port, OTMP_538_port, 
      OTMP_537_port, OTMP_536_port, OTMP_535_port, OTMP_534_port, OTMP_533_port
      , OTMP_532_port, OTMP_531_port, OTMP_530_port, OTMP_529_port, 
      OTMP_528_port, OTMP_527_port, OTMP_526_port, OTMP_525_port, OTMP_524_port
      , OTMP_523_port, OTMP_522_port, OTMP_521_port, OTMP_520_port, 
      OTMP_519_port, OTMP_518_port, OTMP_517_port, OTMP_516_port, OTMP_515_port
      , OTMP_514_port, OTMP_513_port, OTMP_512_port, PTMP_895_port, 
      PTMP_894_port, PTMP_893_port, PTMP_892_port, PTMP_891_port, PTMP_890_port
      , PTMP_889_port, PTMP_888_port, PTMP_887_port, PTMP_886_port, 
      PTMP_885_port, PTMP_884_port, PTMP_883_port, PTMP_882_port, PTMP_881_port
      , PTMP_880_port, PTMP_879_port, PTMP_878_port, PTMP_877_port, 
      PTMP_876_port, PTMP_875_port, PTMP_874_port, PTMP_873_port, PTMP_872_port
      , PTMP_871_port, PTMP_870_port, PTMP_869_port, PTMP_868_port, 
      PTMP_867_port, PTMP_866_port, PTMP_865_port, PTMP_864_port, PTMP_863_port
      , PTMP_862_port, PTMP_861_port, PTMP_860_port, PTMP_859_port, 
      PTMP_858_port, PTMP_857_port, PTMP_856_port, PTMP_855_port, PTMP_854_port
      , PTMP_853_port, PTMP_852_port, PTMP_851_port, PTMP_850_port, 
      PTMP_849_port, PTMP_848_port, PTMP_847_port, PTMP_846_port, PTMP_845_port
      , PTMP_844_port, PTMP_843_port, PTMP_842_port, PTMP_841_port, 
      PTMP_840_port, PTMP_839_port, PTMP_838_port, PTMP_837_port, PTMP_836_port
      , PTMP_835_port, PTMP_834_port, PTMP_833_port, PTMP_832_port, 
      PTMP_831_port, PTMP_830_port, PTMP_829_port, PTMP_828_port, PTMP_827_port
      , PTMP_826_port, PTMP_825_port, PTMP_824_port, PTMP_823_port, 
      PTMP_822_port, PTMP_821_port, PTMP_820_port, PTMP_819_port, PTMP_818_port
      , PTMP_817_port, PTMP_816_port, PTMP_815_port, PTMP_814_port, 
      PTMP_813_port, PTMP_812_port, PTMP_811_port, PTMP_810_port, PTMP_809_port
      , PTMP_808_port, PTMP_807_port, PTMP_806_port, PTMP_805_port, 
      PTMP_804_port, PTMP_803_port, PTMP_802_port, PTMP_801_port, PTMP_800_port
      , PTMP_799_port, PTMP_798_port, PTMP_797_port, PTMP_796_port, 
      PTMP_795_port, PTMP_794_port, PTMP_793_port, PTMP_792_port, PTMP_791_port
      , PTMP_790_port, PTMP_789_port, PTMP_788_port, PTMP_787_port, 
      PTMP_786_port, PTMP_785_port, PTMP_784_port, PTMP_783_port, PTMP_782_port
      , PTMP_781_port, PTMP_780_port, PTMP_779_port, PTMP_778_port, 
      PTMP_777_port, PTMP_776_port, PTMP_775_port, PTMP_774_port, PTMP_773_port
      , PTMP_772_port, PTMP_771_port, PTMP_770_port, PTMP_769_port, 
      PTMP_768_port, PTMP_767_port, PTMP_766_port, PTMP_765_port, PTMP_764_port
      , PTMP_763_port, PTMP_762_port, PTMP_761_port, PTMP_760_port, 
      PTMP_759_port, PTMP_758_port, PTMP_757_port, PTMP_756_port, PTMP_755_port
      , PTMP_754_port, PTMP_753_port, PTMP_752_port, PTMP_751_port, 
      PTMP_750_port, PTMP_749_port, PTMP_748_port, PTMP_747_port, PTMP_746_port
      , PTMP_745_port, PTMP_744_port, PTMP_743_port, PTMP_742_port, 
      PTMP_741_port, PTMP_740_port, PTMP_739_port, PTMP_738_port, PTMP_737_port
      , PTMP_736_port, PTMP_735_port, PTMP_734_port, PTMP_733_port, 
      PTMP_732_port, PTMP_731_port, PTMP_730_port, PTMP_729_port, PTMP_728_port
      , PTMP_727_port, PTMP_726_port, PTMP_725_port, PTMP_724_port, 
      PTMP_723_port, PTMP_722_port, PTMP_721_port, PTMP_720_port, PTMP_719_port
      , PTMP_718_port, PTMP_717_port, PTMP_716_port, PTMP_715_port, 
      PTMP_714_port, PTMP_713_port, PTMP_712_port, PTMP_711_port, PTMP_710_port
      , PTMP_709_port, PTMP_708_port, PTMP_707_port, PTMP_706_port, 
      PTMP_705_port, PTMP_704_port, PTMP_703_port, PTMP_702_port, PTMP_701_port
      , PTMP_700_port, PTMP_699_port, PTMP_698_port, PTMP_697_port, 
      PTMP_696_port, PTMP_695_port, PTMP_694_port, PTMP_693_port, PTMP_692_port
      , PTMP_691_port, PTMP_690_port, PTMP_689_port, PTMP_688_port, 
      PTMP_687_port, PTMP_686_port, PTMP_685_port, PTMP_684_port, PTMP_683_port
      , PTMP_682_port, PTMP_681_port, PTMP_680_port, PTMP_679_port, 
      PTMP_678_port, PTMP_677_port, PTMP_676_port, PTMP_675_port, PTMP_674_port
      , PTMP_673_port, PTMP_672_port, PTMP_671_port, PTMP_670_port, 
      PTMP_669_port, PTMP_668_port, PTMP_667_port, PTMP_666_port, PTMP_665_port
      , PTMP_664_port, PTMP_663_port, PTMP_662_port, PTMP_661_port, 
      PTMP_660_port, PTMP_659_port, PTMP_658_port, PTMP_657_port, PTMP_656_port
      , PTMP_655_port, PTMP_654_port, PTMP_653_port, PTMP_652_port, 
      PTMP_651_port, PTMP_650_port, PTMP_649_port, PTMP_648_port, PTMP_647_port
      , PTMP_646_port, PTMP_645_port, PTMP_644_port, PTMP_643_port, 
      PTMP_642_port, PTMP_641_port, PTMP_640_port, PTMP_639_port, PTMP_638_port
      , PTMP_637_port, PTMP_636_port, PTMP_635_port, PTMP_634_port, 
      PTMP_633_port, PTMP_632_port, PTMP_631_port, PTMP_630_port, PTMP_629_port
      , PTMP_628_port, PTMP_627_port, PTMP_626_port, PTMP_625_port, 
      PTMP_624_port, PTMP_623_port, PTMP_622_port, PTMP_621_port, PTMP_620_port
      , PTMP_619_port, PTMP_618_port, PTMP_617_port, PTMP_616_port, 
      PTMP_615_port, PTMP_614_port, PTMP_613_port, PTMP_612_port, PTMP_611_port
      , PTMP_610_port, PTMP_609_port, PTMP_608_port, PTMP_607_port, 
      PTMP_606_port, PTMP_605_port, PTMP_604_port, PTMP_603_port, PTMP_602_port
      , PTMP_601_port, PTMP_600_port, PTMP_599_port, PTMP_598_port, 
      PTMP_597_port, PTMP_596_port, PTMP_595_port, PTMP_594_port, PTMP_593_port
      , PTMP_592_port, PTMP_591_port, PTMP_590_port, PTMP_589_port, 
      PTMP_588_port, PTMP_587_port, PTMP_586_port, PTMP_585_port, PTMP_584_port
      , PTMP_583_port, PTMP_582_port, PTMP_581_port, PTMP_580_port, 
      PTMP_579_port, PTMP_578_port, PTMP_577_port, PTMP_576_port, PTMP_575_port
      , PTMP_574_port, PTMP_573_port, PTMP_572_port, PTMP_571_port, 
      PTMP_570_port, PTMP_569_port, PTMP_568_port, PTMP_567_port, PTMP_566_port
      , PTMP_565_port, PTMP_564_port, PTMP_563_port, PTMP_562_port, 
      PTMP_561_port, PTMP_560_port, PTMP_559_port, PTMP_558_port, PTMP_557_port
      , PTMP_556_port, PTMP_555_port, PTMP_554_port, PTMP_553_port, 
      PTMP_552_port, PTMP_551_port, PTMP_550_port, PTMP_549_port, PTMP_548_port
      , PTMP_547_port, PTMP_546_port, PTMP_545_port, PTMP_544_port, 
      PTMP_543_port, PTMP_542_port, PTMP_541_port, PTMP_540_port, PTMP_539_port
      , PTMP_538_port, PTMP_537_port, PTMP_536_port, PTMP_535_port, 
      PTMP_534_port, PTMP_533_port, PTMP_532_port, PTMP_531_port, PTMP_530_port
      , PTMP_529_port, PTMP_528_port, PTMP_527_port, PTMP_526_port, 
      PTMP_525_port, PTMP_524_port, PTMP_523_port, PTMP_522_port, PTMP_521_port
      , PTMP_520_port, PTMP_519_port, PTMP_518_port, PTMP_517_port, 
      PTMP_516_port, PTMP_515_port, PTMP_514_port, PTMP_513_port, PTMP_512_port
      , PTMP_511_port, PTMP_510_port, PTMP_509_port, PTMP_508_port, 
      PTMP_507_port, PTMP_506_port, PTMP_505_port, PTMP_504_port, PTMP_503_port
      , PTMP_502_port, PTMP_501_port, PTMP_500_port, PTMP_499_port, 
      PTMP_498_port, PTMP_497_port, PTMP_496_port, PTMP_495_port, PTMP_494_port
      , PTMP_493_port, PTMP_492_port, PTMP_491_port, PTMP_490_port, 
      PTMP_489_port, PTMP_488_port, PTMP_487_port, PTMP_486_port, PTMP_485_port
      , PTMP_484_port, PTMP_483_port, PTMP_482_port, PTMP_481_port, 
      PTMP_480_port, PTMP_479_port, PTMP_478_port, PTMP_477_port, PTMP_476_port
      , PTMP_475_port, PTMP_474_port, PTMP_473_port, PTMP_472_port, 
      PTMP_471_port, PTMP_470_port, PTMP_469_port, PTMP_468_port, PTMP_467_port
      , PTMP_466_port, PTMP_465_port, PTMP_464_port, PTMP_463_port, 
      PTMP_462_port, PTMP_461_port, PTMP_460_port, PTMP_459_port, PTMP_458_port
      , PTMP_457_port, PTMP_456_port, PTMP_455_port, PTMP_454_port, 
      PTMP_453_port, PTMP_452_port, PTMP_451_port, PTMP_450_port, PTMP_449_port
      , PTMP_448_port, PTMP_447_port, PTMP_446_port, PTMP_445_port, 
      PTMP_444_port, PTMP_443_port, PTMP_442_port, PTMP_441_port, PTMP_440_port
      , PTMP_439_port, PTMP_438_port, PTMP_437_port, PTMP_436_port, 
      PTMP_435_port, PTMP_434_port, PTMP_433_port, PTMP_432_port, PTMP_431_port
      , PTMP_430_port, PTMP_429_port, PTMP_428_port, PTMP_427_port, 
      PTMP_426_port, PTMP_425_port, PTMP_424_port, PTMP_423_port, PTMP_422_port
      , PTMP_421_port, PTMP_420_port, PTMP_419_port, PTMP_418_port, 
      PTMP_417_port, PTMP_416_port, PTMP_415_port, PTMP_414_port, PTMP_413_port
      , PTMP_412_port, PTMP_411_port, PTMP_410_port, PTMP_409_port, 
      PTMP_408_port, PTMP_407_port, PTMP_406_port, PTMP_405_port, PTMP_404_port
      , PTMP_403_port, PTMP_402_port, PTMP_401_port, PTMP_400_port, 
      PTMP_399_port, PTMP_398_port, PTMP_397_port, PTMP_396_port, PTMP_395_port
      , PTMP_394_port, PTMP_393_port, PTMP_392_port, PTMP_391_port, 
      PTMP_390_port, PTMP_389_port, PTMP_388_port, PTMP_387_port, PTMP_386_port
      , PTMP_385_port, PTMP_384_port, PTMP_383_port, PTMP_382_port, 
      PTMP_381_port, PTMP_380_port, PTMP_379_port, PTMP_378_port, PTMP_377_port
      , PTMP_376_port, PTMP_375_port, PTMP_374_port, PTMP_373_port, 
      PTMP_372_port, PTMP_371_port, PTMP_370_port, PTMP_369_port, PTMP_368_port
      , PTMP_367_port, PTMP_366_port, PTMP_365_port, PTMP_364_port, 
      PTMP_363_port, PTMP_362_port, PTMP_361_port, PTMP_360_port, PTMP_359_port
      , PTMP_358_port, PTMP_357_port, PTMP_356_port, PTMP_355_port, 
      PTMP_354_port, PTMP_353_port, PTMP_352_port, PTMP_351_port, PTMP_350_port
      , PTMP_349_port, PTMP_348_port, PTMP_347_port, PTMP_346_port, 
      PTMP_345_port, PTMP_344_port, PTMP_343_port, PTMP_342_port, PTMP_341_port
      , PTMP_340_port, PTMP_339_port, PTMP_338_port, PTMP_337_port, 
      PTMP_336_port, PTMP_335_port, PTMP_334_port, PTMP_333_port, PTMP_332_port
      , PTMP_331_port, PTMP_330_port, PTMP_329_port, PTMP_328_port, 
      PTMP_327_port, PTMP_326_port, PTMP_325_port, PTMP_324_port, PTMP_323_port
      , PTMP_322_port, PTMP_321_port, PTMP_320_port, PTMP_319_port, 
      PTMP_318_port, PTMP_317_port, PTMP_316_port, PTMP_315_port, PTMP_314_port
      , PTMP_313_port, PTMP_312_port, PTMP_311_port, PTMP_310_port, 
      PTMP_309_port, PTMP_308_port, PTMP_307_port, PTMP_306_port, PTMP_305_port
      , PTMP_304_port, PTMP_303_port, PTMP_302_port, PTMP_301_port, 
      PTMP_300_port, PTMP_299_port, PTMP_298_port, PTMP_297_port, PTMP_296_port
      , PTMP_295_port, PTMP_294_port, PTMP_293_port, PTMP_292_port, 
      PTMP_291_port, PTMP_290_port, PTMP_289_port, PTMP_288_port, PTMP_287_port
      , PTMP_286_port, PTMP_285_port, PTMP_284_port, PTMP_283_port, 
      PTMP_282_port, PTMP_281_port, PTMP_280_port, PTMP_279_port, PTMP_278_port
      , PTMP_277_port, PTMP_276_port, PTMP_275_port, PTMP_274_port, 
      PTMP_273_port, PTMP_272_port, PTMP_271_port, PTMP_270_port, PTMP_269_port
      , PTMP_268_port, PTMP_267_port, PTMP_266_port, PTMP_265_port, 
      PTMP_264_port, PTMP_263_port, PTMP_262_port, PTMP_261_port, PTMP_260_port
      , PTMP_259_port, PTMP_258_port, PTMP_257_port, PTMP_256_port, 
      PTMP_255_port, PTMP_254_port, PTMP_253_port, PTMP_252_port, PTMP_251_port
      , PTMP_250_port, PTMP_249_port, PTMP_248_port, PTMP_247_port, 
      PTMP_246_port, PTMP_245_port, PTMP_244_port, PTMP_243_port, PTMP_242_port
      , PTMP_241_port, PTMP_240_port, PTMP_239_port, PTMP_238_port, 
      PTMP_237_port, PTMP_236_port, PTMP_235_port, PTMP_234_port, PTMP_233_port
      , PTMP_232_port, PTMP_231_port, PTMP_230_port, PTMP_229_port, 
      PTMP_228_port, PTMP_227_port, PTMP_226_port, PTMP_225_port, PTMP_224_port
      , PTMP_223_port, PTMP_222_port, PTMP_221_port, PTMP_220_port, 
      PTMP_219_port, PTMP_218_port, PTMP_217_port, PTMP_216_port, PTMP_215_port
      , PTMP_214_port, PTMP_213_port, PTMP_212_port, PTMP_211_port, 
      PTMP_210_port, PTMP_209_port, PTMP_208_port, PTMP_207_port, PTMP_206_port
      , PTMP_205_port, PTMP_204_port, PTMP_203_port, PTMP_202_port, 
      PTMP_201_port, PTMP_200_port, PTMP_199_port, PTMP_198_port, PTMP_197_port
      , PTMP_196_port, PTMP_195_port, PTMP_194_port, PTMP_193_port, 
      PTMP_192_port, PTMP_191_port, PTMP_190_port, PTMP_189_port, PTMP_188_port
      , PTMP_187_port, PTMP_186_port, PTMP_185_port, PTMP_184_port, 
      PTMP_183_port, PTMP_182_port, PTMP_181_port, PTMP_180_port, PTMP_179_port
      , PTMP_178_port, PTMP_177_port, PTMP_176_port, PTMP_175_port, 
      PTMP_174_port, PTMP_173_port, PTMP_172_port, PTMP_171_port, PTMP_170_port
      , PTMP_169_port, PTMP_168_port, PTMP_167_port, PTMP_166_port, 
      PTMP_165_port, PTMP_164_port, PTMP_163_port, PTMP_162_port, PTMP_161_port
      , PTMP_160_port, PTMP_159_port, PTMP_158_port, PTMP_157_port, 
      PTMP_156_port, PTMP_155_port, PTMP_154_port, PTMP_153_port, PTMP_152_port
      , PTMP_151_port, PTMP_150_port, PTMP_149_port, PTMP_148_port, 
      PTMP_147_port, PTMP_146_port, PTMP_145_port, PTMP_144_port, PTMP_143_port
      , PTMP_142_port, PTMP_141_port, PTMP_140_port, PTMP_139_port, 
      PTMP_138_port, PTMP_137_port, PTMP_136_port, PTMP_135_port, PTMP_134_port
      , PTMP_133_port, PTMP_132_port, PTMP_131_port, PTMP_130_port, 
      PTMP_129_port, PTMP_128_port, PTMP_127_port, PTMP_126_port, PTMP_125_port
      , PTMP_124_port, PTMP_123_port, PTMP_122_port, PTMP_121_port, 
      PTMP_120_port, PTMP_119_port, PTMP_118_port, PTMP_117_port, PTMP_116_port
      , PTMP_115_port, PTMP_114_port, PTMP_113_port, PTMP_112_port, 
      PTMP_111_port, PTMP_110_port, PTMP_109_port, PTMP_108_port, PTMP_107_port
      , PTMP_106_port, PTMP_105_port, PTMP_104_port, PTMP_103_port, 
      PTMP_102_port, PTMP_101_port, PTMP_100_port, PTMP_99_port, PTMP_98_port, 
      PTMP_97_port, PTMP_96_port, PTMP_95_port, PTMP_94_port, PTMP_93_port, 
      PTMP_92_port, PTMP_91_port, PTMP_90_port, PTMP_89_port, PTMP_88_port, 
      PTMP_87_port, PTMP_86_port, PTMP_85_port, PTMP_84_port, PTMP_83_port, 
      PTMP_82_port, PTMP_81_port, PTMP_80_port, PTMP_79_port, PTMP_78_port, 
      PTMP_77_port, PTMP_76_port, PTMP_75_port, PTMP_74_port, PTMP_73_port, 
      PTMP_72_port, PTMP_71_port, PTMP_70_port, PTMP_69_port, PTMP_68_port, 
      PTMP_67_port, PTMP_66_port, PTMP_65_port, PTMP_64_port, PTMP_63_port, 
      PTMP_62_port, PTMP_61_port, PTMP_60_port, PTMP_59_port, PTMP_58_port, 
      PTMP_57_port, PTMP_56_port, PTMP_55_port, PTMP_54_port, PTMP_53_port, 
      PTMP_52_port, PTMP_51_port, PTMP_50_port, PTMP_49_port, PTMP_48_port, 
      PTMP_47_port, PTMP_46_port, PTMP_45_port, PTMP_44_port, PTMP_43_port, 
      PTMP_42_port, PTMP_41_port, PTMP_40_port, PTMP_39_port, PTMP_38_port, 
      PTMP_37_port, PTMP_36_port, PTMP_35_port, PTMP_34_port, PTMP_33_port, 
      PTMP_32_port, PTMP_31_port, PTMP_30_port, PTMP_29_port, PTMP_28_port, 
      PTMP_27_port, PTMP_26_port, PTMP_25_port, PTMP_24_port, PTMP_23_port, 
      PTMP_22_port, PTMP_21_port, PTMP_20_port, PTMP_19_port, PTMP_18_port, 
      PTMP_17_port, PTMP_16_port, PTMP_15_port, PTMP_14_port, PTMP_13_port, 
      PTMP_12_port, PTMP_11_port, PTMP_10_port, PTMP_9_port, PTMP_8_port, 
      PTMP_7_port, PTMP_6_port, PTMP_5_port, PTMP_4_port, PTMP_3_port, 
      PTMP_2_port, PTMP_1_port, PTMP_0_port, net46772, net46773, net46774, 
      net46775, net46776, net46777, net46778, net46779, net46780, net46781, 
      net46782, net46783, net46784, net46785, net46786, net46787, net46788, 
      net46789, net46790, net46791, net46792, net46793, net46794, net46795, 
      net46796, net46797, net46798, net46799, net46800, net46801, net46802, 
      net46803, net46804, net46805, net46806, net46807, net46808, net46809, 
      net46810, net46811, net46812, net46813, net46814, net46815, net46816, 
      net46817, net46818, net46819, net46820, net46821, net46822, net46823, 
      net46824, net46825, net46826, net46827, net46828, net46829, net46830, 
      net46831, net46832, net46833, net46834, net46835, net46836, net46837, 
      net46838, net46839, net46840, net46841, net46842, net46843, net46844, 
      net46845, net46846, net46847, net46848, net46849, net46850, net46851, 
      net46852, net46853, net46854, net46855, net46856, net46857, net46858, 
      net46859, net46860, net46861, net46862, net46863, net46864, net46865, 
      net46866, net46867, net46868, net46869, net46870, net46871, net46872, 
      net46873, net46874, net46875, net46876, net46877, net46878, net46879, 
      net46880, net46881, net46882, net46883, net46884, net46885, net46886, 
      net46887, net46888, net46889, net46890, net46891, net46892, net46893, 
      net46894, net46895, net46896, net46897, net46898, net46899, net46900, 
      net46901, net46902, net46903, net46904, net46905, net46906, net46907, 
      net46908, net46909, net46910, net46911, net46912, net46913, net46914, 
      net46915, net46916, net46917, net46918, net46919, net46920, net46921, 
      net46922, net46923, net46924, net46925, net46926, net46927, net46928, 
      net46929, net46930, net46931, net46932, net46933, net46934, net46935, 
      net46936, net46937, net46938, net46939, net46940, net46941, net46942, 
      net46943, net46944, net46945, net46946, net46947, net46948, net46949, 
      net46950, net46951, net46952, net46953, net46954, net46955, net46956, 
      net46957, net46958, net46959, net46960, net46961, net46962, net46963, 
      net46964, net46965, net46966, net46967, net46968, net46969, net46970, 
      net46971, net46972, net46973, net46974, net46975, net46976, net46977, 
      net46978, net46979, net46980, net46981, net46982, net46983, net46984, 
      net46985, net46986, net46987, net46988, net46989, net46990, net46991, 
      net46992, net46993, net46994, net46995, net46996, net46997, net46998, 
      net46999, net47000, net47001, net47002, net47003, net47004, net47005, 
      net47006, net47007, net47008, net47009, net47010, net47011, net47012, 
      net47013, net47014, net47015, net47016, net47017, net47018, net47019, 
      net47020, net47021, net47022, net47023, net47024, net47025, net47026, 
      net47027, net47028, net47029, net47030, net47031, net47032, net47033, 
      net47034, net47035, net47036, net47037, net47038, net47039, net47040, 
      net47041, net47042, net47043, net47044, net47045, net47046, net47047, 
      net47048, net47049, net47050, net47051, net47052, net47053, net47054, 
      net47055, net47056, net47057, net47058, net47059, net47060, net47061, 
      net47062, net47063, net47064, net47065, net47066, net47067, net47068, 
      net47069, net47070, net47071, net47072, net47073, net47074, net47075, 
      net47076, net47077, net47078, net47079, net47080, net47081, net47082, 
      net47083, net47084, net47085, net47086, net47087, net47088, net47089, 
      net47090, net47091, net47092, net47093, net47094, net47095, net47096, 
      net47097, net47098, net47099, net47100, net47101, net47102, net47103, 
      net47104, net47105, net47106, net47107, net47108, net47109, net47110, 
      net47111, net47112, net47113, net47114, net47115, net47116, net47117, 
      net47118, net47119, net47120, net47121, net47122, net47123, net47124, 
      net47125, net47126, net47127, net47128, net47129, net47130, net47131, 
      net47132, net47133, net47134, net47135, net47136, net47137, net47138, 
      net47139, net47140, net47141, net47142, net47143, net47144, net47145, 
      net47146, net47147, net47148, net47149, net47150, net47151, net47152, 
      net47153, net47154, net47155, net47156, net47157, net47158, net47159, 
      net47160, net47161, net47162, net47163, net47164, net47165, net47166, 
      net47167, net47168, net47169, net47170, net47171, net47172, net47173, 
      net47174, net47175, net47176, net47177, net47178, net47179, net47180, 
      net47181, net47182, net47183, net47184, net47185, net47186, net47187, 
      net47188, net47189, net47190, net47191, net47192, net47193, net47194, 
      net47195, net47196, net47197, net47198, net47199, net47200, net47201, 
      net47202, net47203, net47204, net47205, net47206, net47207, net47208, 
      net47209, net47210, net47211, net47212, net47213, net47214, net47215, 
      net47216, net47217, net47218, net47219, net47220, net47221, net47222, 
      net47223, net47224, net47225, net47226, net47227, net47228, net47229, 
      net47230, net47231, net47232, net47233, net47234, net47235, net47236, 
      net47237, net47238, net47239, net47240, net47241, net47242, net47243, 
      net47244, net47245, net47246, net47247, net47248, net47249, net47250, 
      net47251, net47252, net47253, net47254, net47255, net47256, net47257, 
      net47258, net47259, net47260, net47261, net47262, net47263, net47264, 
      net47265, net47266, net47267, net47268, net47269, net47270, net47271, 
      net47272, net47273, net47274, net47275, net47276, net47277, net47278, 
      net47279, net47280, net47281, net47282, net47283, net47284, net47285, 
      net47286, net47287, net47288, net47289, net47290, net47291, net47292, 
      net47293, net47294, net47295, net47296, net47297, net47298, net47299, 
      net47300, net47301, net47302, net47303, net47304, net47305, net47306, 
      net47307, net47308, net47309, net47310, net47311, net47312, net47313, 
      net47314, net47315, net47316, net47317, net47318, net47319, net47320, 
      net47321, net47322, net47323, net47324, net47325, net47326, net47327, 
      net47328, net47329, net47330, net47331, net47332, net47333, net47334, 
      net47335, net47336, net47337, net47338, net47339, net47340, net47341, 
      net47342, net47343, net47344, net47345, net47346, net47347, net47348, 
      net47349, net47350, net47351, net47352, net47353, net47354, net47355, 
      net47356, net47357, net47358, net47359, net47360, net47361, net47362, 
      net47363, net47364, net47365, net47366, net47367, net47368, net47369, 
      net47370, net47371, net47372, net47373, net47374, net47375, net47376, 
      net47377, net47378, net47379, net47380, net47381, net47382, net47383, 
      net47384, net47385, net47386, net47387, net47388, net47389, net47390, 
      net47391, net47392, net47393, net47394, net47395, net47396, net47397, 
      net47398, net47399, net47400, net47401, net47402, net47403, net47404, 
      net47405, net47406, net47407, net47408, net47409, net47410, net47411, 
      net47412, net47413, net47414, net47415, net47416, net47417, net47418, 
      net47419, net47420, net47421, net47422, net47423, net47424, net47425, 
      net47426, net47427, net47428, net47429, net47430, net47431, net47432, 
      net47433, net47434, net47435, net47436, net47437, net47438, net47439, 
      net47440, net47441, net47442, net47443, net47444, net47445, net47446, 
      net47447, net47448, net47449, net47450, net47451, net47452, net47453, 
      net47454, net47455, net47456, net47457, net47458, net47459, net47460, 
      net47461, net47462, net47463, net47464, net47465, net47466, net47467, 
      net47468, net47469, net47470, net47471, net47472, net47473, net47474, 
      net47475, net47476, net47477, net47478, net47479, net47480, net47481, 
      net47482, net47483, net47484, net47485, net47486, net47487, net47488, 
      net47489, net47490, net47491, net47492, net47493, net47494, net47495, 
      net47496, net47497, net47498, net47499, net47500, net47501, net47502, 
      net47503, net47504, net47505, net47506, net47507, net47508, net47509, 
      net47510, net47511, net47512, net47513, net47514, net47515, net47516, 
      net47517, net47518, net47519, net47520, net47521, net47522, net47523, 
      net47524, net47525, net47526, net47527, net47528, net47529, net47530, 
      net47531, net47532, net47533, net47534, net47535, net47536, net47537, 
      net47538, net47539, net47540, net47541, net47542, net47543, net47544, 
      net47545, net47546, net47547, net47548, net47549, net47550, net47551, 
      net47552, net47553, net47554, net47555, net47556, net47557, net47558, 
      net47559, net47560, net47561, net47562, net47563, net47564, net47565, 
      net47566, net47567, net47568, net47569, net47570, net47571, net47572, 
      net47573, net47574, net47575, net47576, net47577, net47578, net47579, 
      net47580, net47581, net47582, net47583, net47584, net47585, net47586, 
      net47587, net47588, net47589, net47590, net47591, net47592, net47593, 
      net47594, net47595, net47596, net47597, net47598, net47599, net47600, 
      net47601, net47602, net47603, net47604, net47605, net47606, net47607, 
      net47608, net47609, net47610, net47611, net47612, net47613, net47614, 
      net47615, net47616, net47617, net47618, net47619, net47620, net47621, 
      net47622, net47623, net47624, net47625, net47626, net47627, net47628, 
      net47629, net47630, net47631, net47632, net47633, net47634, net47635, 
      net47636, net47637, net47638, net47639, net47640, net47641, net47642, 
      net47643, net47644, net47645, net47646, net47647, net47648, net47649, 
      net47650, net47651, net47652, net47653, net47654, net47655, net47656, 
      net47657, net47658, net47659, net47660, net47661, net47662, net47663, 
      net47664, net47665, net47666, net47667, net47668, net47669, net47670, 
      net47671, net47672, net47673, net47674, net47675, net47676, net47677, 
      net47678, net47679, net47680, net47681, net47682, net47683, net47684, 
      net47685, net47686, net47687, net47688, net47689, net47690, net47691, 
      net47692, net47693, net47694, net47695, net47696, net47697, net47698, 
      net47699, net47700, net47701, net47702, net47703, net47704, net47705, 
      net47706, net47707, net47708, net47709, net47710, net47711, net47712, 
      net47713, net47714, net47715, net47716, net47717, net47718, net47719, 
      net47720, net47721, net47722, net47723, net47724, net47725, net47726, 
      net47727, net47728, net47729, net47730, net47731, net47732, net47733, 
      net47734, net47735, net47736, net47737, net47738, net47739, net47740, 
      net47741, net47742, net47743, net47744, net47745, net47746, net47747, 
      net47748, net47749, net47750, net47751, net47752, net47753, net47754, 
      net47755, net47756, net47757, net47758, net47759, net47760, net47761, 
      net47762, net47763, net47764, net47765, net47766, net47767, net47768, 
      net47769, net47770, net47771, net47772, net47773, net47774, net47775, 
      net47776, net47777, net47778, net47779, net47780, net47781, net47782, 
      net47783, net47784, net47785, net47786, net47787, net47788, net47789, 
      net47790, net47791, net47792, net47793, net47794, net47795, net47796, 
      net47797, net47798, net47799, net47800, net47801, net47802, net47803, 
      net47804, net47805, net47806, net47807, net47808, net47809, net47810, 
      net47811, net47812, net47813, net47814, net47815, net47816, net47817, 
      net47818, net47819, net47820, net47821, net47822, net47823, net47824, 
      net47825, net47826, net47827, net47828, net47829, net47830, net47831, 
      net47832, net47833, net47834, net47835, net47836, net47837, net47838, 
      net47839, net47840, net47841, net47842, net47843, net47844, net47845, 
      net47846, net47847, net47848, net47849, net47850, net47851, net47852, 
      net47853, net47854, net47855, net47856, net47857, net47858, net47859, 
      net47860, net47861, net47862, net47863, net47864, net47865, net47866, 
      net47867, net47868, net47869, net47870, net47871, net47872, net47873, 
      net47874, net47875, net47876, net47877, net47878, net47879, net47880, 
      net47881, net47882, net47883, net47884, net47885, net47886, net47887, 
      net47888, net47889, net47890, net47891, net47892, net47893, net47894, 
      net47895, net47896, net47897, net47898, net47899, net47900, net47901, 
      net47902, net47903, net47904, net47905, net47906, net47907, net47908, 
      net47909, net47910, net47911, net47912, net47913, net47914, net47915, 
      net47916, net47917, net47918, net47919, net47920, net47921, net47922, 
      net47923, net47924, net47925, net47926, net47927, net47928, net47929, 
      net47930, net47931, net47932, net47933, net47934, net47935, net47936, 
      net47937, net47938, net47939, net47940, net47941, net47942, net47943, 
      net47944, net47945, net47946, net47947, net47948, net47949, net47950, 
      net47951, net47952, net47953, net47954, net47955, net47956, net47957, 
      net47958, net47959, net47960, net47961, net47962, net47963, net47964, 
      net47965, net47966, net47967, net47968, net47969, net47970, net47971, 
      net47972, net47973, net47974, net47975, net47976, net47977, net47978, 
      net47979, net47980, net47981, net47982, net47983, net47984, net47985, 
      net47986, net47987, net47988, net47989, net47990, net47991, net47992, 
      net47993, net47994, net47995, net47996, net47997, net47998, net47999, 
      net48000, net48001, net48002, net48003, net48004, net48005, net48006, 
      net48007, net48008, net48009, net48010, net48011, net48012, net48013, 
      net48014, net48015, net48016, net48017, net48018, net48019, net48020, 
      net48021, net48022, net48023, net48024, net48025, net48026, net48027, 
      net48028, net48029, net48030, net48031, net48032, net48033, net48034, 
      net48035, net48036, net48037, net48038, net48039, net48040, net48041, 
      net48042, net48043, net48044, net48045, net48046, net48047, net48048, 
      net48049, net48050, net48051, net48052, net48053, net48054, net48055, 
      net48056, net48057, net48058, net48059, net48060, net48061, net48062, 
      net48063, net48064, net48065, net48066, net48067, net48068, net48069, 
      net48070, net48071, net48072, net48073, net48074, net48075, net48076, 
      net48077, net48078, net48079, net48080, net48081, net48082, net48083, 
      net48084, net48085, net48086, net48087, net48088, net48089, net48090, 
      net48091, net48092, net48093, net48094, net48095, net48096, net48097, 
      net48098, net48099, net48100, net48101, net48102, net48103, net48104, 
      net48105, net48106, net48107, net48108, net48109, net48110, net48111, 
      net48112, net48113, net48114, net48115, net48116, net48117, net48118, 
      net48119, net48120, net48121, net48122, net48123, net48124, net48125, 
      net48126, net48127, net48128, net48129, net48130, net48131, net48132, 
      net48133, net48134, net48135, net48136, net48137, net48138, net48139, 
      net48140, net48141, net48142, net48143, net48144, net48145, net48146, 
      net48147, net48148, net48149, net48150, net48151, net48152, net48153, 
      net48154, net48155, net48156, net48157, net48158, net48159, net48160, 
      net48161, net48162, net48163, net48164, net48165, net48166, net48167, 
      net48168, net48169, net48170, net48171, net48172, net48173, net48174, 
      net48175, net48176, net48177, net48178, net48179, net48180, net48181, 
      net48182, net48183, net48184, net48185, net48186, net48187, net48188, 
      net48189, net48190, net48191, net48192, net48193, net48194, net48195, 
      net48196, net48197, net48198, net48199, net48200, net48201, net48202, 
      net48203, net48204, net48205, net48206, net48207, net48208, net48209, 
      net48210, net48211, net48212, net48213, net48214, net48215, net48216, 
      net48217, net48218, net48219, net48220, net48221, net48222, net48223, 
      net48224, net48225, net48226, net48227, net48228, net48229, net48230, 
      net48231, net48232, net48233, net48234, net48235, net48236, net48237, 
      net48238, net48239, net48240, net48241, net48242, net48243, net48244, 
      net48245, net48246, net48247, net48248, net48249, net48250, net48251, 
      net48252, net48253, net48254, net48255, net48256, net48257, net48258, 
      net48259, net48260, net48261, net48262, net48263, net48264, net48265, 
      net48266, net48267, net48268, net48269, net48270, net48271, net48272, 
      net48273, net48274, net48275, net48276, net48277, net48278, net48279, 
      net48280, net48281, net48282, net48283, net48284, net48285, net48286, 
      net48287, net48288, net48289, net48290, net48291, net48292, net48293, 
      net48294, net48295, net48296, net48297, net48298, net48299, net48300, 
      net48301, net48302, net48303, net48304, net48305, net48306, net48307, 
      net48308, net48309, net48310, net48311, net48312, net48313, net48314, 
      net48315, net48316, net48317, net48318, net48319, net48320, net48321, 
      net48322, net48323, net48324, net48325, net48326, net48327, net48328, 
      net48329, net48330, net48331, net48332, net48333, net48334, net48335, 
      net48336, net48337, net48338, net48339, net48340, net48341, net48342, 
      net48343, net48344, net48345, net48346, net48347, net48348, net48349, 
      net48350, net48351, net48352, net48353, net48354, net48355, net48356, 
      net48357, net48358, net48359, net48360, net48361, net48362, net48363, 
      net48364, net48365, net48366, net48367, net48368, net48369, net48370, 
      net48371, net48372, net48373, net48374, net48375, net48376, net48377, 
      net48378, net48379, net48380, net48381, net48382, net48383, net48384, 
      net48385, net48386, net48387, net48388, net48389, net48390, net48391, 
      net48392, net48393, net48394, net48395, net48396, net48397, net48398, 
      net48399, net48400, net48401, net48402, net48403, net48404, net48405, 
      net48406, net48407, net48408, net48409, net48410, net48411, net48412, 
      net48413, net48414, net48415, net48416, net48417, net48418, net48419, 
      net48420, net48421, net48422, net48423, net48424, net48425, net48426, 
      net48427, net48428, net48429, net48430, net48431, net48432, net48433, 
      net48434, net48435, net48436, net48437, net48438, net48439, net48440, 
      net48441, net48442, net48443, net48444, net48445, net48446, net48447, 
      net48448, net48449, net48450, net48451, net48452, net48453, net48454, 
      net48455, net48456, net48457, net48458, net48459, net48460, net48461, 
      net48462, net48463, net48464, net48465, net48466, net48467, net48468, 
      net48469, net48470, net48471, net48472, net48473, net48474, net48475, 
      net48476, net48477, net48478, net48479, net48480, net48481, net48482, 
      net48483, net48484, net48485, net48486, net48487, net48488, net48489, 
      net48490, net48491, net48492, net48493, net48494, net48495, net48496, 
      net48497, net48498, net48499, net48500, net48501, net48502, net48503, 
      net48504, net48505, net48506, net48507, net48508, net48509, net48510, 
      net48511, net48512, net48513, net48514, net48515, net48516, net48517, 
      net48518, net48519, net48520, net48521, net48522, net48523, net48524, 
      net48525, net48526, net48527, net48528, net48529, net48530, net48531, 
      net48532, net48533, net48534, net48535, net48536, net48537, net48538, 
      net48539, net48540, net48541, net48542, net48543, net48544, net48545, 
      net48546, net48547, net48548, net48549, net48550, net48551, net48552, 
      net48553, net48554, net48555, net48556, net48557, net48558, net48559, 
      net48560, net48561, net48562, net48563, net48564, net48565, net48566, 
      net48567, net48568, net48569, net48570, net48571, net48572, net48573, 
      net48574, net48575, net48576, net48577, net48578, net48579, net48580, 
      net48581, net48582, net48583, net48584, net48585, net48586, net48587, 
      net48588, net48589, net48590, net48591, net48592, net48593, net48594, 
      net48595, net48596, net48597, net48598, net48599, net48600, net48601, 
      net48602, net48603, net48604, net48605, net48606, net48607, net48608, 
      net48609, net48610, net48611, net48612, net48613, net48614, net48615, 
      net48616, net48617, net48618, net48619, net48620, net48621, net48622, 
      net48623, net48624, net48625, net48626, net48627, net48628, net48629, 
      net48630, net48631, net48632, net48633, net48634, net48635, net48636, 
      net48637, net48638, net48639, net48640, net48641, net48642, net48643, 
      net48644, net48645, net48646, net48647, net48648, net48649, net48650, 
      net48651, net48652, net48653, net48654, net48655, net48656, net48657, 
      net48658, net48659, net48660, net48661, net48662, net48663, net48664, 
      net48665, net48666, net48667, net48668, net48669, net48670, net48671, 
      net48672, net48673, net48674, net48675, net48676, net48677, net48678, 
      net48679, net48680, net48681, net48682, net48683, net48684, net48685, 
      net48686, net48687, net48688, net48689, net48690, net48691, net48692, 
      net48693, net48694, net48695, net48696, net48697, net48698, net48699, 
      net48700, net48701, net48702, net48703, net48704, net48705, net48706, 
      net48707, net48708, net48709, net48710, net48711, net48712, net48713, 
      net48714, net48715, net48716, net48717, net48718, net48719, net48720, 
      net48721, net48722, net48723, net48724, net48725, net48726, net48727, 
      net48728, net48729, net48730, net48731, net48732, net48733, net48734, 
      net48735, net48736, net48737, net48738, net48739, net48740, net48741, 
      net48742, net48743, net48744, net48745, net48746, net48747, net48748, 
      net48749, net48750, net48751, net48752, net48753, net48754, net48755, 
      net48756, net48757, net48758, net48759, net48760, net48761, net48762, 
      net48763, net48764, net48765, net48766, net48767, net48768, net48769, 
      net48770, net48771, net48772, net48773, net48774, net48775, net48776, 
      net48777, net48778, net48779, net48780, net48781, net48782, net48783, 
      net48784, net48785, net48786, net48787, net48788, net48789, net48790, 
      net48791, net48792, net48793, net48794, net48795, net48796, net48797, 
      net48798, net48799, net48800, net48801, net48802, net48803, net48804, 
      net48805, net48806, net48807, net48808, net48809, net48810, net48811, 
      net48812, net48813, net48814, net48815, net48816, net48817, net48818, 
      net48819, n4, n5, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100,
      n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, 
      n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, 
      n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, 
      n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, 
      n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, 
      n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, 
      n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, 
      n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, 
      n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, 
      n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, 
      n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, 
      n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, 
      n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, 
      n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, 
      n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, 
      n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, 
      n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, 
      n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, 
      n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, 
      n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, 
      n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, 
      n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, 
      n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, 
      n_1308, n_1309, n_1310 : std_logic;

begin
   
   X_Logic0_port <= '0';
   net46772 <= '0';
   net46773 <= '0';
   net46774 <= '0';
   net46775 <= '0';
   net46776 <= '0';
   net46777 <= '0';
   net46778 <= '0';
   net46779 <= '0';
   net46780 <= '0';
   net46781 <= '0';
   net46782 <= '0';
   net46783 <= '0';
   net46784 <= '0';
   net46785 <= '0';
   net46786 <= '0';
   net46787 <= '0';
   net46788 <= '0';
   net46789 <= '0';
   net46790 <= '0';
   net46791 <= '0';
   net46792 <= '0';
   net46793 <= '0';
   net46794 <= '0';
   net46795 <= '0';
   net46796 <= '0';
   net46797 <= '0';
   net46798 <= '0';
   net46799 <= '0';
   net46800 <= '0';
   net46801 <= '0';
   net46802 <= '0';
   net46803 <= '0';
   net46804 <= '0';
   net46805 <= '0';
   net46806 <= '0';
   net46807 <= '0';
   net46808 <= '0';
   net46809 <= '0';
   net46810 <= '0';
   net46811 <= '0';
   net46812 <= '0';
   net46813 <= '0';
   net46814 <= '0';
   net46815 <= '0';
   net46816 <= '0';
   net46817 <= '0';
   net46818 <= '0';
   net46819 <= '0';
   net46820 <= '0';
   net46821 <= '0';
   net46822 <= '0';
   net46823 <= '0';
   net46824 <= '0';
   net46825 <= '0';
   net46826 <= '0';
   net46827 <= '0';
   net46828 <= '0';
   net46829 <= '0';
   net46830 <= '0';
   net46831 <= '0';
   net46832 <= '0';
   net46833 <= '0';
   net46834 <= '0';
   net46835 <= '0';
   net46836 <= '0';
   net46837 <= '0';
   net46838 <= '0';
   net46839 <= '0';
   net46840 <= '0';
   net46841 <= '0';
   net46842 <= '0';
   net46843 <= '0';
   net46844 <= '0';
   net46845 <= '0';
   net46846 <= '0';
   net46847 <= '0';
   net46848 <= '0';
   net46849 <= '0';
   net46850 <= '0';
   net46851 <= '0';
   net46852 <= '0';
   net46853 <= '0';
   net46854 <= '0';
   net46855 <= '0';
   net46856 <= '0';
   net46857 <= '0';
   net46858 <= '0';
   net46859 <= '0';
   net46860 <= '0';
   net46861 <= '0';
   net46862 <= '0';
   net46863 <= '0';
   net46864 <= '0';
   net46865 <= '0';
   net46866 <= '0';
   net46867 <= '0';
   net46868 <= '0';
   net46869 <= '0';
   net46870 <= '0';
   net46871 <= '0';
   net46872 <= '0';
   net46873 <= '0';
   net46874 <= '0';
   net46875 <= '0';
   net46876 <= '0';
   net46877 <= '0';
   net46878 <= '0';
   net46879 <= '0';
   net46880 <= '0';
   net46881 <= '0';
   net46882 <= '0';
   net46883 <= '0';
   net46884 <= '0';
   net46885 <= '0';
   net46886 <= '0';
   net46887 <= '0';
   net46888 <= '0';
   net46889 <= '0';
   net46890 <= '0';
   net46891 <= '0';
   net46892 <= '0';
   net46893 <= '0';
   net46894 <= '0';
   net46895 <= '0';
   net46896 <= '0';
   net46897 <= '0';
   net46898 <= '0';
   net46899 <= '0';
   net46900 <= '0';
   net46901 <= '0';
   net46902 <= '0';
   net46903 <= '0';
   net46904 <= '0';
   net46905 <= '0';
   net46906 <= '0';
   net46907 <= '0';
   net46908 <= '0';
   net46909 <= '0';
   net46910 <= '0';
   net46911 <= '0';
   net46912 <= '0';
   net46913 <= '0';
   net46914 <= '0';
   net46915 <= '0';
   net46916 <= '0';
   net46917 <= '0';
   net46918 <= '0';
   net46919 <= '0';
   net46920 <= '0';
   net46921 <= '0';
   net46922 <= '0';
   net46923 <= '0';
   net46924 <= '0';
   net46925 <= '0';
   net46926 <= '0';
   net46927 <= '0';
   net46928 <= '0';
   net46929 <= '0';
   net46930 <= '0';
   net46931 <= '0';
   net46932 <= '0';
   net46933 <= '0';
   net46934 <= '0';
   net46935 <= '0';
   net46936 <= '0';
   net46937 <= '0';
   net46938 <= '0';
   net46939 <= '0';
   net46940 <= '0';
   net46941 <= '0';
   net46942 <= '0';
   net46943 <= '0';
   net46944 <= '0';
   net46945 <= '0';
   net46946 <= '0';
   net46947 <= '0';
   net46948 <= '0';
   net46949 <= '0';
   net46950 <= '0';
   net46951 <= '0';
   net46952 <= '0';
   net46953 <= '0';
   net46954 <= '0';
   net46955 <= '0';
   net46956 <= '0';
   net46957 <= '0';
   net46958 <= '0';
   net46959 <= '0';
   net46960 <= '0';
   net46961 <= '0';
   net46962 <= '0';
   net46963 <= '0';
   net46964 <= '0';
   net46965 <= '0';
   net46966 <= '0';
   net46967 <= '0';
   net46968 <= '0';
   net46969 <= '0';
   net46970 <= '0';
   net46971 <= '0';
   net46972 <= '0';
   net46973 <= '0';
   net46974 <= '0';
   net46975 <= '0';
   net46976 <= '0';
   net46977 <= '0';
   net46978 <= '0';
   net46979 <= '0';
   net46980 <= '0';
   net46981 <= '0';
   net46982 <= '0';
   net46983 <= '0';
   net46984 <= '0';
   net46985 <= '0';
   net46986 <= '0';
   net46987 <= '0';
   net46988 <= '0';
   net46989 <= '0';
   net46990 <= '0';
   net46991 <= '0';
   net46992 <= '0';
   net46993 <= '0';
   net46994 <= '0';
   net46995 <= '0';
   net46996 <= '0';
   net46997 <= '0';
   net46998 <= '0';
   net46999 <= '0';
   net47000 <= '0';
   net47001 <= '0';
   net47002 <= '0';
   net47003 <= '0';
   net47004 <= '0';
   net47005 <= '0';
   net47006 <= '0';
   net47007 <= '0';
   net47008 <= '0';
   net47009 <= '0';
   net47010 <= '0';
   net47011 <= '0';
   net47012 <= '0';
   net47013 <= '0';
   net47014 <= '0';
   net47015 <= '0';
   net47016 <= '0';
   net47017 <= '0';
   net47018 <= '0';
   net47019 <= '0';
   net47020 <= '0';
   net47021 <= '0';
   net47022 <= '0';
   net47023 <= '0';
   net47024 <= '0';
   net47025 <= '0';
   net47026 <= '0';
   net47027 <= '0';
   net47028 <= '0';
   net47029 <= '0';
   net47030 <= '0';
   net47031 <= '0';
   net47032 <= '0';
   net47033 <= '0';
   net47034 <= '0';
   net47035 <= '0';
   net47036 <= '0';
   net47037 <= '0';
   net47038 <= '0';
   net47039 <= '0';
   net47040 <= '0';
   net47041 <= '0';
   net47042 <= '0';
   net47043 <= '0';
   net47044 <= '0';
   net47045 <= '0';
   net47046 <= '0';
   net47047 <= '0';
   net47048 <= '0';
   net47049 <= '0';
   net47050 <= '0';
   net47051 <= '0';
   net47052 <= '0';
   net47053 <= '0';
   net47054 <= '0';
   net47055 <= '0';
   net47056 <= '0';
   net47057 <= '0';
   net47058 <= '0';
   net47059 <= '0';
   net47060 <= '0';
   net47061 <= '0';
   net47062 <= '0';
   net47063 <= '0';
   net47064 <= '0';
   net47065 <= '0';
   net47066 <= '0';
   net47067 <= '0';
   net47068 <= '0';
   net47069 <= '0';
   net47070 <= '0';
   net47071 <= '0';
   net47072 <= '0';
   net47073 <= '0';
   net47074 <= '0';
   net47075 <= '0';
   net47076 <= '0';
   net47077 <= '0';
   net47078 <= '0';
   net47079 <= '0';
   net47080 <= '0';
   net47081 <= '0';
   net47082 <= '0';
   net47083 <= '0';
   net47084 <= '0';
   net47085 <= '0';
   net47086 <= '0';
   net47087 <= '0';
   net47088 <= '0';
   net47089 <= '0';
   net47090 <= '0';
   net47091 <= '0';
   net47092 <= '0';
   net47093 <= '0';
   net47094 <= '0';
   net47095 <= '0';
   net47096 <= '0';
   net47097 <= '0';
   net47098 <= '0';
   net47099 <= '0';
   net47100 <= '0';
   net47101 <= '0';
   net47102 <= '0';
   net47103 <= '0';
   net47104 <= '0';
   net47105 <= '0';
   net47106 <= '0';
   net47107 <= '0';
   net47108 <= '0';
   net47109 <= '0';
   net47110 <= '0';
   net47111 <= '0';
   net47112 <= '0';
   net47113 <= '0';
   net47114 <= '0';
   net47115 <= '0';
   net47116 <= '0';
   net47117 <= '0';
   net47118 <= '0';
   net47119 <= '0';
   net47120 <= '0';
   net47121 <= '0';
   net47122 <= '0';
   net47123 <= '0';
   net47124 <= '0';
   net47125 <= '0';
   net47126 <= '0';
   net47127 <= '0';
   net47128 <= '0';
   net47129 <= '0';
   net47130 <= '0';
   net47131 <= '0';
   net47132 <= '0';
   net47133 <= '0';
   net47134 <= '0';
   net47135 <= '0';
   net47136 <= '0';
   net47137 <= '0';
   net47138 <= '0';
   net47139 <= '0';
   net47140 <= '0';
   net47141 <= '0';
   net47142 <= '0';
   net47143 <= '0';
   net47144 <= '0';
   net47145 <= '0';
   net47146 <= '0';
   net47147 <= '0';
   net47148 <= '0';
   net47149 <= '0';
   net47150 <= '0';
   net47151 <= '0';
   net47152 <= '0';
   net47153 <= '0';
   net47154 <= '0';
   net47155 <= '0';
   net47156 <= '0';
   net47157 <= '0';
   net47158 <= '0';
   net47159 <= '0';
   net47160 <= '0';
   net47161 <= '0';
   net47162 <= '0';
   net47163 <= '0';
   net47164 <= '0';
   net47165 <= '0';
   net47166 <= '0';
   net47167 <= '0';
   net47168 <= '0';
   net47169 <= '0';
   net47170 <= '0';
   net47171 <= '0';
   net47172 <= '0';
   net47173 <= '0';
   net47174 <= '0';
   net47175 <= '0';
   net47176 <= '0';
   net47177 <= '0';
   net47178 <= '0';
   net47179 <= '0';
   net47180 <= '0';
   net47181 <= '0';
   net47182 <= '0';
   net47183 <= '0';
   net47184 <= '0';
   net47185 <= '0';
   net47186 <= '0';
   net47187 <= '0';
   net47188 <= '0';
   net47189 <= '0';
   net47190 <= '0';
   net47191 <= '0';
   net47192 <= '0';
   net47193 <= '0';
   net47194 <= '0';
   net47195 <= '0';
   net47196 <= '0';
   net47197 <= '0';
   net47198 <= '0';
   net47199 <= '0';
   net47200 <= '0';
   net47201 <= '0';
   net47202 <= '0';
   net47203 <= '0';
   net47204 <= '0';
   net47205 <= '0';
   net47206 <= '0';
   net47207 <= '0';
   net47208 <= '0';
   net47209 <= '0';
   net47210 <= '0';
   net47211 <= '0';
   net47212 <= '0';
   net47213 <= '0';
   net47214 <= '0';
   net47215 <= '0';
   net47216 <= '0';
   net47217 <= '0';
   net47218 <= '0';
   net47219 <= '0';
   net47220 <= '0';
   net47221 <= '0';
   net47222 <= '0';
   net47223 <= '0';
   net47224 <= '0';
   net47225 <= '0';
   net47226 <= '0';
   net47227 <= '0';
   net47228 <= '0';
   net47229 <= '0';
   net47230 <= '0';
   net47231 <= '0';
   net47232 <= '0';
   net47233 <= '0';
   net47234 <= '0';
   net47235 <= '0';
   net47236 <= '0';
   net47237 <= '0';
   net47238 <= '0';
   net47239 <= '0';
   net47240 <= '0';
   net47241 <= '0';
   net47242 <= '0';
   net47243 <= '0';
   net47244 <= '0';
   net47245 <= '0';
   net47246 <= '0';
   net47247 <= '0';
   net47248 <= '0';
   net47249 <= '0';
   net47250 <= '0';
   net47251 <= '0';
   net47252 <= '0';
   net47253 <= '0';
   net47254 <= '0';
   net47255 <= '0';
   net47256 <= '0';
   net47257 <= '0';
   net47258 <= '0';
   net47259 <= '0';
   net47260 <= '0';
   net47261 <= '0';
   net47262 <= '0';
   net47263 <= '0';
   net47264 <= '0';
   net47265 <= '0';
   net47266 <= '0';
   net47267 <= '0';
   net47268 <= '0';
   net47269 <= '0';
   net47270 <= '0';
   net47271 <= '0';
   net47272 <= '0';
   net47273 <= '0';
   net47274 <= '0';
   net47275 <= '0';
   net47276 <= '0';
   net47277 <= '0';
   net47278 <= '0';
   net47279 <= '0';
   net47280 <= '0';
   net47281 <= '0';
   net47282 <= '0';
   net47283 <= '0';
   net47284 <= '0';
   net47285 <= '0';
   net47286 <= '0';
   net47287 <= '0';
   net47288 <= '0';
   net47289 <= '0';
   net47290 <= '0';
   net47291 <= '0';
   net47292 <= '0';
   net47293 <= '0';
   net47294 <= '0';
   net47295 <= '0';
   net47296 <= '0';
   net47297 <= '0';
   net47298 <= '0';
   net47299 <= '0';
   net47300 <= '0';
   net47301 <= '0';
   net47302 <= '0';
   net47303 <= '0';
   net47304 <= '0';
   net47305 <= '0';
   net47306 <= '0';
   net47307 <= '0';
   net47308 <= '0';
   net47309 <= '0';
   net47310 <= '0';
   net47311 <= '0';
   net47312 <= '0';
   net47313 <= '0';
   net47314 <= '0';
   net47315 <= '0';
   net47316 <= '0';
   net47317 <= '0';
   net47318 <= '0';
   net47319 <= '0';
   net47320 <= '0';
   net47321 <= '0';
   net47322 <= '0';
   net47323 <= '0';
   net47324 <= '0';
   net47325 <= '0';
   net47326 <= '0';
   net47327 <= '0';
   net47328 <= '0';
   net47329 <= '0';
   net47330 <= '0';
   net47331 <= '0';
   net47332 <= '0';
   net47333 <= '0';
   net47334 <= '0';
   net47335 <= '0';
   net47336 <= '0';
   net47337 <= '0';
   net47338 <= '0';
   net47339 <= '0';
   net47340 <= '0';
   net47341 <= '0';
   net47342 <= '0';
   net47343 <= '0';
   net47344 <= '0';
   net47345 <= '0';
   net47346 <= '0';
   net47347 <= '0';
   net47348 <= '0';
   net47349 <= '0';
   net47350 <= '0';
   net47351 <= '0';
   net47352 <= '0';
   net47353 <= '0';
   net47354 <= '0';
   net47355 <= '0';
   net47356 <= '0';
   net47357 <= '0';
   net47358 <= '0';
   net47359 <= '0';
   net47360 <= '0';
   net47361 <= '0';
   net47362 <= '0';
   net47363 <= '0';
   net47364 <= '0';
   net47365 <= '0';
   net47366 <= '0';
   net47367 <= '0';
   net47368 <= '0';
   net47369 <= '0';
   net47370 <= '0';
   net47371 <= '0';
   net47372 <= '0';
   net47373 <= '0';
   net47374 <= '0';
   net47375 <= '0';
   net47376 <= '0';
   net47377 <= '0';
   net47378 <= '0';
   net47379 <= '0';
   net47380 <= '0';
   net47381 <= '0';
   net47382 <= '0';
   net47383 <= '0';
   net47384 <= '0';
   net47385 <= '0';
   net47386 <= '0';
   net47387 <= '0';
   net47388 <= '0';
   net47389 <= '0';
   net47390 <= '0';
   net47391 <= '0';
   net47392 <= '0';
   net47393 <= '0';
   net47394 <= '0';
   net47395 <= '0';
   net47396 <= '0';
   net47397 <= '0';
   net47398 <= '0';
   net47399 <= '0';
   net47400 <= '0';
   net47401 <= '0';
   net47402 <= '0';
   net47403 <= '0';
   net47404 <= '0';
   net47405 <= '0';
   net47406 <= '0';
   net47407 <= '0';
   net47408 <= '0';
   net47409 <= '0';
   net47410 <= '0';
   net47411 <= '0';
   net47412 <= '0';
   net47413 <= '0';
   net47414 <= '0';
   net47415 <= '0';
   net47416 <= '0';
   net47417 <= '0';
   net47418 <= '0';
   net47419 <= '0';
   net47420 <= '0';
   net47421 <= '0';
   net47422 <= '0';
   net47423 <= '0';
   net47424 <= '0';
   net47425 <= '0';
   net47426 <= '0';
   net47427 <= '0';
   net47428 <= '0';
   net47429 <= '0';
   net47430 <= '0';
   net47431 <= '0';
   net47432 <= '0';
   net47433 <= '0';
   net47434 <= '0';
   net47435 <= '0';
   net47436 <= '0';
   net47437 <= '0';
   net47438 <= '0';
   net47439 <= '0';
   net47440 <= '0';
   net47441 <= '0';
   net47442 <= '0';
   net47443 <= '0';
   net47444 <= '0';
   net47445 <= '0';
   net47446 <= '0';
   net47447 <= '0';
   net47448 <= '0';
   net47449 <= '0';
   net47450 <= '0';
   net47451 <= '0';
   net47452 <= '0';
   net47453 <= '0';
   net47454 <= '0';
   net47455 <= '0';
   net47456 <= '0';
   net47457 <= '0';
   net47458 <= '0';
   net47459 <= '0';
   net47460 <= '0';
   net47461 <= '0';
   net47462 <= '0';
   net47463 <= '0';
   net47464 <= '0';
   net47465 <= '0';
   net47466 <= '0';
   net47467 <= '0';
   net47468 <= '0';
   net47469 <= '0';
   net47470 <= '0';
   net47471 <= '0';
   net47472 <= '0';
   net47473 <= '0';
   net47474 <= '0';
   net47475 <= '0';
   net47476 <= '0';
   net47477 <= '0';
   net47478 <= '0';
   net47479 <= '0';
   net47480 <= '0';
   net47481 <= '0';
   net47482 <= '0';
   net47483 <= '0';
   net47484 <= '0';
   net47485 <= '0';
   net47486 <= '0';
   net47487 <= '0';
   net47488 <= '0';
   net47489 <= '0';
   net47490 <= '0';
   net47491 <= '0';
   net47492 <= '0';
   net47493 <= '0';
   net47494 <= '0';
   net47495 <= '0';
   net47496 <= '0';
   net47497 <= '0';
   net47498 <= '0';
   net47499 <= '0';
   net47500 <= '0';
   net47501 <= '0';
   net47502 <= '0';
   net47503 <= '0';
   net47504 <= '0';
   net47505 <= '0';
   net47506 <= '0';
   net47507 <= '0';
   net47508 <= '0';
   net47509 <= '0';
   net47510 <= '0';
   net47511 <= '0';
   net47512 <= '0';
   net47513 <= '0';
   net47514 <= '0';
   net47515 <= '0';
   net47516 <= '0';
   net47517 <= '0';
   net47518 <= '0';
   net47519 <= '0';
   net47520 <= '0';
   net47521 <= '0';
   net47522 <= '0';
   net47523 <= '0';
   net47524 <= '0';
   net47525 <= '0';
   net47526 <= '0';
   net47527 <= '0';
   net47528 <= '0';
   net47529 <= '0';
   net47530 <= '0';
   net47531 <= '0';
   net47532 <= '0';
   net47533 <= '0';
   net47534 <= '0';
   net47535 <= '0';
   net47536 <= '0';
   net47537 <= '0';
   net47538 <= '0';
   net47539 <= '0';
   net47540 <= '0';
   net47541 <= '0';
   net47542 <= '0';
   net47543 <= '0';
   net47544 <= '0';
   net47545 <= '0';
   net47546 <= '0';
   net47547 <= '0';
   net47548 <= '0';
   net47549 <= '0';
   net47550 <= '0';
   net47551 <= '0';
   net47552 <= '0';
   net47553 <= '0';
   net47554 <= '0';
   net47555 <= '0';
   net47556 <= '0';
   net47557 <= '0';
   net47558 <= '0';
   net47559 <= '0';
   net47560 <= '0';
   net47561 <= '0';
   net47562 <= '0';
   net47563 <= '0';
   net47564 <= '0';
   net47565 <= '0';
   net47566 <= '0';
   net47567 <= '0';
   net47568 <= '0';
   net47569 <= '0';
   net47570 <= '0';
   net47571 <= '0';
   net47572 <= '0';
   net47573 <= '0';
   net47574 <= '0';
   net47575 <= '0';
   net47576 <= '0';
   net47577 <= '0';
   net47578 <= '0';
   net47579 <= '0';
   net47580 <= '0';
   net47581 <= '0';
   net47582 <= '0';
   net47583 <= '0';
   net47584 <= '0';
   net47585 <= '0';
   net47586 <= '0';
   net47587 <= '0';
   net47588 <= '0';
   net47589 <= '0';
   net47590 <= '0';
   net47591 <= '0';
   net47592 <= '0';
   net47593 <= '0';
   net47594 <= '0';
   net47595 <= '0';
   net47596 <= '0';
   net47597 <= '0';
   net47598 <= '0';
   net47599 <= '0';
   net47600 <= '0';
   net47601 <= '0';
   net47602 <= '0';
   net47603 <= '0';
   net47604 <= '0';
   net47605 <= '0';
   net47606 <= '0';
   net47607 <= '0';
   net47608 <= '0';
   net47609 <= '0';
   net47610 <= '0';
   net47611 <= '0';
   net47612 <= '0';
   net47613 <= '0';
   net47614 <= '0';
   net47615 <= '0';
   net47616 <= '0';
   net47617 <= '0';
   net47618 <= '0';
   net47619 <= '0';
   net47620 <= '0';
   net47621 <= '0';
   net47622 <= '0';
   net47623 <= '0';
   net47624 <= '0';
   net47625 <= '0';
   net47626 <= '0';
   net47627 <= '0';
   net47628 <= '0';
   net47629 <= '0';
   net47630 <= '0';
   net47631 <= '0';
   net47632 <= '0';
   net47633 <= '0';
   net47634 <= '0';
   net47635 <= '0';
   net47636 <= '0';
   net47637 <= '0';
   net47638 <= '0';
   net47639 <= '0';
   net47640 <= '0';
   net47641 <= '0';
   net47642 <= '0';
   net47643 <= '0';
   net47644 <= '0';
   net47645 <= '0';
   net47646 <= '0';
   net47647 <= '0';
   net47648 <= '0';
   net47649 <= '0';
   net47650 <= '0';
   net47651 <= '0';
   net47652 <= '0';
   net47653 <= '0';
   net47654 <= '0';
   net47655 <= '0';
   net47656 <= '0';
   net47657 <= '0';
   net47658 <= '0';
   net47659 <= '0';
   net47660 <= '0';
   net47661 <= '0';
   net47662 <= '0';
   net47663 <= '0';
   net47664 <= '0';
   net47665 <= '0';
   net47666 <= '0';
   net47667 <= '0';
   net47668 <= '0';
   net47669 <= '0';
   net47670 <= '0';
   net47671 <= '0';
   net47672 <= '0';
   net47673 <= '0';
   net47674 <= '0';
   net47675 <= '0';
   net47676 <= '0';
   net47677 <= '0';
   net47678 <= '0';
   net47679 <= '0';
   net47680 <= '0';
   net47681 <= '0';
   net47682 <= '0';
   net47683 <= '0';
   net47684 <= '0';
   net47685 <= '0';
   net47686 <= '0';
   net47687 <= '0';
   net47688 <= '0';
   net47689 <= '0';
   net47690 <= '0';
   net47691 <= '0';
   net47692 <= '0';
   net47693 <= '0';
   net47694 <= '0';
   net47695 <= '0';
   net47696 <= '0';
   net47697 <= '0';
   net47698 <= '0';
   net47699 <= '0';
   net47700 <= '0';
   net47701 <= '0';
   net47702 <= '0';
   net47703 <= '0';
   net47704 <= '0';
   net47705 <= '0';
   net47706 <= '0';
   net47707 <= '0';
   net47708 <= '0';
   net47709 <= '0';
   net47710 <= '0';
   net47711 <= '0';
   net47712 <= '0';
   net47713 <= '0';
   net47714 <= '0';
   net47715 <= '0';
   net47716 <= '0';
   net47717 <= '0';
   net47718 <= '0';
   net47719 <= '0';
   net47720 <= '0';
   net47721 <= '0';
   net47722 <= '0';
   net47723 <= '0';
   net47724 <= '0';
   net47725 <= '0';
   net47726 <= '0';
   net47727 <= '0';
   net47728 <= '0';
   net47729 <= '0';
   net47730 <= '0';
   net47731 <= '0';
   net47732 <= '0';
   net47733 <= '0';
   net47734 <= '0';
   net47735 <= '0';
   net47736 <= '0';
   net47737 <= '0';
   net47738 <= '0';
   net47739 <= '0';
   net47740 <= '0';
   net47741 <= '0';
   net47742 <= '0';
   net47743 <= '0';
   net47744 <= '0';
   net47745 <= '0';
   net47746 <= '0';
   net47747 <= '0';
   net47748 <= '0';
   net47749 <= '0';
   net47750 <= '0';
   net47751 <= '0';
   net47752 <= '0';
   net47753 <= '0';
   net47754 <= '0';
   net47755 <= '0';
   net47756 <= '0';
   net47757 <= '0';
   net47758 <= '0';
   net47759 <= '0';
   net47760 <= '0';
   net47761 <= '0';
   net47762 <= '0';
   net47763 <= '0';
   net47764 <= '0';
   net47765 <= '0';
   net47766 <= '0';
   net47767 <= '0';
   net47768 <= '0';
   net47769 <= '0';
   net47770 <= '0';
   net47771 <= '0';
   net47772 <= '0';
   net47773 <= '0';
   net47774 <= '0';
   net47775 <= '0';
   net47776 <= '0';
   net47777 <= '0';
   net47778 <= '0';
   net47779 <= '0';
   net47780 <= '0';
   net47781 <= '0';
   net47782 <= '0';
   net47783 <= '0';
   net47784 <= '0';
   net47785 <= '0';
   net47786 <= '0';
   net47787 <= '0';
   net47788 <= '0';
   net47789 <= '0';
   net47790 <= '0';
   net47791 <= '0';
   net47792 <= '0';
   net47793 <= '0';
   net47794 <= '0';
   net47795 <= '0';
   net47796 <= '0';
   net47797 <= '0';
   net47798 <= '0';
   net47799 <= '0';
   net47800 <= '0';
   net47801 <= '0';
   net47802 <= '0';
   net47803 <= '0';
   net47804 <= '0';
   net47805 <= '0';
   net47806 <= '0';
   net47807 <= '0';
   net47808 <= '0';
   net47809 <= '0';
   net47810 <= '0';
   net47811 <= '0';
   net47812 <= '0';
   net47813 <= '0';
   net47814 <= '0';
   net47815 <= '0';
   net47816 <= '0';
   net47817 <= '0';
   net47818 <= '0';
   net47819 <= '0';
   net47820 <= '0';
   net47821 <= '0';
   net47822 <= '0';
   net47823 <= '0';
   net47824 <= '0';
   net47825 <= '0';
   net47826 <= '0';
   net47827 <= '0';
   net47828 <= '0';
   net47829 <= '0';
   net47830 <= '0';
   net47831 <= '0';
   net47832 <= '0';
   net47833 <= '0';
   net47834 <= '0';
   net47835 <= '0';
   net47836 <= '0';
   net47837 <= '0';
   net47838 <= '0';
   net47839 <= '0';
   net47840 <= '0';
   net47841 <= '0';
   net47842 <= '0';
   net47843 <= '0';
   net47844 <= '0';
   net47845 <= '0';
   net47846 <= '0';
   net47847 <= '0';
   net47848 <= '0';
   net47849 <= '0';
   net47850 <= '0';
   net47851 <= '0';
   net47852 <= '0';
   net47853 <= '0';
   net47854 <= '0';
   net47855 <= '0';
   net47856 <= '0';
   net47857 <= '0';
   net47858 <= '0';
   net47859 <= '0';
   net47860 <= '0';
   net47861 <= '0';
   net47862 <= '0';
   net47863 <= '0';
   net47864 <= '0';
   net47865 <= '0';
   net47866 <= '0';
   net47867 <= '0';
   net47868 <= '0';
   net47869 <= '0';
   net47870 <= '0';
   net47871 <= '0';
   net47872 <= '0';
   net47873 <= '0';
   net47874 <= '0';
   net47875 <= '0';
   net47876 <= '0';
   net47877 <= '0';
   net47878 <= '0';
   net47879 <= '0';
   net47880 <= '0';
   net47881 <= '0';
   net47882 <= '0';
   net47883 <= '0';
   net47884 <= '0';
   net47885 <= '0';
   net47886 <= '0';
   net47887 <= '0';
   net47888 <= '0';
   net47889 <= '0';
   net47890 <= '0';
   net47891 <= '0';
   net47892 <= '0';
   net47893 <= '0';
   net47894 <= '0';
   net47895 <= '0';
   net47896 <= '0';
   net47897 <= '0';
   net47898 <= '0';
   net47899 <= '0';
   net47900 <= '0';
   net47901 <= '0';
   net47902 <= '0';
   net47903 <= '0';
   net47904 <= '0';
   net47905 <= '0';
   net47906 <= '0';
   net47907 <= '0';
   net47908 <= '0';
   net47909 <= '0';
   net47910 <= '0';
   net47911 <= '0';
   net47912 <= '0';
   net47913 <= '0';
   net47914 <= '0';
   net47915 <= '0';
   net47916 <= '0';
   net47917 <= '0';
   net47918 <= '0';
   net47919 <= '0';
   net47920 <= '0';
   net47921 <= '0';
   net47922 <= '0';
   net47923 <= '0';
   net47924 <= '0';
   net47925 <= '0';
   net47926 <= '0';
   net47927 <= '0';
   net47928 <= '0';
   net47929 <= '0';
   net47930 <= '0';
   net47931 <= '0';
   net47932 <= '0';
   net47933 <= '0';
   net47934 <= '0';
   net47935 <= '0';
   net47936 <= '0';
   net47937 <= '0';
   net47938 <= '0';
   net47939 <= '0';
   net47940 <= '0';
   net47941 <= '0';
   net47942 <= '0';
   net47943 <= '0';
   net47944 <= '0';
   net47945 <= '0';
   net47946 <= '0';
   net47947 <= '0';
   net47948 <= '0';
   net47949 <= '0';
   net47950 <= '0';
   net47951 <= '0';
   net47952 <= '0';
   net47953 <= '0';
   net47954 <= '0';
   net47955 <= '0';
   net47956 <= '0';
   net47957 <= '0';
   net47958 <= '0';
   net47959 <= '0';
   net47960 <= '0';
   net47961 <= '0';
   net47962 <= '0';
   net47963 <= '0';
   net47964 <= '0';
   net47965 <= '0';
   net47966 <= '0';
   net47967 <= '0';
   net47968 <= '0';
   net47969 <= '0';
   net47970 <= '0';
   net47971 <= '0';
   net47972 <= '0';
   net47973 <= '0';
   net47974 <= '0';
   net47975 <= '0';
   net47976 <= '0';
   net47977 <= '0';
   net47978 <= '0';
   net47979 <= '0';
   net47980 <= '0';
   net47981 <= '0';
   net47982 <= '0';
   net47983 <= '0';
   net47984 <= '0';
   net47985 <= '0';
   net47986 <= '0';
   net47987 <= '0';
   net47988 <= '0';
   net47989 <= '0';
   net47990 <= '0';
   net47991 <= '0';
   net47992 <= '0';
   net47993 <= '0';
   net47994 <= '0';
   net47995 <= '0';
   net47996 <= '0';
   net47997 <= '0';
   net47998 <= '0';
   net47999 <= '0';
   net48000 <= '0';
   net48001 <= '0';
   net48002 <= '0';
   net48003 <= '0';
   net48004 <= '0';
   net48005 <= '0';
   net48006 <= '0';
   net48007 <= '0';
   net48008 <= '0';
   net48009 <= '0';
   net48010 <= '0';
   net48011 <= '0';
   net48012 <= '0';
   net48013 <= '0';
   net48014 <= '0';
   net48015 <= '0';
   net48016 <= '0';
   net48017 <= '0';
   net48018 <= '0';
   net48019 <= '0';
   net48020 <= '0';
   net48021 <= '0';
   net48022 <= '0';
   net48023 <= '0';
   net48024 <= '0';
   net48025 <= '0';
   net48026 <= '0';
   net48027 <= '0';
   net48028 <= '0';
   net48029 <= '0';
   net48030 <= '0';
   net48031 <= '0';
   net48032 <= '0';
   net48033 <= '0';
   net48034 <= '0';
   net48035 <= '0';
   net48036 <= '0';
   net48037 <= '0';
   net48038 <= '0';
   net48039 <= '0';
   net48040 <= '0';
   net48041 <= '0';
   net48042 <= '0';
   net48043 <= '0';
   net48044 <= '0';
   net48045 <= '0';
   net48046 <= '0';
   net48047 <= '0';
   net48048 <= '0';
   net48049 <= '0';
   net48050 <= '0';
   net48051 <= '0';
   net48052 <= '0';
   net48053 <= '0';
   net48054 <= '0';
   net48055 <= '0';
   net48056 <= '0';
   net48057 <= '0';
   net48058 <= '0';
   net48059 <= '0';
   net48060 <= '0';
   net48061 <= '0';
   net48062 <= '0';
   net48063 <= '0';
   net48064 <= '0';
   net48065 <= '0';
   net48066 <= '0';
   net48067 <= '0';
   net48068 <= '0';
   net48069 <= '0';
   net48070 <= '0';
   net48071 <= '0';
   net48072 <= '0';
   net48073 <= '0';
   net48074 <= '0';
   net48075 <= '0';
   net48076 <= '0';
   net48077 <= '0';
   net48078 <= '0';
   net48079 <= '0';
   net48080 <= '0';
   net48081 <= '0';
   net48082 <= '0';
   net48083 <= '0';
   net48084 <= '0';
   net48085 <= '0';
   net48086 <= '0';
   net48087 <= '0';
   net48088 <= '0';
   net48089 <= '0';
   net48090 <= '0';
   net48091 <= '0';
   net48092 <= '0';
   net48093 <= '0';
   net48094 <= '0';
   net48095 <= '0';
   net48096 <= '0';
   net48097 <= '0';
   net48098 <= '0';
   net48099 <= '0';
   net48100 <= '0';
   net48101 <= '0';
   net48102 <= '0';
   net48103 <= '0';
   net48104 <= '0';
   net48105 <= '0';
   net48106 <= '0';
   net48107 <= '0';
   net48108 <= '0';
   net48109 <= '0';
   net48110 <= '0';
   net48111 <= '0';
   net48112 <= '0';
   net48113 <= '0';
   net48114 <= '0';
   net48115 <= '0';
   net48116 <= '0';
   net48117 <= '0';
   net48118 <= '0';
   net48119 <= '0';
   net48120 <= '0';
   net48121 <= '0';
   net48122 <= '0';
   net48123 <= '0';
   net48124 <= '0';
   net48125 <= '0';
   net48126 <= '0';
   net48127 <= '0';
   net48128 <= '0';
   net48129 <= '0';
   net48130 <= '0';
   net48131 <= '0';
   net48132 <= '0';
   net48133 <= '0';
   net48134 <= '0';
   net48135 <= '0';
   net48136 <= '0';
   net48137 <= '0';
   net48138 <= '0';
   net48139 <= '0';
   net48140 <= '0';
   net48141 <= '0';
   net48142 <= '0';
   net48143 <= '0';
   net48144 <= '0';
   net48145 <= '0';
   net48146 <= '0';
   net48147 <= '0';
   net48148 <= '0';
   net48149 <= '0';
   net48150 <= '0';
   net48151 <= '0';
   net48152 <= '0';
   net48153 <= '0';
   net48154 <= '0';
   net48155 <= '0';
   net48156 <= '0';
   net48157 <= '0';
   net48158 <= '0';
   net48159 <= '0';
   net48160 <= '0';
   net48161 <= '0';
   net48162 <= '0';
   net48163 <= '0';
   net48164 <= '0';
   net48165 <= '0';
   net48166 <= '0';
   net48167 <= '0';
   net48168 <= '0';
   net48169 <= '0';
   net48170 <= '0';
   net48171 <= '0';
   net48172 <= '0';
   net48173 <= '0';
   net48174 <= '0';
   net48175 <= '0';
   net48176 <= '0';
   net48177 <= '0';
   net48178 <= '0';
   net48179 <= '0';
   net48180 <= '0';
   net48181 <= '0';
   net48182 <= '0';
   net48183 <= '0';
   net48184 <= '0';
   net48185 <= '0';
   net48186 <= '0';
   net48187 <= '0';
   net48188 <= '0';
   net48189 <= '0';
   net48190 <= '0';
   net48191 <= '0';
   net48192 <= '0';
   net48193 <= '0';
   net48194 <= '0';
   net48195 <= '0';
   net48196 <= '0';
   net48197 <= '0';
   net48198 <= '0';
   net48199 <= '0';
   net48200 <= '0';
   net48201 <= '0';
   net48202 <= '0';
   net48203 <= '0';
   net48204 <= '0';
   net48205 <= '0';
   net48206 <= '0';
   net48207 <= '0';
   net48208 <= '0';
   net48209 <= '0';
   net48210 <= '0';
   net48211 <= '0';
   net48212 <= '0';
   net48213 <= '0';
   net48214 <= '0';
   net48215 <= '0';
   net48216 <= '0';
   net48217 <= '0';
   net48218 <= '0';
   net48219 <= '0';
   net48220 <= '0';
   net48221 <= '0';
   net48222 <= '0';
   net48223 <= '0';
   net48224 <= '0';
   net48225 <= '0';
   net48226 <= '0';
   net48227 <= '0';
   net48228 <= '0';
   net48229 <= '0';
   net48230 <= '0';
   net48231 <= '0';
   net48232 <= '0';
   net48233 <= '0';
   net48234 <= '0';
   net48235 <= '0';
   net48236 <= '0';
   net48237 <= '0';
   net48238 <= '0';
   net48239 <= '0';
   net48240 <= '0';
   net48241 <= '0';
   net48242 <= '0';
   net48243 <= '0';
   net48244 <= '0';
   net48245 <= '0';
   net48246 <= '0';
   net48247 <= '0';
   net48248 <= '0';
   net48249 <= '0';
   net48250 <= '0';
   net48251 <= '0';
   net48252 <= '0';
   net48253 <= '0';
   net48254 <= '0';
   net48255 <= '0';
   net48256 <= '0';
   net48257 <= '0';
   net48258 <= '0';
   net48259 <= '0';
   net48260 <= '0';
   net48261 <= '0';
   net48262 <= '0';
   net48263 <= '0';
   net48264 <= '0';
   net48265 <= '0';
   net48266 <= '0';
   net48267 <= '0';
   net48268 <= '0';
   net48269 <= '0';
   net48270 <= '0';
   net48271 <= '0';
   net48272 <= '0';
   net48273 <= '0';
   net48274 <= '0';
   net48275 <= '0';
   net48276 <= '0';
   net48277 <= '0';
   net48278 <= '0';
   net48279 <= '0';
   net48280 <= '0';
   net48281 <= '0';
   net48282 <= '0';
   net48283 <= '0';
   net48284 <= '0';
   net48285 <= '0';
   net48286 <= '0';
   net48287 <= '0';
   net48288 <= '0';
   net48289 <= '0';
   net48290 <= '0';
   net48291 <= '0';
   net48292 <= '0';
   net48293 <= '0';
   net48294 <= '0';
   net48295 <= '0';
   net48296 <= '0';
   net48297 <= '0';
   net48298 <= '0';
   net48299 <= '0';
   net48300 <= '0';
   net48301 <= '0';
   net48302 <= '0';
   net48303 <= '0';
   net48304 <= '0';
   net48305 <= '0';
   net48306 <= '0';
   net48307 <= '0';
   net48308 <= '0';
   net48309 <= '0';
   net48310 <= '0';
   net48311 <= '0';
   net48312 <= '0';
   net48313 <= '0';
   net48314 <= '0';
   net48315 <= '0';
   net48316 <= '0';
   net48317 <= '0';
   net48318 <= '0';
   net48319 <= '0';
   net48320 <= '0';
   net48321 <= '0';
   net48322 <= '0';
   net48323 <= '0';
   net48324 <= '0';
   net48325 <= '0';
   net48326 <= '0';
   net48327 <= '0';
   net48328 <= '0';
   net48329 <= '0';
   net48330 <= '0';
   net48331 <= '0';
   net48332 <= '0';
   net48333 <= '0';
   net48334 <= '0';
   net48335 <= '0';
   net48336 <= '0';
   net48337 <= '0';
   net48338 <= '0';
   net48339 <= '0';
   net48340 <= '0';
   net48341 <= '0';
   net48342 <= '0';
   net48343 <= '0';
   net48344 <= '0';
   net48345 <= '0';
   net48346 <= '0';
   net48347 <= '0';
   net48348 <= '0';
   net48349 <= '0';
   net48350 <= '0';
   net48351 <= '0';
   net48352 <= '0';
   net48353 <= '0';
   net48354 <= '0';
   net48355 <= '0';
   net48356 <= '0';
   net48357 <= '0';
   net48358 <= '0';
   net48359 <= '0';
   net48360 <= '0';
   net48361 <= '0';
   net48362 <= '0';
   net48363 <= '0';
   net48364 <= '0';
   net48365 <= '0';
   net48366 <= '0';
   net48367 <= '0';
   net48368 <= '0';
   net48369 <= '0';
   net48370 <= '0';
   net48371 <= '0';
   net48372 <= '0';
   net48373 <= '0';
   net48374 <= '0';
   net48375 <= '0';
   net48376 <= '0';
   net48377 <= '0';
   net48378 <= '0';
   net48379 <= '0';
   net48380 <= '0';
   net48381 <= '0';
   net48382 <= '0';
   net48383 <= '0';
   net48384 <= '0';
   net48385 <= '0';
   net48386 <= '0';
   net48387 <= '0';
   net48388 <= '0';
   net48389 <= '0';
   net48390 <= '0';
   net48391 <= '0';
   net48392 <= '0';
   net48393 <= '0';
   net48394 <= '0';
   net48395 <= '0';
   net48396 <= '0';
   net48397 <= '0';
   net48398 <= '0';
   net48399 <= '0';
   net48400 <= '0';
   net48401 <= '0';
   net48402 <= '0';
   net48403 <= '0';
   net48404 <= '0';
   net48405 <= '0';
   net48406 <= '0';
   net48407 <= '0';
   net48408 <= '0';
   net48409 <= '0';
   net48410 <= '0';
   net48411 <= '0';
   net48412 <= '0';
   net48413 <= '0';
   net48414 <= '0';
   net48415 <= '0';
   net48416 <= '0';
   net48417 <= '0';
   net48418 <= '0';
   net48419 <= '0';
   net48420 <= '0';
   net48421 <= '0';
   net48422 <= '0';
   net48423 <= '0';
   net48424 <= '0';
   net48425 <= '0';
   net48426 <= '0';
   net48427 <= '0';
   net48428 <= '0';
   net48429 <= '0';
   net48430 <= '0';
   net48431 <= '0';
   net48432 <= '0';
   net48433 <= '0';
   net48434 <= '0';
   net48435 <= '0';
   net48436 <= '0';
   net48437 <= '0';
   net48438 <= '0';
   net48439 <= '0';
   net48440 <= '0';
   net48441 <= '0';
   net48442 <= '0';
   net48443 <= '0';
   net48444 <= '0';
   net48445 <= '0';
   net48446 <= '0';
   net48447 <= '0';
   net48448 <= '0';
   net48449 <= '0';
   net48450 <= '0';
   net48451 <= '0';
   net48452 <= '0';
   net48453 <= '0';
   net48454 <= '0';
   net48455 <= '0';
   net48456 <= '0';
   net48457 <= '0';
   net48458 <= '0';
   net48459 <= '0';
   net48460 <= '0';
   net48461 <= '0';
   net48462 <= '0';
   net48463 <= '0';
   net48464 <= '0';
   net48465 <= '0';
   net48466 <= '0';
   net48467 <= '0';
   net48468 <= '0';
   net48469 <= '0';
   net48470 <= '0';
   net48471 <= '0';
   net48472 <= '0';
   net48473 <= '0';
   net48474 <= '0';
   net48475 <= '0';
   net48476 <= '0';
   net48477 <= '0';
   net48478 <= '0';
   net48479 <= '0';
   net48480 <= '0';
   net48481 <= '0';
   net48482 <= '0';
   net48483 <= '0';
   net48484 <= '0';
   net48485 <= '0';
   net48486 <= '0';
   net48487 <= '0';
   net48488 <= '0';
   net48489 <= '0';
   net48490 <= '0';
   net48491 <= '0';
   net48492 <= '0';
   net48493 <= '0';
   net48494 <= '0';
   net48495 <= '0';
   net48496 <= '0';
   net48497 <= '0';
   net48498 <= '0';
   net48499 <= '0';
   net48500 <= '0';
   net48501 <= '0';
   net48502 <= '0';
   net48503 <= '0';
   net48504 <= '0';
   net48505 <= '0';
   net48506 <= '0';
   net48507 <= '0';
   net48508 <= '0';
   net48509 <= '0';
   net48510 <= '0';
   net48511 <= '0';
   net48512 <= '0';
   net48513 <= '0';
   net48514 <= '0';
   net48515 <= '0';
   net48516 <= '0';
   net48517 <= '0';
   net48518 <= '0';
   net48519 <= '0';
   net48520 <= '0';
   net48521 <= '0';
   net48522 <= '0';
   net48523 <= '0';
   net48524 <= '0';
   net48525 <= '0';
   net48526 <= '0';
   net48527 <= '0';
   net48528 <= '0';
   net48529 <= '0';
   net48530 <= '0';
   net48531 <= '0';
   net48532 <= '0';
   net48533 <= '0';
   net48534 <= '0';
   net48535 <= '0';
   net48536 <= '0';
   net48537 <= '0';
   net48538 <= '0';
   net48539 <= '0';
   net48540 <= '0';
   net48541 <= '0';
   net48542 <= '0';
   net48543 <= '0';
   net48544 <= '0';
   net48545 <= '0';
   net48546 <= '0';
   net48547 <= '0';
   net48548 <= '0';
   net48549 <= '0';
   net48550 <= '0';
   net48551 <= '0';
   net48552 <= '0';
   net48553 <= '0';
   net48554 <= '0';
   net48555 <= '0';
   net48556 <= '0';
   net48557 <= '0';
   net48558 <= '0';
   net48559 <= '0';
   net48560 <= '0';
   net48561 <= '0';
   net48562 <= '0';
   net48563 <= '0';
   net48564 <= '0';
   net48565 <= '0';
   net48566 <= '0';
   net48567 <= '0';
   net48568 <= '0';
   net48569 <= '0';
   net48570 <= '0';
   net48571 <= '0';
   net48572 <= '0';
   net48573 <= '0';
   net48574 <= '0';
   net48575 <= '0';
   net48576 <= '0';
   net48577 <= '0';
   net48578 <= '0';
   net48579 <= '0';
   net48580 <= '0';
   net48581 <= '0';
   net48582 <= '0';
   net48583 <= '0';
   net48584 <= '0';
   net48585 <= '0';
   net48586 <= '0';
   net48587 <= '0';
   net48588 <= '0';
   net48589 <= '0';
   net48590 <= '0';
   net48591 <= '0';
   net48592 <= '0';
   net48593 <= '0';
   net48594 <= '0';
   net48595 <= '0';
   net48596 <= '0';
   net48597 <= '0';
   net48598 <= '0';
   net48599 <= '0';
   net48600 <= '0';
   net48601 <= '0';
   net48602 <= '0';
   net48603 <= '0';
   net48604 <= '0';
   net48605 <= '0';
   net48606 <= '0';
   net48607 <= '0';
   net48608 <= '0';
   net48609 <= '0';
   net48610 <= '0';
   net48611 <= '0';
   net48612 <= '0';
   net48613 <= '0';
   net48614 <= '0';
   net48615 <= '0';
   net48616 <= '0';
   net48617 <= '0';
   net48618 <= '0';
   net48619 <= '0';
   net48620 <= '0';
   net48621 <= '0';
   net48622 <= '0';
   net48623 <= '0';
   net48624 <= '0';
   net48625 <= '0';
   net48626 <= '0';
   net48627 <= '0';
   net48628 <= '0';
   net48629 <= '0';
   net48630 <= '0';
   net48631 <= '0';
   net48632 <= '0';
   net48633 <= '0';
   net48634 <= '0';
   net48635 <= '0';
   net48636 <= '0';
   net48637 <= '0';
   net48638 <= '0';
   net48639 <= '0';
   net48640 <= '0';
   net48641 <= '0';
   net48642 <= '0';
   net48643 <= '0';
   net48644 <= '0';
   net48645 <= '0';
   net48646 <= '0';
   net48647 <= '0';
   net48648 <= '0';
   net48649 <= '0';
   net48650 <= '0';
   net48651 <= '0';
   net48652 <= '0';
   net48653 <= '0';
   net48654 <= '0';
   net48655 <= '0';
   net48656 <= '0';
   net48657 <= '0';
   net48658 <= '0';
   net48659 <= '0';
   net48660 <= '0';
   net48661 <= '0';
   net48662 <= '0';
   net48663 <= '0';
   net48664 <= '0';
   net48665 <= '0';
   net48666 <= '0';
   net48667 <= '0';
   net48668 <= '0';
   net48669 <= '0';
   net48670 <= '0';
   net48671 <= '0';
   net48672 <= '0';
   net48673 <= '0';
   net48674 <= '0';
   net48675 <= '0';
   net48676 <= '0';
   net48677 <= '0';
   net48678 <= '0';
   net48679 <= '0';
   net48680 <= '0';
   net48681 <= '0';
   net48682 <= '0';
   net48683 <= '0';
   net48684 <= '0';
   net48685 <= '0';
   net48686 <= '0';
   net48687 <= '0';
   net48688 <= '0';
   net48689 <= '0';
   net48690 <= '0';
   net48691 <= '0';
   net48692 <= '0';
   net48693 <= '0';
   net48694 <= '0';
   net48695 <= '0';
   net48696 <= '0';
   net48697 <= '0';
   net48698 <= '0';
   net48699 <= '0';
   net48700 <= '0';
   net48701 <= '0';
   net48702 <= '0';
   net48703 <= '0';
   net48704 <= '0';
   net48705 <= '0';
   net48706 <= '0';
   net48707 <= '0';
   net48708 <= '0';
   net48709 <= '0';
   net48710 <= '0';
   net48711 <= '0';
   net48712 <= '0';
   net48713 <= '0';
   net48714 <= '0';
   net48715 <= '0';
   net48716 <= '0';
   net48717 <= '0';
   net48718 <= '0';
   net48719 <= '0';
   net48720 <= '0';
   net48721 <= '0';
   net48722 <= '0';
   net48723 <= '0';
   net48724 <= '0';
   net48725 <= '0';
   net48726 <= '0';
   net48727 <= '0';
   net48728 <= '0';
   net48729 <= '0';
   net48730 <= '0';
   net48731 <= '0';
   net48732 <= '0';
   net48733 <= '0';
   net48734 <= '0';
   net48735 <= '0';
   net48736 <= '0';
   net48737 <= '0';
   net48738 <= '0';
   net48739 <= '0';
   net48740 <= '0';
   net48741 <= '0';
   net48742 <= '0';
   net48743 <= '0';
   net48744 <= '0';
   net48745 <= '0';
   net48746 <= '0';
   net48747 <= '0';
   net48748 <= '0';
   net48749 <= '0';
   net48750 <= '0';
   net48751 <= '0';
   net48752 <= '0';
   net48753 <= '0';
   net48754 <= '0';
   net48755 <= '0';
   net48756 <= '0';
   net48757 <= '0';
   net48758 <= '0';
   net48759 <= '0';
   net48760 <= '0';
   net48761 <= '0';
   net48762 <= '0';
   net48763 <= '0';
   net48764 <= '0';
   net48765 <= '0';
   net48766 <= '0';
   net48767 <= '0';
   net48768 <= '0';
   net48769 <= '0';
   net48770 <= '0';
   net48771 <= '0';
   net48772 <= '0';
   net48773 <= '0';
   net48774 <= '0';
   net48775 <= '0';
   net48776 <= '0';
   net48777 <= '0';
   net48778 <= '0';
   net48779 <= '0';
   net48780 <= '0';
   net48781 <= '0';
   net48782 <= '0';
   net48783 <= '0';
   net48784 <= '0';
   net48785 <= '0';
   net48786 <= '0';
   net48787 <= '0';
   net48788 <= '0';
   net48789 <= '0';
   net48790 <= '0';
   net48791 <= '0';
   net48792 <= '0';
   net48793 <= '0';
   net48794 <= '0';
   net48795 <= '0';
   net48796 <= '0';
   net48797 <= '0';
   net48798 <= '0';
   net48799 <= '0';
   net48800 <= '0';
   net48801 <= '0';
   net48802 <= '0';
   net48803 <= '0';
   net48804 <= '0';
   net48805 <= '0';
   net48806 <= '0';
   net48807 <= '0';
   net48808 <= '0';
   net48809 <= '0';
   net48810 <= '0';
   net48811 <= '0';
   net48812 <= '0';
   net48813 <= '0';
   net48814 <= '0';
   net48815 <= '0';
   net48816 <= '0';
   net48817 <= '0';
   net48818 <= '0';
   net48819 <= '0';
   OTMP_960_port <= '0';
   SHIFT_n_960_port <= '0';
   SHIFT_n_961_port <= '0';
   SHIFT_960_port <= '0';
   SHIFT_961_port <= '0';
   OTMP_896_port <= '0';
   SHIFT_n_896_port <= '0';
   SHIFT_n_897_port <= '0';
   SHIFT_896_port <= '0';
   SHIFT_897_port <= '0';
   OTMP_832_port <= '0';
   SHIFT_n_832_port <= '0';
   SHIFT_n_833_port <= '0';
   SHIFT_832_port <= '0';
   SHIFT_833_port <= '0';
   OTMP_768_port <= '0';
   SHIFT_n_768_port <= '0';
   SHIFT_n_769_port <= '0';
   SHIFT_768_port <= '0';
   SHIFT_769_port <= '0';
   OTMP_704_port <= '0';
   SHIFT_n_704_port <= '0';
   SHIFT_n_705_port <= '0';
   SHIFT_704_port <= '0';
   SHIFT_705_port <= '0';
   OTMP_640_port <= '0';
   SHIFT_n_640_port <= '0';
   SHIFT_n_641_port <= '0';
   SHIFT_640_port <= '0';
   SHIFT_641_port <= '0';
   OTMP_576_port <= '0';
   SHIFT_n_576_port <= '0';
   SHIFT_n_577_port <= '0';
   SHIFT_576_port <= '0';
   SHIFT_577_port <= '0';
   OTMP_512_port <= '0';
   SHIFT_n_512_port <= '0';
   SHIFT_n_513_port <= '0';
   SHIFT_512_port <= '0';
   SHIFT_513_port <= '0';
   OTMP_448_port <= '0';
   SHIFT_n_448_port <= '0';
   SHIFT_n_449_port <= '0';
   SHIFT_448_port <= '0';
   SHIFT_449_port <= '0';
   OTMP_384_port <= '0';
   SHIFT_n_384_port <= '0';
   SHIFT_n_385_port <= '0';
   SHIFT_384_port <= '0';
   SHIFT_385_port <= '0';
   OTMP_320_port <= '0';
   SHIFT_n_320_port <= '0';
   SHIFT_n_321_port <= '0';
   SHIFT_320_port <= '0';
   SHIFT_321_port <= '0';
   OTMP_256_port <= '0';
   SHIFT_n_256_port <= '0';
   SHIFT_n_257_port <= '0';
   SHIFT_256_port <= '0';
   SHIFT_257_port <= '0';
   OTMP_192_port <= '0';
   SHIFT_n_192_port <= '0';
   SHIFT_n_193_port <= '0';
   SHIFT_192_port <= '0';
   SHIFT_193_port <= '0';
   OTMP_128_port <= '0';
   SHIFT_n_128_port <= '0';
   SHIFT_n_129_port <= '0';
   SHIFT_128_port <= '0';
   SHIFT_129_port <= '0';
   OTMP_64_port <= '0';
   SHIFT_n_64_port <= '0';
   SHIFT_64_port <= '0';
   n4 <= '0';
   n5 <= '0';
   BOOTHENC_I_1 : BOOTHENC_NBIT64_i0 port map( A(63) => net48692, A(62) => 
                           net48693, A(61) => net48694, A(60) => net48695, 
                           A(59) => net48696, A(58) => net48697, A(57) => 
                           net48698, A(56) => net48699, A(55) => net48700, 
                           A(54) => net48701, A(53) => net48702, A(52) => 
                           net48703, A(51) => net48704, A(50) => net48705, 
                           A(49) => net48706, A(48) => net48707, A(47) => 
                           net48708, A(46) => net48709, A(45) => net48710, 
                           A(44) => net48711, A(43) => net48712, A(42) => 
                           net48713, A(41) => net48714, A(40) => net48715, 
                           A(39) => net48716, A(38) => net48717, A(37) => 
                           net48718, A(36) => net48719, A(35) => net48720, 
                           A(34) => net48721, A(33) => net48722, A(32) => 
                           net48723, A(31) => net48724, A(30) => net48725, 
                           A(29) => net48726, A(28) => net48727, A(27) => 
                           net48728, A(26) => net48729, A(25) => net48730, 
                           A(24) => net48731, A(23) => net48732, A(22) => 
                           net48733, A(21) => net48734, A(20) => net48735, 
                           A(19) => net48736, A(18) => net48737, A(17) => 
                           net48738, A(16) => net48739, A(15) => net48740, 
                           A(14) => net48741, A(13) => net48742, A(12) => 
                           net48743, A(11) => net48744, A(10) => net48745, A(9)
                           => net48746, A(8) => net48747, A(7) => net48748, 
                           A(6) => net48749, A(5) => net48750, A(4) => net48751
                           , A(3) => net48752, A(2) => net48753, A(1) => 
                           net48754, A(0) => net48755, A_n(63) => net48756, 
                           A_n(62) => net48757, A_n(61) => net48758, A_n(60) =>
                           net48759, A_n(59) => net48760, A_n(58) => net48761, 
                           A_n(57) => net48762, A_n(56) => net48763, A_n(55) =>
                           net48764, A_n(54) => net48765, A_n(53) => net48766, 
                           A_n(52) => net48767, A_n(51) => net48768, A_n(50) =>
                           net48769, A_n(49) => net48770, A_n(48) => net48771, 
                           A_n(47) => net48772, A_n(46) => net48773, A_n(45) =>
                           net48774, A_n(44) => net48775, A_n(43) => net48776, 
                           A_n(42) => net48777, A_n(41) => net48778, A_n(40) =>
                           net48779, A_n(39) => net48780, A_n(38) => net48781, 
                           A_n(37) => net48782, A_n(36) => net48783, A_n(35) =>
                           net48784, A_n(34) => net48785, A_n(33) => net48786, 
                           A_n(32) => net48787, A_n(31) => net48788, A_n(30) =>
                           net48789, A_n(29) => net48790, A_n(28) => net48791, 
                           A_n(27) => net48792, A_n(26) => net48793, A_n(25) =>
                           net48794, A_n(24) => net48795, A_n(23) => net48796, 
                           A_n(22) => net48797, A_n(21) => net48798, A_n(20) =>
                           net48799, A_n(19) => net48800, A_n(18) => net48801, 
                           A_n(17) => net48802, A_n(16) => net48803, A_n(15) =>
                           net48804, A_n(14) => net48805, A_n(13) => net48806, 
                           A_n(12) => net48807, A_n(11) => net48808, A_n(10) =>
                           net48809, A_n(9) => net48810, A_n(8) => net48811, 
                           A_n(7) => net48812, A_n(6) => net48813, A_n(5) => 
                           net48814, A_n(4) => net48815, A_n(3) => net48816, 
                           A_n(2) => net48817, A_n(1) => net48818, A_n(0) => 
                           net48819, A_ns(63) => A_n_63, A_ns(62) => A_n_63, 
                           A_ns(61) => A_n_63, A_ns(60) => A_n_63, A_ns(59) => 
                           A_n_63, A_ns(58) => A_n_63, A_ns(57) => A_n_63, 
                           A_ns(56) => A_n_63, A_ns(55) => A_n_63, A_ns(54) => 
                           A_n_63, A_ns(53) => A_n_63, A_ns(52) => A_n_63, 
                           A_ns(51) => A_n_63, A_ns(50) => A_n_63, A_ns(49) => 
                           A_n_63, A_ns(48) => A_n_63, A_ns(47) => A_n_63, 
                           A_ns(46) => A_n_63, A_ns(45) => A_n_63, A_ns(44) => 
                           A_n_63, A_ns(43) => A_n_63, A_ns(42) => A_n_63, 
                           A_ns(41) => A_n_63, A_ns(40) => A_n_63, A_ns(39) => 
                           A_n_63, A_ns(38) => A_n_63, A_ns(37) => A_n_63, 
                           A_ns(36) => A_n_63, A_ns(35) => A_n_63, A_ns(34) => 
                           A_n_63, A_ns(33) => A_n_63, A_ns(32) => A_n_63, 
                           A_ns(31) => A_n_63, A_ns(30) => A_n_30_port, 
                           A_ns(29) => A_n_29_port, A_ns(28) => A_n_28_port, 
                           A_ns(27) => A_n_27_port, A_ns(26) => A_n_26_port, 
                           A_ns(25) => A_n_25_port, A_ns(24) => A_n_24_port, 
                           A_ns(23) => A_n_23_port, A_ns(22) => A_n_22_port, 
                           A_ns(21) => A_n_21_port, A_ns(20) => A_n_20_port, 
                           A_ns(19) => A_n_19_port, A_ns(18) => A_n_18_port, 
                           A_ns(17) => A_n_17_port, A_ns(16) => A_n_16_port, 
                           A_ns(15) => A_n_15_port, A_ns(14) => A_n_14_port, 
                           A_ns(13) => A_n_13_port, A_ns(12) => A_n_12_port, 
                           A_ns(11) => A_n_11_port, A_ns(10) => A_n_10_port, 
                           A_ns(9) => A_n_9_port, A_ns(8) => A_n_8_port, 
                           A_ns(7) => A_n_7_port, A_ns(6) => A_n_6_port, 
                           A_ns(5) => A_n_5_port, A_ns(4) => A_n_4_port, 
                           A_ns(3) => A_n_3_port, A_ns(2) => A_n_2_port, 
                           A_ns(1) => A_n_1_port, A_ns(0) => A_n_0_port, 
                           A_s(63) => A(31), A_s(62) => A(31), A_s(61) => A(31)
                           , A_s(60) => A(31), A_s(59) => A(31), A_s(58) => 
                           A(31), A_s(57) => A(31), A_s(56) => A(31), A_s(55) 
                           => A(31), A_s(54) => A(31), A_s(53) => A(31), 
                           A_s(52) => A(31), A_s(51) => A(31), A_s(50) => A(31)
                           , A_s(49) => A(31), A_s(48) => A(31), A_s(47) => 
                           A(31), A_s(46) => A(31), A_s(45) => A(31), A_s(44) 
                           => A(31), A_s(43) => A(31), A_s(42) => A(31), 
                           A_s(41) => A(31), A_s(40) => A(31), A_s(39) => A(31)
                           , A_s(38) => A(31), A_s(37) => A(31), A_s(36) => 
                           A(31), A_s(35) => A(31), A_s(34) => A(31), A_s(33) 
                           => A(31), A_s(32) => A(31), A_s(31) => A(31), 
                           A_s(30) => A(30), A_s(29) => A(29), A_s(28) => A(28)
                           , A_s(27) => A(27), A_s(26) => A(26), A_s(25) => 
                           A(25), A_s(24) => A(24), A_s(23) => A(23), A_s(22) 
                           => A(22), A_s(21) => A(21), A_s(20) => A(20), 
                           A_s(19) => A(19), A_s(18) => A(18), A_s(17) => A(17)
                           , A_s(16) => A(16), A_s(15) => A(15), A_s(14) => 
                           A(14), A_s(13) => A(13), A_s(12) => A(12), A_s(11) 
                           => A(11), A_s(10) => A(10), A_s(9) => A(9), A_s(8) 
                           => A(8), A_s(7) => A(7), A_s(6) => A(6), A_s(5) => 
                           A(5), A_s(4) => A(4), A_s(3) => A(3), A_s(2) => A(2)
                           , A_s(1) => A(1), A_s(0) => A(0), B(63) => B(31), 
                           B(62) => B(31), B(61) => B(31), B(60) => B(31), 
                           B(59) => B(31), B(58) => B(31), B(57) => B(31), 
                           B(56) => B(31), B(55) => B(31), B(54) => B(31), 
                           B(53) => B(31), B(52) => B(31), B(51) => B(31), 
                           B(50) => B(31), B(49) => B(31), B(48) => B(31), 
                           B(47) => B(31), B(46) => B(31), B(45) => B(31), 
                           B(44) => B(31), B(43) => B(31), B(42) => B(31), 
                           B(41) => B(31), B(40) => B(31), B(39) => B(31), 
                           B(38) => B(31), B(37) => B(31), B(36) => B(31), 
                           B(35) => B(31), B(34) => B(31), B(33) => B(31), 
                           B(32) => B(31), B(31) => B(31), B(30) => B(30), 
                           B(29) => B(29), B(28) => B(28), B(27) => B(27), 
                           B(26) => B(26), B(25) => B(25), B(24) => B(24), 
                           B(23) => B(23), B(22) => B(22), B(21) => B(21), 
                           B(20) => B(20), B(19) => B(19), B(18) => B(18), 
                           B(17) => B(17), B(16) => B(16), B(15) => B(15), 
                           B(14) => B(14), B(13) => B(13), B(12) => B(12), 
                           B(11) => B(11), B(10) => B(10), B(9) => B(9), B(8) 
                           => B(8), B(7) => B(7), B(6) => B(6), B(5) => B(5), 
                           B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), O(63) => OTMP_63_port, O(62) => 
                           OTMP_62_port, O(61) => OTMP_61_port, O(60) => 
                           OTMP_60_port, O(59) => OTMP_59_port, O(58) => 
                           OTMP_58_port, O(57) => OTMP_57_port, O(56) => 
                           OTMP_56_port, O(55) => OTMP_55_port, O(54) => 
                           OTMP_54_port, O(53) => OTMP_53_port, O(52) => 
                           OTMP_52_port, O(51) => OTMP_51_port, O(50) => 
                           OTMP_50_port, O(49) => OTMP_49_port, O(48) => 
                           OTMP_48_port, O(47) => OTMP_47_port, O(46) => 
                           OTMP_46_port, O(45) => OTMP_45_port, O(44) => 
                           OTMP_44_port, O(43) => OTMP_43_port, O(42) => 
                           OTMP_42_port, O(41) => OTMP_41_port, O(40) => 
                           OTMP_40_port, O(39) => OTMP_39_port, O(38) => 
                           OTMP_38_port, O(37) => OTMP_37_port, O(36) => 
                           OTMP_36_port, O(35) => OTMP_35_port, O(34) => 
                           OTMP_34_port, O(33) => OTMP_33_port, O(32) => 
                           OTMP_32_port, O(31) => OTMP_31_port, O(30) => 
                           OTMP_30_port, O(29) => OTMP_29_port, O(28) => 
                           OTMP_28_port, O(27) => OTMP_27_port, O(26) => 
                           OTMP_26_port, O(25) => OTMP_25_port, O(24) => 
                           OTMP_24_port, O(23) => OTMP_23_port, O(22) => 
                           OTMP_22_port, O(21) => OTMP_21_port, O(20) => 
                           OTMP_20_port, O(19) => OTMP_19_port, O(18) => 
                           OTMP_18_port, O(17) => OTMP_17_port, O(16) => 
                           OTMP_16_port, O(15) => OTMP_15_port, O(14) => 
                           OTMP_14_port, O(13) => OTMP_13_port, O(12) => 
                           OTMP_12_port, O(11) => OTMP_11_port, O(10) => 
                           OTMP_10_port, O(9) => OTMP_9_port, O(8) => 
                           OTMP_8_port, O(7) => OTMP_7_port, O(6) => 
                           OTMP_6_port, O(5) => OTMP_5_port, O(4) => 
                           OTMP_4_port, O(3) => OTMP_3_port, O(2) => 
                           OTMP_2_port, O(1) => OTMP_1_port, O(0) => 
                           OTMP_0_port, A_so(63) => SHIFT_127_port, A_so(62) =>
                           SHIFT_126_port, A_so(61) => SHIFT_125_port, A_so(60)
                           => SHIFT_124_port, A_so(59) => SHIFT_123_port, 
                           A_so(58) => SHIFT_122_port, A_so(57) => 
                           SHIFT_121_port, A_so(56) => SHIFT_120_port, A_so(55)
                           => SHIFT_119_port, A_so(54) => SHIFT_118_port, 
                           A_so(53) => SHIFT_117_port, A_so(52) => 
                           SHIFT_116_port, A_so(51) => SHIFT_115_port, A_so(50)
                           => SHIFT_114_port, A_so(49) => SHIFT_113_port, 
                           A_so(48) => SHIFT_112_port, A_so(47) => 
                           SHIFT_111_port, A_so(46) => SHIFT_110_port, A_so(45)
                           => SHIFT_109_port, A_so(44) => SHIFT_108_port, 
                           A_so(43) => SHIFT_107_port, A_so(42) => 
                           SHIFT_106_port, A_so(41) => SHIFT_105_port, A_so(40)
                           => SHIFT_104_port, A_so(39) => SHIFT_103_port, 
                           A_so(38) => SHIFT_102_port, A_so(37) => 
                           SHIFT_101_port, A_so(36) => SHIFT_100_port, A_so(35)
                           => SHIFT_99_port, A_so(34) => SHIFT_98_port, 
                           A_so(33) => SHIFT_97_port, A_so(32) => SHIFT_96_port
                           , A_so(31) => SHIFT_95_port, A_so(30) => 
                           SHIFT_94_port, A_so(29) => SHIFT_93_port, A_so(28) 
                           => SHIFT_92_port, A_so(27) => SHIFT_91_port, 
                           A_so(26) => SHIFT_90_port, A_so(25) => SHIFT_89_port
                           , A_so(24) => SHIFT_88_port, A_so(23) => 
                           SHIFT_87_port, A_so(22) => SHIFT_86_port, A_so(21) 
                           => SHIFT_85_port, A_so(20) => SHIFT_84_port, 
                           A_so(19) => SHIFT_83_port, A_so(18) => SHIFT_82_port
                           , A_so(17) => SHIFT_81_port, A_so(16) => 
                           SHIFT_80_port, A_so(15) => SHIFT_79_port, A_so(14) 
                           => SHIFT_78_port, A_so(13) => SHIFT_77_port, 
                           A_so(12) => SHIFT_76_port, A_so(11) => SHIFT_75_port
                           , A_so(10) => SHIFT_74_port, A_so(9) => 
                           SHIFT_73_port, A_so(8) => SHIFT_72_port, A_so(7) => 
                           SHIFT_71_port, A_so(6) => SHIFT_70_port, A_so(5) => 
                           SHIFT_69_port, A_so(4) => SHIFT_68_port, A_so(3) => 
                           SHIFT_67_port, A_so(2) => SHIFT_66_port, A_so(1) => 
                           SHIFT_65_port, A_so(0) => n_1094, A_nso(63) => 
                           SHIFT_n_127_port, A_nso(62) => SHIFT_n_126_port, 
                           A_nso(61) => SHIFT_n_125_port, A_nso(60) => 
                           SHIFT_n_124_port, A_nso(59) => SHIFT_n_123_port, 
                           A_nso(58) => SHIFT_n_122_port, A_nso(57) => 
                           SHIFT_n_121_port, A_nso(56) => SHIFT_n_120_port, 
                           A_nso(55) => SHIFT_n_119_port, A_nso(54) => 
                           SHIFT_n_118_port, A_nso(53) => SHIFT_n_117_port, 
                           A_nso(52) => SHIFT_n_116_port, A_nso(51) => 
                           SHIFT_n_115_port, A_nso(50) => SHIFT_n_114_port, 
                           A_nso(49) => SHIFT_n_113_port, A_nso(48) => 
                           SHIFT_n_112_port, A_nso(47) => SHIFT_n_111_port, 
                           A_nso(46) => SHIFT_n_110_port, A_nso(45) => 
                           SHIFT_n_109_port, A_nso(44) => SHIFT_n_108_port, 
                           A_nso(43) => SHIFT_n_107_port, A_nso(42) => 
                           SHIFT_n_106_port, A_nso(41) => SHIFT_n_105_port, 
                           A_nso(40) => SHIFT_n_104_port, A_nso(39) => 
                           SHIFT_n_103_port, A_nso(38) => SHIFT_n_102_port, 
                           A_nso(37) => SHIFT_n_101_port, A_nso(36) => 
                           SHIFT_n_100_port, A_nso(35) => SHIFT_n_99_port, 
                           A_nso(34) => SHIFT_n_98_port, A_nso(33) => 
                           SHIFT_n_97_port, A_nso(32) => SHIFT_n_96_port, 
                           A_nso(31) => SHIFT_n_95_port, A_nso(30) => 
                           SHIFT_n_94_port, A_nso(29) => SHIFT_n_93_port, 
                           A_nso(28) => SHIFT_n_92_port, A_nso(27) => 
                           SHIFT_n_91_port, A_nso(26) => SHIFT_n_90_port, 
                           A_nso(25) => SHIFT_n_89_port, A_nso(24) => 
                           SHIFT_n_88_port, A_nso(23) => SHIFT_n_87_port, 
                           A_nso(22) => SHIFT_n_86_port, A_nso(21) => 
                           SHIFT_n_85_port, A_nso(20) => SHIFT_n_84_port, 
                           A_nso(19) => SHIFT_n_83_port, A_nso(18) => 
                           SHIFT_n_82_port, A_nso(17) => SHIFT_n_81_port, 
                           A_nso(16) => SHIFT_n_80_port, A_nso(15) => 
                           SHIFT_n_79_port, A_nso(14) => SHIFT_n_78_port, 
                           A_nso(13) => SHIFT_n_77_port, A_nso(12) => 
                           SHIFT_n_76_port, A_nso(11) => SHIFT_n_75_port, 
                           A_nso(10) => SHIFT_n_74_port, A_nso(9) => 
                           SHIFT_n_73_port, A_nso(8) => SHIFT_n_72_port, 
                           A_nso(7) => SHIFT_n_71_port, A_nso(6) => 
                           SHIFT_n_70_port, A_nso(5) => SHIFT_n_69_port, 
                           A_nso(4) => SHIFT_n_68_port, A_nso(3) => 
                           SHIFT_n_67_port, A_nso(2) => SHIFT_n_66_port, 
                           A_nso(1) => SHIFT_n_65_port, A_nso(0) => n_1095);
   BOOTHENC_I_2 : BOOTHENC_NBIT64_i2 port map( A(63) => net48564, A(62) => 
                           net48565, A(61) => net48566, A(60) => net48567, 
                           A(59) => net48568, A(58) => net48569, A(57) => 
                           net48570, A(56) => net48571, A(55) => net48572, 
                           A(54) => net48573, A(53) => net48574, A(52) => 
                           net48575, A(51) => net48576, A(50) => net48577, 
                           A(49) => net48578, A(48) => net48579, A(47) => 
                           net48580, A(46) => net48581, A(45) => net48582, 
                           A(44) => net48583, A(43) => net48584, A(42) => 
                           net48585, A(41) => net48586, A(40) => net48587, 
                           A(39) => net48588, A(38) => net48589, A(37) => 
                           net48590, A(36) => net48591, A(35) => net48592, 
                           A(34) => net48593, A(33) => net48594, A(32) => 
                           net48595, A(31) => net48596, A(30) => net48597, 
                           A(29) => net48598, A(28) => net48599, A(27) => 
                           net48600, A(26) => net48601, A(25) => net48602, 
                           A(24) => net48603, A(23) => net48604, A(22) => 
                           net48605, A(21) => net48606, A(20) => net48607, 
                           A(19) => net48608, A(18) => net48609, A(17) => 
                           net48610, A(16) => net48611, A(15) => net48612, 
                           A(14) => net48613, A(13) => net48614, A(12) => 
                           net48615, A(11) => net48616, A(10) => net48617, A(9)
                           => net48618, A(8) => net48619, A(7) => net48620, 
                           A(6) => net48621, A(5) => net48622, A(4) => net48623
                           , A(3) => net48624, A(2) => net48625, A(1) => 
                           net48626, A(0) => net48627, A_n(63) => net48628, 
                           A_n(62) => net48629, A_n(61) => net48630, A_n(60) =>
                           net48631, A_n(59) => net48632, A_n(58) => net48633, 
                           A_n(57) => net48634, A_n(56) => net48635, A_n(55) =>
                           net48636, A_n(54) => net48637, A_n(53) => net48638, 
                           A_n(52) => net48639, A_n(51) => net48640, A_n(50) =>
                           net48641, A_n(49) => net48642, A_n(48) => net48643, 
                           A_n(47) => net48644, A_n(46) => net48645, A_n(45) =>
                           net48646, A_n(44) => net48647, A_n(43) => net48648, 
                           A_n(42) => net48649, A_n(41) => net48650, A_n(40) =>
                           net48651, A_n(39) => net48652, A_n(38) => net48653, 
                           A_n(37) => net48654, A_n(36) => net48655, A_n(35) =>
                           net48656, A_n(34) => net48657, A_n(33) => net48658, 
                           A_n(32) => net48659, A_n(31) => net48660, A_n(30) =>
                           net48661, A_n(29) => net48662, A_n(28) => net48663, 
                           A_n(27) => net48664, A_n(26) => net48665, A_n(25) =>
                           net48666, A_n(24) => net48667, A_n(23) => net48668, 
                           A_n(22) => net48669, A_n(21) => net48670, A_n(20) =>
                           net48671, A_n(19) => net48672, A_n(18) => net48673, 
                           A_n(17) => net48674, A_n(16) => net48675, A_n(15) =>
                           net48676, A_n(14) => net48677, A_n(13) => net48678, 
                           A_n(12) => net48679, A_n(11) => net48680, A_n(10) =>
                           net48681, A_n(9) => net48682, A_n(8) => net48683, 
                           A_n(7) => net48684, A_n(6) => net48685, A_n(5) => 
                           net48686, A_n(4) => net48687, A_n(3) => net48688, 
                           A_n(2) => net48689, A_n(1) => net48690, A_n(0) => 
                           net48691, A_ns(63) => SHIFT_n_127_port, A_ns(62) => 
                           SHIFT_n_126_port, A_ns(61) => SHIFT_n_125_port, 
                           A_ns(60) => SHIFT_n_124_port, A_ns(59) => 
                           SHIFT_n_123_port, A_ns(58) => SHIFT_n_122_port, 
                           A_ns(57) => SHIFT_n_121_port, A_ns(56) => 
                           SHIFT_n_120_port, A_ns(55) => SHIFT_n_119_port, 
                           A_ns(54) => SHIFT_n_118_port, A_ns(53) => 
                           SHIFT_n_117_port, A_ns(52) => SHIFT_n_116_port, 
                           A_ns(51) => SHIFT_n_115_port, A_ns(50) => 
                           SHIFT_n_114_port, A_ns(49) => SHIFT_n_113_port, 
                           A_ns(48) => SHIFT_n_112_port, A_ns(47) => 
                           SHIFT_n_111_port, A_ns(46) => SHIFT_n_110_port, 
                           A_ns(45) => SHIFT_n_109_port, A_ns(44) => 
                           SHIFT_n_108_port, A_ns(43) => SHIFT_n_107_port, 
                           A_ns(42) => SHIFT_n_106_port, A_ns(41) => 
                           SHIFT_n_105_port, A_ns(40) => SHIFT_n_104_port, 
                           A_ns(39) => SHIFT_n_103_port, A_ns(38) => 
                           SHIFT_n_102_port, A_ns(37) => SHIFT_n_101_port, 
                           A_ns(36) => SHIFT_n_100_port, A_ns(35) => 
                           SHIFT_n_99_port, A_ns(34) => SHIFT_n_98_port, 
                           A_ns(33) => SHIFT_n_97_port, A_ns(32) => 
                           SHIFT_n_96_port, A_ns(31) => SHIFT_n_95_port, 
                           A_ns(30) => SHIFT_n_94_port, A_ns(29) => 
                           SHIFT_n_93_port, A_ns(28) => SHIFT_n_92_port, 
                           A_ns(27) => SHIFT_n_91_port, A_ns(26) => 
                           SHIFT_n_90_port, A_ns(25) => SHIFT_n_89_port, 
                           A_ns(24) => SHIFT_n_88_port, A_ns(23) => 
                           SHIFT_n_87_port, A_ns(22) => SHIFT_n_86_port, 
                           A_ns(21) => SHIFT_n_85_port, A_ns(20) => 
                           SHIFT_n_84_port, A_ns(19) => SHIFT_n_83_port, 
                           A_ns(18) => SHIFT_n_82_port, A_ns(17) => 
                           SHIFT_n_81_port, A_ns(16) => SHIFT_n_80_port, 
                           A_ns(15) => SHIFT_n_79_port, A_ns(14) => 
                           SHIFT_n_78_port, A_ns(13) => SHIFT_n_77_port, 
                           A_ns(12) => SHIFT_n_76_port, A_ns(11) => 
                           SHIFT_n_75_port, A_ns(10) => SHIFT_n_74_port, 
                           A_ns(9) => SHIFT_n_73_port, A_ns(8) => 
                           SHIFT_n_72_port, A_ns(7) => SHIFT_n_71_port, A_ns(6)
                           => SHIFT_n_70_port, A_ns(5) => SHIFT_n_69_port, 
                           A_ns(4) => SHIFT_n_68_port, A_ns(3) => 
                           SHIFT_n_67_port, A_ns(2) => SHIFT_n_66_port, A_ns(1)
                           => SHIFT_n_65_port, A_ns(0) => SHIFT_n_64_port, 
                           A_s(63) => SHIFT_127_port, A_s(62) => SHIFT_126_port
                           , A_s(61) => SHIFT_125_port, A_s(60) => 
                           SHIFT_124_port, A_s(59) => SHIFT_123_port, A_s(58) 
                           => SHIFT_122_port, A_s(57) => SHIFT_121_port, 
                           A_s(56) => SHIFT_120_port, A_s(55) => SHIFT_119_port
                           , A_s(54) => SHIFT_118_port, A_s(53) => 
                           SHIFT_117_port, A_s(52) => SHIFT_116_port, A_s(51) 
                           => SHIFT_115_port, A_s(50) => SHIFT_114_port, 
                           A_s(49) => SHIFT_113_port, A_s(48) => SHIFT_112_port
                           , A_s(47) => SHIFT_111_port, A_s(46) => 
                           SHIFT_110_port, A_s(45) => SHIFT_109_port, A_s(44) 
                           => SHIFT_108_port, A_s(43) => SHIFT_107_port, 
                           A_s(42) => SHIFT_106_port, A_s(41) => SHIFT_105_port
                           , A_s(40) => SHIFT_104_port, A_s(39) => 
                           SHIFT_103_port, A_s(38) => SHIFT_102_port, A_s(37) 
                           => SHIFT_101_port, A_s(36) => SHIFT_100_port, 
                           A_s(35) => SHIFT_99_port, A_s(34) => SHIFT_98_port, 
                           A_s(33) => SHIFT_97_port, A_s(32) => SHIFT_96_port, 
                           A_s(31) => SHIFT_95_port, A_s(30) => SHIFT_94_port, 
                           A_s(29) => SHIFT_93_port, A_s(28) => SHIFT_92_port, 
                           A_s(27) => SHIFT_91_port, A_s(26) => SHIFT_90_port, 
                           A_s(25) => SHIFT_89_port, A_s(24) => SHIFT_88_port, 
                           A_s(23) => SHIFT_87_port, A_s(22) => SHIFT_86_port, 
                           A_s(21) => SHIFT_85_port, A_s(20) => SHIFT_84_port, 
                           A_s(19) => SHIFT_83_port, A_s(18) => SHIFT_82_port, 
                           A_s(17) => SHIFT_81_port, A_s(16) => SHIFT_80_port, 
                           A_s(15) => SHIFT_79_port, A_s(14) => SHIFT_78_port, 
                           A_s(13) => SHIFT_77_port, A_s(12) => SHIFT_76_port, 
                           A_s(11) => SHIFT_75_port, A_s(10) => SHIFT_74_port, 
                           A_s(9) => SHIFT_73_port, A_s(8) => SHIFT_72_port, 
                           A_s(7) => SHIFT_71_port, A_s(6) => SHIFT_70_port, 
                           A_s(5) => SHIFT_69_port, A_s(4) => SHIFT_68_port, 
                           A_s(3) => SHIFT_67_port, A_s(2) => SHIFT_66_port, 
                           A_s(1) => SHIFT_65_port, A_s(0) => SHIFT_64_port, 
                           B(63) => B(31), B(62) => B(31), B(61) => B(31), 
                           B(60) => B(31), B(59) => B(31), B(58) => B(31), 
                           B(57) => B(31), B(56) => B(31), B(55) => B(31), 
                           B(54) => B(31), B(53) => B(31), B(52) => B(31), 
                           B(51) => B(31), B(50) => B(31), B(49) => B(31), 
                           B(48) => B(31), B(47) => B(31), B(46) => B(31), 
                           B(45) => B(31), B(44) => B(31), B(43) => B(31), 
                           B(42) => B(31), B(41) => B(31), B(40) => B(31), 
                           B(39) => B(31), B(38) => B(31), B(37) => B(31), 
                           B(36) => B(31), B(35) => B(31), B(34) => B(31), 
                           B(33) => B(31), B(32) => B(31), B(31) => B(31), 
                           B(30) => B(30), B(29) => B(29), B(28) => B(28), 
                           B(27) => B(27), B(26) => B(26), B(25) => B(25), 
                           B(24) => B(24), B(23) => B(23), B(22) => B(22), 
                           B(21) => B(21), B(20) => B(20), B(19) => B(19), 
                           B(18) => B(18), B(17) => B(17), B(16) => B(16), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => B(0), O(63) => 
                           OTMP_127_port, O(62) => OTMP_126_port, O(61) => 
                           OTMP_125_port, O(60) => OTMP_124_port, O(59) => 
                           OTMP_123_port, O(58) => OTMP_122_port, O(57) => 
                           OTMP_121_port, O(56) => OTMP_120_port, O(55) => 
                           OTMP_119_port, O(54) => OTMP_118_port, O(53) => 
                           OTMP_117_port, O(52) => OTMP_116_port, O(51) => 
                           OTMP_115_port, O(50) => OTMP_114_port, O(49) => 
                           OTMP_113_port, O(48) => OTMP_112_port, O(47) => 
                           OTMP_111_port, O(46) => OTMP_110_port, O(45) => 
                           OTMP_109_port, O(44) => OTMP_108_port, O(43) => 
                           OTMP_107_port, O(42) => OTMP_106_port, O(41) => 
                           OTMP_105_port, O(40) => OTMP_104_port, O(39) => 
                           OTMP_103_port, O(38) => OTMP_102_port, O(37) => 
                           OTMP_101_port, O(36) => OTMP_100_port, O(35) => 
                           OTMP_99_port, O(34) => OTMP_98_port, O(33) => 
                           OTMP_97_port, O(32) => OTMP_96_port, O(31) => 
                           OTMP_95_port, O(30) => OTMP_94_port, O(29) => 
                           OTMP_93_port, O(28) => OTMP_92_port, O(27) => 
                           OTMP_91_port, O(26) => OTMP_90_port, O(25) => 
                           OTMP_89_port, O(24) => OTMP_88_port, O(23) => 
                           OTMP_87_port, O(22) => OTMP_86_port, O(21) => 
                           OTMP_85_port, O(20) => OTMP_84_port, O(19) => 
                           OTMP_83_port, O(18) => OTMP_82_port, O(17) => 
                           OTMP_81_port, O(16) => OTMP_80_port, O(15) => 
                           OTMP_79_port, O(14) => OTMP_78_port, O(13) => 
                           OTMP_77_port, O(12) => OTMP_76_port, O(11) => 
                           OTMP_75_port, O(10) => OTMP_74_port, O(9) => 
                           OTMP_73_port, O(8) => OTMP_72_port, O(7) => 
                           OTMP_71_port, O(6) => OTMP_70_port, O(5) => 
                           OTMP_69_port, O(4) => OTMP_68_port, O(3) => 
                           OTMP_67_port, O(2) => OTMP_66_port, O(1) => 
                           OTMP_65_port, O(0) => n_1096, A_so(63) => 
                           SHIFT_191_port, A_so(62) => SHIFT_190_port, A_so(61)
                           => SHIFT_189_port, A_so(60) => SHIFT_188_port, 
                           A_so(59) => SHIFT_187_port, A_so(58) => 
                           SHIFT_186_port, A_so(57) => SHIFT_185_port, A_so(56)
                           => SHIFT_184_port, A_so(55) => SHIFT_183_port, 
                           A_so(54) => SHIFT_182_port, A_so(53) => 
                           SHIFT_181_port, A_so(52) => SHIFT_180_port, A_so(51)
                           => SHIFT_179_port, A_so(50) => SHIFT_178_port, 
                           A_so(49) => SHIFT_177_port, A_so(48) => 
                           SHIFT_176_port, A_so(47) => SHIFT_175_port, A_so(46)
                           => SHIFT_174_port, A_so(45) => SHIFT_173_port, 
                           A_so(44) => SHIFT_172_port, A_so(43) => 
                           SHIFT_171_port, A_so(42) => SHIFT_170_port, A_so(41)
                           => SHIFT_169_port, A_so(40) => SHIFT_168_port, 
                           A_so(39) => SHIFT_167_port, A_so(38) => 
                           SHIFT_166_port, A_so(37) => SHIFT_165_port, A_so(36)
                           => SHIFT_164_port, A_so(35) => SHIFT_163_port, 
                           A_so(34) => SHIFT_162_port, A_so(33) => 
                           SHIFT_161_port, A_so(32) => SHIFT_160_port, A_so(31)
                           => SHIFT_159_port, A_so(30) => SHIFT_158_port, 
                           A_so(29) => SHIFT_157_port, A_so(28) => 
                           SHIFT_156_port, A_so(27) => SHIFT_155_port, A_so(26)
                           => SHIFT_154_port, A_so(25) => SHIFT_153_port, 
                           A_so(24) => SHIFT_152_port, A_so(23) => 
                           SHIFT_151_port, A_so(22) => SHIFT_150_port, A_so(21)
                           => SHIFT_149_port, A_so(20) => SHIFT_148_port, 
                           A_so(19) => SHIFT_147_port, A_so(18) => 
                           SHIFT_146_port, A_so(17) => SHIFT_145_port, A_so(16)
                           => SHIFT_144_port, A_so(15) => SHIFT_143_port, 
                           A_so(14) => SHIFT_142_port, A_so(13) => 
                           SHIFT_141_port, A_so(12) => SHIFT_140_port, A_so(11)
                           => SHIFT_139_port, A_so(10) => SHIFT_138_port, 
                           A_so(9) => SHIFT_137_port, A_so(8) => SHIFT_136_port
                           , A_so(7) => SHIFT_135_port, A_so(6) => 
                           SHIFT_134_port, A_so(5) => SHIFT_133_port, A_so(4) 
                           => SHIFT_132_port, A_so(3) => SHIFT_131_port, 
                           A_so(2) => SHIFT_130_port, A_so(1) => n_1097, 
                           A_so(0) => n_1098, A_nso(63) => SHIFT_n_191_port, 
                           A_nso(62) => SHIFT_n_190_port, A_nso(61) => 
                           SHIFT_n_189_port, A_nso(60) => SHIFT_n_188_port, 
                           A_nso(59) => SHIFT_n_187_port, A_nso(58) => 
                           SHIFT_n_186_port, A_nso(57) => SHIFT_n_185_port, 
                           A_nso(56) => SHIFT_n_184_port, A_nso(55) => 
                           SHIFT_n_183_port, A_nso(54) => SHIFT_n_182_port, 
                           A_nso(53) => SHIFT_n_181_port, A_nso(52) => 
                           SHIFT_n_180_port, A_nso(51) => SHIFT_n_179_port, 
                           A_nso(50) => SHIFT_n_178_port, A_nso(49) => 
                           SHIFT_n_177_port, A_nso(48) => SHIFT_n_176_port, 
                           A_nso(47) => SHIFT_n_175_port, A_nso(46) => 
                           SHIFT_n_174_port, A_nso(45) => SHIFT_n_173_port, 
                           A_nso(44) => SHIFT_n_172_port, A_nso(43) => 
                           SHIFT_n_171_port, A_nso(42) => SHIFT_n_170_port, 
                           A_nso(41) => SHIFT_n_169_port, A_nso(40) => 
                           SHIFT_n_168_port, A_nso(39) => SHIFT_n_167_port, 
                           A_nso(38) => SHIFT_n_166_port, A_nso(37) => 
                           SHIFT_n_165_port, A_nso(36) => SHIFT_n_164_port, 
                           A_nso(35) => SHIFT_n_163_port, A_nso(34) => 
                           SHIFT_n_162_port, A_nso(33) => SHIFT_n_161_port, 
                           A_nso(32) => SHIFT_n_160_port, A_nso(31) => 
                           SHIFT_n_159_port, A_nso(30) => SHIFT_n_158_port, 
                           A_nso(29) => SHIFT_n_157_port, A_nso(28) => 
                           SHIFT_n_156_port, A_nso(27) => SHIFT_n_155_port, 
                           A_nso(26) => SHIFT_n_154_port, A_nso(25) => 
                           SHIFT_n_153_port, A_nso(24) => SHIFT_n_152_port, 
                           A_nso(23) => SHIFT_n_151_port, A_nso(22) => 
                           SHIFT_n_150_port, A_nso(21) => SHIFT_n_149_port, 
                           A_nso(20) => SHIFT_n_148_port, A_nso(19) => 
                           SHIFT_n_147_port, A_nso(18) => SHIFT_n_146_port, 
                           A_nso(17) => SHIFT_n_145_port, A_nso(16) => 
                           SHIFT_n_144_port, A_nso(15) => SHIFT_n_143_port, 
                           A_nso(14) => SHIFT_n_142_port, A_nso(13) => 
                           SHIFT_n_141_port, A_nso(12) => SHIFT_n_140_port, 
                           A_nso(11) => SHIFT_n_139_port, A_nso(10) => 
                           SHIFT_n_138_port, A_nso(9) => SHIFT_n_137_port, 
                           A_nso(8) => SHIFT_n_136_port, A_nso(7) => 
                           SHIFT_n_135_port, A_nso(6) => SHIFT_n_134_port, 
                           A_nso(5) => SHIFT_n_133_port, A_nso(4) => 
                           SHIFT_n_132_port, A_nso(3) => SHIFT_n_131_port, 
                           A_nso(2) => SHIFT_n_130_port, A_nso(1) => n_1099, 
                           A_nso(0) => n_1100);
   BOOTHENC_I_3 : BOOTHENC_NBIT64_i4 port map( A(63) => net48436, A(62) => 
                           net48437, A(61) => net48438, A(60) => net48439, 
                           A(59) => net48440, A(58) => net48441, A(57) => 
                           net48442, A(56) => net48443, A(55) => net48444, 
                           A(54) => net48445, A(53) => net48446, A(52) => 
                           net48447, A(51) => net48448, A(50) => net48449, 
                           A(49) => net48450, A(48) => net48451, A(47) => 
                           net48452, A(46) => net48453, A(45) => net48454, 
                           A(44) => net48455, A(43) => net48456, A(42) => 
                           net48457, A(41) => net48458, A(40) => net48459, 
                           A(39) => net48460, A(38) => net48461, A(37) => 
                           net48462, A(36) => net48463, A(35) => net48464, 
                           A(34) => net48465, A(33) => net48466, A(32) => 
                           net48467, A(31) => net48468, A(30) => net48469, 
                           A(29) => net48470, A(28) => net48471, A(27) => 
                           net48472, A(26) => net48473, A(25) => net48474, 
                           A(24) => net48475, A(23) => net48476, A(22) => 
                           net48477, A(21) => net48478, A(20) => net48479, 
                           A(19) => net48480, A(18) => net48481, A(17) => 
                           net48482, A(16) => net48483, A(15) => net48484, 
                           A(14) => net48485, A(13) => net48486, A(12) => 
                           net48487, A(11) => net48488, A(10) => net48489, A(9)
                           => net48490, A(8) => net48491, A(7) => net48492, 
                           A(6) => net48493, A(5) => net48494, A(4) => net48495
                           , A(3) => net48496, A(2) => net48497, A(1) => 
                           net48498, A(0) => net48499, A_n(63) => net48500, 
                           A_n(62) => net48501, A_n(61) => net48502, A_n(60) =>
                           net48503, A_n(59) => net48504, A_n(58) => net48505, 
                           A_n(57) => net48506, A_n(56) => net48507, A_n(55) =>
                           net48508, A_n(54) => net48509, A_n(53) => net48510, 
                           A_n(52) => net48511, A_n(51) => net48512, A_n(50) =>
                           net48513, A_n(49) => net48514, A_n(48) => net48515, 
                           A_n(47) => net48516, A_n(46) => net48517, A_n(45) =>
                           net48518, A_n(44) => net48519, A_n(43) => net48520, 
                           A_n(42) => net48521, A_n(41) => net48522, A_n(40) =>
                           net48523, A_n(39) => net48524, A_n(38) => net48525, 
                           A_n(37) => net48526, A_n(36) => net48527, A_n(35) =>
                           net48528, A_n(34) => net48529, A_n(33) => net48530, 
                           A_n(32) => net48531, A_n(31) => net48532, A_n(30) =>
                           net48533, A_n(29) => net48534, A_n(28) => net48535, 
                           A_n(27) => net48536, A_n(26) => net48537, A_n(25) =>
                           net48538, A_n(24) => net48539, A_n(23) => net48540, 
                           A_n(22) => net48541, A_n(21) => net48542, A_n(20) =>
                           net48543, A_n(19) => net48544, A_n(18) => net48545, 
                           A_n(17) => net48546, A_n(16) => net48547, A_n(15) =>
                           net48548, A_n(14) => net48549, A_n(13) => net48550, 
                           A_n(12) => net48551, A_n(11) => net48552, A_n(10) =>
                           net48553, A_n(9) => net48554, A_n(8) => net48555, 
                           A_n(7) => net48556, A_n(6) => net48557, A_n(5) => 
                           net48558, A_n(4) => net48559, A_n(3) => net48560, 
                           A_n(2) => net48561, A_n(1) => net48562, A_n(0) => 
                           net48563, A_ns(63) => SHIFT_n_191_port, A_ns(62) => 
                           SHIFT_n_190_port, A_ns(61) => SHIFT_n_189_port, 
                           A_ns(60) => SHIFT_n_188_port, A_ns(59) => 
                           SHIFT_n_187_port, A_ns(58) => SHIFT_n_186_port, 
                           A_ns(57) => SHIFT_n_185_port, A_ns(56) => 
                           SHIFT_n_184_port, A_ns(55) => SHIFT_n_183_port, 
                           A_ns(54) => SHIFT_n_182_port, A_ns(53) => 
                           SHIFT_n_181_port, A_ns(52) => SHIFT_n_180_port, 
                           A_ns(51) => SHIFT_n_179_port, A_ns(50) => 
                           SHIFT_n_178_port, A_ns(49) => SHIFT_n_177_port, 
                           A_ns(48) => SHIFT_n_176_port, A_ns(47) => 
                           SHIFT_n_175_port, A_ns(46) => SHIFT_n_174_port, 
                           A_ns(45) => SHIFT_n_173_port, A_ns(44) => 
                           SHIFT_n_172_port, A_ns(43) => SHIFT_n_171_port, 
                           A_ns(42) => SHIFT_n_170_port, A_ns(41) => 
                           SHIFT_n_169_port, A_ns(40) => SHIFT_n_168_port, 
                           A_ns(39) => SHIFT_n_167_port, A_ns(38) => 
                           SHIFT_n_166_port, A_ns(37) => SHIFT_n_165_port, 
                           A_ns(36) => SHIFT_n_164_port, A_ns(35) => 
                           SHIFT_n_163_port, A_ns(34) => SHIFT_n_162_port, 
                           A_ns(33) => SHIFT_n_161_port, A_ns(32) => 
                           SHIFT_n_160_port, A_ns(31) => SHIFT_n_159_port, 
                           A_ns(30) => SHIFT_n_158_port, A_ns(29) => 
                           SHIFT_n_157_port, A_ns(28) => SHIFT_n_156_port, 
                           A_ns(27) => SHIFT_n_155_port, A_ns(26) => 
                           SHIFT_n_154_port, A_ns(25) => SHIFT_n_153_port, 
                           A_ns(24) => SHIFT_n_152_port, A_ns(23) => 
                           SHIFT_n_151_port, A_ns(22) => SHIFT_n_150_port, 
                           A_ns(21) => SHIFT_n_149_port, A_ns(20) => 
                           SHIFT_n_148_port, A_ns(19) => SHIFT_n_147_port, 
                           A_ns(18) => SHIFT_n_146_port, A_ns(17) => 
                           SHIFT_n_145_port, A_ns(16) => SHIFT_n_144_port, 
                           A_ns(15) => SHIFT_n_143_port, A_ns(14) => 
                           SHIFT_n_142_port, A_ns(13) => SHIFT_n_141_port, 
                           A_ns(12) => SHIFT_n_140_port, A_ns(11) => 
                           SHIFT_n_139_port, A_ns(10) => SHIFT_n_138_port, 
                           A_ns(9) => SHIFT_n_137_port, A_ns(8) => 
                           SHIFT_n_136_port, A_ns(7) => SHIFT_n_135_port, 
                           A_ns(6) => SHIFT_n_134_port, A_ns(5) => 
                           SHIFT_n_133_port, A_ns(4) => SHIFT_n_132_port, 
                           A_ns(3) => SHIFT_n_131_port, A_ns(2) => 
                           SHIFT_n_130_port, A_ns(1) => SHIFT_n_129_port, 
                           A_ns(0) => SHIFT_n_128_port, A_s(63) => 
                           SHIFT_191_port, A_s(62) => SHIFT_190_port, A_s(61) 
                           => SHIFT_189_port, A_s(60) => SHIFT_188_port, 
                           A_s(59) => SHIFT_187_port, A_s(58) => SHIFT_186_port
                           , A_s(57) => SHIFT_185_port, A_s(56) => 
                           SHIFT_184_port, A_s(55) => SHIFT_183_port, A_s(54) 
                           => SHIFT_182_port, A_s(53) => SHIFT_181_port, 
                           A_s(52) => SHIFT_180_port, A_s(51) => SHIFT_179_port
                           , A_s(50) => SHIFT_178_port, A_s(49) => 
                           SHIFT_177_port, A_s(48) => SHIFT_176_port, A_s(47) 
                           => SHIFT_175_port, A_s(46) => SHIFT_174_port, 
                           A_s(45) => SHIFT_173_port, A_s(44) => SHIFT_172_port
                           , A_s(43) => SHIFT_171_port, A_s(42) => 
                           SHIFT_170_port, A_s(41) => SHIFT_169_port, A_s(40) 
                           => SHIFT_168_port, A_s(39) => SHIFT_167_port, 
                           A_s(38) => SHIFT_166_port, A_s(37) => SHIFT_165_port
                           , A_s(36) => SHIFT_164_port, A_s(35) => 
                           SHIFT_163_port, A_s(34) => SHIFT_162_port, A_s(33) 
                           => SHIFT_161_port, A_s(32) => SHIFT_160_port, 
                           A_s(31) => SHIFT_159_port, A_s(30) => SHIFT_158_port
                           , A_s(29) => SHIFT_157_port, A_s(28) => 
                           SHIFT_156_port, A_s(27) => SHIFT_155_port, A_s(26) 
                           => SHIFT_154_port, A_s(25) => SHIFT_153_port, 
                           A_s(24) => SHIFT_152_port, A_s(23) => SHIFT_151_port
                           , A_s(22) => SHIFT_150_port, A_s(21) => 
                           SHIFT_149_port, A_s(20) => SHIFT_148_port, A_s(19) 
                           => SHIFT_147_port, A_s(18) => SHIFT_146_port, 
                           A_s(17) => SHIFT_145_port, A_s(16) => SHIFT_144_port
                           , A_s(15) => SHIFT_143_port, A_s(14) => 
                           SHIFT_142_port, A_s(13) => SHIFT_141_port, A_s(12) 
                           => SHIFT_140_port, A_s(11) => SHIFT_139_port, 
                           A_s(10) => SHIFT_138_port, A_s(9) => SHIFT_137_port,
                           A_s(8) => SHIFT_136_port, A_s(7) => SHIFT_135_port, 
                           A_s(6) => SHIFT_134_port, A_s(5) => SHIFT_133_port, 
                           A_s(4) => SHIFT_132_port, A_s(3) => SHIFT_131_port, 
                           A_s(2) => SHIFT_130_port, A_s(1) => SHIFT_129_port, 
                           A_s(0) => SHIFT_128_port, B(63) => B(31), B(62) => 
                           B(31), B(61) => B(31), B(60) => B(31), B(59) => 
                           B(31), B(58) => B(31), B(57) => B(31), B(56) => 
                           B(31), B(55) => B(31), B(54) => B(31), B(53) => 
                           B(31), B(52) => B(31), B(51) => B(31), B(50) => 
                           B(31), B(49) => B(31), B(48) => B(31), B(47) => 
                           B(31), B(46) => B(31), B(45) => B(31), B(44) => 
                           B(31), B(43) => B(31), B(42) => B(31), B(41) => 
                           B(31), B(40) => B(31), B(39) => B(31), B(38) => 
                           B(31), B(37) => B(31), B(36) => B(31), B(35) => 
                           B(31), B(34) => B(31), B(33) => B(31), B(32) => 
                           B(31), B(31) => B(31), B(30) => B(30), B(29) => 
                           B(29), B(28) => B(28), B(27) => B(27), B(26) => 
                           B(26), B(25) => B(25), B(24) => B(24), B(23) => 
                           B(23), B(22) => B(22), B(21) => B(21), B(20) => 
                           B(20), B(19) => B(19), B(18) => B(18), B(17) => 
                           B(17), B(16) => B(16), B(15) => B(15), B(14) => 
                           B(14), B(13) => B(13), B(12) => B(12), B(11) => 
                           B(11), B(10) => B(10), B(9) => B(9), B(8) => B(8), 
                           B(7) => B(7), B(6) => B(6), B(5) => B(5), B(4) => 
                           B(4), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), O(63) => OTMP_191_port, O(62) => 
                           OTMP_190_port, O(61) => OTMP_189_port, O(60) => 
                           OTMP_188_port, O(59) => OTMP_187_port, O(58) => 
                           OTMP_186_port, O(57) => OTMP_185_port, O(56) => 
                           OTMP_184_port, O(55) => OTMP_183_port, O(54) => 
                           OTMP_182_port, O(53) => OTMP_181_port, O(52) => 
                           OTMP_180_port, O(51) => OTMP_179_port, O(50) => 
                           OTMP_178_port, O(49) => OTMP_177_port, O(48) => 
                           OTMP_176_port, O(47) => OTMP_175_port, O(46) => 
                           OTMP_174_port, O(45) => OTMP_173_port, O(44) => 
                           OTMP_172_port, O(43) => OTMP_171_port, O(42) => 
                           OTMP_170_port, O(41) => OTMP_169_port, O(40) => 
                           OTMP_168_port, O(39) => OTMP_167_port, O(38) => 
                           OTMP_166_port, O(37) => OTMP_165_port, O(36) => 
                           OTMP_164_port, O(35) => OTMP_163_port, O(34) => 
                           OTMP_162_port, O(33) => OTMP_161_port, O(32) => 
                           OTMP_160_port, O(31) => OTMP_159_port, O(30) => 
                           OTMP_158_port, O(29) => OTMP_157_port, O(28) => 
                           OTMP_156_port, O(27) => OTMP_155_port, O(26) => 
                           OTMP_154_port, O(25) => OTMP_153_port, O(24) => 
                           OTMP_152_port, O(23) => OTMP_151_port, O(22) => 
                           OTMP_150_port, O(21) => OTMP_149_port, O(20) => 
                           OTMP_148_port, O(19) => OTMP_147_port, O(18) => 
                           OTMP_146_port, O(17) => OTMP_145_port, O(16) => 
                           OTMP_144_port, O(15) => OTMP_143_port, O(14) => 
                           OTMP_142_port, O(13) => OTMP_141_port, O(12) => 
                           OTMP_140_port, O(11) => OTMP_139_port, O(10) => 
                           OTMP_138_port, O(9) => OTMP_137_port, O(8) => 
                           OTMP_136_port, O(7) => OTMP_135_port, O(6) => 
                           OTMP_134_port, O(5) => OTMP_133_port, O(4) => 
                           OTMP_132_port, O(3) => OTMP_131_port, O(2) => 
                           OTMP_130_port, O(1) => OTMP_129_port, O(0) => n_1101
                           , A_so(63) => SHIFT_255_port, A_so(62) => 
                           SHIFT_254_port, A_so(61) => SHIFT_253_port, A_so(60)
                           => SHIFT_252_port, A_so(59) => SHIFT_251_port, 
                           A_so(58) => SHIFT_250_port, A_so(57) => 
                           SHIFT_249_port, A_so(56) => SHIFT_248_port, A_so(55)
                           => SHIFT_247_port, A_so(54) => SHIFT_246_port, 
                           A_so(53) => SHIFT_245_port, A_so(52) => 
                           SHIFT_244_port, A_so(51) => SHIFT_243_port, A_so(50)
                           => SHIFT_242_port, A_so(49) => SHIFT_241_port, 
                           A_so(48) => SHIFT_240_port, A_so(47) => 
                           SHIFT_239_port, A_so(46) => SHIFT_238_port, A_so(45)
                           => SHIFT_237_port, A_so(44) => SHIFT_236_port, 
                           A_so(43) => SHIFT_235_port, A_so(42) => 
                           SHIFT_234_port, A_so(41) => SHIFT_233_port, A_so(40)
                           => SHIFT_232_port, A_so(39) => SHIFT_231_port, 
                           A_so(38) => SHIFT_230_port, A_so(37) => 
                           SHIFT_229_port, A_so(36) => SHIFT_228_port, A_so(35)
                           => SHIFT_227_port, A_so(34) => SHIFT_226_port, 
                           A_so(33) => SHIFT_225_port, A_so(32) => 
                           SHIFT_224_port, A_so(31) => SHIFT_223_port, A_so(30)
                           => SHIFT_222_port, A_so(29) => SHIFT_221_port, 
                           A_so(28) => SHIFT_220_port, A_so(27) => 
                           SHIFT_219_port, A_so(26) => SHIFT_218_port, A_so(25)
                           => SHIFT_217_port, A_so(24) => SHIFT_216_port, 
                           A_so(23) => SHIFT_215_port, A_so(22) => 
                           SHIFT_214_port, A_so(21) => SHIFT_213_port, A_so(20)
                           => SHIFT_212_port, A_so(19) => SHIFT_211_port, 
                           A_so(18) => SHIFT_210_port, A_so(17) => 
                           SHIFT_209_port, A_so(16) => SHIFT_208_port, A_so(15)
                           => SHIFT_207_port, A_so(14) => SHIFT_206_port, 
                           A_so(13) => SHIFT_205_port, A_so(12) => 
                           SHIFT_204_port, A_so(11) => SHIFT_203_port, A_so(10)
                           => SHIFT_202_port, A_so(9) => SHIFT_201_port, 
                           A_so(8) => SHIFT_200_port, A_so(7) => SHIFT_199_port
                           , A_so(6) => SHIFT_198_port, A_so(5) => 
                           SHIFT_197_port, A_so(4) => SHIFT_196_port, A_so(3) 
                           => SHIFT_195_port, A_so(2) => SHIFT_194_port, 
                           A_so(1) => n_1102, A_so(0) => n_1103, A_nso(63) => 
                           SHIFT_n_255_port, A_nso(62) => SHIFT_n_254_port, 
                           A_nso(61) => SHIFT_n_253_port, A_nso(60) => 
                           SHIFT_n_252_port, A_nso(59) => SHIFT_n_251_port, 
                           A_nso(58) => SHIFT_n_250_port, A_nso(57) => 
                           SHIFT_n_249_port, A_nso(56) => SHIFT_n_248_port, 
                           A_nso(55) => SHIFT_n_247_port, A_nso(54) => 
                           SHIFT_n_246_port, A_nso(53) => SHIFT_n_245_port, 
                           A_nso(52) => SHIFT_n_244_port, A_nso(51) => 
                           SHIFT_n_243_port, A_nso(50) => SHIFT_n_242_port, 
                           A_nso(49) => SHIFT_n_241_port, A_nso(48) => 
                           SHIFT_n_240_port, A_nso(47) => SHIFT_n_239_port, 
                           A_nso(46) => SHIFT_n_238_port, A_nso(45) => 
                           SHIFT_n_237_port, A_nso(44) => SHIFT_n_236_port, 
                           A_nso(43) => SHIFT_n_235_port, A_nso(42) => 
                           SHIFT_n_234_port, A_nso(41) => SHIFT_n_233_port, 
                           A_nso(40) => SHIFT_n_232_port, A_nso(39) => 
                           SHIFT_n_231_port, A_nso(38) => SHIFT_n_230_port, 
                           A_nso(37) => SHIFT_n_229_port, A_nso(36) => 
                           SHIFT_n_228_port, A_nso(35) => SHIFT_n_227_port, 
                           A_nso(34) => SHIFT_n_226_port, A_nso(33) => 
                           SHIFT_n_225_port, A_nso(32) => SHIFT_n_224_port, 
                           A_nso(31) => SHIFT_n_223_port, A_nso(30) => 
                           SHIFT_n_222_port, A_nso(29) => SHIFT_n_221_port, 
                           A_nso(28) => SHIFT_n_220_port, A_nso(27) => 
                           SHIFT_n_219_port, A_nso(26) => SHIFT_n_218_port, 
                           A_nso(25) => SHIFT_n_217_port, A_nso(24) => 
                           SHIFT_n_216_port, A_nso(23) => SHIFT_n_215_port, 
                           A_nso(22) => SHIFT_n_214_port, A_nso(21) => 
                           SHIFT_n_213_port, A_nso(20) => SHIFT_n_212_port, 
                           A_nso(19) => SHIFT_n_211_port, A_nso(18) => 
                           SHIFT_n_210_port, A_nso(17) => SHIFT_n_209_port, 
                           A_nso(16) => SHIFT_n_208_port, A_nso(15) => 
                           SHIFT_n_207_port, A_nso(14) => SHIFT_n_206_port, 
                           A_nso(13) => SHIFT_n_205_port, A_nso(12) => 
                           SHIFT_n_204_port, A_nso(11) => SHIFT_n_203_port, 
                           A_nso(10) => SHIFT_n_202_port, A_nso(9) => 
                           SHIFT_n_201_port, A_nso(8) => SHIFT_n_200_port, 
                           A_nso(7) => SHIFT_n_199_port, A_nso(6) => 
                           SHIFT_n_198_port, A_nso(5) => SHIFT_n_197_port, 
                           A_nso(4) => SHIFT_n_196_port, A_nso(3) => 
                           SHIFT_n_195_port, A_nso(2) => SHIFT_n_194_port, 
                           A_nso(1) => n_1104, A_nso(0) => n_1105);
   BOOTHENC_I_4 : BOOTHENC_NBIT64_i6 port map( A(63) => net48308, A(62) => 
                           net48309, A(61) => net48310, A(60) => net48311, 
                           A(59) => net48312, A(58) => net48313, A(57) => 
                           net48314, A(56) => net48315, A(55) => net48316, 
                           A(54) => net48317, A(53) => net48318, A(52) => 
                           net48319, A(51) => net48320, A(50) => net48321, 
                           A(49) => net48322, A(48) => net48323, A(47) => 
                           net48324, A(46) => net48325, A(45) => net48326, 
                           A(44) => net48327, A(43) => net48328, A(42) => 
                           net48329, A(41) => net48330, A(40) => net48331, 
                           A(39) => net48332, A(38) => net48333, A(37) => 
                           net48334, A(36) => net48335, A(35) => net48336, 
                           A(34) => net48337, A(33) => net48338, A(32) => 
                           net48339, A(31) => net48340, A(30) => net48341, 
                           A(29) => net48342, A(28) => net48343, A(27) => 
                           net48344, A(26) => net48345, A(25) => net48346, 
                           A(24) => net48347, A(23) => net48348, A(22) => 
                           net48349, A(21) => net48350, A(20) => net48351, 
                           A(19) => net48352, A(18) => net48353, A(17) => 
                           net48354, A(16) => net48355, A(15) => net48356, 
                           A(14) => net48357, A(13) => net48358, A(12) => 
                           net48359, A(11) => net48360, A(10) => net48361, A(9)
                           => net48362, A(8) => net48363, A(7) => net48364, 
                           A(6) => net48365, A(5) => net48366, A(4) => net48367
                           , A(3) => net48368, A(2) => net48369, A(1) => 
                           net48370, A(0) => net48371, A_n(63) => net48372, 
                           A_n(62) => net48373, A_n(61) => net48374, A_n(60) =>
                           net48375, A_n(59) => net48376, A_n(58) => net48377, 
                           A_n(57) => net48378, A_n(56) => net48379, A_n(55) =>
                           net48380, A_n(54) => net48381, A_n(53) => net48382, 
                           A_n(52) => net48383, A_n(51) => net48384, A_n(50) =>
                           net48385, A_n(49) => net48386, A_n(48) => net48387, 
                           A_n(47) => net48388, A_n(46) => net48389, A_n(45) =>
                           net48390, A_n(44) => net48391, A_n(43) => net48392, 
                           A_n(42) => net48393, A_n(41) => net48394, A_n(40) =>
                           net48395, A_n(39) => net48396, A_n(38) => net48397, 
                           A_n(37) => net48398, A_n(36) => net48399, A_n(35) =>
                           net48400, A_n(34) => net48401, A_n(33) => net48402, 
                           A_n(32) => net48403, A_n(31) => net48404, A_n(30) =>
                           net48405, A_n(29) => net48406, A_n(28) => net48407, 
                           A_n(27) => net48408, A_n(26) => net48409, A_n(25) =>
                           net48410, A_n(24) => net48411, A_n(23) => net48412, 
                           A_n(22) => net48413, A_n(21) => net48414, A_n(20) =>
                           net48415, A_n(19) => net48416, A_n(18) => net48417, 
                           A_n(17) => net48418, A_n(16) => net48419, A_n(15) =>
                           net48420, A_n(14) => net48421, A_n(13) => net48422, 
                           A_n(12) => net48423, A_n(11) => net48424, A_n(10) =>
                           net48425, A_n(9) => net48426, A_n(8) => net48427, 
                           A_n(7) => net48428, A_n(6) => net48429, A_n(5) => 
                           net48430, A_n(4) => net48431, A_n(3) => net48432, 
                           A_n(2) => net48433, A_n(1) => net48434, A_n(0) => 
                           net48435, A_ns(63) => SHIFT_n_255_port, A_ns(62) => 
                           SHIFT_n_254_port, A_ns(61) => SHIFT_n_253_port, 
                           A_ns(60) => SHIFT_n_252_port, A_ns(59) => 
                           SHIFT_n_251_port, A_ns(58) => SHIFT_n_250_port, 
                           A_ns(57) => SHIFT_n_249_port, A_ns(56) => 
                           SHIFT_n_248_port, A_ns(55) => SHIFT_n_247_port, 
                           A_ns(54) => SHIFT_n_246_port, A_ns(53) => 
                           SHIFT_n_245_port, A_ns(52) => SHIFT_n_244_port, 
                           A_ns(51) => SHIFT_n_243_port, A_ns(50) => 
                           SHIFT_n_242_port, A_ns(49) => SHIFT_n_241_port, 
                           A_ns(48) => SHIFT_n_240_port, A_ns(47) => 
                           SHIFT_n_239_port, A_ns(46) => SHIFT_n_238_port, 
                           A_ns(45) => SHIFT_n_237_port, A_ns(44) => 
                           SHIFT_n_236_port, A_ns(43) => SHIFT_n_235_port, 
                           A_ns(42) => SHIFT_n_234_port, A_ns(41) => 
                           SHIFT_n_233_port, A_ns(40) => SHIFT_n_232_port, 
                           A_ns(39) => SHIFT_n_231_port, A_ns(38) => 
                           SHIFT_n_230_port, A_ns(37) => SHIFT_n_229_port, 
                           A_ns(36) => SHIFT_n_228_port, A_ns(35) => 
                           SHIFT_n_227_port, A_ns(34) => SHIFT_n_226_port, 
                           A_ns(33) => SHIFT_n_225_port, A_ns(32) => 
                           SHIFT_n_224_port, A_ns(31) => SHIFT_n_223_port, 
                           A_ns(30) => SHIFT_n_222_port, A_ns(29) => 
                           SHIFT_n_221_port, A_ns(28) => SHIFT_n_220_port, 
                           A_ns(27) => SHIFT_n_219_port, A_ns(26) => 
                           SHIFT_n_218_port, A_ns(25) => SHIFT_n_217_port, 
                           A_ns(24) => SHIFT_n_216_port, A_ns(23) => 
                           SHIFT_n_215_port, A_ns(22) => SHIFT_n_214_port, 
                           A_ns(21) => SHIFT_n_213_port, A_ns(20) => 
                           SHIFT_n_212_port, A_ns(19) => SHIFT_n_211_port, 
                           A_ns(18) => SHIFT_n_210_port, A_ns(17) => 
                           SHIFT_n_209_port, A_ns(16) => SHIFT_n_208_port, 
                           A_ns(15) => SHIFT_n_207_port, A_ns(14) => 
                           SHIFT_n_206_port, A_ns(13) => SHIFT_n_205_port, 
                           A_ns(12) => SHIFT_n_204_port, A_ns(11) => 
                           SHIFT_n_203_port, A_ns(10) => SHIFT_n_202_port, 
                           A_ns(9) => SHIFT_n_201_port, A_ns(8) => 
                           SHIFT_n_200_port, A_ns(7) => SHIFT_n_199_port, 
                           A_ns(6) => SHIFT_n_198_port, A_ns(5) => 
                           SHIFT_n_197_port, A_ns(4) => SHIFT_n_196_port, 
                           A_ns(3) => SHIFT_n_195_port, A_ns(2) => 
                           SHIFT_n_194_port, A_ns(1) => SHIFT_n_193_port, 
                           A_ns(0) => SHIFT_n_192_port, A_s(63) => 
                           SHIFT_255_port, A_s(62) => SHIFT_254_port, A_s(61) 
                           => SHIFT_253_port, A_s(60) => SHIFT_252_port, 
                           A_s(59) => SHIFT_251_port, A_s(58) => SHIFT_250_port
                           , A_s(57) => SHIFT_249_port, A_s(56) => 
                           SHIFT_248_port, A_s(55) => SHIFT_247_port, A_s(54) 
                           => SHIFT_246_port, A_s(53) => SHIFT_245_port, 
                           A_s(52) => SHIFT_244_port, A_s(51) => SHIFT_243_port
                           , A_s(50) => SHIFT_242_port, A_s(49) => 
                           SHIFT_241_port, A_s(48) => SHIFT_240_port, A_s(47) 
                           => SHIFT_239_port, A_s(46) => SHIFT_238_port, 
                           A_s(45) => SHIFT_237_port, A_s(44) => SHIFT_236_port
                           , A_s(43) => SHIFT_235_port, A_s(42) => 
                           SHIFT_234_port, A_s(41) => SHIFT_233_port, A_s(40) 
                           => SHIFT_232_port, A_s(39) => SHIFT_231_port, 
                           A_s(38) => SHIFT_230_port, A_s(37) => SHIFT_229_port
                           , A_s(36) => SHIFT_228_port, A_s(35) => 
                           SHIFT_227_port, A_s(34) => SHIFT_226_port, A_s(33) 
                           => SHIFT_225_port, A_s(32) => SHIFT_224_port, 
                           A_s(31) => SHIFT_223_port, A_s(30) => SHIFT_222_port
                           , A_s(29) => SHIFT_221_port, A_s(28) => 
                           SHIFT_220_port, A_s(27) => SHIFT_219_port, A_s(26) 
                           => SHIFT_218_port, A_s(25) => SHIFT_217_port, 
                           A_s(24) => SHIFT_216_port, A_s(23) => SHIFT_215_port
                           , A_s(22) => SHIFT_214_port, A_s(21) => 
                           SHIFT_213_port, A_s(20) => SHIFT_212_port, A_s(19) 
                           => SHIFT_211_port, A_s(18) => SHIFT_210_port, 
                           A_s(17) => SHIFT_209_port, A_s(16) => SHIFT_208_port
                           , A_s(15) => SHIFT_207_port, A_s(14) => 
                           SHIFT_206_port, A_s(13) => SHIFT_205_port, A_s(12) 
                           => SHIFT_204_port, A_s(11) => SHIFT_203_port, 
                           A_s(10) => SHIFT_202_port, A_s(9) => SHIFT_201_port,
                           A_s(8) => SHIFT_200_port, A_s(7) => SHIFT_199_port, 
                           A_s(6) => SHIFT_198_port, A_s(5) => SHIFT_197_port, 
                           A_s(4) => SHIFT_196_port, A_s(3) => SHIFT_195_port, 
                           A_s(2) => SHIFT_194_port, A_s(1) => SHIFT_193_port, 
                           A_s(0) => SHIFT_192_port, B(63) => B(31), B(62) => 
                           B(31), B(61) => B(31), B(60) => B(31), B(59) => 
                           B(31), B(58) => B(31), B(57) => B(31), B(56) => 
                           B(31), B(55) => B(31), B(54) => B(31), B(53) => 
                           B(31), B(52) => B(31), B(51) => B(31), B(50) => 
                           B(31), B(49) => B(31), B(48) => B(31), B(47) => 
                           B(31), B(46) => B(31), B(45) => B(31), B(44) => 
                           B(31), B(43) => B(31), B(42) => B(31), B(41) => 
                           B(31), B(40) => B(31), B(39) => B(31), B(38) => 
                           B(31), B(37) => B(31), B(36) => B(31), B(35) => 
                           B(31), B(34) => B(31), B(33) => B(31), B(32) => 
                           B(31), B(31) => B(31), B(30) => B(30), B(29) => 
                           B(29), B(28) => B(28), B(27) => B(27), B(26) => 
                           B(26), B(25) => B(25), B(24) => B(24), B(23) => 
                           B(23), B(22) => B(22), B(21) => B(21), B(20) => 
                           B(20), B(19) => B(19), B(18) => B(18), B(17) => 
                           B(17), B(16) => B(16), B(15) => B(15), B(14) => 
                           B(14), B(13) => B(13), B(12) => B(12), B(11) => 
                           B(11), B(10) => B(10), B(9) => B(9), B(8) => B(8), 
                           B(7) => B(7), B(6) => B(6), B(5) => B(5), B(4) => 
                           B(4), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), O(63) => OTMP_255_port, O(62) => 
                           OTMP_254_port, O(61) => OTMP_253_port, O(60) => 
                           OTMP_252_port, O(59) => OTMP_251_port, O(58) => 
                           OTMP_250_port, O(57) => OTMP_249_port, O(56) => 
                           OTMP_248_port, O(55) => OTMP_247_port, O(54) => 
                           OTMP_246_port, O(53) => OTMP_245_port, O(52) => 
                           OTMP_244_port, O(51) => OTMP_243_port, O(50) => 
                           OTMP_242_port, O(49) => OTMP_241_port, O(48) => 
                           OTMP_240_port, O(47) => OTMP_239_port, O(46) => 
                           OTMP_238_port, O(45) => OTMP_237_port, O(44) => 
                           OTMP_236_port, O(43) => OTMP_235_port, O(42) => 
                           OTMP_234_port, O(41) => OTMP_233_port, O(40) => 
                           OTMP_232_port, O(39) => OTMP_231_port, O(38) => 
                           OTMP_230_port, O(37) => OTMP_229_port, O(36) => 
                           OTMP_228_port, O(35) => OTMP_227_port, O(34) => 
                           OTMP_226_port, O(33) => OTMP_225_port, O(32) => 
                           OTMP_224_port, O(31) => OTMP_223_port, O(30) => 
                           OTMP_222_port, O(29) => OTMP_221_port, O(28) => 
                           OTMP_220_port, O(27) => OTMP_219_port, O(26) => 
                           OTMP_218_port, O(25) => OTMP_217_port, O(24) => 
                           OTMP_216_port, O(23) => OTMP_215_port, O(22) => 
                           OTMP_214_port, O(21) => OTMP_213_port, O(20) => 
                           OTMP_212_port, O(19) => OTMP_211_port, O(18) => 
                           OTMP_210_port, O(17) => OTMP_209_port, O(16) => 
                           OTMP_208_port, O(15) => OTMP_207_port, O(14) => 
                           OTMP_206_port, O(13) => OTMP_205_port, O(12) => 
                           OTMP_204_port, O(11) => OTMP_203_port, O(10) => 
                           OTMP_202_port, O(9) => OTMP_201_port, O(8) => 
                           OTMP_200_port, O(7) => OTMP_199_port, O(6) => 
                           OTMP_198_port, O(5) => OTMP_197_port, O(4) => 
                           OTMP_196_port, O(3) => OTMP_195_port, O(2) => 
                           OTMP_194_port, O(1) => OTMP_193_port, O(0) => n_1106
                           , A_so(63) => SHIFT_319_port, A_so(62) => 
                           SHIFT_318_port, A_so(61) => SHIFT_317_port, A_so(60)
                           => SHIFT_316_port, A_so(59) => SHIFT_315_port, 
                           A_so(58) => SHIFT_314_port, A_so(57) => 
                           SHIFT_313_port, A_so(56) => SHIFT_312_port, A_so(55)
                           => SHIFT_311_port, A_so(54) => SHIFT_310_port, 
                           A_so(53) => SHIFT_309_port, A_so(52) => 
                           SHIFT_308_port, A_so(51) => SHIFT_307_port, A_so(50)
                           => SHIFT_306_port, A_so(49) => SHIFT_305_port, 
                           A_so(48) => SHIFT_304_port, A_so(47) => 
                           SHIFT_303_port, A_so(46) => SHIFT_302_port, A_so(45)
                           => SHIFT_301_port, A_so(44) => SHIFT_300_port, 
                           A_so(43) => SHIFT_299_port, A_so(42) => 
                           SHIFT_298_port, A_so(41) => SHIFT_297_port, A_so(40)
                           => SHIFT_296_port, A_so(39) => SHIFT_295_port, 
                           A_so(38) => SHIFT_294_port, A_so(37) => 
                           SHIFT_293_port, A_so(36) => SHIFT_292_port, A_so(35)
                           => SHIFT_291_port, A_so(34) => SHIFT_290_port, 
                           A_so(33) => SHIFT_289_port, A_so(32) => 
                           SHIFT_288_port, A_so(31) => SHIFT_287_port, A_so(30)
                           => SHIFT_286_port, A_so(29) => SHIFT_285_port, 
                           A_so(28) => SHIFT_284_port, A_so(27) => 
                           SHIFT_283_port, A_so(26) => SHIFT_282_port, A_so(25)
                           => SHIFT_281_port, A_so(24) => SHIFT_280_port, 
                           A_so(23) => SHIFT_279_port, A_so(22) => 
                           SHIFT_278_port, A_so(21) => SHIFT_277_port, A_so(20)
                           => SHIFT_276_port, A_so(19) => SHIFT_275_port, 
                           A_so(18) => SHIFT_274_port, A_so(17) => 
                           SHIFT_273_port, A_so(16) => SHIFT_272_port, A_so(15)
                           => SHIFT_271_port, A_so(14) => SHIFT_270_port, 
                           A_so(13) => SHIFT_269_port, A_so(12) => 
                           SHIFT_268_port, A_so(11) => SHIFT_267_port, A_so(10)
                           => SHIFT_266_port, A_so(9) => SHIFT_265_port, 
                           A_so(8) => SHIFT_264_port, A_so(7) => SHIFT_263_port
                           , A_so(6) => SHIFT_262_port, A_so(5) => 
                           SHIFT_261_port, A_so(4) => SHIFT_260_port, A_so(3) 
                           => SHIFT_259_port, A_so(2) => SHIFT_258_port, 
                           A_so(1) => n_1107, A_so(0) => n_1108, A_nso(63) => 
                           SHIFT_n_319_port, A_nso(62) => SHIFT_n_318_port, 
                           A_nso(61) => SHIFT_n_317_port, A_nso(60) => 
                           SHIFT_n_316_port, A_nso(59) => SHIFT_n_315_port, 
                           A_nso(58) => SHIFT_n_314_port, A_nso(57) => 
                           SHIFT_n_313_port, A_nso(56) => SHIFT_n_312_port, 
                           A_nso(55) => SHIFT_n_311_port, A_nso(54) => 
                           SHIFT_n_310_port, A_nso(53) => SHIFT_n_309_port, 
                           A_nso(52) => SHIFT_n_308_port, A_nso(51) => 
                           SHIFT_n_307_port, A_nso(50) => SHIFT_n_306_port, 
                           A_nso(49) => SHIFT_n_305_port, A_nso(48) => 
                           SHIFT_n_304_port, A_nso(47) => SHIFT_n_303_port, 
                           A_nso(46) => SHIFT_n_302_port, A_nso(45) => 
                           SHIFT_n_301_port, A_nso(44) => SHIFT_n_300_port, 
                           A_nso(43) => SHIFT_n_299_port, A_nso(42) => 
                           SHIFT_n_298_port, A_nso(41) => SHIFT_n_297_port, 
                           A_nso(40) => SHIFT_n_296_port, A_nso(39) => 
                           SHIFT_n_295_port, A_nso(38) => SHIFT_n_294_port, 
                           A_nso(37) => SHIFT_n_293_port, A_nso(36) => 
                           SHIFT_n_292_port, A_nso(35) => SHIFT_n_291_port, 
                           A_nso(34) => SHIFT_n_290_port, A_nso(33) => 
                           SHIFT_n_289_port, A_nso(32) => SHIFT_n_288_port, 
                           A_nso(31) => SHIFT_n_287_port, A_nso(30) => 
                           SHIFT_n_286_port, A_nso(29) => SHIFT_n_285_port, 
                           A_nso(28) => SHIFT_n_284_port, A_nso(27) => 
                           SHIFT_n_283_port, A_nso(26) => SHIFT_n_282_port, 
                           A_nso(25) => SHIFT_n_281_port, A_nso(24) => 
                           SHIFT_n_280_port, A_nso(23) => SHIFT_n_279_port, 
                           A_nso(22) => SHIFT_n_278_port, A_nso(21) => 
                           SHIFT_n_277_port, A_nso(20) => SHIFT_n_276_port, 
                           A_nso(19) => SHIFT_n_275_port, A_nso(18) => 
                           SHIFT_n_274_port, A_nso(17) => SHIFT_n_273_port, 
                           A_nso(16) => SHIFT_n_272_port, A_nso(15) => 
                           SHIFT_n_271_port, A_nso(14) => SHIFT_n_270_port, 
                           A_nso(13) => SHIFT_n_269_port, A_nso(12) => 
                           SHIFT_n_268_port, A_nso(11) => SHIFT_n_267_port, 
                           A_nso(10) => SHIFT_n_266_port, A_nso(9) => 
                           SHIFT_n_265_port, A_nso(8) => SHIFT_n_264_port, 
                           A_nso(7) => SHIFT_n_263_port, A_nso(6) => 
                           SHIFT_n_262_port, A_nso(5) => SHIFT_n_261_port, 
                           A_nso(4) => SHIFT_n_260_port, A_nso(3) => 
                           SHIFT_n_259_port, A_nso(2) => SHIFT_n_258_port, 
                           A_nso(1) => n_1109, A_nso(0) => n_1110);
   BOOTHENC_I_5 : BOOTHENC_NBIT64_i8 port map( A(63) => net48180, A(62) => 
                           net48181, A(61) => net48182, A(60) => net48183, 
                           A(59) => net48184, A(58) => net48185, A(57) => 
                           net48186, A(56) => net48187, A(55) => net48188, 
                           A(54) => net48189, A(53) => net48190, A(52) => 
                           net48191, A(51) => net48192, A(50) => net48193, 
                           A(49) => net48194, A(48) => net48195, A(47) => 
                           net48196, A(46) => net48197, A(45) => net48198, 
                           A(44) => net48199, A(43) => net48200, A(42) => 
                           net48201, A(41) => net48202, A(40) => net48203, 
                           A(39) => net48204, A(38) => net48205, A(37) => 
                           net48206, A(36) => net48207, A(35) => net48208, 
                           A(34) => net48209, A(33) => net48210, A(32) => 
                           net48211, A(31) => net48212, A(30) => net48213, 
                           A(29) => net48214, A(28) => net48215, A(27) => 
                           net48216, A(26) => net48217, A(25) => net48218, 
                           A(24) => net48219, A(23) => net48220, A(22) => 
                           net48221, A(21) => net48222, A(20) => net48223, 
                           A(19) => net48224, A(18) => net48225, A(17) => 
                           net48226, A(16) => net48227, A(15) => net48228, 
                           A(14) => net48229, A(13) => net48230, A(12) => 
                           net48231, A(11) => net48232, A(10) => net48233, A(9)
                           => net48234, A(8) => net48235, A(7) => net48236, 
                           A(6) => net48237, A(5) => net48238, A(4) => net48239
                           , A(3) => net48240, A(2) => net48241, A(1) => 
                           net48242, A(0) => net48243, A_n(63) => net48244, 
                           A_n(62) => net48245, A_n(61) => net48246, A_n(60) =>
                           net48247, A_n(59) => net48248, A_n(58) => net48249, 
                           A_n(57) => net48250, A_n(56) => net48251, A_n(55) =>
                           net48252, A_n(54) => net48253, A_n(53) => net48254, 
                           A_n(52) => net48255, A_n(51) => net48256, A_n(50) =>
                           net48257, A_n(49) => net48258, A_n(48) => net48259, 
                           A_n(47) => net48260, A_n(46) => net48261, A_n(45) =>
                           net48262, A_n(44) => net48263, A_n(43) => net48264, 
                           A_n(42) => net48265, A_n(41) => net48266, A_n(40) =>
                           net48267, A_n(39) => net48268, A_n(38) => net48269, 
                           A_n(37) => net48270, A_n(36) => net48271, A_n(35) =>
                           net48272, A_n(34) => net48273, A_n(33) => net48274, 
                           A_n(32) => net48275, A_n(31) => net48276, A_n(30) =>
                           net48277, A_n(29) => net48278, A_n(28) => net48279, 
                           A_n(27) => net48280, A_n(26) => net48281, A_n(25) =>
                           net48282, A_n(24) => net48283, A_n(23) => net48284, 
                           A_n(22) => net48285, A_n(21) => net48286, A_n(20) =>
                           net48287, A_n(19) => net48288, A_n(18) => net48289, 
                           A_n(17) => net48290, A_n(16) => net48291, A_n(15) =>
                           net48292, A_n(14) => net48293, A_n(13) => net48294, 
                           A_n(12) => net48295, A_n(11) => net48296, A_n(10) =>
                           net48297, A_n(9) => net48298, A_n(8) => net48299, 
                           A_n(7) => net48300, A_n(6) => net48301, A_n(5) => 
                           net48302, A_n(4) => net48303, A_n(3) => net48304, 
                           A_n(2) => net48305, A_n(1) => net48306, A_n(0) => 
                           net48307, A_ns(63) => SHIFT_n_319_port, A_ns(62) => 
                           SHIFT_n_318_port, A_ns(61) => SHIFT_n_317_port, 
                           A_ns(60) => SHIFT_n_316_port, A_ns(59) => 
                           SHIFT_n_315_port, A_ns(58) => SHIFT_n_314_port, 
                           A_ns(57) => SHIFT_n_313_port, A_ns(56) => 
                           SHIFT_n_312_port, A_ns(55) => SHIFT_n_311_port, 
                           A_ns(54) => SHIFT_n_310_port, A_ns(53) => 
                           SHIFT_n_309_port, A_ns(52) => SHIFT_n_308_port, 
                           A_ns(51) => SHIFT_n_307_port, A_ns(50) => 
                           SHIFT_n_306_port, A_ns(49) => SHIFT_n_305_port, 
                           A_ns(48) => SHIFT_n_304_port, A_ns(47) => 
                           SHIFT_n_303_port, A_ns(46) => SHIFT_n_302_port, 
                           A_ns(45) => SHIFT_n_301_port, A_ns(44) => 
                           SHIFT_n_300_port, A_ns(43) => SHIFT_n_299_port, 
                           A_ns(42) => SHIFT_n_298_port, A_ns(41) => 
                           SHIFT_n_297_port, A_ns(40) => SHIFT_n_296_port, 
                           A_ns(39) => SHIFT_n_295_port, A_ns(38) => 
                           SHIFT_n_294_port, A_ns(37) => SHIFT_n_293_port, 
                           A_ns(36) => SHIFT_n_292_port, A_ns(35) => 
                           SHIFT_n_291_port, A_ns(34) => SHIFT_n_290_port, 
                           A_ns(33) => SHIFT_n_289_port, A_ns(32) => 
                           SHIFT_n_288_port, A_ns(31) => SHIFT_n_287_port, 
                           A_ns(30) => SHIFT_n_286_port, A_ns(29) => 
                           SHIFT_n_285_port, A_ns(28) => SHIFT_n_284_port, 
                           A_ns(27) => SHIFT_n_283_port, A_ns(26) => 
                           SHIFT_n_282_port, A_ns(25) => SHIFT_n_281_port, 
                           A_ns(24) => SHIFT_n_280_port, A_ns(23) => 
                           SHIFT_n_279_port, A_ns(22) => SHIFT_n_278_port, 
                           A_ns(21) => SHIFT_n_277_port, A_ns(20) => 
                           SHIFT_n_276_port, A_ns(19) => SHIFT_n_275_port, 
                           A_ns(18) => SHIFT_n_274_port, A_ns(17) => 
                           SHIFT_n_273_port, A_ns(16) => SHIFT_n_272_port, 
                           A_ns(15) => SHIFT_n_271_port, A_ns(14) => 
                           SHIFT_n_270_port, A_ns(13) => SHIFT_n_269_port, 
                           A_ns(12) => SHIFT_n_268_port, A_ns(11) => 
                           SHIFT_n_267_port, A_ns(10) => SHIFT_n_266_port, 
                           A_ns(9) => SHIFT_n_265_port, A_ns(8) => 
                           SHIFT_n_264_port, A_ns(7) => SHIFT_n_263_port, 
                           A_ns(6) => SHIFT_n_262_port, A_ns(5) => 
                           SHIFT_n_261_port, A_ns(4) => SHIFT_n_260_port, 
                           A_ns(3) => SHIFT_n_259_port, A_ns(2) => 
                           SHIFT_n_258_port, A_ns(1) => SHIFT_n_257_port, 
                           A_ns(0) => SHIFT_n_256_port, A_s(63) => 
                           SHIFT_319_port, A_s(62) => SHIFT_318_port, A_s(61) 
                           => SHIFT_317_port, A_s(60) => SHIFT_316_port, 
                           A_s(59) => SHIFT_315_port, A_s(58) => SHIFT_314_port
                           , A_s(57) => SHIFT_313_port, A_s(56) => 
                           SHIFT_312_port, A_s(55) => SHIFT_311_port, A_s(54) 
                           => SHIFT_310_port, A_s(53) => SHIFT_309_port, 
                           A_s(52) => SHIFT_308_port, A_s(51) => SHIFT_307_port
                           , A_s(50) => SHIFT_306_port, A_s(49) => 
                           SHIFT_305_port, A_s(48) => SHIFT_304_port, A_s(47) 
                           => SHIFT_303_port, A_s(46) => SHIFT_302_port, 
                           A_s(45) => SHIFT_301_port, A_s(44) => SHIFT_300_port
                           , A_s(43) => SHIFT_299_port, A_s(42) => 
                           SHIFT_298_port, A_s(41) => SHIFT_297_port, A_s(40) 
                           => SHIFT_296_port, A_s(39) => SHIFT_295_port, 
                           A_s(38) => SHIFT_294_port, A_s(37) => SHIFT_293_port
                           , A_s(36) => SHIFT_292_port, A_s(35) => 
                           SHIFT_291_port, A_s(34) => SHIFT_290_port, A_s(33) 
                           => SHIFT_289_port, A_s(32) => SHIFT_288_port, 
                           A_s(31) => SHIFT_287_port, A_s(30) => SHIFT_286_port
                           , A_s(29) => SHIFT_285_port, A_s(28) => 
                           SHIFT_284_port, A_s(27) => SHIFT_283_port, A_s(26) 
                           => SHIFT_282_port, A_s(25) => SHIFT_281_port, 
                           A_s(24) => SHIFT_280_port, A_s(23) => SHIFT_279_port
                           , A_s(22) => SHIFT_278_port, A_s(21) => 
                           SHIFT_277_port, A_s(20) => SHIFT_276_port, A_s(19) 
                           => SHIFT_275_port, A_s(18) => SHIFT_274_port, 
                           A_s(17) => SHIFT_273_port, A_s(16) => SHIFT_272_port
                           , A_s(15) => SHIFT_271_port, A_s(14) => 
                           SHIFT_270_port, A_s(13) => SHIFT_269_port, A_s(12) 
                           => SHIFT_268_port, A_s(11) => SHIFT_267_port, 
                           A_s(10) => SHIFT_266_port, A_s(9) => SHIFT_265_port,
                           A_s(8) => SHIFT_264_port, A_s(7) => SHIFT_263_port, 
                           A_s(6) => SHIFT_262_port, A_s(5) => SHIFT_261_port, 
                           A_s(4) => SHIFT_260_port, A_s(3) => SHIFT_259_port, 
                           A_s(2) => SHIFT_258_port, A_s(1) => SHIFT_257_port, 
                           A_s(0) => SHIFT_256_port, B(63) => B(31), B(62) => 
                           B(31), B(61) => B(31), B(60) => B(31), B(59) => 
                           B(31), B(58) => B(31), B(57) => B(31), B(56) => 
                           B(31), B(55) => B(31), B(54) => B(31), B(53) => 
                           B(31), B(52) => B(31), B(51) => B(31), B(50) => 
                           B(31), B(49) => B(31), B(48) => B(31), B(47) => 
                           B(31), B(46) => B(31), B(45) => B(31), B(44) => 
                           B(31), B(43) => B(31), B(42) => B(31), B(41) => 
                           B(31), B(40) => B(31), B(39) => B(31), B(38) => 
                           B(31), B(37) => B(31), B(36) => B(31), B(35) => 
                           B(31), B(34) => B(31), B(33) => B(31), B(32) => 
                           B(31), B(31) => B(31), B(30) => B(30), B(29) => 
                           B(29), B(28) => B(28), B(27) => B(27), B(26) => 
                           B(26), B(25) => B(25), B(24) => B(24), B(23) => 
                           B(23), B(22) => B(22), B(21) => B(21), B(20) => 
                           B(20), B(19) => B(19), B(18) => B(18), B(17) => 
                           B(17), B(16) => B(16), B(15) => B(15), B(14) => 
                           B(14), B(13) => B(13), B(12) => B(12), B(11) => 
                           B(11), B(10) => B(10), B(9) => B(9), B(8) => B(8), 
                           B(7) => B(7), B(6) => B(6), B(5) => B(5), B(4) => 
                           B(4), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), O(63) => OTMP_319_port, O(62) => 
                           OTMP_318_port, O(61) => OTMP_317_port, O(60) => 
                           OTMP_316_port, O(59) => OTMP_315_port, O(58) => 
                           OTMP_314_port, O(57) => OTMP_313_port, O(56) => 
                           OTMP_312_port, O(55) => OTMP_311_port, O(54) => 
                           OTMP_310_port, O(53) => OTMP_309_port, O(52) => 
                           OTMP_308_port, O(51) => OTMP_307_port, O(50) => 
                           OTMP_306_port, O(49) => OTMP_305_port, O(48) => 
                           OTMP_304_port, O(47) => OTMP_303_port, O(46) => 
                           OTMP_302_port, O(45) => OTMP_301_port, O(44) => 
                           OTMP_300_port, O(43) => OTMP_299_port, O(42) => 
                           OTMP_298_port, O(41) => OTMP_297_port, O(40) => 
                           OTMP_296_port, O(39) => OTMP_295_port, O(38) => 
                           OTMP_294_port, O(37) => OTMP_293_port, O(36) => 
                           OTMP_292_port, O(35) => OTMP_291_port, O(34) => 
                           OTMP_290_port, O(33) => OTMP_289_port, O(32) => 
                           OTMP_288_port, O(31) => OTMP_287_port, O(30) => 
                           OTMP_286_port, O(29) => OTMP_285_port, O(28) => 
                           OTMP_284_port, O(27) => OTMP_283_port, O(26) => 
                           OTMP_282_port, O(25) => OTMP_281_port, O(24) => 
                           OTMP_280_port, O(23) => OTMP_279_port, O(22) => 
                           OTMP_278_port, O(21) => OTMP_277_port, O(20) => 
                           OTMP_276_port, O(19) => OTMP_275_port, O(18) => 
                           OTMP_274_port, O(17) => OTMP_273_port, O(16) => 
                           OTMP_272_port, O(15) => OTMP_271_port, O(14) => 
                           OTMP_270_port, O(13) => OTMP_269_port, O(12) => 
                           OTMP_268_port, O(11) => OTMP_267_port, O(10) => 
                           OTMP_266_port, O(9) => OTMP_265_port, O(8) => 
                           OTMP_264_port, O(7) => OTMP_263_port, O(6) => 
                           OTMP_262_port, O(5) => OTMP_261_port, O(4) => 
                           OTMP_260_port, O(3) => OTMP_259_port, O(2) => 
                           OTMP_258_port, O(1) => OTMP_257_port, O(0) => n_1111
                           , A_so(63) => SHIFT_383_port, A_so(62) => 
                           SHIFT_382_port, A_so(61) => SHIFT_381_port, A_so(60)
                           => SHIFT_380_port, A_so(59) => SHIFT_379_port, 
                           A_so(58) => SHIFT_378_port, A_so(57) => 
                           SHIFT_377_port, A_so(56) => SHIFT_376_port, A_so(55)
                           => SHIFT_375_port, A_so(54) => SHIFT_374_port, 
                           A_so(53) => SHIFT_373_port, A_so(52) => 
                           SHIFT_372_port, A_so(51) => SHIFT_371_port, A_so(50)
                           => SHIFT_370_port, A_so(49) => SHIFT_369_port, 
                           A_so(48) => SHIFT_368_port, A_so(47) => 
                           SHIFT_367_port, A_so(46) => SHIFT_366_port, A_so(45)
                           => SHIFT_365_port, A_so(44) => SHIFT_364_port, 
                           A_so(43) => SHIFT_363_port, A_so(42) => 
                           SHIFT_362_port, A_so(41) => SHIFT_361_port, A_so(40)
                           => SHIFT_360_port, A_so(39) => SHIFT_359_port, 
                           A_so(38) => SHIFT_358_port, A_so(37) => 
                           SHIFT_357_port, A_so(36) => SHIFT_356_port, A_so(35)
                           => SHIFT_355_port, A_so(34) => SHIFT_354_port, 
                           A_so(33) => SHIFT_353_port, A_so(32) => 
                           SHIFT_352_port, A_so(31) => SHIFT_351_port, A_so(30)
                           => SHIFT_350_port, A_so(29) => SHIFT_349_port, 
                           A_so(28) => SHIFT_348_port, A_so(27) => 
                           SHIFT_347_port, A_so(26) => SHIFT_346_port, A_so(25)
                           => SHIFT_345_port, A_so(24) => SHIFT_344_port, 
                           A_so(23) => SHIFT_343_port, A_so(22) => 
                           SHIFT_342_port, A_so(21) => SHIFT_341_port, A_so(20)
                           => SHIFT_340_port, A_so(19) => SHIFT_339_port, 
                           A_so(18) => SHIFT_338_port, A_so(17) => 
                           SHIFT_337_port, A_so(16) => SHIFT_336_port, A_so(15)
                           => SHIFT_335_port, A_so(14) => SHIFT_334_port, 
                           A_so(13) => SHIFT_333_port, A_so(12) => 
                           SHIFT_332_port, A_so(11) => SHIFT_331_port, A_so(10)
                           => SHIFT_330_port, A_so(9) => SHIFT_329_port, 
                           A_so(8) => SHIFT_328_port, A_so(7) => SHIFT_327_port
                           , A_so(6) => SHIFT_326_port, A_so(5) => 
                           SHIFT_325_port, A_so(4) => SHIFT_324_port, A_so(3) 
                           => SHIFT_323_port, A_so(2) => SHIFT_322_port, 
                           A_so(1) => n_1112, A_so(0) => n_1113, A_nso(63) => 
                           SHIFT_n_383_port, A_nso(62) => SHIFT_n_382_port, 
                           A_nso(61) => SHIFT_n_381_port, A_nso(60) => 
                           SHIFT_n_380_port, A_nso(59) => SHIFT_n_379_port, 
                           A_nso(58) => SHIFT_n_378_port, A_nso(57) => 
                           SHIFT_n_377_port, A_nso(56) => SHIFT_n_376_port, 
                           A_nso(55) => SHIFT_n_375_port, A_nso(54) => 
                           SHIFT_n_374_port, A_nso(53) => SHIFT_n_373_port, 
                           A_nso(52) => SHIFT_n_372_port, A_nso(51) => 
                           SHIFT_n_371_port, A_nso(50) => SHIFT_n_370_port, 
                           A_nso(49) => SHIFT_n_369_port, A_nso(48) => 
                           SHIFT_n_368_port, A_nso(47) => SHIFT_n_367_port, 
                           A_nso(46) => SHIFT_n_366_port, A_nso(45) => 
                           SHIFT_n_365_port, A_nso(44) => SHIFT_n_364_port, 
                           A_nso(43) => SHIFT_n_363_port, A_nso(42) => 
                           SHIFT_n_362_port, A_nso(41) => SHIFT_n_361_port, 
                           A_nso(40) => SHIFT_n_360_port, A_nso(39) => 
                           SHIFT_n_359_port, A_nso(38) => SHIFT_n_358_port, 
                           A_nso(37) => SHIFT_n_357_port, A_nso(36) => 
                           SHIFT_n_356_port, A_nso(35) => SHIFT_n_355_port, 
                           A_nso(34) => SHIFT_n_354_port, A_nso(33) => 
                           SHIFT_n_353_port, A_nso(32) => SHIFT_n_352_port, 
                           A_nso(31) => SHIFT_n_351_port, A_nso(30) => 
                           SHIFT_n_350_port, A_nso(29) => SHIFT_n_349_port, 
                           A_nso(28) => SHIFT_n_348_port, A_nso(27) => 
                           SHIFT_n_347_port, A_nso(26) => SHIFT_n_346_port, 
                           A_nso(25) => SHIFT_n_345_port, A_nso(24) => 
                           SHIFT_n_344_port, A_nso(23) => SHIFT_n_343_port, 
                           A_nso(22) => SHIFT_n_342_port, A_nso(21) => 
                           SHIFT_n_341_port, A_nso(20) => SHIFT_n_340_port, 
                           A_nso(19) => SHIFT_n_339_port, A_nso(18) => 
                           SHIFT_n_338_port, A_nso(17) => SHIFT_n_337_port, 
                           A_nso(16) => SHIFT_n_336_port, A_nso(15) => 
                           SHIFT_n_335_port, A_nso(14) => SHIFT_n_334_port, 
                           A_nso(13) => SHIFT_n_333_port, A_nso(12) => 
                           SHIFT_n_332_port, A_nso(11) => SHIFT_n_331_port, 
                           A_nso(10) => SHIFT_n_330_port, A_nso(9) => 
                           SHIFT_n_329_port, A_nso(8) => SHIFT_n_328_port, 
                           A_nso(7) => SHIFT_n_327_port, A_nso(6) => 
                           SHIFT_n_326_port, A_nso(5) => SHIFT_n_325_port, 
                           A_nso(4) => SHIFT_n_324_port, A_nso(3) => 
                           SHIFT_n_323_port, A_nso(2) => SHIFT_n_322_port, 
                           A_nso(1) => n_1114, A_nso(0) => n_1115);
   BOOTHENC_I_6 : BOOTHENC_NBIT64_i10 port map( A(63) => net48052, A(62) => 
                           net48053, A(61) => net48054, A(60) => net48055, 
                           A(59) => net48056, A(58) => net48057, A(57) => 
                           net48058, A(56) => net48059, A(55) => net48060, 
                           A(54) => net48061, A(53) => net48062, A(52) => 
                           net48063, A(51) => net48064, A(50) => net48065, 
                           A(49) => net48066, A(48) => net48067, A(47) => 
                           net48068, A(46) => net48069, A(45) => net48070, 
                           A(44) => net48071, A(43) => net48072, A(42) => 
                           net48073, A(41) => net48074, A(40) => net48075, 
                           A(39) => net48076, A(38) => net48077, A(37) => 
                           net48078, A(36) => net48079, A(35) => net48080, 
                           A(34) => net48081, A(33) => net48082, A(32) => 
                           net48083, A(31) => net48084, A(30) => net48085, 
                           A(29) => net48086, A(28) => net48087, A(27) => 
                           net48088, A(26) => net48089, A(25) => net48090, 
                           A(24) => net48091, A(23) => net48092, A(22) => 
                           net48093, A(21) => net48094, A(20) => net48095, 
                           A(19) => net48096, A(18) => net48097, A(17) => 
                           net48098, A(16) => net48099, A(15) => net48100, 
                           A(14) => net48101, A(13) => net48102, A(12) => 
                           net48103, A(11) => net48104, A(10) => net48105, A(9)
                           => net48106, A(8) => net48107, A(7) => net48108, 
                           A(6) => net48109, A(5) => net48110, A(4) => net48111
                           , A(3) => net48112, A(2) => net48113, A(1) => 
                           net48114, A(0) => net48115, A_n(63) => net48116, 
                           A_n(62) => net48117, A_n(61) => net48118, A_n(60) =>
                           net48119, A_n(59) => net48120, A_n(58) => net48121, 
                           A_n(57) => net48122, A_n(56) => net48123, A_n(55) =>
                           net48124, A_n(54) => net48125, A_n(53) => net48126, 
                           A_n(52) => net48127, A_n(51) => net48128, A_n(50) =>
                           net48129, A_n(49) => net48130, A_n(48) => net48131, 
                           A_n(47) => net48132, A_n(46) => net48133, A_n(45) =>
                           net48134, A_n(44) => net48135, A_n(43) => net48136, 
                           A_n(42) => net48137, A_n(41) => net48138, A_n(40) =>
                           net48139, A_n(39) => net48140, A_n(38) => net48141, 
                           A_n(37) => net48142, A_n(36) => net48143, A_n(35) =>
                           net48144, A_n(34) => net48145, A_n(33) => net48146, 
                           A_n(32) => net48147, A_n(31) => net48148, A_n(30) =>
                           net48149, A_n(29) => net48150, A_n(28) => net48151, 
                           A_n(27) => net48152, A_n(26) => net48153, A_n(25) =>
                           net48154, A_n(24) => net48155, A_n(23) => net48156, 
                           A_n(22) => net48157, A_n(21) => net48158, A_n(20) =>
                           net48159, A_n(19) => net48160, A_n(18) => net48161, 
                           A_n(17) => net48162, A_n(16) => net48163, A_n(15) =>
                           net48164, A_n(14) => net48165, A_n(13) => net48166, 
                           A_n(12) => net48167, A_n(11) => net48168, A_n(10) =>
                           net48169, A_n(9) => net48170, A_n(8) => net48171, 
                           A_n(7) => net48172, A_n(6) => net48173, A_n(5) => 
                           net48174, A_n(4) => net48175, A_n(3) => net48176, 
                           A_n(2) => net48177, A_n(1) => net48178, A_n(0) => 
                           net48179, A_ns(63) => SHIFT_n_383_port, A_ns(62) => 
                           SHIFT_n_382_port, A_ns(61) => SHIFT_n_381_port, 
                           A_ns(60) => SHIFT_n_380_port, A_ns(59) => 
                           SHIFT_n_379_port, A_ns(58) => SHIFT_n_378_port, 
                           A_ns(57) => SHIFT_n_377_port, A_ns(56) => 
                           SHIFT_n_376_port, A_ns(55) => SHIFT_n_375_port, 
                           A_ns(54) => SHIFT_n_374_port, A_ns(53) => 
                           SHIFT_n_373_port, A_ns(52) => SHIFT_n_372_port, 
                           A_ns(51) => SHIFT_n_371_port, A_ns(50) => 
                           SHIFT_n_370_port, A_ns(49) => SHIFT_n_369_port, 
                           A_ns(48) => SHIFT_n_368_port, A_ns(47) => 
                           SHIFT_n_367_port, A_ns(46) => SHIFT_n_366_port, 
                           A_ns(45) => SHIFT_n_365_port, A_ns(44) => 
                           SHIFT_n_364_port, A_ns(43) => SHIFT_n_363_port, 
                           A_ns(42) => SHIFT_n_362_port, A_ns(41) => 
                           SHIFT_n_361_port, A_ns(40) => SHIFT_n_360_port, 
                           A_ns(39) => SHIFT_n_359_port, A_ns(38) => 
                           SHIFT_n_358_port, A_ns(37) => SHIFT_n_357_port, 
                           A_ns(36) => SHIFT_n_356_port, A_ns(35) => 
                           SHIFT_n_355_port, A_ns(34) => SHIFT_n_354_port, 
                           A_ns(33) => SHIFT_n_353_port, A_ns(32) => 
                           SHIFT_n_352_port, A_ns(31) => SHIFT_n_351_port, 
                           A_ns(30) => SHIFT_n_350_port, A_ns(29) => 
                           SHIFT_n_349_port, A_ns(28) => SHIFT_n_348_port, 
                           A_ns(27) => SHIFT_n_347_port, A_ns(26) => 
                           SHIFT_n_346_port, A_ns(25) => SHIFT_n_345_port, 
                           A_ns(24) => SHIFT_n_344_port, A_ns(23) => 
                           SHIFT_n_343_port, A_ns(22) => SHIFT_n_342_port, 
                           A_ns(21) => SHIFT_n_341_port, A_ns(20) => 
                           SHIFT_n_340_port, A_ns(19) => SHIFT_n_339_port, 
                           A_ns(18) => SHIFT_n_338_port, A_ns(17) => 
                           SHIFT_n_337_port, A_ns(16) => SHIFT_n_336_port, 
                           A_ns(15) => SHIFT_n_335_port, A_ns(14) => 
                           SHIFT_n_334_port, A_ns(13) => SHIFT_n_333_port, 
                           A_ns(12) => SHIFT_n_332_port, A_ns(11) => 
                           SHIFT_n_331_port, A_ns(10) => SHIFT_n_330_port, 
                           A_ns(9) => SHIFT_n_329_port, A_ns(8) => 
                           SHIFT_n_328_port, A_ns(7) => SHIFT_n_327_port, 
                           A_ns(6) => SHIFT_n_326_port, A_ns(5) => 
                           SHIFT_n_325_port, A_ns(4) => SHIFT_n_324_port, 
                           A_ns(3) => SHIFT_n_323_port, A_ns(2) => 
                           SHIFT_n_322_port, A_ns(1) => SHIFT_n_321_port, 
                           A_ns(0) => SHIFT_n_320_port, A_s(63) => 
                           SHIFT_383_port, A_s(62) => SHIFT_382_port, A_s(61) 
                           => SHIFT_381_port, A_s(60) => SHIFT_380_port, 
                           A_s(59) => SHIFT_379_port, A_s(58) => SHIFT_378_port
                           , A_s(57) => SHIFT_377_port, A_s(56) => 
                           SHIFT_376_port, A_s(55) => SHIFT_375_port, A_s(54) 
                           => SHIFT_374_port, A_s(53) => SHIFT_373_port, 
                           A_s(52) => SHIFT_372_port, A_s(51) => SHIFT_371_port
                           , A_s(50) => SHIFT_370_port, A_s(49) => 
                           SHIFT_369_port, A_s(48) => SHIFT_368_port, A_s(47) 
                           => SHIFT_367_port, A_s(46) => SHIFT_366_port, 
                           A_s(45) => SHIFT_365_port, A_s(44) => SHIFT_364_port
                           , A_s(43) => SHIFT_363_port, A_s(42) => 
                           SHIFT_362_port, A_s(41) => SHIFT_361_port, A_s(40) 
                           => SHIFT_360_port, A_s(39) => SHIFT_359_port, 
                           A_s(38) => SHIFT_358_port, A_s(37) => SHIFT_357_port
                           , A_s(36) => SHIFT_356_port, A_s(35) => 
                           SHIFT_355_port, A_s(34) => SHIFT_354_port, A_s(33) 
                           => SHIFT_353_port, A_s(32) => SHIFT_352_port, 
                           A_s(31) => SHIFT_351_port, A_s(30) => SHIFT_350_port
                           , A_s(29) => SHIFT_349_port, A_s(28) => 
                           SHIFT_348_port, A_s(27) => SHIFT_347_port, A_s(26) 
                           => SHIFT_346_port, A_s(25) => SHIFT_345_port, 
                           A_s(24) => SHIFT_344_port, A_s(23) => SHIFT_343_port
                           , A_s(22) => SHIFT_342_port, A_s(21) => 
                           SHIFT_341_port, A_s(20) => SHIFT_340_port, A_s(19) 
                           => SHIFT_339_port, A_s(18) => SHIFT_338_port, 
                           A_s(17) => SHIFT_337_port, A_s(16) => SHIFT_336_port
                           , A_s(15) => SHIFT_335_port, A_s(14) => 
                           SHIFT_334_port, A_s(13) => SHIFT_333_port, A_s(12) 
                           => SHIFT_332_port, A_s(11) => SHIFT_331_port, 
                           A_s(10) => SHIFT_330_port, A_s(9) => SHIFT_329_port,
                           A_s(8) => SHIFT_328_port, A_s(7) => SHIFT_327_port, 
                           A_s(6) => SHIFT_326_port, A_s(5) => SHIFT_325_port, 
                           A_s(4) => SHIFT_324_port, A_s(3) => SHIFT_323_port, 
                           A_s(2) => SHIFT_322_port, A_s(1) => SHIFT_321_port, 
                           A_s(0) => SHIFT_320_port, B(63) => B(31), B(62) => 
                           B(31), B(61) => B(31), B(60) => B(31), B(59) => 
                           B(31), B(58) => B(31), B(57) => B(31), B(56) => 
                           B(31), B(55) => B(31), B(54) => B(31), B(53) => 
                           B(31), B(52) => B(31), B(51) => B(31), B(50) => 
                           B(31), B(49) => B(31), B(48) => B(31), B(47) => 
                           B(31), B(46) => B(31), B(45) => B(31), B(44) => 
                           B(31), B(43) => B(31), B(42) => B(31), B(41) => 
                           B(31), B(40) => B(31), B(39) => B(31), B(38) => 
                           B(31), B(37) => B(31), B(36) => B(31), B(35) => 
                           B(31), B(34) => B(31), B(33) => B(31), B(32) => 
                           B(31), B(31) => B(31), B(30) => B(30), B(29) => 
                           B(29), B(28) => B(28), B(27) => B(27), B(26) => 
                           B(26), B(25) => B(25), B(24) => B(24), B(23) => 
                           B(23), B(22) => B(22), B(21) => B(21), B(20) => 
                           B(20), B(19) => B(19), B(18) => B(18), B(17) => 
                           B(17), B(16) => B(16), B(15) => B(15), B(14) => 
                           B(14), B(13) => B(13), B(12) => B(12), B(11) => 
                           B(11), B(10) => B(10), B(9) => B(9), B(8) => B(8), 
                           B(7) => B(7), B(6) => B(6), B(5) => B(5), B(4) => 
                           B(4), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), O(63) => OTMP_383_port, O(62) => 
                           OTMP_382_port, O(61) => OTMP_381_port, O(60) => 
                           OTMP_380_port, O(59) => OTMP_379_port, O(58) => 
                           OTMP_378_port, O(57) => OTMP_377_port, O(56) => 
                           OTMP_376_port, O(55) => OTMP_375_port, O(54) => 
                           OTMP_374_port, O(53) => OTMP_373_port, O(52) => 
                           OTMP_372_port, O(51) => OTMP_371_port, O(50) => 
                           OTMP_370_port, O(49) => OTMP_369_port, O(48) => 
                           OTMP_368_port, O(47) => OTMP_367_port, O(46) => 
                           OTMP_366_port, O(45) => OTMP_365_port, O(44) => 
                           OTMP_364_port, O(43) => OTMP_363_port, O(42) => 
                           OTMP_362_port, O(41) => OTMP_361_port, O(40) => 
                           OTMP_360_port, O(39) => OTMP_359_port, O(38) => 
                           OTMP_358_port, O(37) => OTMP_357_port, O(36) => 
                           OTMP_356_port, O(35) => OTMP_355_port, O(34) => 
                           OTMP_354_port, O(33) => OTMP_353_port, O(32) => 
                           OTMP_352_port, O(31) => OTMP_351_port, O(30) => 
                           OTMP_350_port, O(29) => OTMP_349_port, O(28) => 
                           OTMP_348_port, O(27) => OTMP_347_port, O(26) => 
                           OTMP_346_port, O(25) => OTMP_345_port, O(24) => 
                           OTMP_344_port, O(23) => OTMP_343_port, O(22) => 
                           OTMP_342_port, O(21) => OTMP_341_port, O(20) => 
                           OTMP_340_port, O(19) => OTMP_339_port, O(18) => 
                           OTMP_338_port, O(17) => OTMP_337_port, O(16) => 
                           OTMP_336_port, O(15) => OTMP_335_port, O(14) => 
                           OTMP_334_port, O(13) => OTMP_333_port, O(12) => 
                           OTMP_332_port, O(11) => OTMP_331_port, O(10) => 
                           OTMP_330_port, O(9) => OTMP_329_port, O(8) => 
                           OTMP_328_port, O(7) => OTMP_327_port, O(6) => 
                           OTMP_326_port, O(5) => OTMP_325_port, O(4) => 
                           OTMP_324_port, O(3) => OTMP_323_port, O(2) => 
                           OTMP_322_port, O(1) => OTMP_321_port, O(0) => n_1116
                           , A_so(63) => SHIFT_447_port, A_so(62) => 
                           SHIFT_446_port, A_so(61) => SHIFT_445_port, A_so(60)
                           => SHIFT_444_port, A_so(59) => SHIFT_443_port, 
                           A_so(58) => SHIFT_442_port, A_so(57) => 
                           SHIFT_441_port, A_so(56) => SHIFT_440_port, A_so(55)
                           => SHIFT_439_port, A_so(54) => SHIFT_438_port, 
                           A_so(53) => SHIFT_437_port, A_so(52) => 
                           SHIFT_436_port, A_so(51) => SHIFT_435_port, A_so(50)
                           => SHIFT_434_port, A_so(49) => SHIFT_433_port, 
                           A_so(48) => SHIFT_432_port, A_so(47) => 
                           SHIFT_431_port, A_so(46) => SHIFT_430_port, A_so(45)
                           => SHIFT_429_port, A_so(44) => SHIFT_428_port, 
                           A_so(43) => SHIFT_427_port, A_so(42) => 
                           SHIFT_426_port, A_so(41) => SHIFT_425_port, A_so(40)
                           => SHIFT_424_port, A_so(39) => SHIFT_423_port, 
                           A_so(38) => SHIFT_422_port, A_so(37) => 
                           SHIFT_421_port, A_so(36) => SHIFT_420_port, A_so(35)
                           => SHIFT_419_port, A_so(34) => SHIFT_418_port, 
                           A_so(33) => SHIFT_417_port, A_so(32) => 
                           SHIFT_416_port, A_so(31) => SHIFT_415_port, A_so(30)
                           => SHIFT_414_port, A_so(29) => SHIFT_413_port, 
                           A_so(28) => SHIFT_412_port, A_so(27) => 
                           SHIFT_411_port, A_so(26) => SHIFT_410_port, A_so(25)
                           => SHIFT_409_port, A_so(24) => SHIFT_408_port, 
                           A_so(23) => SHIFT_407_port, A_so(22) => 
                           SHIFT_406_port, A_so(21) => SHIFT_405_port, A_so(20)
                           => SHIFT_404_port, A_so(19) => SHIFT_403_port, 
                           A_so(18) => SHIFT_402_port, A_so(17) => 
                           SHIFT_401_port, A_so(16) => SHIFT_400_port, A_so(15)
                           => SHIFT_399_port, A_so(14) => SHIFT_398_port, 
                           A_so(13) => SHIFT_397_port, A_so(12) => 
                           SHIFT_396_port, A_so(11) => SHIFT_395_port, A_so(10)
                           => SHIFT_394_port, A_so(9) => SHIFT_393_port, 
                           A_so(8) => SHIFT_392_port, A_so(7) => SHIFT_391_port
                           , A_so(6) => SHIFT_390_port, A_so(5) => 
                           SHIFT_389_port, A_so(4) => SHIFT_388_port, A_so(3) 
                           => SHIFT_387_port, A_so(2) => SHIFT_386_port, 
                           A_so(1) => n_1117, A_so(0) => n_1118, A_nso(63) => 
                           SHIFT_n_447_port, A_nso(62) => SHIFT_n_446_port, 
                           A_nso(61) => SHIFT_n_445_port, A_nso(60) => 
                           SHIFT_n_444_port, A_nso(59) => SHIFT_n_443_port, 
                           A_nso(58) => SHIFT_n_442_port, A_nso(57) => 
                           SHIFT_n_441_port, A_nso(56) => SHIFT_n_440_port, 
                           A_nso(55) => SHIFT_n_439_port, A_nso(54) => 
                           SHIFT_n_438_port, A_nso(53) => SHIFT_n_437_port, 
                           A_nso(52) => SHIFT_n_436_port, A_nso(51) => 
                           SHIFT_n_435_port, A_nso(50) => SHIFT_n_434_port, 
                           A_nso(49) => SHIFT_n_433_port, A_nso(48) => 
                           SHIFT_n_432_port, A_nso(47) => SHIFT_n_431_port, 
                           A_nso(46) => SHIFT_n_430_port, A_nso(45) => 
                           SHIFT_n_429_port, A_nso(44) => SHIFT_n_428_port, 
                           A_nso(43) => SHIFT_n_427_port, A_nso(42) => 
                           SHIFT_n_426_port, A_nso(41) => SHIFT_n_425_port, 
                           A_nso(40) => SHIFT_n_424_port, A_nso(39) => 
                           SHIFT_n_423_port, A_nso(38) => SHIFT_n_422_port, 
                           A_nso(37) => SHIFT_n_421_port, A_nso(36) => 
                           SHIFT_n_420_port, A_nso(35) => SHIFT_n_419_port, 
                           A_nso(34) => SHIFT_n_418_port, A_nso(33) => 
                           SHIFT_n_417_port, A_nso(32) => SHIFT_n_416_port, 
                           A_nso(31) => SHIFT_n_415_port, A_nso(30) => 
                           SHIFT_n_414_port, A_nso(29) => SHIFT_n_413_port, 
                           A_nso(28) => SHIFT_n_412_port, A_nso(27) => 
                           SHIFT_n_411_port, A_nso(26) => SHIFT_n_410_port, 
                           A_nso(25) => SHIFT_n_409_port, A_nso(24) => 
                           SHIFT_n_408_port, A_nso(23) => SHIFT_n_407_port, 
                           A_nso(22) => SHIFT_n_406_port, A_nso(21) => 
                           SHIFT_n_405_port, A_nso(20) => SHIFT_n_404_port, 
                           A_nso(19) => SHIFT_n_403_port, A_nso(18) => 
                           SHIFT_n_402_port, A_nso(17) => SHIFT_n_401_port, 
                           A_nso(16) => SHIFT_n_400_port, A_nso(15) => 
                           SHIFT_n_399_port, A_nso(14) => SHIFT_n_398_port, 
                           A_nso(13) => SHIFT_n_397_port, A_nso(12) => 
                           SHIFT_n_396_port, A_nso(11) => SHIFT_n_395_port, 
                           A_nso(10) => SHIFT_n_394_port, A_nso(9) => 
                           SHIFT_n_393_port, A_nso(8) => SHIFT_n_392_port, 
                           A_nso(7) => SHIFT_n_391_port, A_nso(6) => 
                           SHIFT_n_390_port, A_nso(5) => SHIFT_n_389_port, 
                           A_nso(4) => SHIFT_n_388_port, A_nso(3) => 
                           SHIFT_n_387_port, A_nso(2) => SHIFT_n_386_port, 
                           A_nso(1) => n_1119, A_nso(0) => n_1120);
   BOOTHENC_I_7 : BOOTHENC_NBIT64_i12 port map( A(63) => net47924, A(62) => 
                           net47925, A(61) => net47926, A(60) => net47927, 
                           A(59) => net47928, A(58) => net47929, A(57) => 
                           net47930, A(56) => net47931, A(55) => net47932, 
                           A(54) => net47933, A(53) => net47934, A(52) => 
                           net47935, A(51) => net47936, A(50) => net47937, 
                           A(49) => net47938, A(48) => net47939, A(47) => 
                           net47940, A(46) => net47941, A(45) => net47942, 
                           A(44) => net47943, A(43) => net47944, A(42) => 
                           net47945, A(41) => net47946, A(40) => net47947, 
                           A(39) => net47948, A(38) => net47949, A(37) => 
                           net47950, A(36) => net47951, A(35) => net47952, 
                           A(34) => net47953, A(33) => net47954, A(32) => 
                           net47955, A(31) => net47956, A(30) => net47957, 
                           A(29) => net47958, A(28) => net47959, A(27) => 
                           net47960, A(26) => net47961, A(25) => net47962, 
                           A(24) => net47963, A(23) => net47964, A(22) => 
                           net47965, A(21) => net47966, A(20) => net47967, 
                           A(19) => net47968, A(18) => net47969, A(17) => 
                           net47970, A(16) => net47971, A(15) => net47972, 
                           A(14) => net47973, A(13) => net47974, A(12) => 
                           net47975, A(11) => net47976, A(10) => net47977, A(9)
                           => net47978, A(8) => net47979, A(7) => net47980, 
                           A(6) => net47981, A(5) => net47982, A(4) => net47983
                           , A(3) => net47984, A(2) => net47985, A(1) => 
                           net47986, A(0) => net47987, A_n(63) => net47988, 
                           A_n(62) => net47989, A_n(61) => net47990, A_n(60) =>
                           net47991, A_n(59) => net47992, A_n(58) => net47993, 
                           A_n(57) => net47994, A_n(56) => net47995, A_n(55) =>
                           net47996, A_n(54) => net47997, A_n(53) => net47998, 
                           A_n(52) => net47999, A_n(51) => net48000, A_n(50) =>
                           net48001, A_n(49) => net48002, A_n(48) => net48003, 
                           A_n(47) => net48004, A_n(46) => net48005, A_n(45) =>
                           net48006, A_n(44) => net48007, A_n(43) => net48008, 
                           A_n(42) => net48009, A_n(41) => net48010, A_n(40) =>
                           net48011, A_n(39) => net48012, A_n(38) => net48013, 
                           A_n(37) => net48014, A_n(36) => net48015, A_n(35) =>
                           net48016, A_n(34) => net48017, A_n(33) => net48018, 
                           A_n(32) => net48019, A_n(31) => net48020, A_n(30) =>
                           net48021, A_n(29) => net48022, A_n(28) => net48023, 
                           A_n(27) => net48024, A_n(26) => net48025, A_n(25) =>
                           net48026, A_n(24) => net48027, A_n(23) => net48028, 
                           A_n(22) => net48029, A_n(21) => net48030, A_n(20) =>
                           net48031, A_n(19) => net48032, A_n(18) => net48033, 
                           A_n(17) => net48034, A_n(16) => net48035, A_n(15) =>
                           net48036, A_n(14) => net48037, A_n(13) => net48038, 
                           A_n(12) => net48039, A_n(11) => net48040, A_n(10) =>
                           net48041, A_n(9) => net48042, A_n(8) => net48043, 
                           A_n(7) => net48044, A_n(6) => net48045, A_n(5) => 
                           net48046, A_n(4) => net48047, A_n(3) => net48048, 
                           A_n(2) => net48049, A_n(1) => net48050, A_n(0) => 
                           net48051, A_ns(63) => SHIFT_n_447_port, A_ns(62) => 
                           SHIFT_n_446_port, A_ns(61) => SHIFT_n_445_port, 
                           A_ns(60) => SHIFT_n_444_port, A_ns(59) => 
                           SHIFT_n_443_port, A_ns(58) => SHIFT_n_442_port, 
                           A_ns(57) => SHIFT_n_441_port, A_ns(56) => 
                           SHIFT_n_440_port, A_ns(55) => SHIFT_n_439_port, 
                           A_ns(54) => SHIFT_n_438_port, A_ns(53) => 
                           SHIFT_n_437_port, A_ns(52) => SHIFT_n_436_port, 
                           A_ns(51) => SHIFT_n_435_port, A_ns(50) => 
                           SHIFT_n_434_port, A_ns(49) => SHIFT_n_433_port, 
                           A_ns(48) => SHIFT_n_432_port, A_ns(47) => 
                           SHIFT_n_431_port, A_ns(46) => SHIFT_n_430_port, 
                           A_ns(45) => SHIFT_n_429_port, A_ns(44) => 
                           SHIFT_n_428_port, A_ns(43) => SHIFT_n_427_port, 
                           A_ns(42) => SHIFT_n_426_port, A_ns(41) => 
                           SHIFT_n_425_port, A_ns(40) => SHIFT_n_424_port, 
                           A_ns(39) => SHIFT_n_423_port, A_ns(38) => 
                           SHIFT_n_422_port, A_ns(37) => SHIFT_n_421_port, 
                           A_ns(36) => SHIFT_n_420_port, A_ns(35) => 
                           SHIFT_n_419_port, A_ns(34) => SHIFT_n_418_port, 
                           A_ns(33) => SHIFT_n_417_port, A_ns(32) => 
                           SHIFT_n_416_port, A_ns(31) => SHIFT_n_415_port, 
                           A_ns(30) => SHIFT_n_414_port, A_ns(29) => 
                           SHIFT_n_413_port, A_ns(28) => SHIFT_n_412_port, 
                           A_ns(27) => SHIFT_n_411_port, A_ns(26) => 
                           SHIFT_n_410_port, A_ns(25) => SHIFT_n_409_port, 
                           A_ns(24) => SHIFT_n_408_port, A_ns(23) => 
                           SHIFT_n_407_port, A_ns(22) => SHIFT_n_406_port, 
                           A_ns(21) => SHIFT_n_405_port, A_ns(20) => 
                           SHIFT_n_404_port, A_ns(19) => SHIFT_n_403_port, 
                           A_ns(18) => SHIFT_n_402_port, A_ns(17) => 
                           SHIFT_n_401_port, A_ns(16) => SHIFT_n_400_port, 
                           A_ns(15) => SHIFT_n_399_port, A_ns(14) => 
                           SHIFT_n_398_port, A_ns(13) => SHIFT_n_397_port, 
                           A_ns(12) => SHIFT_n_396_port, A_ns(11) => 
                           SHIFT_n_395_port, A_ns(10) => SHIFT_n_394_port, 
                           A_ns(9) => SHIFT_n_393_port, A_ns(8) => 
                           SHIFT_n_392_port, A_ns(7) => SHIFT_n_391_port, 
                           A_ns(6) => SHIFT_n_390_port, A_ns(5) => 
                           SHIFT_n_389_port, A_ns(4) => SHIFT_n_388_port, 
                           A_ns(3) => SHIFT_n_387_port, A_ns(2) => 
                           SHIFT_n_386_port, A_ns(1) => SHIFT_n_385_port, 
                           A_ns(0) => SHIFT_n_384_port, A_s(63) => 
                           SHIFT_447_port, A_s(62) => SHIFT_446_port, A_s(61) 
                           => SHIFT_445_port, A_s(60) => SHIFT_444_port, 
                           A_s(59) => SHIFT_443_port, A_s(58) => SHIFT_442_port
                           , A_s(57) => SHIFT_441_port, A_s(56) => 
                           SHIFT_440_port, A_s(55) => SHIFT_439_port, A_s(54) 
                           => SHIFT_438_port, A_s(53) => SHIFT_437_port, 
                           A_s(52) => SHIFT_436_port, A_s(51) => SHIFT_435_port
                           , A_s(50) => SHIFT_434_port, A_s(49) => 
                           SHIFT_433_port, A_s(48) => SHIFT_432_port, A_s(47) 
                           => SHIFT_431_port, A_s(46) => SHIFT_430_port, 
                           A_s(45) => SHIFT_429_port, A_s(44) => SHIFT_428_port
                           , A_s(43) => SHIFT_427_port, A_s(42) => 
                           SHIFT_426_port, A_s(41) => SHIFT_425_port, A_s(40) 
                           => SHIFT_424_port, A_s(39) => SHIFT_423_port, 
                           A_s(38) => SHIFT_422_port, A_s(37) => SHIFT_421_port
                           , A_s(36) => SHIFT_420_port, A_s(35) => 
                           SHIFT_419_port, A_s(34) => SHIFT_418_port, A_s(33) 
                           => SHIFT_417_port, A_s(32) => SHIFT_416_port, 
                           A_s(31) => SHIFT_415_port, A_s(30) => SHIFT_414_port
                           , A_s(29) => SHIFT_413_port, A_s(28) => 
                           SHIFT_412_port, A_s(27) => SHIFT_411_port, A_s(26) 
                           => SHIFT_410_port, A_s(25) => SHIFT_409_port, 
                           A_s(24) => SHIFT_408_port, A_s(23) => SHIFT_407_port
                           , A_s(22) => SHIFT_406_port, A_s(21) => 
                           SHIFT_405_port, A_s(20) => SHIFT_404_port, A_s(19) 
                           => SHIFT_403_port, A_s(18) => SHIFT_402_port, 
                           A_s(17) => SHIFT_401_port, A_s(16) => SHIFT_400_port
                           , A_s(15) => SHIFT_399_port, A_s(14) => 
                           SHIFT_398_port, A_s(13) => SHIFT_397_port, A_s(12) 
                           => SHIFT_396_port, A_s(11) => SHIFT_395_port, 
                           A_s(10) => SHIFT_394_port, A_s(9) => SHIFT_393_port,
                           A_s(8) => SHIFT_392_port, A_s(7) => SHIFT_391_port, 
                           A_s(6) => SHIFT_390_port, A_s(5) => SHIFT_389_port, 
                           A_s(4) => SHIFT_388_port, A_s(3) => SHIFT_387_port, 
                           A_s(2) => SHIFT_386_port, A_s(1) => SHIFT_385_port, 
                           A_s(0) => SHIFT_384_port, B(63) => B(31), B(62) => 
                           B(31), B(61) => B(31), B(60) => B(31), B(59) => 
                           B(31), B(58) => B(31), B(57) => B(31), B(56) => 
                           B(31), B(55) => B(31), B(54) => B(31), B(53) => 
                           B(31), B(52) => B(31), B(51) => B(31), B(50) => 
                           B(31), B(49) => B(31), B(48) => B(31), B(47) => 
                           B(31), B(46) => B(31), B(45) => B(31), B(44) => 
                           B(31), B(43) => B(31), B(42) => B(31), B(41) => 
                           B(31), B(40) => B(31), B(39) => B(31), B(38) => 
                           B(31), B(37) => B(31), B(36) => B(31), B(35) => 
                           B(31), B(34) => B(31), B(33) => B(31), B(32) => 
                           B(31), B(31) => B(31), B(30) => B(30), B(29) => 
                           B(29), B(28) => B(28), B(27) => B(27), B(26) => 
                           B(26), B(25) => B(25), B(24) => B(24), B(23) => 
                           B(23), B(22) => B(22), B(21) => B(21), B(20) => 
                           B(20), B(19) => B(19), B(18) => B(18), B(17) => 
                           B(17), B(16) => B(16), B(15) => B(15), B(14) => 
                           B(14), B(13) => B(13), B(12) => B(12), B(11) => 
                           B(11), B(10) => B(10), B(9) => B(9), B(8) => B(8), 
                           B(7) => B(7), B(6) => B(6), B(5) => B(5), B(4) => 
                           B(4), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), O(63) => OTMP_447_port, O(62) => 
                           OTMP_446_port, O(61) => OTMP_445_port, O(60) => 
                           OTMP_444_port, O(59) => OTMP_443_port, O(58) => 
                           OTMP_442_port, O(57) => OTMP_441_port, O(56) => 
                           OTMP_440_port, O(55) => OTMP_439_port, O(54) => 
                           OTMP_438_port, O(53) => OTMP_437_port, O(52) => 
                           OTMP_436_port, O(51) => OTMP_435_port, O(50) => 
                           OTMP_434_port, O(49) => OTMP_433_port, O(48) => 
                           OTMP_432_port, O(47) => OTMP_431_port, O(46) => 
                           OTMP_430_port, O(45) => OTMP_429_port, O(44) => 
                           OTMP_428_port, O(43) => OTMP_427_port, O(42) => 
                           OTMP_426_port, O(41) => OTMP_425_port, O(40) => 
                           OTMP_424_port, O(39) => OTMP_423_port, O(38) => 
                           OTMP_422_port, O(37) => OTMP_421_port, O(36) => 
                           OTMP_420_port, O(35) => OTMP_419_port, O(34) => 
                           OTMP_418_port, O(33) => OTMP_417_port, O(32) => 
                           OTMP_416_port, O(31) => OTMP_415_port, O(30) => 
                           OTMP_414_port, O(29) => OTMP_413_port, O(28) => 
                           OTMP_412_port, O(27) => OTMP_411_port, O(26) => 
                           OTMP_410_port, O(25) => OTMP_409_port, O(24) => 
                           OTMP_408_port, O(23) => OTMP_407_port, O(22) => 
                           OTMP_406_port, O(21) => OTMP_405_port, O(20) => 
                           OTMP_404_port, O(19) => OTMP_403_port, O(18) => 
                           OTMP_402_port, O(17) => OTMP_401_port, O(16) => 
                           OTMP_400_port, O(15) => OTMP_399_port, O(14) => 
                           OTMP_398_port, O(13) => OTMP_397_port, O(12) => 
                           OTMP_396_port, O(11) => OTMP_395_port, O(10) => 
                           OTMP_394_port, O(9) => OTMP_393_port, O(8) => 
                           OTMP_392_port, O(7) => OTMP_391_port, O(6) => 
                           OTMP_390_port, O(5) => OTMP_389_port, O(4) => 
                           OTMP_388_port, O(3) => OTMP_387_port, O(2) => 
                           OTMP_386_port, O(1) => OTMP_385_port, O(0) => n_1121
                           , A_so(63) => SHIFT_511_port, A_so(62) => 
                           SHIFT_510_port, A_so(61) => SHIFT_509_port, A_so(60)
                           => SHIFT_508_port, A_so(59) => SHIFT_507_port, 
                           A_so(58) => SHIFT_506_port, A_so(57) => 
                           SHIFT_505_port, A_so(56) => SHIFT_504_port, A_so(55)
                           => SHIFT_503_port, A_so(54) => SHIFT_502_port, 
                           A_so(53) => SHIFT_501_port, A_so(52) => 
                           SHIFT_500_port, A_so(51) => SHIFT_499_port, A_so(50)
                           => SHIFT_498_port, A_so(49) => SHIFT_497_port, 
                           A_so(48) => SHIFT_496_port, A_so(47) => 
                           SHIFT_495_port, A_so(46) => SHIFT_494_port, A_so(45)
                           => SHIFT_493_port, A_so(44) => SHIFT_492_port, 
                           A_so(43) => SHIFT_491_port, A_so(42) => 
                           SHIFT_490_port, A_so(41) => SHIFT_489_port, A_so(40)
                           => SHIFT_488_port, A_so(39) => SHIFT_487_port, 
                           A_so(38) => SHIFT_486_port, A_so(37) => 
                           SHIFT_485_port, A_so(36) => SHIFT_484_port, A_so(35)
                           => SHIFT_483_port, A_so(34) => SHIFT_482_port, 
                           A_so(33) => SHIFT_481_port, A_so(32) => 
                           SHIFT_480_port, A_so(31) => SHIFT_479_port, A_so(30)
                           => SHIFT_478_port, A_so(29) => SHIFT_477_port, 
                           A_so(28) => SHIFT_476_port, A_so(27) => 
                           SHIFT_475_port, A_so(26) => SHIFT_474_port, A_so(25)
                           => SHIFT_473_port, A_so(24) => SHIFT_472_port, 
                           A_so(23) => SHIFT_471_port, A_so(22) => 
                           SHIFT_470_port, A_so(21) => SHIFT_469_port, A_so(20)
                           => SHIFT_468_port, A_so(19) => SHIFT_467_port, 
                           A_so(18) => SHIFT_466_port, A_so(17) => 
                           SHIFT_465_port, A_so(16) => SHIFT_464_port, A_so(15)
                           => SHIFT_463_port, A_so(14) => SHIFT_462_port, 
                           A_so(13) => SHIFT_461_port, A_so(12) => 
                           SHIFT_460_port, A_so(11) => SHIFT_459_port, A_so(10)
                           => SHIFT_458_port, A_so(9) => SHIFT_457_port, 
                           A_so(8) => SHIFT_456_port, A_so(7) => SHIFT_455_port
                           , A_so(6) => SHIFT_454_port, A_so(5) => 
                           SHIFT_453_port, A_so(4) => SHIFT_452_port, A_so(3) 
                           => SHIFT_451_port, A_so(2) => SHIFT_450_port, 
                           A_so(1) => n_1122, A_so(0) => n_1123, A_nso(63) => 
                           SHIFT_n_511_port, A_nso(62) => SHIFT_n_510_port, 
                           A_nso(61) => SHIFT_n_509_port, A_nso(60) => 
                           SHIFT_n_508_port, A_nso(59) => SHIFT_n_507_port, 
                           A_nso(58) => SHIFT_n_506_port, A_nso(57) => 
                           SHIFT_n_505_port, A_nso(56) => SHIFT_n_504_port, 
                           A_nso(55) => SHIFT_n_503_port, A_nso(54) => 
                           SHIFT_n_502_port, A_nso(53) => SHIFT_n_501_port, 
                           A_nso(52) => SHIFT_n_500_port, A_nso(51) => 
                           SHIFT_n_499_port, A_nso(50) => SHIFT_n_498_port, 
                           A_nso(49) => SHIFT_n_497_port, A_nso(48) => 
                           SHIFT_n_496_port, A_nso(47) => SHIFT_n_495_port, 
                           A_nso(46) => SHIFT_n_494_port, A_nso(45) => 
                           SHIFT_n_493_port, A_nso(44) => SHIFT_n_492_port, 
                           A_nso(43) => SHIFT_n_491_port, A_nso(42) => 
                           SHIFT_n_490_port, A_nso(41) => SHIFT_n_489_port, 
                           A_nso(40) => SHIFT_n_488_port, A_nso(39) => 
                           SHIFT_n_487_port, A_nso(38) => SHIFT_n_486_port, 
                           A_nso(37) => SHIFT_n_485_port, A_nso(36) => 
                           SHIFT_n_484_port, A_nso(35) => SHIFT_n_483_port, 
                           A_nso(34) => SHIFT_n_482_port, A_nso(33) => 
                           SHIFT_n_481_port, A_nso(32) => SHIFT_n_480_port, 
                           A_nso(31) => SHIFT_n_479_port, A_nso(30) => 
                           SHIFT_n_478_port, A_nso(29) => SHIFT_n_477_port, 
                           A_nso(28) => SHIFT_n_476_port, A_nso(27) => 
                           SHIFT_n_475_port, A_nso(26) => SHIFT_n_474_port, 
                           A_nso(25) => SHIFT_n_473_port, A_nso(24) => 
                           SHIFT_n_472_port, A_nso(23) => SHIFT_n_471_port, 
                           A_nso(22) => SHIFT_n_470_port, A_nso(21) => 
                           SHIFT_n_469_port, A_nso(20) => SHIFT_n_468_port, 
                           A_nso(19) => SHIFT_n_467_port, A_nso(18) => 
                           SHIFT_n_466_port, A_nso(17) => SHIFT_n_465_port, 
                           A_nso(16) => SHIFT_n_464_port, A_nso(15) => 
                           SHIFT_n_463_port, A_nso(14) => SHIFT_n_462_port, 
                           A_nso(13) => SHIFT_n_461_port, A_nso(12) => 
                           SHIFT_n_460_port, A_nso(11) => SHIFT_n_459_port, 
                           A_nso(10) => SHIFT_n_458_port, A_nso(9) => 
                           SHIFT_n_457_port, A_nso(8) => SHIFT_n_456_port, 
                           A_nso(7) => SHIFT_n_455_port, A_nso(6) => 
                           SHIFT_n_454_port, A_nso(5) => SHIFT_n_453_port, 
                           A_nso(4) => SHIFT_n_452_port, A_nso(3) => 
                           SHIFT_n_451_port, A_nso(2) => SHIFT_n_450_port, 
                           A_nso(1) => n_1124, A_nso(0) => n_1125);
   BOOTHENC_I_8 : BOOTHENC_NBIT64_i14 port map( A(63) => net47796, A(62) => 
                           net47797, A(61) => net47798, A(60) => net47799, 
                           A(59) => net47800, A(58) => net47801, A(57) => 
                           net47802, A(56) => net47803, A(55) => net47804, 
                           A(54) => net47805, A(53) => net47806, A(52) => 
                           net47807, A(51) => net47808, A(50) => net47809, 
                           A(49) => net47810, A(48) => net47811, A(47) => 
                           net47812, A(46) => net47813, A(45) => net47814, 
                           A(44) => net47815, A(43) => net47816, A(42) => 
                           net47817, A(41) => net47818, A(40) => net47819, 
                           A(39) => net47820, A(38) => net47821, A(37) => 
                           net47822, A(36) => net47823, A(35) => net47824, 
                           A(34) => net47825, A(33) => net47826, A(32) => 
                           net47827, A(31) => net47828, A(30) => net47829, 
                           A(29) => net47830, A(28) => net47831, A(27) => 
                           net47832, A(26) => net47833, A(25) => net47834, 
                           A(24) => net47835, A(23) => net47836, A(22) => 
                           net47837, A(21) => net47838, A(20) => net47839, 
                           A(19) => net47840, A(18) => net47841, A(17) => 
                           net47842, A(16) => net47843, A(15) => net47844, 
                           A(14) => net47845, A(13) => net47846, A(12) => 
                           net47847, A(11) => net47848, A(10) => net47849, A(9)
                           => net47850, A(8) => net47851, A(7) => net47852, 
                           A(6) => net47853, A(5) => net47854, A(4) => net47855
                           , A(3) => net47856, A(2) => net47857, A(1) => 
                           net47858, A(0) => net47859, A_n(63) => net47860, 
                           A_n(62) => net47861, A_n(61) => net47862, A_n(60) =>
                           net47863, A_n(59) => net47864, A_n(58) => net47865, 
                           A_n(57) => net47866, A_n(56) => net47867, A_n(55) =>
                           net47868, A_n(54) => net47869, A_n(53) => net47870, 
                           A_n(52) => net47871, A_n(51) => net47872, A_n(50) =>
                           net47873, A_n(49) => net47874, A_n(48) => net47875, 
                           A_n(47) => net47876, A_n(46) => net47877, A_n(45) =>
                           net47878, A_n(44) => net47879, A_n(43) => net47880, 
                           A_n(42) => net47881, A_n(41) => net47882, A_n(40) =>
                           net47883, A_n(39) => net47884, A_n(38) => net47885, 
                           A_n(37) => net47886, A_n(36) => net47887, A_n(35) =>
                           net47888, A_n(34) => net47889, A_n(33) => net47890, 
                           A_n(32) => net47891, A_n(31) => net47892, A_n(30) =>
                           net47893, A_n(29) => net47894, A_n(28) => net47895, 
                           A_n(27) => net47896, A_n(26) => net47897, A_n(25) =>
                           net47898, A_n(24) => net47899, A_n(23) => net47900, 
                           A_n(22) => net47901, A_n(21) => net47902, A_n(20) =>
                           net47903, A_n(19) => net47904, A_n(18) => net47905, 
                           A_n(17) => net47906, A_n(16) => net47907, A_n(15) =>
                           net47908, A_n(14) => net47909, A_n(13) => net47910, 
                           A_n(12) => net47911, A_n(11) => net47912, A_n(10) =>
                           net47913, A_n(9) => net47914, A_n(8) => net47915, 
                           A_n(7) => net47916, A_n(6) => net47917, A_n(5) => 
                           net47918, A_n(4) => net47919, A_n(3) => net47920, 
                           A_n(2) => net47921, A_n(1) => net47922, A_n(0) => 
                           net47923, A_ns(63) => SHIFT_n_511_port, A_ns(62) => 
                           SHIFT_n_510_port, A_ns(61) => SHIFT_n_509_port, 
                           A_ns(60) => SHIFT_n_508_port, A_ns(59) => 
                           SHIFT_n_507_port, A_ns(58) => SHIFT_n_506_port, 
                           A_ns(57) => SHIFT_n_505_port, A_ns(56) => 
                           SHIFT_n_504_port, A_ns(55) => SHIFT_n_503_port, 
                           A_ns(54) => SHIFT_n_502_port, A_ns(53) => 
                           SHIFT_n_501_port, A_ns(52) => SHIFT_n_500_port, 
                           A_ns(51) => SHIFT_n_499_port, A_ns(50) => 
                           SHIFT_n_498_port, A_ns(49) => SHIFT_n_497_port, 
                           A_ns(48) => SHIFT_n_496_port, A_ns(47) => 
                           SHIFT_n_495_port, A_ns(46) => SHIFT_n_494_port, 
                           A_ns(45) => SHIFT_n_493_port, A_ns(44) => 
                           SHIFT_n_492_port, A_ns(43) => SHIFT_n_491_port, 
                           A_ns(42) => SHIFT_n_490_port, A_ns(41) => 
                           SHIFT_n_489_port, A_ns(40) => SHIFT_n_488_port, 
                           A_ns(39) => SHIFT_n_487_port, A_ns(38) => 
                           SHIFT_n_486_port, A_ns(37) => SHIFT_n_485_port, 
                           A_ns(36) => SHIFT_n_484_port, A_ns(35) => 
                           SHIFT_n_483_port, A_ns(34) => SHIFT_n_482_port, 
                           A_ns(33) => SHIFT_n_481_port, A_ns(32) => 
                           SHIFT_n_480_port, A_ns(31) => SHIFT_n_479_port, 
                           A_ns(30) => SHIFT_n_478_port, A_ns(29) => 
                           SHIFT_n_477_port, A_ns(28) => SHIFT_n_476_port, 
                           A_ns(27) => SHIFT_n_475_port, A_ns(26) => 
                           SHIFT_n_474_port, A_ns(25) => SHIFT_n_473_port, 
                           A_ns(24) => SHIFT_n_472_port, A_ns(23) => 
                           SHIFT_n_471_port, A_ns(22) => SHIFT_n_470_port, 
                           A_ns(21) => SHIFT_n_469_port, A_ns(20) => 
                           SHIFT_n_468_port, A_ns(19) => SHIFT_n_467_port, 
                           A_ns(18) => SHIFT_n_466_port, A_ns(17) => 
                           SHIFT_n_465_port, A_ns(16) => SHIFT_n_464_port, 
                           A_ns(15) => SHIFT_n_463_port, A_ns(14) => 
                           SHIFT_n_462_port, A_ns(13) => SHIFT_n_461_port, 
                           A_ns(12) => SHIFT_n_460_port, A_ns(11) => 
                           SHIFT_n_459_port, A_ns(10) => SHIFT_n_458_port, 
                           A_ns(9) => SHIFT_n_457_port, A_ns(8) => 
                           SHIFT_n_456_port, A_ns(7) => SHIFT_n_455_port, 
                           A_ns(6) => SHIFT_n_454_port, A_ns(5) => 
                           SHIFT_n_453_port, A_ns(4) => SHIFT_n_452_port, 
                           A_ns(3) => SHIFT_n_451_port, A_ns(2) => 
                           SHIFT_n_450_port, A_ns(1) => SHIFT_n_449_port, 
                           A_ns(0) => SHIFT_n_448_port, A_s(63) => 
                           SHIFT_511_port, A_s(62) => SHIFT_510_port, A_s(61) 
                           => SHIFT_509_port, A_s(60) => SHIFT_508_port, 
                           A_s(59) => SHIFT_507_port, A_s(58) => SHIFT_506_port
                           , A_s(57) => SHIFT_505_port, A_s(56) => 
                           SHIFT_504_port, A_s(55) => SHIFT_503_port, A_s(54) 
                           => SHIFT_502_port, A_s(53) => SHIFT_501_port, 
                           A_s(52) => SHIFT_500_port, A_s(51) => SHIFT_499_port
                           , A_s(50) => SHIFT_498_port, A_s(49) => 
                           SHIFT_497_port, A_s(48) => SHIFT_496_port, A_s(47) 
                           => SHIFT_495_port, A_s(46) => SHIFT_494_port, 
                           A_s(45) => SHIFT_493_port, A_s(44) => SHIFT_492_port
                           , A_s(43) => SHIFT_491_port, A_s(42) => 
                           SHIFT_490_port, A_s(41) => SHIFT_489_port, A_s(40) 
                           => SHIFT_488_port, A_s(39) => SHIFT_487_port, 
                           A_s(38) => SHIFT_486_port, A_s(37) => SHIFT_485_port
                           , A_s(36) => SHIFT_484_port, A_s(35) => 
                           SHIFT_483_port, A_s(34) => SHIFT_482_port, A_s(33) 
                           => SHIFT_481_port, A_s(32) => SHIFT_480_port, 
                           A_s(31) => SHIFT_479_port, A_s(30) => SHIFT_478_port
                           , A_s(29) => SHIFT_477_port, A_s(28) => 
                           SHIFT_476_port, A_s(27) => SHIFT_475_port, A_s(26) 
                           => SHIFT_474_port, A_s(25) => SHIFT_473_port, 
                           A_s(24) => SHIFT_472_port, A_s(23) => SHIFT_471_port
                           , A_s(22) => SHIFT_470_port, A_s(21) => 
                           SHIFT_469_port, A_s(20) => SHIFT_468_port, A_s(19) 
                           => SHIFT_467_port, A_s(18) => SHIFT_466_port, 
                           A_s(17) => SHIFT_465_port, A_s(16) => SHIFT_464_port
                           , A_s(15) => SHIFT_463_port, A_s(14) => 
                           SHIFT_462_port, A_s(13) => SHIFT_461_port, A_s(12) 
                           => SHIFT_460_port, A_s(11) => SHIFT_459_port, 
                           A_s(10) => SHIFT_458_port, A_s(9) => SHIFT_457_port,
                           A_s(8) => SHIFT_456_port, A_s(7) => SHIFT_455_port, 
                           A_s(6) => SHIFT_454_port, A_s(5) => SHIFT_453_port, 
                           A_s(4) => SHIFT_452_port, A_s(3) => SHIFT_451_port, 
                           A_s(2) => SHIFT_450_port, A_s(1) => SHIFT_449_port, 
                           A_s(0) => SHIFT_448_port, B(63) => B(31), B(62) => 
                           B(31), B(61) => B(31), B(60) => B(31), B(59) => 
                           B(31), B(58) => B(31), B(57) => B(31), B(56) => 
                           B(31), B(55) => B(31), B(54) => B(31), B(53) => 
                           B(31), B(52) => B(31), B(51) => B(31), B(50) => 
                           B(31), B(49) => B(31), B(48) => B(31), B(47) => 
                           B(31), B(46) => B(31), B(45) => B(31), B(44) => 
                           B(31), B(43) => B(31), B(42) => B(31), B(41) => 
                           B(31), B(40) => B(31), B(39) => B(31), B(38) => 
                           B(31), B(37) => B(31), B(36) => B(31), B(35) => 
                           B(31), B(34) => B(31), B(33) => B(31), B(32) => 
                           B(31), B(31) => B(31), B(30) => B(30), B(29) => 
                           B(29), B(28) => B(28), B(27) => B(27), B(26) => 
                           B(26), B(25) => B(25), B(24) => B(24), B(23) => 
                           B(23), B(22) => B(22), B(21) => B(21), B(20) => 
                           B(20), B(19) => B(19), B(18) => B(18), B(17) => 
                           B(17), B(16) => B(16), B(15) => B(15), B(14) => 
                           B(14), B(13) => B(13), B(12) => B(12), B(11) => 
                           B(11), B(10) => B(10), B(9) => B(9), B(8) => B(8), 
                           B(7) => B(7), B(6) => B(6), B(5) => B(5), B(4) => 
                           B(4), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), O(63) => OTMP_511_port, O(62) => 
                           OTMP_510_port, O(61) => OTMP_509_port, O(60) => 
                           OTMP_508_port, O(59) => OTMP_507_port, O(58) => 
                           OTMP_506_port, O(57) => OTMP_505_port, O(56) => 
                           OTMP_504_port, O(55) => OTMP_503_port, O(54) => 
                           OTMP_502_port, O(53) => OTMP_501_port, O(52) => 
                           OTMP_500_port, O(51) => OTMP_499_port, O(50) => 
                           OTMP_498_port, O(49) => OTMP_497_port, O(48) => 
                           OTMP_496_port, O(47) => OTMP_495_port, O(46) => 
                           OTMP_494_port, O(45) => OTMP_493_port, O(44) => 
                           OTMP_492_port, O(43) => OTMP_491_port, O(42) => 
                           OTMP_490_port, O(41) => OTMP_489_port, O(40) => 
                           OTMP_488_port, O(39) => OTMP_487_port, O(38) => 
                           OTMP_486_port, O(37) => OTMP_485_port, O(36) => 
                           OTMP_484_port, O(35) => OTMP_483_port, O(34) => 
                           OTMP_482_port, O(33) => OTMP_481_port, O(32) => 
                           OTMP_480_port, O(31) => OTMP_479_port, O(30) => 
                           OTMP_478_port, O(29) => OTMP_477_port, O(28) => 
                           OTMP_476_port, O(27) => OTMP_475_port, O(26) => 
                           OTMP_474_port, O(25) => OTMP_473_port, O(24) => 
                           OTMP_472_port, O(23) => OTMP_471_port, O(22) => 
                           OTMP_470_port, O(21) => OTMP_469_port, O(20) => 
                           OTMP_468_port, O(19) => OTMP_467_port, O(18) => 
                           OTMP_466_port, O(17) => OTMP_465_port, O(16) => 
                           OTMP_464_port, O(15) => OTMP_463_port, O(14) => 
                           OTMP_462_port, O(13) => OTMP_461_port, O(12) => 
                           OTMP_460_port, O(11) => OTMP_459_port, O(10) => 
                           OTMP_458_port, O(9) => OTMP_457_port, O(8) => 
                           OTMP_456_port, O(7) => OTMP_455_port, O(6) => 
                           OTMP_454_port, O(5) => OTMP_453_port, O(4) => 
                           OTMP_452_port, O(3) => OTMP_451_port, O(2) => 
                           OTMP_450_port, O(1) => OTMP_449_port, O(0) => n_1126
                           , A_so(63) => SHIFT_575_port, A_so(62) => 
                           SHIFT_574_port, A_so(61) => SHIFT_573_port, A_so(60)
                           => SHIFT_572_port, A_so(59) => SHIFT_571_port, 
                           A_so(58) => SHIFT_570_port, A_so(57) => 
                           SHIFT_569_port, A_so(56) => SHIFT_568_port, A_so(55)
                           => SHIFT_567_port, A_so(54) => SHIFT_566_port, 
                           A_so(53) => SHIFT_565_port, A_so(52) => 
                           SHIFT_564_port, A_so(51) => SHIFT_563_port, A_so(50)
                           => SHIFT_562_port, A_so(49) => SHIFT_561_port, 
                           A_so(48) => SHIFT_560_port, A_so(47) => 
                           SHIFT_559_port, A_so(46) => SHIFT_558_port, A_so(45)
                           => SHIFT_557_port, A_so(44) => SHIFT_556_port, 
                           A_so(43) => SHIFT_555_port, A_so(42) => 
                           SHIFT_554_port, A_so(41) => SHIFT_553_port, A_so(40)
                           => SHIFT_552_port, A_so(39) => SHIFT_551_port, 
                           A_so(38) => SHIFT_550_port, A_so(37) => 
                           SHIFT_549_port, A_so(36) => SHIFT_548_port, A_so(35)
                           => SHIFT_547_port, A_so(34) => SHIFT_546_port, 
                           A_so(33) => SHIFT_545_port, A_so(32) => 
                           SHIFT_544_port, A_so(31) => SHIFT_543_port, A_so(30)
                           => SHIFT_542_port, A_so(29) => SHIFT_541_port, 
                           A_so(28) => SHIFT_540_port, A_so(27) => 
                           SHIFT_539_port, A_so(26) => SHIFT_538_port, A_so(25)
                           => SHIFT_537_port, A_so(24) => SHIFT_536_port, 
                           A_so(23) => SHIFT_535_port, A_so(22) => 
                           SHIFT_534_port, A_so(21) => SHIFT_533_port, A_so(20)
                           => SHIFT_532_port, A_so(19) => SHIFT_531_port, 
                           A_so(18) => SHIFT_530_port, A_so(17) => 
                           SHIFT_529_port, A_so(16) => SHIFT_528_port, A_so(15)
                           => SHIFT_527_port, A_so(14) => SHIFT_526_port, 
                           A_so(13) => SHIFT_525_port, A_so(12) => 
                           SHIFT_524_port, A_so(11) => SHIFT_523_port, A_so(10)
                           => SHIFT_522_port, A_so(9) => SHIFT_521_port, 
                           A_so(8) => SHIFT_520_port, A_so(7) => SHIFT_519_port
                           , A_so(6) => SHIFT_518_port, A_so(5) => 
                           SHIFT_517_port, A_so(4) => SHIFT_516_port, A_so(3) 
                           => SHIFT_515_port, A_so(2) => SHIFT_514_port, 
                           A_so(1) => n_1127, A_so(0) => n_1128, A_nso(63) => 
                           SHIFT_n_575_port, A_nso(62) => SHIFT_n_574_port, 
                           A_nso(61) => SHIFT_n_573_port, A_nso(60) => 
                           SHIFT_n_572_port, A_nso(59) => SHIFT_n_571_port, 
                           A_nso(58) => SHIFT_n_570_port, A_nso(57) => 
                           SHIFT_n_569_port, A_nso(56) => SHIFT_n_568_port, 
                           A_nso(55) => SHIFT_n_567_port, A_nso(54) => 
                           SHIFT_n_566_port, A_nso(53) => SHIFT_n_565_port, 
                           A_nso(52) => SHIFT_n_564_port, A_nso(51) => 
                           SHIFT_n_563_port, A_nso(50) => SHIFT_n_562_port, 
                           A_nso(49) => SHIFT_n_561_port, A_nso(48) => 
                           SHIFT_n_560_port, A_nso(47) => SHIFT_n_559_port, 
                           A_nso(46) => SHIFT_n_558_port, A_nso(45) => 
                           SHIFT_n_557_port, A_nso(44) => SHIFT_n_556_port, 
                           A_nso(43) => SHIFT_n_555_port, A_nso(42) => 
                           SHIFT_n_554_port, A_nso(41) => SHIFT_n_553_port, 
                           A_nso(40) => SHIFT_n_552_port, A_nso(39) => 
                           SHIFT_n_551_port, A_nso(38) => SHIFT_n_550_port, 
                           A_nso(37) => SHIFT_n_549_port, A_nso(36) => 
                           SHIFT_n_548_port, A_nso(35) => SHIFT_n_547_port, 
                           A_nso(34) => SHIFT_n_546_port, A_nso(33) => 
                           SHIFT_n_545_port, A_nso(32) => SHIFT_n_544_port, 
                           A_nso(31) => SHIFT_n_543_port, A_nso(30) => 
                           SHIFT_n_542_port, A_nso(29) => SHIFT_n_541_port, 
                           A_nso(28) => SHIFT_n_540_port, A_nso(27) => 
                           SHIFT_n_539_port, A_nso(26) => SHIFT_n_538_port, 
                           A_nso(25) => SHIFT_n_537_port, A_nso(24) => 
                           SHIFT_n_536_port, A_nso(23) => SHIFT_n_535_port, 
                           A_nso(22) => SHIFT_n_534_port, A_nso(21) => 
                           SHIFT_n_533_port, A_nso(20) => SHIFT_n_532_port, 
                           A_nso(19) => SHIFT_n_531_port, A_nso(18) => 
                           SHIFT_n_530_port, A_nso(17) => SHIFT_n_529_port, 
                           A_nso(16) => SHIFT_n_528_port, A_nso(15) => 
                           SHIFT_n_527_port, A_nso(14) => SHIFT_n_526_port, 
                           A_nso(13) => SHIFT_n_525_port, A_nso(12) => 
                           SHIFT_n_524_port, A_nso(11) => SHIFT_n_523_port, 
                           A_nso(10) => SHIFT_n_522_port, A_nso(9) => 
                           SHIFT_n_521_port, A_nso(8) => SHIFT_n_520_port, 
                           A_nso(7) => SHIFT_n_519_port, A_nso(6) => 
                           SHIFT_n_518_port, A_nso(5) => SHIFT_n_517_port, 
                           A_nso(4) => SHIFT_n_516_port, A_nso(3) => 
                           SHIFT_n_515_port, A_nso(2) => SHIFT_n_514_port, 
                           A_nso(1) => n_1129, A_nso(0) => n_1130);
   BOOTHENC_I_9 : BOOTHENC_NBIT64_i16 port map( A(63) => net47668, A(62) => 
                           net47669, A(61) => net47670, A(60) => net47671, 
                           A(59) => net47672, A(58) => net47673, A(57) => 
                           net47674, A(56) => net47675, A(55) => net47676, 
                           A(54) => net47677, A(53) => net47678, A(52) => 
                           net47679, A(51) => net47680, A(50) => net47681, 
                           A(49) => net47682, A(48) => net47683, A(47) => 
                           net47684, A(46) => net47685, A(45) => net47686, 
                           A(44) => net47687, A(43) => net47688, A(42) => 
                           net47689, A(41) => net47690, A(40) => net47691, 
                           A(39) => net47692, A(38) => net47693, A(37) => 
                           net47694, A(36) => net47695, A(35) => net47696, 
                           A(34) => net47697, A(33) => net47698, A(32) => 
                           net47699, A(31) => net47700, A(30) => net47701, 
                           A(29) => net47702, A(28) => net47703, A(27) => 
                           net47704, A(26) => net47705, A(25) => net47706, 
                           A(24) => net47707, A(23) => net47708, A(22) => 
                           net47709, A(21) => net47710, A(20) => net47711, 
                           A(19) => net47712, A(18) => net47713, A(17) => 
                           net47714, A(16) => net47715, A(15) => net47716, 
                           A(14) => net47717, A(13) => net47718, A(12) => 
                           net47719, A(11) => net47720, A(10) => net47721, A(9)
                           => net47722, A(8) => net47723, A(7) => net47724, 
                           A(6) => net47725, A(5) => net47726, A(4) => net47727
                           , A(3) => net47728, A(2) => net47729, A(1) => 
                           net47730, A(0) => net47731, A_n(63) => net47732, 
                           A_n(62) => net47733, A_n(61) => net47734, A_n(60) =>
                           net47735, A_n(59) => net47736, A_n(58) => net47737, 
                           A_n(57) => net47738, A_n(56) => net47739, A_n(55) =>
                           net47740, A_n(54) => net47741, A_n(53) => net47742, 
                           A_n(52) => net47743, A_n(51) => net47744, A_n(50) =>
                           net47745, A_n(49) => net47746, A_n(48) => net47747, 
                           A_n(47) => net47748, A_n(46) => net47749, A_n(45) =>
                           net47750, A_n(44) => net47751, A_n(43) => net47752, 
                           A_n(42) => net47753, A_n(41) => net47754, A_n(40) =>
                           net47755, A_n(39) => net47756, A_n(38) => net47757, 
                           A_n(37) => net47758, A_n(36) => net47759, A_n(35) =>
                           net47760, A_n(34) => net47761, A_n(33) => net47762, 
                           A_n(32) => net47763, A_n(31) => net47764, A_n(30) =>
                           net47765, A_n(29) => net47766, A_n(28) => net47767, 
                           A_n(27) => net47768, A_n(26) => net47769, A_n(25) =>
                           net47770, A_n(24) => net47771, A_n(23) => net47772, 
                           A_n(22) => net47773, A_n(21) => net47774, A_n(20) =>
                           net47775, A_n(19) => net47776, A_n(18) => net47777, 
                           A_n(17) => net47778, A_n(16) => net47779, A_n(15) =>
                           net47780, A_n(14) => net47781, A_n(13) => net47782, 
                           A_n(12) => net47783, A_n(11) => net47784, A_n(10) =>
                           net47785, A_n(9) => net47786, A_n(8) => net47787, 
                           A_n(7) => net47788, A_n(6) => net47789, A_n(5) => 
                           net47790, A_n(4) => net47791, A_n(3) => net47792, 
                           A_n(2) => net47793, A_n(1) => net47794, A_n(0) => 
                           net47795, A_ns(63) => SHIFT_n_575_port, A_ns(62) => 
                           SHIFT_n_574_port, A_ns(61) => SHIFT_n_573_port, 
                           A_ns(60) => SHIFT_n_572_port, A_ns(59) => 
                           SHIFT_n_571_port, A_ns(58) => SHIFT_n_570_port, 
                           A_ns(57) => SHIFT_n_569_port, A_ns(56) => 
                           SHIFT_n_568_port, A_ns(55) => SHIFT_n_567_port, 
                           A_ns(54) => SHIFT_n_566_port, A_ns(53) => 
                           SHIFT_n_565_port, A_ns(52) => SHIFT_n_564_port, 
                           A_ns(51) => SHIFT_n_563_port, A_ns(50) => 
                           SHIFT_n_562_port, A_ns(49) => SHIFT_n_561_port, 
                           A_ns(48) => SHIFT_n_560_port, A_ns(47) => 
                           SHIFT_n_559_port, A_ns(46) => SHIFT_n_558_port, 
                           A_ns(45) => SHIFT_n_557_port, A_ns(44) => 
                           SHIFT_n_556_port, A_ns(43) => SHIFT_n_555_port, 
                           A_ns(42) => SHIFT_n_554_port, A_ns(41) => 
                           SHIFT_n_553_port, A_ns(40) => SHIFT_n_552_port, 
                           A_ns(39) => SHIFT_n_551_port, A_ns(38) => 
                           SHIFT_n_550_port, A_ns(37) => SHIFT_n_549_port, 
                           A_ns(36) => SHIFT_n_548_port, A_ns(35) => 
                           SHIFT_n_547_port, A_ns(34) => SHIFT_n_546_port, 
                           A_ns(33) => SHIFT_n_545_port, A_ns(32) => 
                           SHIFT_n_544_port, A_ns(31) => SHIFT_n_543_port, 
                           A_ns(30) => SHIFT_n_542_port, A_ns(29) => 
                           SHIFT_n_541_port, A_ns(28) => SHIFT_n_540_port, 
                           A_ns(27) => SHIFT_n_539_port, A_ns(26) => 
                           SHIFT_n_538_port, A_ns(25) => SHIFT_n_537_port, 
                           A_ns(24) => SHIFT_n_536_port, A_ns(23) => 
                           SHIFT_n_535_port, A_ns(22) => SHIFT_n_534_port, 
                           A_ns(21) => SHIFT_n_533_port, A_ns(20) => 
                           SHIFT_n_532_port, A_ns(19) => SHIFT_n_531_port, 
                           A_ns(18) => SHIFT_n_530_port, A_ns(17) => 
                           SHIFT_n_529_port, A_ns(16) => SHIFT_n_528_port, 
                           A_ns(15) => SHIFT_n_527_port, A_ns(14) => 
                           SHIFT_n_526_port, A_ns(13) => SHIFT_n_525_port, 
                           A_ns(12) => SHIFT_n_524_port, A_ns(11) => 
                           SHIFT_n_523_port, A_ns(10) => SHIFT_n_522_port, 
                           A_ns(9) => SHIFT_n_521_port, A_ns(8) => 
                           SHIFT_n_520_port, A_ns(7) => SHIFT_n_519_port, 
                           A_ns(6) => SHIFT_n_518_port, A_ns(5) => 
                           SHIFT_n_517_port, A_ns(4) => SHIFT_n_516_port, 
                           A_ns(3) => SHIFT_n_515_port, A_ns(2) => 
                           SHIFT_n_514_port, A_ns(1) => SHIFT_n_513_port, 
                           A_ns(0) => SHIFT_n_512_port, A_s(63) => 
                           SHIFT_575_port, A_s(62) => SHIFT_574_port, A_s(61) 
                           => SHIFT_573_port, A_s(60) => SHIFT_572_port, 
                           A_s(59) => SHIFT_571_port, A_s(58) => SHIFT_570_port
                           , A_s(57) => SHIFT_569_port, A_s(56) => 
                           SHIFT_568_port, A_s(55) => SHIFT_567_port, A_s(54) 
                           => SHIFT_566_port, A_s(53) => SHIFT_565_port, 
                           A_s(52) => SHIFT_564_port, A_s(51) => SHIFT_563_port
                           , A_s(50) => SHIFT_562_port, A_s(49) => 
                           SHIFT_561_port, A_s(48) => SHIFT_560_port, A_s(47) 
                           => SHIFT_559_port, A_s(46) => SHIFT_558_port, 
                           A_s(45) => SHIFT_557_port, A_s(44) => SHIFT_556_port
                           , A_s(43) => SHIFT_555_port, A_s(42) => 
                           SHIFT_554_port, A_s(41) => SHIFT_553_port, A_s(40) 
                           => SHIFT_552_port, A_s(39) => SHIFT_551_port, 
                           A_s(38) => SHIFT_550_port, A_s(37) => SHIFT_549_port
                           , A_s(36) => SHIFT_548_port, A_s(35) => 
                           SHIFT_547_port, A_s(34) => SHIFT_546_port, A_s(33) 
                           => SHIFT_545_port, A_s(32) => SHIFT_544_port, 
                           A_s(31) => SHIFT_543_port, A_s(30) => SHIFT_542_port
                           , A_s(29) => SHIFT_541_port, A_s(28) => 
                           SHIFT_540_port, A_s(27) => SHIFT_539_port, A_s(26) 
                           => SHIFT_538_port, A_s(25) => SHIFT_537_port, 
                           A_s(24) => SHIFT_536_port, A_s(23) => SHIFT_535_port
                           , A_s(22) => SHIFT_534_port, A_s(21) => 
                           SHIFT_533_port, A_s(20) => SHIFT_532_port, A_s(19) 
                           => SHIFT_531_port, A_s(18) => SHIFT_530_port, 
                           A_s(17) => SHIFT_529_port, A_s(16) => SHIFT_528_port
                           , A_s(15) => SHIFT_527_port, A_s(14) => 
                           SHIFT_526_port, A_s(13) => SHIFT_525_port, A_s(12) 
                           => SHIFT_524_port, A_s(11) => SHIFT_523_port, 
                           A_s(10) => SHIFT_522_port, A_s(9) => SHIFT_521_port,
                           A_s(8) => SHIFT_520_port, A_s(7) => SHIFT_519_port, 
                           A_s(6) => SHIFT_518_port, A_s(5) => SHIFT_517_port, 
                           A_s(4) => SHIFT_516_port, A_s(3) => SHIFT_515_port, 
                           A_s(2) => SHIFT_514_port, A_s(1) => SHIFT_513_port, 
                           A_s(0) => SHIFT_512_port, B(63) => B(31), B(62) => 
                           B(31), B(61) => B(31), B(60) => B(31), B(59) => 
                           B(31), B(58) => B(31), B(57) => B(31), B(56) => 
                           B(31), B(55) => B(31), B(54) => B(31), B(53) => 
                           B(31), B(52) => B(31), B(51) => B(31), B(50) => 
                           B(31), B(49) => B(31), B(48) => B(31), B(47) => 
                           B(31), B(46) => B(31), B(45) => B(31), B(44) => 
                           B(31), B(43) => B(31), B(42) => B(31), B(41) => 
                           B(31), B(40) => B(31), B(39) => B(31), B(38) => 
                           B(31), B(37) => B(31), B(36) => B(31), B(35) => 
                           B(31), B(34) => B(31), B(33) => B(31), B(32) => 
                           B(31), B(31) => B(31), B(30) => B(30), B(29) => 
                           B(29), B(28) => B(28), B(27) => B(27), B(26) => 
                           B(26), B(25) => B(25), B(24) => B(24), B(23) => 
                           B(23), B(22) => B(22), B(21) => B(21), B(20) => 
                           B(20), B(19) => B(19), B(18) => B(18), B(17) => 
                           B(17), B(16) => B(16), B(15) => B(15), B(14) => 
                           B(14), B(13) => B(13), B(12) => B(12), B(11) => 
                           B(11), B(10) => B(10), B(9) => B(9), B(8) => B(8), 
                           B(7) => B(7), B(6) => B(6), B(5) => B(5), B(4) => 
                           B(4), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), O(63) => OTMP_575_port, O(62) => 
                           OTMP_574_port, O(61) => OTMP_573_port, O(60) => 
                           OTMP_572_port, O(59) => OTMP_571_port, O(58) => 
                           OTMP_570_port, O(57) => OTMP_569_port, O(56) => 
                           OTMP_568_port, O(55) => OTMP_567_port, O(54) => 
                           OTMP_566_port, O(53) => OTMP_565_port, O(52) => 
                           OTMP_564_port, O(51) => OTMP_563_port, O(50) => 
                           OTMP_562_port, O(49) => OTMP_561_port, O(48) => 
                           OTMP_560_port, O(47) => OTMP_559_port, O(46) => 
                           OTMP_558_port, O(45) => OTMP_557_port, O(44) => 
                           OTMP_556_port, O(43) => OTMP_555_port, O(42) => 
                           OTMP_554_port, O(41) => OTMP_553_port, O(40) => 
                           OTMP_552_port, O(39) => OTMP_551_port, O(38) => 
                           OTMP_550_port, O(37) => OTMP_549_port, O(36) => 
                           OTMP_548_port, O(35) => OTMP_547_port, O(34) => 
                           OTMP_546_port, O(33) => OTMP_545_port, O(32) => 
                           OTMP_544_port, O(31) => OTMP_543_port, O(30) => 
                           OTMP_542_port, O(29) => OTMP_541_port, O(28) => 
                           OTMP_540_port, O(27) => OTMP_539_port, O(26) => 
                           OTMP_538_port, O(25) => OTMP_537_port, O(24) => 
                           OTMP_536_port, O(23) => OTMP_535_port, O(22) => 
                           OTMP_534_port, O(21) => OTMP_533_port, O(20) => 
                           OTMP_532_port, O(19) => OTMP_531_port, O(18) => 
                           OTMP_530_port, O(17) => OTMP_529_port, O(16) => 
                           OTMP_528_port, O(15) => OTMP_527_port, O(14) => 
                           OTMP_526_port, O(13) => OTMP_525_port, O(12) => 
                           OTMP_524_port, O(11) => OTMP_523_port, O(10) => 
                           OTMP_522_port, O(9) => OTMP_521_port, O(8) => 
                           OTMP_520_port, O(7) => OTMP_519_port, O(6) => 
                           OTMP_518_port, O(5) => OTMP_517_port, O(4) => 
                           OTMP_516_port, O(3) => OTMP_515_port, O(2) => 
                           OTMP_514_port, O(1) => OTMP_513_port, O(0) => n_1131
                           , A_so(63) => SHIFT_639_port, A_so(62) => 
                           SHIFT_638_port, A_so(61) => SHIFT_637_port, A_so(60)
                           => SHIFT_636_port, A_so(59) => SHIFT_635_port, 
                           A_so(58) => SHIFT_634_port, A_so(57) => 
                           SHIFT_633_port, A_so(56) => SHIFT_632_port, A_so(55)
                           => SHIFT_631_port, A_so(54) => SHIFT_630_port, 
                           A_so(53) => SHIFT_629_port, A_so(52) => 
                           SHIFT_628_port, A_so(51) => SHIFT_627_port, A_so(50)
                           => SHIFT_626_port, A_so(49) => SHIFT_625_port, 
                           A_so(48) => SHIFT_624_port, A_so(47) => 
                           SHIFT_623_port, A_so(46) => SHIFT_622_port, A_so(45)
                           => SHIFT_621_port, A_so(44) => SHIFT_620_port, 
                           A_so(43) => SHIFT_619_port, A_so(42) => 
                           SHIFT_618_port, A_so(41) => SHIFT_617_port, A_so(40)
                           => SHIFT_616_port, A_so(39) => SHIFT_615_port, 
                           A_so(38) => SHIFT_614_port, A_so(37) => 
                           SHIFT_613_port, A_so(36) => SHIFT_612_port, A_so(35)
                           => SHIFT_611_port, A_so(34) => SHIFT_610_port, 
                           A_so(33) => SHIFT_609_port, A_so(32) => 
                           SHIFT_608_port, A_so(31) => SHIFT_607_port, A_so(30)
                           => SHIFT_606_port, A_so(29) => SHIFT_605_port, 
                           A_so(28) => SHIFT_604_port, A_so(27) => 
                           SHIFT_603_port, A_so(26) => SHIFT_602_port, A_so(25)
                           => SHIFT_601_port, A_so(24) => SHIFT_600_port, 
                           A_so(23) => SHIFT_599_port, A_so(22) => 
                           SHIFT_598_port, A_so(21) => SHIFT_597_port, A_so(20)
                           => SHIFT_596_port, A_so(19) => SHIFT_595_port, 
                           A_so(18) => SHIFT_594_port, A_so(17) => 
                           SHIFT_593_port, A_so(16) => SHIFT_592_port, A_so(15)
                           => SHIFT_591_port, A_so(14) => SHIFT_590_port, 
                           A_so(13) => SHIFT_589_port, A_so(12) => 
                           SHIFT_588_port, A_so(11) => SHIFT_587_port, A_so(10)
                           => SHIFT_586_port, A_so(9) => SHIFT_585_port, 
                           A_so(8) => SHIFT_584_port, A_so(7) => SHIFT_583_port
                           , A_so(6) => SHIFT_582_port, A_so(5) => 
                           SHIFT_581_port, A_so(4) => SHIFT_580_port, A_so(3) 
                           => SHIFT_579_port, A_so(2) => SHIFT_578_port, 
                           A_so(1) => n_1132, A_so(0) => n_1133, A_nso(63) => 
                           SHIFT_n_639_port, A_nso(62) => SHIFT_n_638_port, 
                           A_nso(61) => SHIFT_n_637_port, A_nso(60) => 
                           SHIFT_n_636_port, A_nso(59) => SHIFT_n_635_port, 
                           A_nso(58) => SHIFT_n_634_port, A_nso(57) => 
                           SHIFT_n_633_port, A_nso(56) => SHIFT_n_632_port, 
                           A_nso(55) => SHIFT_n_631_port, A_nso(54) => 
                           SHIFT_n_630_port, A_nso(53) => SHIFT_n_629_port, 
                           A_nso(52) => SHIFT_n_628_port, A_nso(51) => 
                           SHIFT_n_627_port, A_nso(50) => SHIFT_n_626_port, 
                           A_nso(49) => SHIFT_n_625_port, A_nso(48) => 
                           SHIFT_n_624_port, A_nso(47) => SHIFT_n_623_port, 
                           A_nso(46) => SHIFT_n_622_port, A_nso(45) => 
                           SHIFT_n_621_port, A_nso(44) => SHIFT_n_620_port, 
                           A_nso(43) => SHIFT_n_619_port, A_nso(42) => 
                           SHIFT_n_618_port, A_nso(41) => SHIFT_n_617_port, 
                           A_nso(40) => SHIFT_n_616_port, A_nso(39) => 
                           SHIFT_n_615_port, A_nso(38) => SHIFT_n_614_port, 
                           A_nso(37) => SHIFT_n_613_port, A_nso(36) => 
                           SHIFT_n_612_port, A_nso(35) => SHIFT_n_611_port, 
                           A_nso(34) => SHIFT_n_610_port, A_nso(33) => 
                           SHIFT_n_609_port, A_nso(32) => SHIFT_n_608_port, 
                           A_nso(31) => SHIFT_n_607_port, A_nso(30) => 
                           SHIFT_n_606_port, A_nso(29) => SHIFT_n_605_port, 
                           A_nso(28) => SHIFT_n_604_port, A_nso(27) => 
                           SHIFT_n_603_port, A_nso(26) => SHIFT_n_602_port, 
                           A_nso(25) => SHIFT_n_601_port, A_nso(24) => 
                           SHIFT_n_600_port, A_nso(23) => SHIFT_n_599_port, 
                           A_nso(22) => SHIFT_n_598_port, A_nso(21) => 
                           SHIFT_n_597_port, A_nso(20) => SHIFT_n_596_port, 
                           A_nso(19) => SHIFT_n_595_port, A_nso(18) => 
                           SHIFT_n_594_port, A_nso(17) => SHIFT_n_593_port, 
                           A_nso(16) => SHIFT_n_592_port, A_nso(15) => 
                           SHIFT_n_591_port, A_nso(14) => SHIFT_n_590_port, 
                           A_nso(13) => SHIFT_n_589_port, A_nso(12) => 
                           SHIFT_n_588_port, A_nso(11) => SHIFT_n_587_port, 
                           A_nso(10) => SHIFT_n_586_port, A_nso(9) => 
                           SHIFT_n_585_port, A_nso(8) => SHIFT_n_584_port, 
                           A_nso(7) => SHIFT_n_583_port, A_nso(6) => 
                           SHIFT_n_582_port, A_nso(5) => SHIFT_n_581_port, 
                           A_nso(4) => SHIFT_n_580_port, A_nso(3) => 
                           SHIFT_n_579_port, A_nso(2) => SHIFT_n_578_port, 
                           A_nso(1) => n_1134, A_nso(0) => n_1135);
   BOOTHENC_I_10 : BOOTHENC_NBIT64_i18 port map( A(63) => net47540, A(62) => 
                           net47541, A(61) => net47542, A(60) => net47543, 
                           A(59) => net47544, A(58) => net47545, A(57) => 
                           net47546, A(56) => net47547, A(55) => net47548, 
                           A(54) => net47549, A(53) => net47550, A(52) => 
                           net47551, A(51) => net47552, A(50) => net47553, 
                           A(49) => net47554, A(48) => net47555, A(47) => 
                           net47556, A(46) => net47557, A(45) => net47558, 
                           A(44) => net47559, A(43) => net47560, A(42) => 
                           net47561, A(41) => net47562, A(40) => net47563, 
                           A(39) => net47564, A(38) => net47565, A(37) => 
                           net47566, A(36) => net47567, A(35) => net47568, 
                           A(34) => net47569, A(33) => net47570, A(32) => 
                           net47571, A(31) => net47572, A(30) => net47573, 
                           A(29) => net47574, A(28) => net47575, A(27) => 
                           net47576, A(26) => net47577, A(25) => net47578, 
                           A(24) => net47579, A(23) => net47580, A(22) => 
                           net47581, A(21) => net47582, A(20) => net47583, 
                           A(19) => net47584, A(18) => net47585, A(17) => 
                           net47586, A(16) => net47587, A(15) => net47588, 
                           A(14) => net47589, A(13) => net47590, A(12) => 
                           net47591, A(11) => net47592, A(10) => net47593, A(9)
                           => net47594, A(8) => net47595, A(7) => net47596, 
                           A(6) => net47597, A(5) => net47598, A(4) => net47599
                           , A(3) => net47600, A(2) => net47601, A(1) => 
                           net47602, A(0) => net47603, A_n(63) => net47604, 
                           A_n(62) => net47605, A_n(61) => net47606, A_n(60) =>
                           net47607, A_n(59) => net47608, A_n(58) => net47609, 
                           A_n(57) => net47610, A_n(56) => net47611, A_n(55) =>
                           net47612, A_n(54) => net47613, A_n(53) => net47614, 
                           A_n(52) => net47615, A_n(51) => net47616, A_n(50) =>
                           net47617, A_n(49) => net47618, A_n(48) => net47619, 
                           A_n(47) => net47620, A_n(46) => net47621, A_n(45) =>
                           net47622, A_n(44) => net47623, A_n(43) => net47624, 
                           A_n(42) => net47625, A_n(41) => net47626, A_n(40) =>
                           net47627, A_n(39) => net47628, A_n(38) => net47629, 
                           A_n(37) => net47630, A_n(36) => net47631, A_n(35) =>
                           net47632, A_n(34) => net47633, A_n(33) => net47634, 
                           A_n(32) => net47635, A_n(31) => net47636, A_n(30) =>
                           net47637, A_n(29) => net47638, A_n(28) => net47639, 
                           A_n(27) => net47640, A_n(26) => net47641, A_n(25) =>
                           net47642, A_n(24) => net47643, A_n(23) => net47644, 
                           A_n(22) => net47645, A_n(21) => net47646, A_n(20) =>
                           net47647, A_n(19) => net47648, A_n(18) => net47649, 
                           A_n(17) => net47650, A_n(16) => net47651, A_n(15) =>
                           net47652, A_n(14) => net47653, A_n(13) => net47654, 
                           A_n(12) => net47655, A_n(11) => net47656, A_n(10) =>
                           net47657, A_n(9) => net47658, A_n(8) => net47659, 
                           A_n(7) => net47660, A_n(6) => net47661, A_n(5) => 
                           net47662, A_n(4) => net47663, A_n(3) => net47664, 
                           A_n(2) => net47665, A_n(1) => net47666, A_n(0) => 
                           net47667, A_ns(63) => SHIFT_n_639_port, A_ns(62) => 
                           SHIFT_n_638_port, A_ns(61) => SHIFT_n_637_port, 
                           A_ns(60) => SHIFT_n_636_port, A_ns(59) => 
                           SHIFT_n_635_port, A_ns(58) => SHIFT_n_634_port, 
                           A_ns(57) => SHIFT_n_633_port, A_ns(56) => 
                           SHIFT_n_632_port, A_ns(55) => SHIFT_n_631_port, 
                           A_ns(54) => SHIFT_n_630_port, A_ns(53) => 
                           SHIFT_n_629_port, A_ns(52) => SHIFT_n_628_port, 
                           A_ns(51) => SHIFT_n_627_port, A_ns(50) => 
                           SHIFT_n_626_port, A_ns(49) => SHIFT_n_625_port, 
                           A_ns(48) => SHIFT_n_624_port, A_ns(47) => 
                           SHIFT_n_623_port, A_ns(46) => SHIFT_n_622_port, 
                           A_ns(45) => SHIFT_n_621_port, A_ns(44) => 
                           SHIFT_n_620_port, A_ns(43) => SHIFT_n_619_port, 
                           A_ns(42) => SHIFT_n_618_port, A_ns(41) => 
                           SHIFT_n_617_port, A_ns(40) => SHIFT_n_616_port, 
                           A_ns(39) => SHIFT_n_615_port, A_ns(38) => 
                           SHIFT_n_614_port, A_ns(37) => SHIFT_n_613_port, 
                           A_ns(36) => SHIFT_n_612_port, A_ns(35) => 
                           SHIFT_n_611_port, A_ns(34) => SHIFT_n_610_port, 
                           A_ns(33) => SHIFT_n_609_port, A_ns(32) => 
                           SHIFT_n_608_port, A_ns(31) => SHIFT_n_607_port, 
                           A_ns(30) => SHIFT_n_606_port, A_ns(29) => 
                           SHIFT_n_605_port, A_ns(28) => SHIFT_n_604_port, 
                           A_ns(27) => SHIFT_n_603_port, A_ns(26) => 
                           SHIFT_n_602_port, A_ns(25) => SHIFT_n_601_port, 
                           A_ns(24) => SHIFT_n_600_port, A_ns(23) => 
                           SHIFT_n_599_port, A_ns(22) => SHIFT_n_598_port, 
                           A_ns(21) => SHIFT_n_597_port, A_ns(20) => 
                           SHIFT_n_596_port, A_ns(19) => SHIFT_n_595_port, 
                           A_ns(18) => SHIFT_n_594_port, A_ns(17) => 
                           SHIFT_n_593_port, A_ns(16) => SHIFT_n_592_port, 
                           A_ns(15) => SHIFT_n_591_port, A_ns(14) => 
                           SHIFT_n_590_port, A_ns(13) => SHIFT_n_589_port, 
                           A_ns(12) => SHIFT_n_588_port, A_ns(11) => 
                           SHIFT_n_587_port, A_ns(10) => SHIFT_n_586_port, 
                           A_ns(9) => SHIFT_n_585_port, A_ns(8) => 
                           SHIFT_n_584_port, A_ns(7) => SHIFT_n_583_port, 
                           A_ns(6) => SHIFT_n_582_port, A_ns(5) => 
                           SHIFT_n_581_port, A_ns(4) => SHIFT_n_580_port, 
                           A_ns(3) => SHIFT_n_579_port, A_ns(2) => 
                           SHIFT_n_578_port, A_ns(1) => SHIFT_n_577_port, 
                           A_ns(0) => SHIFT_n_576_port, A_s(63) => 
                           SHIFT_639_port, A_s(62) => SHIFT_638_port, A_s(61) 
                           => SHIFT_637_port, A_s(60) => SHIFT_636_port, 
                           A_s(59) => SHIFT_635_port, A_s(58) => SHIFT_634_port
                           , A_s(57) => SHIFT_633_port, A_s(56) => 
                           SHIFT_632_port, A_s(55) => SHIFT_631_port, A_s(54) 
                           => SHIFT_630_port, A_s(53) => SHIFT_629_port, 
                           A_s(52) => SHIFT_628_port, A_s(51) => SHIFT_627_port
                           , A_s(50) => SHIFT_626_port, A_s(49) => 
                           SHIFT_625_port, A_s(48) => SHIFT_624_port, A_s(47) 
                           => SHIFT_623_port, A_s(46) => SHIFT_622_port, 
                           A_s(45) => SHIFT_621_port, A_s(44) => SHIFT_620_port
                           , A_s(43) => SHIFT_619_port, A_s(42) => 
                           SHIFT_618_port, A_s(41) => SHIFT_617_port, A_s(40) 
                           => SHIFT_616_port, A_s(39) => SHIFT_615_port, 
                           A_s(38) => SHIFT_614_port, A_s(37) => SHIFT_613_port
                           , A_s(36) => SHIFT_612_port, A_s(35) => 
                           SHIFT_611_port, A_s(34) => SHIFT_610_port, A_s(33) 
                           => SHIFT_609_port, A_s(32) => SHIFT_608_port, 
                           A_s(31) => SHIFT_607_port, A_s(30) => SHIFT_606_port
                           , A_s(29) => SHIFT_605_port, A_s(28) => 
                           SHIFT_604_port, A_s(27) => SHIFT_603_port, A_s(26) 
                           => SHIFT_602_port, A_s(25) => SHIFT_601_port, 
                           A_s(24) => SHIFT_600_port, A_s(23) => SHIFT_599_port
                           , A_s(22) => SHIFT_598_port, A_s(21) => 
                           SHIFT_597_port, A_s(20) => SHIFT_596_port, A_s(19) 
                           => SHIFT_595_port, A_s(18) => SHIFT_594_port, 
                           A_s(17) => SHIFT_593_port, A_s(16) => SHIFT_592_port
                           , A_s(15) => SHIFT_591_port, A_s(14) => 
                           SHIFT_590_port, A_s(13) => SHIFT_589_port, A_s(12) 
                           => SHIFT_588_port, A_s(11) => SHIFT_587_port, 
                           A_s(10) => SHIFT_586_port, A_s(9) => SHIFT_585_port,
                           A_s(8) => SHIFT_584_port, A_s(7) => SHIFT_583_port, 
                           A_s(6) => SHIFT_582_port, A_s(5) => SHIFT_581_port, 
                           A_s(4) => SHIFT_580_port, A_s(3) => SHIFT_579_port, 
                           A_s(2) => SHIFT_578_port, A_s(1) => SHIFT_577_port, 
                           A_s(0) => SHIFT_576_port, B(63) => B(31), B(62) => 
                           B(31), B(61) => B(31), B(60) => B(31), B(59) => 
                           B(31), B(58) => B(31), B(57) => B(31), B(56) => 
                           B(31), B(55) => B(31), B(54) => B(31), B(53) => 
                           B(31), B(52) => B(31), B(51) => B(31), B(50) => 
                           B(31), B(49) => B(31), B(48) => B(31), B(47) => 
                           B(31), B(46) => B(31), B(45) => B(31), B(44) => 
                           B(31), B(43) => B(31), B(42) => B(31), B(41) => 
                           B(31), B(40) => B(31), B(39) => B(31), B(38) => 
                           B(31), B(37) => B(31), B(36) => B(31), B(35) => 
                           B(31), B(34) => B(31), B(33) => B(31), B(32) => 
                           B(31), B(31) => B(31), B(30) => B(30), B(29) => 
                           B(29), B(28) => B(28), B(27) => B(27), B(26) => 
                           B(26), B(25) => B(25), B(24) => B(24), B(23) => 
                           B(23), B(22) => B(22), B(21) => B(21), B(20) => 
                           B(20), B(19) => B(19), B(18) => B(18), B(17) => 
                           B(17), B(16) => B(16), B(15) => B(15), B(14) => 
                           B(14), B(13) => B(13), B(12) => B(12), B(11) => 
                           B(11), B(10) => B(10), B(9) => B(9), B(8) => B(8), 
                           B(7) => B(7), B(6) => B(6), B(5) => B(5), B(4) => 
                           B(4), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), O(63) => OTMP_639_port, O(62) => 
                           OTMP_638_port, O(61) => OTMP_637_port, O(60) => 
                           OTMP_636_port, O(59) => OTMP_635_port, O(58) => 
                           OTMP_634_port, O(57) => OTMP_633_port, O(56) => 
                           OTMP_632_port, O(55) => OTMP_631_port, O(54) => 
                           OTMP_630_port, O(53) => OTMP_629_port, O(52) => 
                           OTMP_628_port, O(51) => OTMP_627_port, O(50) => 
                           OTMP_626_port, O(49) => OTMP_625_port, O(48) => 
                           OTMP_624_port, O(47) => OTMP_623_port, O(46) => 
                           OTMP_622_port, O(45) => OTMP_621_port, O(44) => 
                           OTMP_620_port, O(43) => OTMP_619_port, O(42) => 
                           OTMP_618_port, O(41) => OTMP_617_port, O(40) => 
                           OTMP_616_port, O(39) => OTMP_615_port, O(38) => 
                           OTMP_614_port, O(37) => OTMP_613_port, O(36) => 
                           OTMP_612_port, O(35) => OTMP_611_port, O(34) => 
                           OTMP_610_port, O(33) => OTMP_609_port, O(32) => 
                           OTMP_608_port, O(31) => OTMP_607_port, O(30) => 
                           OTMP_606_port, O(29) => OTMP_605_port, O(28) => 
                           OTMP_604_port, O(27) => OTMP_603_port, O(26) => 
                           OTMP_602_port, O(25) => OTMP_601_port, O(24) => 
                           OTMP_600_port, O(23) => OTMP_599_port, O(22) => 
                           OTMP_598_port, O(21) => OTMP_597_port, O(20) => 
                           OTMP_596_port, O(19) => OTMP_595_port, O(18) => 
                           OTMP_594_port, O(17) => OTMP_593_port, O(16) => 
                           OTMP_592_port, O(15) => OTMP_591_port, O(14) => 
                           OTMP_590_port, O(13) => OTMP_589_port, O(12) => 
                           OTMP_588_port, O(11) => OTMP_587_port, O(10) => 
                           OTMP_586_port, O(9) => OTMP_585_port, O(8) => 
                           OTMP_584_port, O(7) => OTMP_583_port, O(6) => 
                           OTMP_582_port, O(5) => OTMP_581_port, O(4) => 
                           OTMP_580_port, O(3) => OTMP_579_port, O(2) => 
                           OTMP_578_port, O(1) => OTMP_577_port, O(0) => n_1136
                           , A_so(63) => SHIFT_703_port, A_so(62) => 
                           SHIFT_702_port, A_so(61) => SHIFT_701_port, A_so(60)
                           => SHIFT_700_port, A_so(59) => SHIFT_699_port, 
                           A_so(58) => SHIFT_698_port, A_so(57) => 
                           SHIFT_697_port, A_so(56) => SHIFT_696_port, A_so(55)
                           => SHIFT_695_port, A_so(54) => SHIFT_694_port, 
                           A_so(53) => SHIFT_693_port, A_so(52) => 
                           SHIFT_692_port, A_so(51) => SHIFT_691_port, A_so(50)
                           => SHIFT_690_port, A_so(49) => SHIFT_689_port, 
                           A_so(48) => SHIFT_688_port, A_so(47) => 
                           SHIFT_687_port, A_so(46) => SHIFT_686_port, A_so(45)
                           => SHIFT_685_port, A_so(44) => SHIFT_684_port, 
                           A_so(43) => SHIFT_683_port, A_so(42) => 
                           SHIFT_682_port, A_so(41) => SHIFT_681_port, A_so(40)
                           => SHIFT_680_port, A_so(39) => SHIFT_679_port, 
                           A_so(38) => SHIFT_678_port, A_so(37) => 
                           SHIFT_677_port, A_so(36) => SHIFT_676_port, A_so(35)
                           => SHIFT_675_port, A_so(34) => SHIFT_674_port, 
                           A_so(33) => SHIFT_673_port, A_so(32) => 
                           SHIFT_672_port, A_so(31) => SHIFT_671_port, A_so(30)
                           => SHIFT_670_port, A_so(29) => SHIFT_669_port, 
                           A_so(28) => SHIFT_668_port, A_so(27) => 
                           SHIFT_667_port, A_so(26) => SHIFT_666_port, A_so(25)
                           => SHIFT_665_port, A_so(24) => SHIFT_664_port, 
                           A_so(23) => SHIFT_663_port, A_so(22) => 
                           SHIFT_662_port, A_so(21) => SHIFT_661_port, A_so(20)
                           => SHIFT_660_port, A_so(19) => SHIFT_659_port, 
                           A_so(18) => SHIFT_658_port, A_so(17) => 
                           SHIFT_657_port, A_so(16) => SHIFT_656_port, A_so(15)
                           => SHIFT_655_port, A_so(14) => SHIFT_654_port, 
                           A_so(13) => SHIFT_653_port, A_so(12) => 
                           SHIFT_652_port, A_so(11) => SHIFT_651_port, A_so(10)
                           => SHIFT_650_port, A_so(9) => SHIFT_649_port, 
                           A_so(8) => SHIFT_648_port, A_so(7) => SHIFT_647_port
                           , A_so(6) => SHIFT_646_port, A_so(5) => 
                           SHIFT_645_port, A_so(4) => SHIFT_644_port, A_so(3) 
                           => SHIFT_643_port, A_so(2) => SHIFT_642_port, 
                           A_so(1) => n_1137, A_so(0) => n_1138, A_nso(63) => 
                           SHIFT_n_703_port, A_nso(62) => SHIFT_n_702_port, 
                           A_nso(61) => SHIFT_n_701_port, A_nso(60) => 
                           SHIFT_n_700_port, A_nso(59) => SHIFT_n_699_port, 
                           A_nso(58) => SHIFT_n_698_port, A_nso(57) => 
                           SHIFT_n_697_port, A_nso(56) => SHIFT_n_696_port, 
                           A_nso(55) => SHIFT_n_695_port, A_nso(54) => 
                           SHIFT_n_694_port, A_nso(53) => SHIFT_n_693_port, 
                           A_nso(52) => SHIFT_n_692_port, A_nso(51) => 
                           SHIFT_n_691_port, A_nso(50) => SHIFT_n_690_port, 
                           A_nso(49) => SHIFT_n_689_port, A_nso(48) => 
                           SHIFT_n_688_port, A_nso(47) => SHIFT_n_687_port, 
                           A_nso(46) => SHIFT_n_686_port, A_nso(45) => 
                           SHIFT_n_685_port, A_nso(44) => SHIFT_n_684_port, 
                           A_nso(43) => SHIFT_n_683_port, A_nso(42) => 
                           SHIFT_n_682_port, A_nso(41) => SHIFT_n_681_port, 
                           A_nso(40) => SHIFT_n_680_port, A_nso(39) => 
                           SHIFT_n_679_port, A_nso(38) => SHIFT_n_678_port, 
                           A_nso(37) => SHIFT_n_677_port, A_nso(36) => 
                           SHIFT_n_676_port, A_nso(35) => SHIFT_n_675_port, 
                           A_nso(34) => SHIFT_n_674_port, A_nso(33) => 
                           SHIFT_n_673_port, A_nso(32) => SHIFT_n_672_port, 
                           A_nso(31) => SHIFT_n_671_port, A_nso(30) => 
                           SHIFT_n_670_port, A_nso(29) => SHIFT_n_669_port, 
                           A_nso(28) => SHIFT_n_668_port, A_nso(27) => 
                           SHIFT_n_667_port, A_nso(26) => SHIFT_n_666_port, 
                           A_nso(25) => SHIFT_n_665_port, A_nso(24) => 
                           SHIFT_n_664_port, A_nso(23) => SHIFT_n_663_port, 
                           A_nso(22) => SHIFT_n_662_port, A_nso(21) => 
                           SHIFT_n_661_port, A_nso(20) => SHIFT_n_660_port, 
                           A_nso(19) => SHIFT_n_659_port, A_nso(18) => 
                           SHIFT_n_658_port, A_nso(17) => SHIFT_n_657_port, 
                           A_nso(16) => SHIFT_n_656_port, A_nso(15) => 
                           SHIFT_n_655_port, A_nso(14) => SHIFT_n_654_port, 
                           A_nso(13) => SHIFT_n_653_port, A_nso(12) => 
                           SHIFT_n_652_port, A_nso(11) => SHIFT_n_651_port, 
                           A_nso(10) => SHIFT_n_650_port, A_nso(9) => 
                           SHIFT_n_649_port, A_nso(8) => SHIFT_n_648_port, 
                           A_nso(7) => SHIFT_n_647_port, A_nso(6) => 
                           SHIFT_n_646_port, A_nso(5) => SHIFT_n_645_port, 
                           A_nso(4) => SHIFT_n_644_port, A_nso(3) => 
                           SHIFT_n_643_port, A_nso(2) => SHIFT_n_642_port, 
                           A_nso(1) => n_1139, A_nso(0) => n_1140);
   BOOTHENC_I_11 : BOOTHENC_NBIT64_i20 port map( A(63) => net47412, A(62) => 
                           net47413, A(61) => net47414, A(60) => net47415, 
                           A(59) => net47416, A(58) => net47417, A(57) => 
                           net47418, A(56) => net47419, A(55) => net47420, 
                           A(54) => net47421, A(53) => net47422, A(52) => 
                           net47423, A(51) => net47424, A(50) => net47425, 
                           A(49) => net47426, A(48) => net47427, A(47) => 
                           net47428, A(46) => net47429, A(45) => net47430, 
                           A(44) => net47431, A(43) => net47432, A(42) => 
                           net47433, A(41) => net47434, A(40) => net47435, 
                           A(39) => net47436, A(38) => net47437, A(37) => 
                           net47438, A(36) => net47439, A(35) => net47440, 
                           A(34) => net47441, A(33) => net47442, A(32) => 
                           net47443, A(31) => net47444, A(30) => net47445, 
                           A(29) => net47446, A(28) => net47447, A(27) => 
                           net47448, A(26) => net47449, A(25) => net47450, 
                           A(24) => net47451, A(23) => net47452, A(22) => 
                           net47453, A(21) => net47454, A(20) => net47455, 
                           A(19) => net47456, A(18) => net47457, A(17) => 
                           net47458, A(16) => net47459, A(15) => net47460, 
                           A(14) => net47461, A(13) => net47462, A(12) => 
                           net47463, A(11) => net47464, A(10) => net47465, A(9)
                           => net47466, A(8) => net47467, A(7) => net47468, 
                           A(6) => net47469, A(5) => net47470, A(4) => net47471
                           , A(3) => net47472, A(2) => net47473, A(1) => 
                           net47474, A(0) => net47475, A_n(63) => net47476, 
                           A_n(62) => net47477, A_n(61) => net47478, A_n(60) =>
                           net47479, A_n(59) => net47480, A_n(58) => net47481, 
                           A_n(57) => net47482, A_n(56) => net47483, A_n(55) =>
                           net47484, A_n(54) => net47485, A_n(53) => net47486, 
                           A_n(52) => net47487, A_n(51) => net47488, A_n(50) =>
                           net47489, A_n(49) => net47490, A_n(48) => net47491, 
                           A_n(47) => net47492, A_n(46) => net47493, A_n(45) =>
                           net47494, A_n(44) => net47495, A_n(43) => net47496, 
                           A_n(42) => net47497, A_n(41) => net47498, A_n(40) =>
                           net47499, A_n(39) => net47500, A_n(38) => net47501, 
                           A_n(37) => net47502, A_n(36) => net47503, A_n(35) =>
                           net47504, A_n(34) => net47505, A_n(33) => net47506, 
                           A_n(32) => net47507, A_n(31) => net47508, A_n(30) =>
                           net47509, A_n(29) => net47510, A_n(28) => net47511, 
                           A_n(27) => net47512, A_n(26) => net47513, A_n(25) =>
                           net47514, A_n(24) => net47515, A_n(23) => net47516, 
                           A_n(22) => net47517, A_n(21) => net47518, A_n(20) =>
                           net47519, A_n(19) => net47520, A_n(18) => net47521, 
                           A_n(17) => net47522, A_n(16) => net47523, A_n(15) =>
                           net47524, A_n(14) => net47525, A_n(13) => net47526, 
                           A_n(12) => net47527, A_n(11) => net47528, A_n(10) =>
                           net47529, A_n(9) => net47530, A_n(8) => net47531, 
                           A_n(7) => net47532, A_n(6) => net47533, A_n(5) => 
                           net47534, A_n(4) => net47535, A_n(3) => net47536, 
                           A_n(2) => net47537, A_n(1) => net47538, A_n(0) => 
                           net47539, A_ns(63) => SHIFT_n_703_port, A_ns(62) => 
                           SHIFT_n_702_port, A_ns(61) => SHIFT_n_701_port, 
                           A_ns(60) => SHIFT_n_700_port, A_ns(59) => 
                           SHIFT_n_699_port, A_ns(58) => SHIFT_n_698_port, 
                           A_ns(57) => SHIFT_n_697_port, A_ns(56) => 
                           SHIFT_n_696_port, A_ns(55) => SHIFT_n_695_port, 
                           A_ns(54) => SHIFT_n_694_port, A_ns(53) => 
                           SHIFT_n_693_port, A_ns(52) => SHIFT_n_692_port, 
                           A_ns(51) => SHIFT_n_691_port, A_ns(50) => 
                           SHIFT_n_690_port, A_ns(49) => SHIFT_n_689_port, 
                           A_ns(48) => SHIFT_n_688_port, A_ns(47) => 
                           SHIFT_n_687_port, A_ns(46) => SHIFT_n_686_port, 
                           A_ns(45) => SHIFT_n_685_port, A_ns(44) => 
                           SHIFT_n_684_port, A_ns(43) => SHIFT_n_683_port, 
                           A_ns(42) => SHIFT_n_682_port, A_ns(41) => 
                           SHIFT_n_681_port, A_ns(40) => SHIFT_n_680_port, 
                           A_ns(39) => SHIFT_n_679_port, A_ns(38) => 
                           SHIFT_n_678_port, A_ns(37) => SHIFT_n_677_port, 
                           A_ns(36) => SHIFT_n_676_port, A_ns(35) => 
                           SHIFT_n_675_port, A_ns(34) => SHIFT_n_674_port, 
                           A_ns(33) => SHIFT_n_673_port, A_ns(32) => 
                           SHIFT_n_672_port, A_ns(31) => SHIFT_n_671_port, 
                           A_ns(30) => SHIFT_n_670_port, A_ns(29) => 
                           SHIFT_n_669_port, A_ns(28) => SHIFT_n_668_port, 
                           A_ns(27) => SHIFT_n_667_port, A_ns(26) => 
                           SHIFT_n_666_port, A_ns(25) => SHIFT_n_665_port, 
                           A_ns(24) => SHIFT_n_664_port, A_ns(23) => 
                           SHIFT_n_663_port, A_ns(22) => SHIFT_n_662_port, 
                           A_ns(21) => SHIFT_n_661_port, A_ns(20) => 
                           SHIFT_n_660_port, A_ns(19) => SHIFT_n_659_port, 
                           A_ns(18) => SHIFT_n_658_port, A_ns(17) => 
                           SHIFT_n_657_port, A_ns(16) => SHIFT_n_656_port, 
                           A_ns(15) => SHIFT_n_655_port, A_ns(14) => 
                           SHIFT_n_654_port, A_ns(13) => SHIFT_n_653_port, 
                           A_ns(12) => SHIFT_n_652_port, A_ns(11) => 
                           SHIFT_n_651_port, A_ns(10) => SHIFT_n_650_port, 
                           A_ns(9) => SHIFT_n_649_port, A_ns(8) => 
                           SHIFT_n_648_port, A_ns(7) => SHIFT_n_647_port, 
                           A_ns(6) => SHIFT_n_646_port, A_ns(5) => 
                           SHIFT_n_645_port, A_ns(4) => SHIFT_n_644_port, 
                           A_ns(3) => SHIFT_n_643_port, A_ns(2) => 
                           SHIFT_n_642_port, A_ns(1) => SHIFT_n_641_port, 
                           A_ns(0) => SHIFT_n_640_port, A_s(63) => 
                           SHIFT_703_port, A_s(62) => SHIFT_702_port, A_s(61) 
                           => SHIFT_701_port, A_s(60) => SHIFT_700_port, 
                           A_s(59) => SHIFT_699_port, A_s(58) => SHIFT_698_port
                           , A_s(57) => SHIFT_697_port, A_s(56) => 
                           SHIFT_696_port, A_s(55) => SHIFT_695_port, A_s(54) 
                           => SHIFT_694_port, A_s(53) => SHIFT_693_port, 
                           A_s(52) => SHIFT_692_port, A_s(51) => SHIFT_691_port
                           , A_s(50) => SHIFT_690_port, A_s(49) => 
                           SHIFT_689_port, A_s(48) => SHIFT_688_port, A_s(47) 
                           => SHIFT_687_port, A_s(46) => SHIFT_686_port, 
                           A_s(45) => SHIFT_685_port, A_s(44) => SHIFT_684_port
                           , A_s(43) => SHIFT_683_port, A_s(42) => 
                           SHIFT_682_port, A_s(41) => SHIFT_681_port, A_s(40) 
                           => SHIFT_680_port, A_s(39) => SHIFT_679_port, 
                           A_s(38) => SHIFT_678_port, A_s(37) => SHIFT_677_port
                           , A_s(36) => SHIFT_676_port, A_s(35) => 
                           SHIFT_675_port, A_s(34) => SHIFT_674_port, A_s(33) 
                           => SHIFT_673_port, A_s(32) => SHIFT_672_port, 
                           A_s(31) => SHIFT_671_port, A_s(30) => SHIFT_670_port
                           , A_s(29) => SHIFT_669_port, A_s(28) => 
                           SHIFT_668_port, A_s(27) => SHIFT_667_port, A_s(26) 
                           => SHIFT_666_port, A_s(25) => SHIFT_665_port, 
                           A_s(24) => SHIFT_664_port, A_s(23) => SHIFT_663_port
                           , A_s(22) => SHIFT_662_port, A_s(21) => 
                           SHIFT_661_port, A_s(20) => SHIFT_660_port, A_s(19) 
                           => SHIFT_659_port, A_s(18) => SHIFT_658_port, 
                           A_s(17) => SHIFT_657_port, A_s(16) => SHIFT_656_port
                           , A_s(15) => SHIFT_655_port, A_s(14) => 
                           SHIFT_654_port, A_s(13) => SHIFT_653_port, A_s(12) 
                           => SHIFT_652_port, A_s(11) => SHIFT_651_port, 
                           A_s(10) => SHIFT_650_port, A_s(9) => SHIFT_649_port,
                           A_s(8) => SHIFT_648_port, A_s(7) => SHIFT_647_port, 
                           A_s(6) => SHIFT_646_port, A_s(5) => SHIFT_645_port, 
                           A_s(4) => SHIFT_644_port, A_s(3) => SHIFT_643_port, 
                           A_s(2) => SHIFT_642_port, A_s(1) => SHIFT_641_port, 
                           A_s(0) => SHIFT_640_port, B(63) => B(31), B(62) => 
                           B(31), B(61) => B(31), B(60) => B(31), B(59) => 
                           B(31), B(58) => B(31), B(57) => B(31), B(56) => 
                           B(31), B(55) => B(31), B(54) => B(31), B(53) => 
                           B(31), B(52) => B(31), B(51) => B(31), B(50) => 
                           B(31), B(49) => B(31), B(48) => B(31), B(47) => 
                           B(31), B(46) => B(31), B(45) => B(31), B(44) => 
                           B(31), B(43) => B(31), B(42) => B(31), B(41) => 
                           B(31), B(40) => B(31), B(39) => B(31), B(38) => 
                           B(31), B(37) => B(31), B(36) => B(31), B(35) => 
                           B(31), B(34) => B(31), B(33) => B(31), B(32) => 
                           B(31), B(31) => B(31), B(30) => B(30), B(29) => 
                           B(29), B(28) => B(28), B(27) => B(27), B(26) => 
                           B(26), B(25) => B(25), B(24) => B(24), B(23) => 
                           B(23), B(22) => B(22), B(21) => B(21), B(20) => 
                           B(20), B(19) => B(19), B(18) => B(18), B(17) => 
                           B(17), B(16) => B(16), B(15) => B(15), B(14) => 
                           B(14), B(13) => B(13), B(12) => B(12), B(11) => 
                           B(11), B(10) => B(10), B(9) => B(9), B(8) => B(8), 
                           B(7) => B(7), B(6) => B(6), B(5) => B(5), B(4) => 
                           B(4), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), O(63) => OTMP_703_port, O(62) => 
                           OTMP_702_port, O(61) => OTMP_701_port, O(60) => 
                           OTMP_700_port, O(59) => OTMP_699_port, O(58) => 
                           OTMP_698_port, O(57) => OTMP_697_port, O(56) => 
                           OTMP_696_port, O(55) => OTMP_695_port, O(54) => 
                           OTMP_694_port, O(53) => OTMP_693_port, O(52) => 
                           OTMP_692_port, O(51) => OTMP_691_port, O(50) => 
                           OTMP_690_port, O(49) => OTMP_689_port, O(48) => 
                           OTMP_688_port, O(47) => OTMP_687_port, O(46) => 
                           OTMP_686_port, O(45) => OTMP_685_port, O(44) => 
                           OTMP_684_port, O(43) => OTMP_683_port, O(42) => 
                           OTMP_682_port, O(41) => OTMP_681_port, O(40) => 
                           OTMP_680_port, O(39) => OTMP_679_port, O(38) => 
                           OTMP_678_port, O(37) => OTMP_677_port, O(36) => 
                           OTMP_676_port, O(35) => OTMP_675_port, O(34) => 
                           OTMP_674_port, O(33) => OTMP_673_port, O(32) => 
                           OTMP_672_port, O(31) => OTMP_671_port, O(30) => 
                           OTMP_670_port, O(29) => OTMP_669_port, O(28) => 
                           OTMP_668_port, O(27) => OTMP_667_port, O(26) => 
                           OTMP_666_port, O(25) => OTMP_665_port, O(24) => 
                           OTMP_664_port, O(23) => OTMP_663_port, O(22) => 
                           OTMP_662_port, O(21) => OTMP_661_port, O(20) => 
                           OTMP_660_port, O(19) => OTMP_659_port, O(18) => 
                           OTMP_658_port, O(17) => OTMP_657_port, O(16) => 
                           OTMP_656_port, O(15) => OTMP_655_port, O(14) => 
                           OTMP_654_port, O(13) => OTMP_653_port, O(12) => 
                           OTMP_652_port, O(11) => OTMP_651_port, O(10) => 
                           OTMP_650_port, O(9) => OTMP_649_port, O(8) => 
                           OTMP_648_port, O(7) => OTMP_647_port, O(6) => 
                           OTMP_646_port, O(5) => OTMP_645_port, O(4) => 
                           OTMP_644_port, O(3) => OTMP_643_port, O(2) => 
                           OTMP_642_port, O(1) => OTMP_641_port, O(0) => n_1141
                           , A_so(63) => SHIFT_767_port, A_so(62) => 
                           SHIFT_766_port, A_so(61) => SHIFT_765_port, A_so(60)
                           => SHIFT_764_port, A_so(59) => SHIFT_763_port, 
                           A_so(58) => SHIFT_762_port, A_so(57) => 
                           SHIFT_761_port, A_so(56) => SHIFT_760_port, A_so(55)
                           => SHIFT_759_port, A_so(54) => SHIFT_758_port, 
                           A_so(53) => SHIFT_757_port, A_so(52) => 
                           SHIFT_756_port, A_so(51) => SHIFT_755_port, A_so(50)
                           => SHIFT_754_port, A_so(49) => SHIFT_753_port, 
                           A_so(48) => SHIFT_752_port, A_so(47) => 
                           SHIFT_751_port, A_so(46) => SHIFT_750_port, A_so(45)
                           => SHIFT_749_port, A_so(44) => SHIFT_748_port, 
                           A_so(43) => SHIFT_747_port, A_so(42) => 
                           SHIFT_746_port, A_so(41) => SHIFT_745_port, A_so(40)
                           => SHIFT_744_port, A_so(39) => SHIFT_743_port, 
                           A_so(38) => SHIFT_742_port, A_so(37) => 
                           SHIFT_741_port, A_so(36) => SHIFT_740_port, A_so(35)
                           => SHIFT_739_port, A_so(34) => SHIFT_738_port, 
                           A_so(33) => SHIFT_737_port, A_so(32) => 
                           SHIFT_736_port, A_so(31) => SHIFT_735_port, A_so(30)
                           => SHIFT_734_port, A_so(29) => SHIFT_733_port, 
                           A_so(28) => SHIFT_732_port, A_so(27) => 
                           SHIFT_731_port, A_so(26) => SHIFT_730_port, A_so(25)
                           => SHIFT_729_port, A_so(24) => SHIFT_728_port, 
                           A_so(23) => SHIFT_727_port, A_so(22) => 
                           SHIFT_726_port, A_so(21) => SHIFT_725_port, A_so(20)
                           => SHIFT_724_port, A_so(19) => SHIFT_723_port, 
                           A_so(18) => SHIFT_722_port, A_so(17) => 
                           SHIFT_721_port, A_so(16) => SHIFT_720_port, A_so(15)
                           => SHIFT_719_port, A_so(14) => SHIFT_718_port, 
                           A_so(13) => SHIFT_717_port, A_so(12) => 
                           SHIFT_716_port, A_so(11) => SHIFT_715_port, A_so(10)
                           => SHIFT_714_port, A_so(9) => SHIFT_713_port, 
                           A_so(8) => SHIFT_712_port, A_so(7) => SHIFT_711_port
                           , A_so(6) => SHIFT_710_port, A_so(5) => 
                           SHIFT_709_port, A_so(4) => SHIFT_708_port, A_so(3) 
                           => SHIFT_707_port, A_so(2) => SHIFT_706_port, 
                           A_so(1) => n_1142, A_so(0) => n_1143, A_nso(63) => 
                           SHIFT_n_767_port, A_nso(62) => SHIFT_n_766_port, 
                           A_nso(61) => SHIFT_n_765_port, A_nso(60) => 
                           SHIFT_n_764_port, A_nso(59) => SHIFT_n_763_port, 
                           A_nso(58) => SHIFT_n_762_port, A_nso(57) => 
                           SHIFT_n_761_port, A_nso(56) => SHIFT_n_760_port, 
                           A_nso(55) => SHIFT_n_759_port, A_nso(54) => 
                           SHIFT_n_758_port, A_nso(53) => SHIFT_n_757_port, 
                           A_nso(52) => SHIFT_n_756_port, A_nso(51) => 
                           SHIFT_n_755_port, A_nso(50) => SHIFT_n_754_port, 
                           A_nso(49) => SHIFT_n_753_port, A_nso(48) => 
                           SHIFT_n_752_port, A_nso(47) => SHIFT_n_751_port, 
                           A_nso(46) => SHIFT_n_750_port, A_nso(45) => 
                           SHIFT_n_749_port, A_nso(44) => SHIFT_n_748_port, 
                           A_nso(43) => SHIFT_n_747_port, A_nso(42) => 
                           SHIFT_n_746_port, A_nso(41) => SHIFT_n_745_port, 
                           A_nso(40) => SHIFT_n_744_port, A_nso(39) => 
                           SHIFT_n_743_port, A_nso(38) => SHIFT_n_742_port, 
                           A_nso(37) => SHIFT_n_741_port, A_nso(36) => 
                           SHIFT_n_740_port, A_nso(35) => SHIFT_n_739_port, 
                           A_nso(34) => SHIFT_n_738_port, A_nso(33) => 
                           SHIFT_n_737_port, A_nso(32) => SHIFT_n_736_port, 
                           A_nso(31) => SHIFT_n_735_port, A_nso(30) => 
                           SHIFT_n_734_port, A_nso(29) => SHIFT_n_733_port, 
                           A_nso(28) => SHIFT_n_732_port, A_nso(27) => 
                           SHIFT_n_731_port, A_nso(26) => SHIFT_n_730_port, 
                           A_nso(25) => SHIFT_n_729_port, A_nso(24) => 
                           SHIFT_n_728_port, A_nso(23) => SHIFT_n_727_port, 
                           A_nso(22) => SHIFT_n_726_port, A_nso(21) => 
                           SHIFT_n_725_port, A_nso(20) => SHIFT_n_724_port, 
                           A_nso(19) => SHIFT_n_723_port, A_nso(18) => 
                           SHIFT_n_722_port, A_nso(17) => SHIFT_n_721_port, 
                           A_nso(16) => SHIFT_n_720_port, A_nso(15) => 
                           SHIFT_n_719_port, A_nso(14) => SHIFT_n_718_port, 
                           A_nso(13) => SHIFT_n_717_port, A_nso(12) => 
                           SHIFT_n_716_port, A_nso(11) => SHIFT_n_715_port, 
                           A_nso(10) => SHIFT_n_714_port, A_nso(9) => 
                           SHIFT_n_713_port, A_nso(8) => SHIFT_n_712_port, 
                           A_nso(7) => SHIFT_n_711_port, A_nso(6) => 
                           SHIFT_n_710_port, A_nso(5) => SHIFT_n_709_port, 
                           A_nso(4) => SHIFT_n_708_port, A_nso(3) => 
                           SHIFT_n_707_port, A_nso(2) => SHIFT_n_706_port, 
                           A_nso(1) => n_1144, A_nso(0) => n_1145);
   BOOTHENC_I_12 : BOOTHENC_NBIT64_i22 port map( A(63) => net47284, A(62) => 
                           net47285, A(61) => net47286, A(60) => net47287, 
                           A(59) => net47288, A(58) => net47289, A(57) => 
                           net47290, A(56) => net47291, A(55) => net47292, 
                           A(54) => net47293, A(53) => net47294, A(52) => 
                           net47295, A(51) => net47296, A(50) => net47297, 
                           A(49) => net47298, A(48) => net47299, A(47) => 
                           net47300, A(46) => net47301, A(45) => net47302, 
                           A(44) => net47303, A(43) => net47304, A(42) => 
                           net47305, A(41) => net47306, A(40) => net47307, 
                           A(39) => net47308, A(38) => net47309, A(37) => 
                           net47310, A(36) => net47311, A(35) => net47312, 
                           A(34) => net47313, A(33) => net47314, A(32) => 
                           net47315, A(31) => net47316, A(30) => net47317, 
                           A(29) => net47318, A(28) => net47319, A(27) => 
                           net47320, A(26) => net47321, A(25) => net47322, 
                           A(24) => net47323, A(23) => net47324, A(22) => 
                           net47325, A(21) => net47326, A(20) => net47327, 
                           A(19) => net47328, A(18) => net47329, A(17) => 
                           net47330, A(16) => net47331, A(15) => net47332, 
                           A(14) => net47333, A(13) => net47334, A(12) => 
                           net47335, A(11) => net47336, A(10) => net47337, A(9)
                           => net47338, A(8) => net47339, A(7) => net47340, 
                           A(6) => net47341, A(5) => net47342, A(4) => net47343
                           , A(3) => net47344, A(2) => net47345, A(1) => 
                           net47346, A(0) => net47347, A_n(63) => net47348, 
                           A_n(62) => net47349, A_n(61) => net47350, A_n(60) =>
                           net47351, A_n(59) => net47352, A_n(58) => net47353, 
                           A_n(57) => net47354, A_n(56) => net47355, A_n(55) =>
                           net47356, A_n(54) => net47357, A_n(53) => net47358, 
                           A_n(52) => net47359, A_n(51) => net47360, A_n(50) =>
                           net47361, A_n(49) => net47362, A_n(48) => net47363, 
                           A_n(47) => net47364, A_n(46) => net47365, A_n(45) =>
                           net47366, A_n(44) => net47367, A_n(43) => net47368, 
                           A_n(42) => net47369, A_n(41) => net47370, A_n(40) =>
                           net47371, A_n(39) => net47372, A_n(38) => net47373, 
                           A_n(37) => net47374, A_n(36) => net47375, A_n(35) =>
                           net47376, A_n(34) => net47377, A_n(33) => net47378, 
                           A_n(32) => net47379, A_n(31) => net47380, A_n(30) =>
                           net47381, A_n(29) => net47382, A_n(28) => net47383, 
                           A_n(27) => net47384, A_n(26) => net47385, A_n(25) =>
                           net47386, A_n(24) => net47387, A_n(23) => net47388, 
                           A_n(22) => net47389, A_n(21) => net47390, A_n(20) =>
                           net47391, A_n(19) => net47392, A_n(18) => net47393, 
                           A_n(17) => net47394, A_n(16) => net47395, A_n(15) =>
                           net47396, A_n(14) => net47397, A_n(13) => net47398, 
                           A_n(12) => net47399, A_n(11) => net47400, A_n(10) =>
                           net47401, A_n(9) => net47402, A_n(8) => net47403, 
                           A_n(7) => net47404, A_n(6) => net47405, A_n(5) => 
                           net47406, A_n(4) => net47407, A_n(3) => net47408, 
                           A_n(2) => net47409, A_n(1) => net47410, A_n(0) => 
                           net47411, A_ns(63) => SHIFT_n_767_port, A_ns(62) => 
                           SHIFT_n_766_port, A_ns(61) => SHIFT_n_765_port, 
                           A_ns(60) => SHIFT_n_764_port, A_ns(59) => 
                           SHIFT_n_763_port, A_ns(58) => SHIFT_n_762_port, 
                           A_ns(57) => SHIFT_n_761_port, A_ns(56) => 
                           SHIFT_n_760_port, A_ns(55) => SHIFT_n_759_port, 
                           A_ns(54) => SHIFT_n_758_port, A_ns(53) => 
                           SHIFT_n_757_port, A_ns(52) => SHIFT_n_756_port, 
                           A_ns(51) => SHIFT_n_755_port, A_ns(50) => 
                           SHIFT_n_754_port, A_ns(49) => SHIFT_n_753_port, 
                           A_ns(48) => SHIFT_n_752_port, A_ns(47) => 
                           SHIFT_n_751_port, A_ns(46) => SHIFT_n_750_port, 
                           A_ns(45) => SHIFT_n_749_port, A_ns(44) => 
                           SHIFT_n_748_port, A_ns(43) => SHIFT_n_747_port, 
                           A_ns(42) => SHIFT_n_746_port, A_ns(41) => 
                           SHIFT_n_745_port, A_ns(40) => SHIFT_n_744_port, 
                           A_ns(39) => SHIFT_n_743_port, A_ns(38) => 
                           SHIFT_n_742_port, A_ns(37) => SHIFT_n_741_port, 
                           A_ns(36) => SHIFT_n_740_port, A_ns(35) => 
                           SHIFT_n_739_port, A_ns(34) => SHIFT_n_738_port, 
                           A_ns(33) => SHIFT_n_737_port, A_ns(32) => 
                           SHIFT_n_736_port, A_ns(31) => SHIFT_n_735_port, 
                           A_ns(30) => SHIFT_n_734_port, A_ns(29) => 
                           SHIFT_n_733_port, A_ns(28) => SHIFT_n_732_port, 
                           A_ns(27) => SHIFT_n_731_port, A_ns(26) => 
                           SHIFT_n_730_port, A_ns(25) => SHIFT_n_729_port, 
                           A_ns(24) => SHIFT_n_728_port, A_ns(23) => 
                           SHIFT_n_727_port, A_ns(22) => SHIFT_n_726_port, 
                           A_ns(21) => SHIFT_n_725_port, A_ns(20) => 
                           SHIFT_n_724_port, A_ns(19) => SHIFT_n_723_port, 
                           A_ns(18) => SHIFT_n_722_port, A_ns(17) => 
                           SHIFT_n_721_port, A_ns(16) => SHIFT_n_720_port, 
                           A_ns(15) => SHIFT_n_719_port, A_ns(14) => 
                           SHIFT_n_718_port, A_ns(13) => SHIFT_n_717_port, 
                           A_ns(12) => SHIFT_n_716_port, A_ns(11) => 
                           SHIFT_n_715_port, A_ns(10) => SHIFT_n_714_port, 
                           A_ns(9) => SHIFT_n_713_port, A_ns(8) => 
                           SHIFT_n_712_port, A_ns(7) => SHIFT_n_711_port, 
                           A_ns(6) => SHIFT_n_710_port, A_ns(5) => 
                           SHIFT_n_709_port, A_ns(4) => SHIFT_n_708_port, 
                           A_ns(3) => SHIFT_n_707_port, A_ns(2) => 
                           SHIFT_n_706_port, A_ns(1) => SHIFT_n_705_port, 
                           A_ns(0) => SHIFT_n_704_port, A_s(63) => 
                           SHIFT_767_port, A_s(62) => SHIFT_766_port, A_s(61) 
                           => SHIFT_765_port, A_s(60) => SHIFT_764_port, 
                           A_s(59) => SHIFT_763_port, A_s(58) => SHIFT_762_port
                           , A_s(57) => SHIFT_761_port, A_s(56) => 
                           SHIFT_760_port, A_s(55) => SHIFT_759_port, A_s(54) 
                           => SHIFT_758_port, A_s(53) => SHIFT_757_port, 
                           A_s(52) => SHIFT_756_port, A_s(51) => SHIFT_755_port
                           , A_s(50) => SHIFT_754_port, A_s(49) => 
                           SHIFT_753_port, A_s(48) => SHIFT_752_port, A_s(47) 
                           => SHIFT_751_port, A_s(46) => SHIFT_750_port, 
                           A_s(45) => SHIFT_749_port, A_s(44) => SHIFT_748_port
                           , A_s(43) => SHIFT_747_port, A_s(42) => 
                           SHIFT_746_port, A_s(41) => SHIFT_745_port, A_s(40) 
                           => SHIFT_744_port, A_s(39) => SHIFT_743_port, 
                           A_s(38) => SHIFT_742_port, A_s(37) => SHIFT_741_port
                           , A_s(36) => SHIFT_740_port, A_s(35) => 
                           SHIFT_739_port, A_s(34) => SHIFT_738_port, A_s(33) 
                           => SHIFT_737_port, A_s(32) => SHIFT_736_port, 
                           A_s(31) => SHIFT_735_port, A_s(30) => SHIFT_734_port
                           , A_s(29) => SHIFT_733_port, A_s(28) => 
                           SHIFT_732_port, A_s(27) => SHIFT_731_port, A_s(26) 
                           => SHIFT_730_port, A_s(25) => SHIFT_729_port, 
                           A_s(24) => SHIFT_728_port, A_s(23) => SHIFT_727_port
                           , A_s(22) => SHIFT_726_port, A_s(21) => 
                           SHIFT_725_port, A_s(20) => SHIFT_724_port, A_s(19) 
                           => SHIFT_723_port, A_s(18) => SHIFT_722_port, 
                           A_s(17) => SHIFT_721_port, A_s(16) => SHIFT_720_port
                           , A_s(15) => SHIFT_719_port, A_s(14) => 
                           SHIFT_718_port, A_s(13) => SHIFT_717_port, A_s(12) 
                           => SHIFT_716_port, A_s(11) => SHIFT_715_port, 
                           A_s(10) => SHIFT_714_port, A_s(9) => SHIFT_713_port,
                           A_s(8) => SHIFT_712_port, A_s(7) => SHIFT_711_port, 
                           A_s(6) => SHIFT_710_port, A_s(5) => SHIFT_709_port, 
                           A_s(4) => SHIFT_708_port, A_s(3) => SHIFT_707_port, 
                           A_s(2) => SHIFT_706_port, A_s(1) => SHIFT_705_port, 
                           A_s(0) => SHIFT_704_port, B(63) => B(31), B(62) => 
                           B(31), B(61) => B(31), B(60) => B(31), B(59) => 
                           B(31), B(58) => B(31), B(57) => B(31), B(56) => 
                           B(31), B(55) => B(31), B(54) => B(31), B(53) => 
                           B(31), B(52) => B(31), B(51) => B(31), B(50) => 
                           B(31), B(49) => B(31), B(48) => B(31), B(47) => 
                           B(31), B(46) => B(31), B(45) => B(31), B(44) => 
                           B(31), B(43) => B(31), B(42) => B(31), B(41) => 
                           B(31), B(40) => B(31), B(39) => B(31), B(38) => 
                           B(31), B(37) => B(31), B(36) => B(31), B(35) => 
                           B(31), B(34) => B(31), B(33) => B(31), B(32) => 
                           B(31), B(31) => B(31), B(30) => B(30), B(29) => 
                           B(29), B(28) => B(28), B(27) => B(27), B(26) => 
                           B(26), B(25) => B(25), B(24) => B(24), B(23) => 
                           B(23), B(22) => B(22), B(21) => B(21), B(20) => 
                           B(20), B(19) => B(19), B(18) => B(18), B(17) => 
                           B(17), B(16) => B(16), B(15) => B(15), B(14) => 
                           B(14), B(13) => B(13), B(12) => B(12), B(11) => 
                           B(11), B(10) => B(10), B(9) => B(9), B(8) => B(8), 
                           B(7) => B(7), B(6) => B(6), B(5) => B(5), B(4) => 
                           B(4), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), O(63) => OTMP_767_port, O(62) => 
                           OTMP_766_port, O(61) => OTMP_765_port, O(60) => 
                           OTMP_764_port, O(59) => OTMP_763_port, O(58) => 
                           OTMP_762_port, O(57) => OTMP_761_port, O(56) => 
                           OTMP_760_port, O(55) => OTMP_759_port, O(54) => 
                           OTMP_758_port, O(53) => OTMP_757_port, O(52) => 
                           OTMP_756_port, O(51) => OTMP_755_port, O(50) => 
                           OTMP_754_port, O(49) => OTMP_753_port, O(48) => 
                           OTMP_752_port, O(47) => OTMP_751_port, O(46) => 
                           OTMP_750_port, O(45) => OTMP_749_port, O(44) => 
                           OTMP_748_port, O(43) => OTMP_747_port, O(42) => 
                           OTMP_746_port, O(41) => OTMP_745_port, O(40) => 
                           OTMP_744_port, O(39) => OTMP_743_port, O(38) => 
                           OTMP_742_port, O(37) => OTMP_741_port, O(36) => 
                           OTMP_740_port, O(35) => OTMP_739_port, O(34) => 
                           OTMP_738_port, O(33) => OTMP_737_port, O(32) => 
                           OTMP_736_port, O(31) => OTMP_735_port, O(30) => 
                           OTMP_734_port, O(29) => OTMP_733_port, O(28) => 
                           OTMP_732_port, O(27) => OTMP_731_port, O(26) => 
                           OTMP_730_port, O(25) => OTMP_729_port, O(24) => 
                           OTMP_728_port, O(23) => OTMP_727_port, O(22) => 
                           OTMP_726_port, O(21) => OTMP_725_port, O(20) => 
                           OTMP_724_port, O(19) => OTMP_723_port, O(18) => 
                           OTMP_722_port, O(17) => OTMP_721_port, O(16) => 
                           OTMP_720_port, O(15) => OTMP_719_port, O(14) => 
                           OTMP_718_port, O(13) => OTMP_717_port, O(12) => 
                           OTMP_716_port, O(11) => OTMP_715_port, O(10) => 
                           OTMP_714_port, O(9) => OTMP_713_port, O(8) => 
                           OTMP_712_port, O(7) => OTMP_711_port, O(6) => 
                           OTMP_710_port, O(5) => OTMP_709_port, O(4) => 
                           OTMP_708_port, O(3) => OTMP_707_port, O(2) => 
                           OTMP_706_port, O(1) => OTMP_705_port, O(0) => n_1146
                           , A_so(63) => SHIFT_831_port, A_so(62) => 
                           SHIFT_830_port, A_so(61) => SHIFT_829_port, A_so(60)
                           => SHIFT_828_port, A_so(59) => SHIFT_827_port, 
                           A_so(58) => SHIFT_826_port, A_so(57) => 
                           SHIFT_825_port, A_so(56) => SHIFT_824_port, A_so(55)
                           => SHIFT_823_port, A_so(54) => SHIFT_822_port, 
                           A_so(53) => SHIFT_821_port, A_so(52) => 
                           SHIFT_820_port, A_so(51) => SHIFT_819_port, A_so(50)
                           => SHIFT_818_port, A_so(49) => SHIFT_817_port, 
                           A_so(48) => SHIFT_816_port, A_so(47) => 
                           SHIFT_815_port, A_so(46) => SHIFT_814_port, A_so(45)
                           => SHIFT_813_port, A_so(44) => SHIFT_812_port, 
                           A_so(43) => SHIFT_811_port, A_so(42) => 
                           SHIFT_810_port, A_so(41) => SHIFT_809_port, A_so(40)
                           => SHIFT_808_port, A_so(39) => SHIFT_807_port, 
                           A_so(38) => SHIFT_806_port, A_so(37) => 
                           SHIFT_805_port, A_so(36) => SHIFT_804_port, A_so(35)
                           => SHIFT_803_port, A_so(34) => SHIFT_802_port, 
                           A_so(33) => SHIFT_801_port, A_so(32) => 
                           SHIFT_800_port, A_so(31) => SHIFT_799_port, A_so(30)
                           => SHIFT_798_port, A_so(29) => SHIFT_797_port, 
                           A_so(28) => SHIFT_796_port, A_so(27) => 
                           SHIFT_795_port, A_so(26) => SHIFT_794_port, A_so(25)
                           => SHIFT_793_port, A_so(24) => SHIFT_792_port, 
                           A_so(23) => SHIFT_791_port, A_so(22) => 
                           SHIFT_790_port, A_so(21) => SHIFT_789_port, A_so(20)
                           => SHIFT_788_port, A_so(19) => SHIFT_787_port, 
                           A_so(18) => SHIFT_786_port, A_so(17) => 
                           SHIFT_785_port, A_so(16) => SHIFT_784_port, A_so(15)
                           => SHIFT_783_port, A_so(14) => SHIFT_782_port, 
                           A_so(13) => SHIFT_781_port, A_so(12) => 
                           SHIFT_780_port, A_so(11) => SHIFT_779_port, A_so(10)
                           => SHIFT_778_port, A_so(9) => SHIFT_777_port, 
                           A_so(8) => SHIFT_776_port, A_so(7) => SHIFT_775_port
                           , A_so(6) => SHIFT_774_port, A_so(5) => 
                           SHIFT_773_port, A_so(4) => SHIFT_772_port, A_so(3) 
                           => SHIFT_771_port, A_so(2) => SHIFT_770_port, 
                           A_so(1) => n_1147, A_so(0) => n_1148, A_nso(63) => 
                           SHIFT_n_831_port, A_nso(62) => SHIFT_n_830_port, 
                           A_nso(61) => SHIFT_n_829_port, A_nso(60) => 
                           SHIFT_n_828_port, A_nso(59) => SHIFT_n_827_port, 
                           A_nso(58) => SHIFT_n_826_port, A_nso(57) => 
                           SHIFT_n_825_port, A_nso(56) => SHIFT_n_824_port, 
                           A_nso(55) => SHIFT_n_823_port, A_nso(54) => 
                           SHIFT_n_822_port, A_nso(53) => SHIFT_n_821_port, 
                           A_nso(52) => SHIFT_n_820_port, A_nso(51) => 
                           SHIFT_n_819_port, A_nso(50) => SHIFT_n_818_port, 
                           A_nso(49) => SHIFT_n_817_port, A_nso(48) => 
                           SHIFT_n_816_port, A_nso(47) => SHIFT_n_815_port, 
                           A_nso(46) => SHIFT_n_814_port, A_nso(45) => 
                           SHIFT_n_813_port, A_nso(44) => SHIFT_n_812_port, 
                           A_nso(43) => SHIFT_n_811_port, A_nso(42) => 
                           SHIFT_n_810_port, A_nso(41) => SHIFT_n_809_port, 
                           A_nso(40) => SHIFT_n_808_port, A_nso(39) => 
                           SHIFT_n_807_port, A_nso(38) => SHIFT_n_806_port, 
                           A_nso(37) => SHIFT_n_805_port, A_nso(36) => 
                           SHIFT_n_804_port, A_nso(35) => SHIFT_n_803_port, 
                           A_nso(34) => SHIFT_n_802_port, A_nso(33) => 
                           SHIFT_n_801_port, A_nso(32) => SHIFT_n_800_port, 
                           A_nso(31) => SHIFT_n_799_port, A_nso(30) => 
                           SHIFT_n_798_port, A_nso(29) => SHIFT_n_797_port, 
                           A_nso(28) => SHIFT_n_796_port, A_nso(27) => 
                           SHIFT_n_795_port, A_nso(26) => SHIFT_n_794_port, 
                           A_nso(25) => SHIFT_n_793_port, A_nso(24) => 
                           SHIFT_n_792_port, A_nso(23) => SHIFT_n_791_port, 
                           A_nso(22) => SHIFT_n_790_port, A_nso(21) => 
                           SHIFT_n_789_port, A_nso(20) => SHIFT_n_788_port, 
                           A_nso(19) => SHIFT_n_787_port, A_nso(18) => 
                           SHIFT_n_786_port, A_nso(17) => SHIFT_n_785_port, 
                           A_nso(16) => SHIFT_n_784_port, A_nso(15) => 
                           SHIFT_n_783_port, A_nso(14) => SHIFT_n_782_port, 
                           A_nso(13) => SHIFT_n_781_port, A_nso(12) => 
                           SHIFT_n_780_port, A_nso(11) => SHIFT_n_779_port, 
                           A_nso(10) => SHIFT_n_778_port, A_nso(9) => 
                           SHIFT_n_777_port, A_nso(8) => SHIFT_n_776_port, 
                           A_nso(7) => SHIFT_n_775_port, A_nso(6) => 
                           SHIFT_n_774_port, A_nso(5) => SHIFT_n_773_port, 
                           A_nso(4) => SHIFT_n_772_port, A_nso(3) => 
                           SHIFT_n_771_port, A_nso(2) => SHIFT_n_770_port, 
                           A_nso(1) => n_1149, A_nso(0) => n_1150);
   BOOTHENC_I_13 : BOOTHENC_NBIT64_i24 port map( A(63) => net47156, A(62) => 
                           net47157, A(61) => net47158, A(60) => net47159, 
                           A(59) => net47160, A(58) => net47161, A(57) => 
                           net47162, A(56) => net47163, A(55) => net47164, 
                           A(54) => net47165, A(53) => net47166, A(52) => 
                           net47167, A(51) => net47168, A(50) => net47169, 
                           A(49) => net47170, A(48) => net47171, A(47) => 
                           net47172, A(46) => net47173, A(45) => net47174, 
                           A(44) => net47175, A(43) => net47176, A(42) => 
                           net47177, A(41) => net47178, A(40) => net47179, 
                           A(39) => net47180, A(38) => net47181, A(37) => 
                           net47182, A(36) => net47183, A(35) => net47184, 
                           A(34) => net47185, A(33) => net47186, A(32) => 
                           net47187, A(31) => net47188, A(30) => net47189, 
                           A(29) => net47190, A(28) => net47191, A(27) => 
                           net47192, A(26) => net47193, A(25) => net47194, 
                           A(24) => net47195, A(23) => net47196, A(22) => 
                           net47197, A(21) => net47198, A(20) => net47199, 
                           A(19) => net47200, A(18) => net47201, A(17) => 
                           net47202, A(16) => net47203, A(15) => net47204, 
                           A(14) => net47205, A(13) => net47206, A(12) => 
                           net47207, A(11) => net47208, A(10) => net47209, A(9)
                           => net47210, A(8) => net47211, A(7) => net47212, 
                           A(6) => net47213, A(5) => net47214, A(4) => net47215
                           , A(3) => net47216, A(2) => net47217, A(1) => 
                           net47218, A(0) => net47219, A_n(63) => net47220, 
                           A_n(62) => net47221, A_n(61) => net47222, A_n(60) =>
                           net47223, A_n(59) => net47224, A_n(58) => net47225, 
                           A_n(57) => net47226, A_n(56) => net47227, A_n(55) =>
                           net47228, A_n(54) => net47229, A_n(53) => net47230, 
                           A_n(52) => net47231, A_n(51) => net47232, A_n(50) =>
                           net47233, A_n(49) => net47234, A_n(48) => net47235, 
                           A_n(47) => net47236, A_n(46) => net47237, A_n(45) =>
                           net47238, A_n(44) => net47239, A_n(43) => net47240, 
                           A_n(42) => net47241, A_n(41) => net47242, A_n(40) =>
                           net47243, A_n(39) => net47244, A_n(38) => net47245, 
                           A_n(37) => net47246, A_n(36) => net47247, A_n(35) =>
                           net47248, A_n(34) => net47249, A_n(33) => net47250, 
                           A_n(32) => net47251, A_n(31) => net47252, A_n(30) =>
                           net47253, A_n(29) => net47254, A_n(28) => net47255, 
                           A_n(27) => net47256, A_n(26) => net47257, A_n(25) =>
                           net47258, A_n(24) => net47259, A_n(23) => net47260, 
                           A_n(22) => net47261, A_n(21) => net47262, A_n(20) =>
                           net47263, A_n(19) => net47264, A_n(18) => net47265, 
                           A_n(17) => net47266, A_n(16) => net47267, A_n(15) =>
                           net47268, A_n(14) => net47269, A_n(13) => net47270, 
                           A_n(12) => net47271, A_n(11) => net47272, A_n(10) =>
                           net47273, A_n(9) => net47274, A_n(8) => net47275, 
                           A_n(7) => net47276, A_n(6) => net47277, A_n(5) => 
                           net47278, A_n(4) => net47279, A_n(3) => net47280, 
                           A_n(2) => net47281, A_n(1) => net47282, A_n(0) => 
                           net47283, A_ns(63) => SHIFT_n_831_port, A_ns(62) => 
                           SHIFT_n_830_port, A_ns(61) => SHIFT_n_829_port, 
                           A_ns(60) => SHIFT_n_828_port, A_ns(59) => 
                           SHIFT_n_827_port, A_ns(58) => SHIFT_n_826_port, 
                           A_ns(57) => SHIFT_n_825_port, A_ns(56) => 
                           SHIFT_n_824_port, A_ns(55) => SHIFT_n_823_port, 
                           A_ns(54) => SHIFT_n_822_port, A_ns(53) => 
                           SHIFT_n_821_port, A_ns(52) => SHIFT_n_820_port, 
                           A_ns(51) => SHIFT_n_819_port, A_ns(50) => 
                           SHIFT_n_818_port, A_ns(49) => SHIFT_n_817_port, 
                           A_ns(48) => SHIFT_n_816_port, A_ns(47) => 
                           SHIFT_n_815_port, A_ns(46) => SHIFT_n_814_port, 
                           A_ns(45) => SHIFT_n_813_port, A_ns(44) => 
                           SHIFT_n_812_port, A_ns(43) => SHIFT_n_811_port, 
                           A_ns(42) => SHIFT_n_810_port, A_ns(41) => 
                           SHIFT_n_809_port, A_ns(40) => SHIFT_n_808_port, 
                           A_ns(39) => SHIFT_n_807_port, A_ns(38) => 
                           SHIFT_n_806_port, A_ns(37) => SHIFT_n_805_port, 
                           A_ns(36) => SHIFT_n_804_port, A_ns(35) => 
                           SHIFT_n_803_port, A_ns(34) => SHIFT_n_802_port, 
                           A_ns(33) => SHIFT_n_801_port, A_ns(32) => 
                           SHIFT_n_800_port, A_ns(31) => SHIFT_n_799_port, 
                           A_ns(30) => SHIFT_n_798_port, A_ns(29) => 
                           SHIFT_n_797_port, A_ns(28) => SHIFT_n_796_port, 
                           A_ns(27) => SHIFT_n_795_port, A_ns(26) => 
                           SHIFT_n_794_port, A_ns(25) => SHIFT_n_793_port, 
                           A_ns(24) => SHIFT_n_792_port, A_ns(23) => 
                           SHIFT_n_791_port, A_ns(22) => SHIFT_n_790_port, 
                           A_ns(21) => SHIFT_n_789_port, A_ns(20) => 
                           SHIFT_n_788_port, A_ns(19) => SHIFT_n_787_port, 
                           A_ns(18) => SHIFT_n_786_port, A_ns(17) => 
                           SHIFT_n_785_port, A_ns(16) => SHIFT_n_784_port, 
                           A_ns(15) => SHIFT_n_783_port, A_ns(14) => 
                           SHIFT_n_782_port, A_ns(13) => SHIFT_n_781_port, 
                           A_ns(12) => SHIFT_n_780_port, A_ns(11) => 
                           SHIFT_n_779_port, A_ns(10) => SHIFT_n_778_port, 
                           A_ns(9) => SHIFT_n_777_port, A_ns(8) => 
                           SHIFT_n_776_port, A_ns(7) => SHIFT_n_775_port, 
                           A_ns(6) => SHIFT_n_774_port, A_ns(5) => 
                           SHIFT_n_773_port, A_ns(4) => SHIFT_n_772_port, 
                           A_ns(3) => SHIFT_n_771_port, A_ns(2) => 
                           SHIFT_n_770_port, A_ns(1) => SHIFT_n_769_port, 
                           A_ns(0) => SHIFT_n_768_port, A_s(63) => 
                           SHIFT_831_port, A_s(62) => SHIFT_830_port, A_s(61) 
                           => SHIFT_829_port, A_s(60) => SHIFT_828_port, 
                           A_s(59) => SHIFT_827_port, A_s(58) => SHIFT_826_port
                           , A_s(57) => SHIFT_825_port, A_s(56) => 
                           SHIFT_824_port, A_s(55) => SHIFT_823_port, A_s(54) 
                           => SHIFT_822_port, A_s(53) => SHIFT_821_port, 
                           A_s(52) => SHIFT_820_port, A_s(51) => SHIFT_819_port
                           , A_s(50) => SHIFT_818_port, A_s(49) => 
                           SHIFT_817_port, A_s(48) => SHIFT_816_port, A_s(47) 
                           => SHIFT_815_port, A_s(46) => SHIFT_814_port, 
                           A_s(45) => SHIFT_813_port, A_s(44) => SHIFT_812_port
                           , A_s(43) => SHIFT_811_port, A_s(42) => 
                           SHIFT_810_port, A_s(41) => SHIFT_809_port, A_s(40) 
                           => SHIFT_808_port, A_s(39) => SHIFT_807_port, 
                           A_s(38) => SHIFT_806_port, A_s(37) => SHIFT_805_port
                           , A_s(36) => SHIFT_804_port, A_s(35) => 
                           SHIFT_803_port, A_s(34) => SHIFT_802_port, A_s(33) 
                           => SHIFT_801_port, A_s(32) => SHIFT_800_port, 
                           A_s(31) => SHIFT_799_port, A_s(30) => SHIFT_798_port
                           , A_s(29) => SHIFT_797_port, A_s(28) => 
                           SHIFT_796_port, A_s(27) => SHIFT_795_port, A_s(26) 
                           => SHIFT_794_port, A_s(25) => SHIFT_793_port, 
                           A_s(24) => SHIFT_792_port, A_s(23) => SHIFT_791_port
                           , A_s(22) => SHIFT_790_port, A_s(21) => 
                           SHIFT_789_port, A_s(20) => SHIFT_788_port, A_s(19) 
                           => SHIFT_787_port, A_s(18) => SHIFT_786_port, 
                           A_s(17) => SHIFT_785_port, A_s(16) => SHIFT_784_port
                           , A_s(15) => SHIFT_783_port, A_s(14) => 
                           SHIFT_782_port, A_s(13) => SHIFT_781_port, A_s(12) 
                           => SHIFT_780_port, A_s(11) => SHIFT_779_port, 
                           A_s(10) => SHIFT_778_port, A_s(9) => SHIFT_777_port,
                           A_s(8) => SHIFT_776_port, A_s(7) => SHIFT_775_port, 
                           A_s(6) => SHIFT_774_port, A_s(5) => SHIFT_773_port, 
                           A_s(4) => SHIFT_772_port, A_s(3) => SHIFT_771_port, 
                           A_s(2) => SHIFT_770_port, A_s(1) => SHIFT_769_port, 
                           A_s(0) => SHIFT_768_port, B(63) => B(31), B(62) => 
                           B(31), B(61) => B(31), B(60) => B(31), B(59) => 
                           B(31), B(58) => B(31), B(57) => B(31), B(56) => 
                           B(31), B(55) => B(31), B(54) => B(31), B(53) => 
                           B(31), B(52) => B(31), B(51) => B(31), B(50) => 
                           B(31), B(49) => B(31), B(48) => B(31), B(47) => 
                           B(31), B(46) => B(31), B(45) => B(31), B(44) => 
                           B(31), B(43) => B(31), B(42) => B(31), B(41) => 
                           B(31), B(40) => B(31), B(39) => B(31), B(38) => 
                           B(31), B(37) => B(31), B(36) => B(31), B(35) => 
                           B(31), B(34) => B(31), B(33) => B(31), B(32) => 
                           B(31), B(31) => B(31), B(30) => B(30), B(29) => 
                           B(29), B(28) => B(28), B(27) => B(27), B(26) => 
                           B(26), B(25) => B(25), B(24) => B(24), B(23) => 
                           B(23), B(22) => B(22), B(21) => B(21), B(20) => 
                           B(20), B(19) => B(19), B(18) => B(18), B(17) => 
                           B(17), B(16) => B(16), B(15) => B(15), B(14) => 
                           B(14), B(13) => B(13), B(12) => B(12), B(11) => 
                           B(11), B(10) => B(10), B(9) => B(9), B(8) => B(8), 
                           B(7) => B(7), B(6) => B(6), B(5) => B(5), B(4) => 
                           B(4), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), O(63) => OTMP_831_port, O(62) => 
                           OTMP_830_port, O(61) => OTMP_829_port, O(60) => 
                           OTMP_828_port, O(59) => OTMP_827_port, O(58) => 
                           OTMP_826_port, O(57) => OTMP_825_port, O(56) => 
                           OTMP_824_port, O(55) => OTMP_823_port, O(54) => 
                           OTMP_822_port, O(53) => OTMP_821_port, O(52) => 
                           OTMP_820_port, O(51) => OTMP_819_port, O(50) => 
                           OTMP_818_port, O(49) => OTMP_817_port, O(48) => 
                           OTMP_816_port, O(47) => OTMP_815_port, O(46) => 
                           OTMP_814_port, O(45) => OTMP_813_port, O(44) => 
                           OTMP_812_port, O(43) => OTMP_811_port, O(42) => 
                           OTMP_810_port, O(41) => OTMP_809_port, O(40) => 
                           OTMP_808_port, O(39) => OTMP_807_port, O(38) => 
                           OTMP_806_port, O(37) => OTMP_805_port, O(36) => 
                           OTMP_804_port, O(35) => OTMP_803_port, O(34) => 
                           OTMP_802_port, O(33) => OTMP_801_port, O(32) => 
                           OTMP_800_port, O(31) => OTMP_799_port, O(30) => 
                           OTMP_798_port, O(29) => OTMP_797_port, O(28) => 
                           OTMP_796_port, O(27) => OTMP_795_port, O(26) => 
                           OTMP_794_port, O(25) => OTMP_793_port, O(24) => 
                           OTMP_792_port, O(23) => OTMP_791_port, O(22) => 
                           OTMP_790_port, O(21) => OTMP_789_port, O(20) => 
                           OTMP_788_port, O(19) => OTMP_787_port, O(18) => 
                           OTMP_786_port, O(17) => OTMP_785_port, O(16) => 
                           OTMP_784_port, O(15) => OTMP_783_port, O(14) => 
                           OTMP_782_port, O(13) => OTMP_781_port, O(12) => 
                           OTMP_780_port, O(11) => OTMP_779_port, O(10) => 
                           OTMP_778_port, O(9) => OTMP_777_port, O(8) => 
                           OTMP_776_port, O(7) => OTMP_775_port, O(6) => 
                           OTMP_774_port, O(5) => OTMP_773_port, O(4) => 
                           OTMP_772_port, O(3) => OTMP_771_port, O(2) => 
                           OTMP_770_port, O(1) => OTMP_769_port, O(0) => n_1151
                           , A_so(63) => SHIFT_895_port, A_so(62) => 
                           SHIFT_894_port, A_so(61) => SHIFT_893_port, A_so(60)
                           => SHIFT_892_port, A_so(59) => SHIFT_891_port, 
                           A_so(58) => SHIFT_890_port, A_so(57) => 
                           SHIFT_889_port, A_so(56) => SHIFT_888_port, A_so(55)
                           => SHIFT_887_port, A_so(54) => SHIFT_886_port, 
                           A_so(53) => SHIFT_885_port, A_so(52) => 
                           SHIFT_884_port, A_so(51) => SHIFT_883_port, A_so(50)
                           => SHIFT_882_port, A_so(49) => SHIFT_881_port, 
                           A_so(48) => SHIFT_880_port, A_so(47) => 
                           SHIFT_879_port, A_so(46) => SHIFT_878_port, A_so(45)
                           => SHIFT_877_port, A_so(44) => SHIFT_876_port, 
                           A_so(43) => SHIFT_875_port, A_so(42) => 
                           SHIFT_874_port, A_so(41) => SHIFT_873_port, A_so(40)
                           => SHIFT_872_port, A_so(39) => SHIFT_871_port, 
                           A_so(38) => SHIFT_870_port, A_so(37) => 
                           SHIFT_869_port, A_so(36) => SHIFT_868_port, A_so(35)
                           => SHIFT_867_port, A_so(34) => SHIFT_866_port, 
                           A_so(33) => SHIFT_865_port, A_so(32) => 
                           SHIFT_864_port, A_so(31) => SHIFT_863_port, A_so(30)
                           => SHIFT_862_port, A_so(29) => SHIFT_861_port, 
                           A_so(28) => SHIFT_860_port, A_so(27) => 
                           SHIFT_859_port, A_so(26) => SHIFT_858_port, A_so(25)
                           => SHIFT_857_port, A_so(24) => SHIFT_856_port, 
                           A_so(23) => SHIFT_855_port, A_so(22) => 
                           SHIFT_854_port, A_so(21) => SHIFT_853_port, A_so(20)
                           => SHIFT_852_port, A_so(19) => SHIFT_851_port, 
                           A_so(18) => SHIFT_850_port, A_so(17) => 
                           SHIFT_849_port, A_so(16) => SHIFT_848_port, A_so(15)
                           => SHIFT_847_port, A_so(14) => SHIFT_846_port, 
                           A_so(13) => SHIFT_845_port, A_so(12) => 
                           SHIFT_844_port, A_so(11) => SHIFT_843_port, A_so(10)
                           => SHIFT_842_port, A_so(9) => SHIFT_841_port, 
                           A_so(8) => SHIFT_840_port, A_so(7) => SHIFT_839_port
                           , A_so(6) => SHIFT_838_port, A_so(5) => 
                           SHIFT_837_port, A_so(4) => SHIFT_836_port, A_so(3) 
                           => SHIFT_835_port, A_so(2) => SHIFT_834_port, 
                           A_so(1) => n_1152, A_so(0) => n_1153, A_nso(63) => 
                           SHIFT_n_895_port, A_nso(62) => SHIFT_n_894_port, 
                           A_nso(61) => SHIFT_n_893_port, A_nso(60) => 
                           SHIFT_n_892_port, A_nso(59) => SHIFT_n_891_port, 
                           A_nso(58) => SHIFT_n_890_port, A_nso(57) => 
                           SHIFT_n_889_port, A_nso(56) => SHIFT_n_888_port, 
                           A_nso(55) => SHIFT_n_887_port, A_nso(54) => 
                           SHIFT_n_886_port, A_nso(53) => SHIFT_n_885_port, 
                           A_nso(52) => SHIFT_n_884_port, A_nso(51) => 
                           SHIFT_n_883_port, A_nso(50) => SHIFT_n_882_port, 
                           A_nso(49) => SHIFT_n_881_port, A_nso(48) => 
                           SHIFT_n_880_port, A_nso(47) => SHIFT_n_879_port, 
                           A_nso(46) => SHIFT_n_878_port, A_nso(45) => 
                           SHIFT_n_877_port, A_nso(44) => SHIFT_n_876_port, 
                           A_nso(43) => SHIFT_n_875_port, A_nso(42) => 
                           SHIFT_n_874_port, A_nso(41) => SHIFT_n_873_port, 
                           A_nso(40) => SHIFT_n_872_port, A_nso(39) => 
                           SHIFT_n_871_port, A_nso(38) => SHIFT_n_870_port, 
                           A_nso(37) => SHIFT_n_869_port, A_nso(36) => 
                           SHIFT_n_868_port, A_nso(35) => SHIFT_n_867_port, 
                           A_nso(34) => SHIFT_n_866_port, A_nso(33) => 
                           SHIFT_n_865_port, A_nso(32) => SHIFT_n_864_port, 
                           A_nso(31) => SHIFT_n_863_port, A_nso(30) => 
                           SHIFT_n_862_port, A_nso(29) => SHIFT_n_861_port, 
                           A_nso(28) => SHIFT_n_860_port, A_nso(27) => 
                           SHIFT_n_859_port, A_nso(26) => SHIFT_n_858_port, 
                           A_nso(25) => SHIFT_n_857_port, A_nso(24) => 
                           SHIFT_n_856_port, A_nso(23) => SHIFT_n_855_port, 
                           A_nso(22) => SHIFT_n_854_port, A_nso(21) => 
                           SHIFT_n_853_port, A_nso(20) => SHIFT_n_852_port, 
                           A_nso(19) => SHIFT_n_851_port, A_nso(18) => 
                           SHIFT_n_850_port, A_nso(17) => SHIFT_n_849_port, 
                           A_nso(16) => SHIFT_n_848_port, A_nso(15) => 
                           SHIFT_n_847_port, A_nso(14) => SHIFT_n_846_port, 
                           A_nso(13) => SHIFT_n_845_port, A_nso(12) => 
                           SHIFT_n_844_port, A_nso(11) => SHIFT_n_843_port, 
                           A_nso(10) => SHIFT_n_842_port, A_nso(9) => 
                           SHIFT_n_841_port, A_nso(8) => SHIFT_n_840_port, 
                           A_nso(7) => SHIFT_n_839_port, A_nso(6) => 
                           SHIFT_n_838_port, A_nso(5) => SHIFT_n_837_port, 
                           A_nso(4) => SHIFT_n_836_port, A_nso(3) => 
                           SHIFT_n_835_port, A_nso(2) => SHIFT_n_834_port, 
                           A_nso(1) => n_1154, A_nso(0) => n_1155);
   BOOTHENC_I_14 : BOOTHENC_NBIT64_i26 port map( A(63) => net47028, A(62) => 
                           net47029, A(61) => net47030, A(60) => net47031, 
                           A(59) => net47032, A(58) => net47033, A(57) => 
                           net47034, A(56) => net47035, A(55) => net47036, 
                           A(54) => net47037, A(53) => net47038, A(52) => 
                           net47039, A(51) => net47040, A(50) => net47041, 
                           A(49) => net47042, A(48) => net47043, A(47) => 
                           net47044, A(46) => net47045, A(45) => net47046, 
                           A(44) => net47047, A(43) => net47048, A(42) => 
                           net47049, A(41) => net47050, A(40) => net47051, 
                           A(39) => net47052, A(38) => net47053, A(37) => 
                           net47054, A(36) => net47055, A(35) => net47056, 
                           A(34) => net47057, A(33) => net47058, A(32) => 
                           net47059, A(31) => net47060, A(30) => net47061, 
                           A(29) => net47062, A(28) => net47063, A(27) => 
                           net47064, A(26) => net47065, A(25) => net47066, 
                           A(24) => net47067, A(23) => net47068, A(22) => 
                           net47069, A(21) => net47070, A(20) => net47071, 
                           A(19) => net47072, A(18) => net47073, A(17) => 
                           net47074, A(16) => net47075, A(15) => net47076, 
                           A(14) => net47077, A(13) => net47078, A(12) => 
                           net47079, A(11) => net47080, A(10) => net47081, A(9)
                           => net47082, A(8) => net47083, A(7) => net47084, 
                           A(6) => net47085, A(5) => net47086, A(4) => net47087
                           , A(3) => net47088, A(2) => net47089, A(1) => 
                           net47090, A(0) => net47091, A_n(63) => net47092, 
                           A_n(62) => net47093, A_n(61) => net47094, A_n(60) =>
                           net47095, A_n(59) => net47096, A_n(58) => net47097, 
                           A_n(57) => net47098, A_n(56) => net47099, A_n(55) =>
                           net47100, A_n(54) => net47101, A_n(53) => net47102, 
                           A_n(52) => net47103, A_n(51) => net47104, A_n(50) =>
                           net47105, A_n(49) => net47106, A_n(48) => net47107, 
                           A_n(47) => net47108, A_n(46) => net47109, A_n(45) =>
                           net47110, A_n(44) => net47111, A_n(43) => net47112, 
                           A_n(42) => net47113, A_n(41) => net47114, A_n(40) =>
                           net47115, A_n(39) => net47116, A_n(38) => net47117, 
                           A_n(37) => net47118, A_n(36) => net47119, A_n(35) =>
                           net47120, A_n(34) => net47121, A_n(33) => net47122, 
                           A_n(32) => net47123, A_n(31) => net47124, A_n(30) =>
                           net47125, A_n(29) => net47126, A_n(28) => net47127, 
                           A_n(27) => net47128, A_n(26) => net47129, A_n(25) =>
                           net47130, A_n(24) => net47131, A_n(23) => net47132, 
                           A_n(22) => net47133, A_n(21) => net47134, A_n(20) =>
                           net47135, A_n(19) => net47136, A_n(18) => net47137, 
                           A_n(17) => net47138, A_n(16) => net47139, A_n(15) =>
                           net47140, A_n(14) => net47141, A_n(13) => net47142, 
                           A_n(12) => net47143, A_n(11) => net47144, A_n(10) =>
                           net47145, A_n(9) => net47146, A_n(8) => net47147, 
                           A_n(7) => net47148, A_n(6) => net47149, A_n(5) => 
                           net47150, A_n(4) => net47151, A_n(3) => net47152, 
                           A_n(2) => net47153, A_n(1) => net47154, A_n(0) => 
                           net47155, A_ns(63) => SHIFT_n_895_port, A_ns(62) => 
                           SHIFT_n_894_port, A_ns(61) => SHIFT_n_893_port, 
                           A_ns(60) => SHIFT_n_892_port, A_ns(59) => 
                           SHIFT_n_891_port, A_ns(58) => SHIFT_n_890_port, 
                           A_ns(57) => SHIFT_n_889_port, A_ns(56) => 
                           SHIFT_n_888_port, A_ns(55) => SHIFT_n_887_port, 
                           A_ns(54) => SHIFT_n_886_port, A_ns(53) => 
                           SHIFT_n_885_port, A_ns(52) => SHIFT_n_884_port, 
                           A_ns(51) => SHIFT_n_883_port, A_ns(50) => 
                           SHIFT_n_882_port, A_ns(49) => SHIFT_n_881_port, 
                           A_ns(48) => SHIFT_n_880_port, A_ns(47) => 
                           SHIFT_n_879_port, A_ns(46) => SHIFT_n_878_port, 
                           A_ns(45) => SHIFT_n_877_port, A_ns(44) => 
                           SHIFT_n_876_port, A_ns(43) => SHIFT_n_875_port, 
                           A_ns(42) => SHIFT_n_874_port, A_ns(41) => 
                           SHIFT_n_873_port, A_ns(40) => SHIFT_n_872_port, 
                           A_ns(39) => SHIFT_n_871_port, A_ns(38) => 
                           SHIFT_n_870_port, A_ns(37) => SHIFT_n_869_port, 
                           A_ns(36) => SHIFT_n_868_port, A_ns(35) => 
                           SHIFT_n_867_port, A_ns(34) => SHIFT_n_866_port, 
                           A_ns(33) => SHIFT_n_865_port, A_ns(32) => 
                           SHIFT_n_864_port, A_ns(31) => SHIFT_n_863_port, 
                           A_ns(30) => SHIFT_n_862_port, A_ns(29) => 
                           SHIFT_n_861_port, A_ns(28) => SHIFT_n_860_port, 
                           A_ns(27) => SHIFT_n_859_port, A_ns(26) => 
                           SHIFT_n_858_port, A_ns(25) => SHIFT_n_857_port, 
                           A_ns(24) => SHIFT_n_856_port, A_ns(23) => 
                           SHIFT_n_855_port, A_ns(22) => SHIFT_n_854_port, 
                           A_ns(21) => SHIFT_n_853_port, A_ns(20) => 
                           SHIFT_n_852_port, A_ns(19) => SHIFT_n_851_port, 
                           A_ns(18) => SHIFT_n_850_port, A_ns(17) => 
                           SHIFT_n_849_port, A_ns(16) => SHIFT_n_848_port, 
                           A_ns(15) => SHIFT_n_847_port, A_ns(14) => 
                           SHIFT_n_846_port, A_ns(13) => SHIFT_n_845_port, 
                           A_ns(12) => SHIFT_n_844_port, A_ns(11) => 
                           SHIFT_n_843_port, A_ns(10) => SHIFT_n_842_port, 
                           A_ns(9) => SHIFT_n_841_port, A_ns(8) => 
                           SHIFT_n_840_port, A_ns(7) => SHIFT_n_839_port, 
                           A_ns(6) => SHIFT_n_838_port, A_ns(5) => 
                           SHIFT_n_837_port, A_ns(4) => SHIFT_n_836_port, 
                           A_ns(3) => SHIFT_n_835_port, A_ns(2) => 
                           SHIFT_n_834_port, A_ns(1) => SHIFT_n_833_port, 
                           A_ns(0) => SHIFT_n_832_port, A_s(63) => 
                           SHIFT_895_port, A_s(62) => SHIFT_894_port, A_s(61) 
                           => SHIFT_893_port, A_s(60) => SHIFT_892_port, 
                           A_s(59) => SHIFT_891_port, A_s(58) => SHIFT_890_port
                           , A_s(57) => SHIFT_889_port, A_s(56) => 
                           SHIFT_888_port, A_s(55) => SHIFT_887_port, A_s(54) 
                           => SHIFT_886_port, A_s(53) => SHIFT_885_port, 
                           A_s(52) => SHIFT_884_port, A_s(51) => SHIFT_883_port
                           , A_s(50) => SHIFT_882_port, A_s(49) => 
                           SHIFT_881_port, A_s(48) => SHIFT_880_port, A_s(47) 
                           => SHIFT_879_port, A_s(46) => SHIFT_878_port, 
                           A_s(45) => SHIFT_877_port, A_s(44) => SHIFT_876_port
                           , A_s(43) => SHIFT_875_port, A_s(42) => 
                           SHIFT_874_port, A_s(41) => SHIFT_873_port, A_s(40) 
                           => SHIFT_872_port, A_s(39) => SHIFT_871_port, 
                           A_s(38) => SHIFT_870_port, A_s(37) => SHIFT_869_port
                           , A_s(36) => SHIFT_868_port, A_s(35) => 
                           SHIFT_867_port, A_s(34) => SHIFT_866_port, A_s(33) 
                           => SHIFT_865_port, A_s(32) => SHIFT_864_port, 
                           A_s(31) => SHIFT_863_port, A_s(30) => SHIFT_862_port
                           , A_s(29) => SHIFT_861_port, A_s(28) => 
                           SHIFT_860_port, A_s(27) => SHIFT_859_port, A_s(26) 
                           => SHIFT_858_port, A_s(25) => SHIFT_857_port, 
                           A_s(24) => SHIFT_856_port, A_s(23) => SHIFT_855_port
                           , A_s(22) => SHIFT_854_port, A_s(21) => 
                           SHIFT_853_port, A_s(20) => SHIFT_852_port, A_s(19) 
                           => SHIFT_851_port, A_s(18) => SHIFT_850_port, 
                           A_s(17) => SHIFT_849_port, A_s(16) => SHIFT_848_port
                           , A_s(15) => SHIFT_847_port, A_s(14) => 
                           SHIFT_846_port, A_s(13) => SHIFT_845_port, A_s(12) 
                           => SHIFT_844_port, A_s(11) => SHIFT_843_port, 
                           A_s(10) => SHIFT_842_port, A_s(9) => SHIFT_841_port,
                           A_s(8) => SHIFT_840_port, A_s(7) => SHIFT_839_port, 
                           A_s(6) => SHIFT_838_port, A_s(5) => SHIFT_837_port, 
                           A_s(4) => SHIFT_836_port, A_s(3) => SHIFT_835_port, 
                           A_s(2) => SHIFT_834_port, A_s(1) => SHIFT_833_port, 
                           A_s(0) => SHIFT_832_port, B(63) => B(31), B(62) => 
                           B(31), B(61) => B(31), B(60) => B(31), B(59) => 
                           B(31), B(58) => B(31), B(57) => B(31), B(56) => 
                           B(31), B(55) => B(31), B(54) => B(31), B(53) => 
                           B(31), B(52) => B(31), B(51) => B(31), B(50) => 
                           B(31), B(49) => B(31), B(48) => B(31), B(47) => 
                           B(31), B(46) => B(31), B(45) => B(31), B(44) => 
                           B(31), B(43) => B(31), B(42) => B(31), B(41) => 
                           B(31), B(40) => B(31), B(39) => B(31), B(38) => 
                           B(31), B(37) => B(31), B(36) => B(31), B(35) => 
                           B(31), B(34) => B(31), B(33) => B(31), B(32) => 
                           B(31), B(31) => B(31), B(30) => B(30), B(29) => 
                           B(29), B(28) => B(28), B(27) => B(27), B(26) => 
                           B(26), B(25) => B(25), B(24) => B(24), B(23) => 
                           B(23), B(22) => B(22), B(21) => B(21), B(20) => 
                           B(20), B(19) => B(19), B(18) => B(18), B(17) => 
                           B(17), B(16) => B(16), B(15) => B(15), B(14) => 
                           B(14), B(13) => B(13), B(12) => B(12), B(11) => 
                           B(11), B(10) => B(10), B(9) => B(9), B(8) => B(8), 
                           B(7) => B(7), B(6) => B(6), B(5) => B(5), B(4) => 
                           B(4), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), O(63) => OTMP_895_port, O(62) => 
                           OTMP_894_port, O(61) => OTMP_893_port, O(60) => 
                           OTMP_892_port, O(59) => OTMP_891_port, O(58) => 
                           OTMP_890_port, O(57) => OTMP_889_port, O(56) => 
                           OTMP_888_port, O(55) => OTMP_887_port, O(54) => 
                           OTMP_886_port, O(53) => OTMP_885_port, O(52) => 
                           OTMP_884_port, O(51) => OTMP_883_port, O(50) => 
                           OTMP_882_port, O(49) => OTMP_881_port, O(48) => 
                           OTMP_880_port, O(47) => OTMP_879_port, O(46) => 
                           OTMP_878_port, O(45) => OTMP_877_port, O(44) => 
                           OTMP_876_port, O(43) => OTMP_875_port, O(42) => 
                           OTMP_874_port, O(41) => OTMP_873_port, O(40) => 
                           OTMP_872_port, O(39) => OTMP_871_port, O(38) => 
                           OTMP_870_port, O(37) => OTMP_869_port, O(36) => 
                           OTMP_868_port, O(35) => OTMP_867_port, O(34) => 
                           OTMP_866_port, O(33) => OTMP_865_port, O(32) => 
                           OTMP_864_port, O(31) => OTMP_863_port, O(30) => 
                           OTMP_862_port, O(29) => OTMP_861_port, O(28) => 
                           OTMP_860_port, O(27) => OTMP_859_port, O(26) => 
                           OTMP_858_port, O(25) => OTMP_857_port, O(24) => 
                           OTMP_856_port, O(23) => OTMP_855_port, O(22) => 
                           OTMP_854_port, O(21) => OTMP_853_port, O(20) => 
                           OTMP_852_port, O(19) => OTMP_851_port, O(18) => 
                           OTMP_850_port, O(17) => OTMP_849_port, O(16) => 
                           OTMP_848_port, O(15) => OTMP_847_port, O(14) => 
                           OTMP_846_port, O(13) => OTMP_845_port, O(12) => 
                           OTMP_844_port, O(11) => OTMP_843_port, O(10) => 
                           OTMP_842_port, O(9) => OTMP_841_port, O(8) => 
                           OTMP_840_port, O(7) => OTMP_839_port, O(6) => 
                           OTMP_838_port, O(5) => OTMP_837_port, O(4) => 
                           OTMP_836_port, O(3) => OTMP_835_port, O(2) => 
                           OTMP_834_port, O(1) => OTMP_833_port, O(0) => n_1156
                           , A_so(63) => SHIFT_959_port, A_so(62) => 
                           SHIFT_958_port, A_so(61) => SHIFT_957_port, A_so(60)
                           => SHIFT_956_port, A_so(59) => SHIFT_955_port, 
                           A_so(58) => SHIFT_954_port, A_so(57) => 
                           SHIFT_953_port, A_so(56) => SHIFT_952_port, A_so(55)
                           => SHIFT_951_port, A_so(54) => SHIFT_950_port, 
                           A_so(53) => SHIFT_949_port, A_so(52) => 
                           SHIFT_948_port, A_so(51) => SHIFT_947_port, A_so(50)
                           => SHIFT_946_port, A_so(49) => SHIFT_945_port, 
                           A_so(48) => SHIFT_944_port, A_so(47) => 
                           SHIFT_943_port, A_so(46) => SHIFT_942_port, A_so(45)
                           => SHIFT_941_port, A_so(44) => SHIFT_940_port, 
                           A_so(43) => SHIFT_939_port, A_so(42) => 
                           SHIFT_938_port, A_so(41) => SHIFT_937_port, A_so(40)
                           => SHIFT_936_port, A_so(39) => SHIFT_935_port, 
                           A_so(38) => SHIFT_934_port, A_so(37) => 
                           SHIFT_933_port, A_so(36) => SHIFT_932_port, A_so(35)
                           => SHIFT_931_port, A_so(34) => SHIFT_930_port, 
                           A_so(33) => SHIFT_929_port, A_so(32) => 
                           SHIFT_928_port, A_so(31) => SHIFT_927_port, A_so(30)
                           => SHIFT_926_port, A_so(29) => SHIFT_925_port, 
                           A_so(28) => SHIFT_924_port, A_so(27) => 
                           SHIFT_923_port, A_so(26) => SHIFT_922_port, A_so(25)
                           => SHIFT_921_port, A_so(24) => SHIFT_920_port, 
                           A_so(23) => SHIFT_919_port, A_so(22) => 
                           SHIFT_918_port, A_so(21) => SHIFT_917_port, A_so(20)
                           => SHIFT_916_port, A_so(19) => SHIFT_915_port, 
                           A_so(18) => SHIFT_914_port, A_so(17) => 
                           SHIFT_913_port, A_so(16) => SHIFT_912_port, A_so(15)
                           => SHIFT_911_port, A_so(14) => SHIFT_910_port, 
                           A_so(13) => SHIFT_909_port, A_so(12) => 
                           SHIFT_908_port, A_so(11) => SHIFT_907_port, A_so(10)
                           => SHIFT_906_port, A_so(9) => SHIFT_905_port, 
                           A_so(8) => SHIFT_904_port, A_so(7) => SHIFT_903_port
                           , A_so(6) => SHIFT_902_port, A_so(5) => 
                           SHIFT_901_port, A_so(4) => SHIFT_900_port, A_so(3) 
                           => SHIFT_899_port, A_so(2) => SHIFT_898_port, 
                           A_so(1) => n_1157, A_so(0) => n_1158, A_nso(63) => 
                           SHIFT_n_959_port, A_nso(62) => SHIFT_n_958_port, 
                           A_nso(61) => SHIFT_n_957_port, A_nso(60) => 
                           SHIFT_n_956_port, A_nso(59) => SHIFT_n_955_port, 
                           A_nso(58) => SHIFT_n_954_port, A_nso(57) => 
                           SHIFT_n_953_port, A_nso(56) => SHIFT_n_952_port, 
                           A_nso(55) => SHIFT_n_951_port, A_nso(54) => 
                           SHIFT_n_950_port, A_nso(53) => SHIFT_n_949_port, 
                           A_nso(52) => SHIFT_n_948_port, A_nso(51) => 
                           SHIFT_n_947_port, A_nso(50) => SHIFT_n_946_port, 
                           A_nso(49) => SHIFT_n_945_port, A_nso(48) => 
                           SHIFT_n_944_port, A_nso(47) => SHIFT_n_943_port, 
                           A_nso(46) => SHIFT_n_942_port, A_nso(45) => 
                           SHIFT_n_941_port, A_nso(44) => SHIFT_n_940_port, 
                           A_nso(43) => SHIFT_n_939_port, A_nso(42) => 
                           SHIFT_n_938_port, A_nso(41) => SHIFT_n_937_port, 
                           A_nso(40) => SHIFT_n_936_port, A_nso(39) => 
                           SHIFT_n_935_port, A_nso(38) => SHIFT_n_934_port, 
                           A_nso(37) => SHIFT_n_933_port, A_nso(36) => 
                           SHIFT_n_932_port, A_nso(35) => SHIFT_n_931_port, 
                           A_nso(34) => SHIFT_n_930_port, A_nso(33) => 
                           SHIFT_n_929_port, A_nso(32) => SHIFT_n_928_port, 
                           A_nso(31) => SHIFT_n_927_port, A_nso(30) => 
                           SHIFT_n_926_port, A_nso(29) => SHIFT_n_925_port, 
                           A_nso(28) => SHIFT_n_924_port, A_nso(27) => 
                           SHIFT_n_923_port, A_nso(26) => SHIFT_n_922_port, 
                           A_nso(25) => SHIFT_n_921_port, A_nso(24) => 
                           SHIFT_n_920_port, A_nso(23) => SHIFT_n_919_port, 
                           A_nso(22) => SHIFT_n_918_port, A_nso(21) => 
                           SHIFT_n_917_port, A_nso(20) => SHIFT_n_916_port, 
                           A_nso(19) => SHIFT_n_915_port, A_nso(18) => 
                           SHIFT_n_914_port, A_nso(17) => SHIFT_n_913_port, 
                           A_nso(16) => SHIFT_n_912_port, A_nso(15) => 
                           SHIFT_n_911_port, A_nso(14) => SHIFT_n_910_port, 
                           A_nso(13) => SHIFT_n_909_port, A_nso(12) => 
                           SHIFT_n_908_port, A_nso(11) => SHIFT_n_907_port, 
                           A_nso(10) => SHIFT_n_906_port, A_nso(9) => 
                           SHIFT_n_905_port, A_nso(8) => SHIFT_n_904_port, 
                           A_nso(7) => SHIFT_n_903_port, A_nso(6) => 
                           SHIFT_n_902_port, A_nso(5) => SHIFT_n_901_port, 
                           A_nso(4) => SHIFT_n_900_port, A_nso(3) => 
                           SHIFT_n_899_port, A_nso(2) => SHIFT_n_898_port, 
                           A_nso(1) => n_1159, A_nso(0) => n_1160);
   BOOTHENC_I_15 : BOOTHENC_NBIT64_i28 port map( A(63) => net46900, A(62) => 
                           net46901, A(61) => net46902, A(60) => net46903, 
                           A(59) => net46904, A(58) => net46905, A(57) => 
                           net46906, A(56) => net46907, A(55) => net46908, 
                           A(54) => net46909, A(53) => net46910, A(52) => 
                           net46911, A(51) => net46912, A(50) => net46913, 
                           A(49) => net46914, A(48) => net46915, A(47) => 
                           net46916, A(46) => net46917, A(45) => net46918, 
                           A(44) => net46919, A(43) => net46920, A(42) => 
                           net46921, A(41) => net46922, A(40) => net46923, 
                           A(39) => net46924, A(38) => net46925, A(37) => 
                           net46926, A(36) => net46927, A(35) => net46928, 
                           A(34) => net46929, A(33) => net46930, A(32) => 
                           net46931, A(31) => net46932, A(30) => net46933, 
                           A(29) => net46934, A(28) => net46935, A(27) => 
                           net46936, A(26) => net46937, A(25) => net46938, 
                           A(24) => net46939, A(23) => net46940, A(22) => 
                           net46941, A(21) => net46942, A(20) => net46943, 
                           A(19) => net46944, A(18) => net46945, A(17) => 
                           net46946, A(16) => net46947, A(15) => net46948, 
                           A(14) => net46949, A(13) => net46950, A(12) => 
                           net46951, A(11) => net46952, A(10) => net46953, A(9)
                           => net46954, A(8) => net46955, A(7) => net46956, 
                           A(6) => net46957, A(5) => net46958, A(4) => net46959
                           , A(3) => net46960, A(2) => net46961, A(1) => 
                           net46962, A(0) => net46963, A_n(63) => net46964, 
                           A_n(62) => net46965, A_n(61) => net46966, A_n(60) =>
                           net46967, A_n(59) => net46968, A_n(58) => net46969, 
                           A_n(57) => net46970, A_n(56) => net46971, A_n(55) =>
                           net46972, A_n(54) => net46973, A_n(53) => net46974, 
                           A_n(52) => net46975, A_n(51) => net46976, A_n(50) =>
                           net46977, A_n(49) => net46978, A_n(48) => net46979, 
                           A_n(47) => net46980, A_n(46) => net46981, A_n(45) =>
                           net46982, A_n(44) => net46983, A_n(43) => net46984, 
                           A_n(42) => net46985, A_n(41) => net46986, A_n(40) =>
                           net46987, A_n(39) => net46988, A_n(38) => net46989, 
                           A_n(37) => net46990, A_n(36) => net46991, A_n(35) =>
                           net46992, A_n(34) => net46993, A_n(33) => net46994, 
                           A_n(32) => net46995, A_n(31) => net46996, A_n(30) =>
                           net46997, A_n(29) => net46998, A_n(28) => net46999, 
                           A_n(27) => net47000, A_n(26) => net47001, A_n(25) =>
                           net47002, A_n(24) => net47003, A_n(23) => net47004, 
                           A_n(22) => net47005, A_n(21) => net47006, A_n(20) =>
                           net47007, A_n(19) => net47008, A_n(18) => net47009, 
                           A_n(17) => net47010, A_n(16) => net47011, A_n(15) =>
                           net47012, A_n(14) => net47013, A_n(13) => net47014, 
                           A_n(12) => net47015, A_n(11) => net47016, A_n(10) =>
                           net47017, A_n(9) => net47018, A_n(8) => net47019, 
                           A_n(7) => net47020, A_n(6) => net47021, A_n(5) => 
                           net47022, A_n(4) => net47023, A_n(3) => net47024, 
                           A_n(2) => net47025, A_n(1) => net47026, A_n(0) => 
                           net47027, A_ns(63) => SHIFT_n_959_port, A_ns(62) => 
                           SHIFT_n_958_port, A_ns(61) => SHIFT_n_957_port, 
                           A_ns(60) => SHIFT_n_956_port, A_ns(59) => 
                           SHIFT_n_955_port, A_ns(58) => SHIFT_n_954_port, 
                           A_ns(57) => SHIFT_n_953_port, A_ns(56) => 
                           SHIFT_n_952_port, A_ns(55) => SHIFT_n_951_port, 
                           A_ns(54) => SHIFT_n_950_port, A_ns(53) => 
                           SHIFT_n_949_port, A_ns(52) => SHIFT_n_948_port, 
                           A_ns(51) => SHIFT_n_947_port, A_ns(50) => 
                           SHIFT_n_946_port, A_ns(49) => SHIFT_n_945_port, 
                           A_ns(48) => SHIFT_n_944_port, A_ns(47) => 
                           SHIFT_n_943_port, A_ns(46) => SHIFT_n_942_port, 
                           A_ns(45) => SHIFT_n_941_port, A_ns(44) => 
                           SHIFT_n_940_port, A_ns(43) => SHIFT_n_939_port, 
                           A_ns(42) => SHIFT_n_938_port, A_ns(41) => 
                           SHIFT_n_937_port, A_ns(40) => SHIFT_n_936_port, 
                           A_ns(39) => SHIFT_n_935_port, A_ns(38) => 
                           SHIFT_n_934_port, A_ns(37) => SHIFT_n_933_port, 
                           A_ns(36) => SHIFT_n_932_port, A_ns(35) => 
                           SHIFT_n_931_port, A_ns(34) => SHIFT_n_930_port, 
                           A_ns(33) => SHIFT_n_929_port, A_ns(32) => 
                           SHIFT_n_928_port, A_ns(31) => SHIFT_n_927_port, 
                           A_ns(30) => SHIFT_n_926_port, A_ns(29) => 
                           SHIFT_n_925_port, A_ns(28) => SHIFT_n_924_port, 
                           A_ns(27) => SHIFT_n_923_port, A_ns(26) => 
                           SHIFT_n_922_port, A_ns(25) => SHIFT_n_921_port, 
                           A_ns(24) => SHIFT_n_920_port, A_ns(23) => 
                           SHIFT_n_919_port, A_ns(22) => SHIFT_n_918_port, 
                           A_ns(21) => SHIFT_n_917_port, A_ns(20) => 
                           SHIFT_n_916_port, A_ns(19) => SHIFT_n_915_port, 
                           A_ns(18) => SHIFT_n_914_port, A_ns(17) => 
                           SHIFT_n_913_port, A_ns(16) => SHIFT_n_912_port, 
                           A_ns(15) => SHIFT_n_911_port, A_ns(14) => 
                           SHIFT_n_910_port, A_ns(13) => SHIFT_n_909_port, 
                           A_ns(12) => SHIFT_n_908_port, A_ns(11) => 
                           SHIFT_n_907_port, A_ns(10) => SHIFT_n_906_port, 
                           A_ns(9) => SHIFT_n_905_port, A_ns(8) => 
                           SHIFT_n_904_port, A_ns(7) => SHIFT_n_903_port, 
                           A_ns(6) => SHIFT_n_902_port, A_ns(5) => 
                           SHIFT_n_901_port, A_ns(4) => SHIFT_n_900_port, 
                           A_ns(3) => SHIFT_n_899_port, A_ns(2) => 
                           SHIFT_n_898_port, A_ns(1) => SHIFT_n_897_port, 
                           A_ns(0) => SHIFT_n_896_port, A_s(63) => 
                           SHIFT_959_port, A_s(62) => SHIFT_958_port, A_s(61) 
                           => SHIFT_957_port, A_s(60) => SHIFT_956_port, 
                           A_s(59) => SHIFT_955_port, A_s(58) => SHIFT_954_port
                           , A_s(57) => SHIFT_953_port, A_s(56) => 
                           SHIFT_952_port, A_s(55) => SHIFT_951_port, A_s(54) 
                           => SHIFT_950_port, A_s(53) => SHIFT_949_port, 
                           A_s(52) => SHIFT_948_port, A_s(51) => SHIFT_947_port
                           , A_s(50) => SHIFT_946_port, A_s(49) => 
                           SHIFT_945_port, A_s(48) => SHIFT_944_port, A_s(47) 
                           => SHIFT_943_port, A_s(46) => SHIFT_942_port, 
                           A_s(45) => SHIFT_941_port, A_s(44) => SHIFT_940_port
                           , A_s(43) => SHIFT_939_port, A_s(42) => 
                           SHIFT_938_port, A_s(41) => SHIFT_937_port, A_s(40) 
                           => SHIFT_936_port, A_s(39) => SHIFT_935_port, 
                           A_s(38) => SHIFT_934_port, A_s(37) => SHIFT_933_port
                           , A_s(36) => SHIFT_932_port, A_s(35) => 
                           SHIFT_931_port, A_s(34) => SHIFT_930_port, A_s(33) 
                           => SHIFT_929_port, A_s(32) => SHIFT_928_port, 
                           A_s(31) => SHIFT_927_port, A_s(30) => SHIFT_926_port
                           , A_s(29) => SHIFT_925_port, A_s(28) => 
                           SHIFT_924_port, A_s(27) => SHIFT_923_port, A_s(26) 
                           => SHIFT_922_port, A_s(25) => SHIFT_921_port, 
                           A_s(24) => SHIFT_920_port, A_s(23) => SHIFT_919_port
                           , A_s(22) => SHIFT_918_port, A_s(21) => 
                           SHIFT_917_port, A_s(20) => SHIFT_916_port, A_s(19) 
                           => SHIFT_915_port, A_s(18) => SHIFT_914_port, 
                           A_s(17) => SHIFT_913_port, A_s(16) => SHIFT_912_port
                           , A_s(15) => SHIFT_911_port, A_s(14) => 
                           SHIFT_910_port, A_s(13) => SHIFT_909_port, A_s(12) 
                           => SHIFT_908_port, A_s(11) => SHIFT_907_port, 
                           A_s(10) => SHIFT_906_port, A_s(9) => SHIFT_905_port,
                           A_s(8) => SHIFT_904_port, A_s(7) => SHIFT_903_port, 
                           A_s(6) => SHIFT_902_port, A_s(5) => SHIFT_901_port, 
                           A_s(4) => SHIFT_900_port, A_s(3) => SHIFT_899_port, 
                           A_s(2) => SHIFT_898_port, A_s(1) => SHIFT_897_port, 
                           A_s(0) => SHIFT_896_port, B(63) => B(31), B(62) => 
                           B(31), B(61) => B(31), B(60) => B(31), B(59) => 
                           B(31), B(58) => B(31), B(57) => B(31), B(56) => 
                           B(31), B(55) => B(31), B(54) => B(31), B(53) => 
                           B(31), B(52) => B(31), B(51) => B(31), B(50) => 
                           B(31), B(49) => B(31), B(48) => B(31), B(47) => 
                           B(31), B(46) => B(31), B(45) => B(31), B(44) => 
                           B(31), B(43) => B(31), B(42) => B(31), B(41) => 
                           B(31), B(40) => B(31), B(39) => B(31), B(38) => 
                           B(31), B(37) => B(31), B(36) => B(31), B(35) => 
                           B(31), B(34) => B(31), B(33) => B(31), B(32) => 
                           B(31), B(31) => B(31), B(30) => B(30), B(29) => 
                           B(29), B(28) => B(28), B(27) => B(27), B(26) => 
                           B(26), B(25) => B(25), B(24) => B(24), B(23) => 
                           B(23), B(22) => B(22), B(21) => B(21), B(20) => 
                           B(20), B(19) => B(19), B(18) => B(18), B(17) => 
                           B(17), B(16) => B(16), B(15) => B(15), B(14) => 
                           B(14), B(13) => B(13), B(12) => B(12), B(11) => 
                           B(11), B(10) => B(10), B(9) => B(9), B(8) => B(8), 
                           B(7) => B(7), B(6) => B(6), B(5) => B(5), B(4) => 
                           B(4), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), O(63) => OTMP_959_port, O(62) => 
                           OTMP_958_port, O(61) => OTMP_957_port, O(60) => 
                           OTMP_956_port, O(59) => OTMP_955_port, O(58) => 
                           OTMP_954_port, O(57) => OTMP_953_port, O(56) => 
                           OTMP_952_port, O(55) => OTMP_951_port, O(54) => 
                           OTMP_950_port, O(53) => OTMP_949_port, O(52) => 
                           OTMP_948_port, O(51) => OTMP_947_port, O(50) => 
                           OTMP_946_port, O(49) => OTMP_945_port, O(48) => 
                           OTMP_944_port, O(47) => OTMP_943_port, O(46) => 
                           OTMP_942_port, O(45) => OTMP_941_port, O(44) => 
                           OTMP_940_port, O(43) => OTMP_939_port, O(42) => 
                           OTMP_938_port, O(41) => OTMP_937_port, O(40) => 
                           OTMP_936_port, O(39) => OTMP_935_port, O(38) => 
                           OTMP_934_port, O(37) => OTMP_933_port, O(36) => 
                           OTMP_932_port, O(35) => OTMP_931_port, O(34) => 
                           OTMP_930_port, O(33) => OTMP_929_port, O(32) => 
                           OTMP_928_port, O(31) => OTMP_927_port, O(30) => 
                           OTMP_926_port, O(29) => OTMP_925_port, O(28) => 
                           OTMP_924_port, O(27) => OTMP_923_port, O(26) => 
                           OTMP_922_port, O(25) => OTMP_921_port, O(24) => 
                           OTMP_920_port, O(23) => OTMP_919_port, O(22) => 
                           OTMP_918_port, O(21) => OTMP_917_port, O(20) => 
                           OTMP_916_port, O(19) => OTMP_915_port, O(18) => 
                           OTMP_914_port, O(17) => OTMP_913_port, O(16) => 
                           OTMP_912_port, O(15) => OTMP_911_port, O(14) => 
                           OTMP_910_port, O(13) => OTMP_909_port, O(12) => 
                           OTMP_908_port, O(11) => OTMP_907_port, O(10) => 
                           OTMP_906_port, O(9) => OTMP_905_port, O(8) => 
                           OTMP_904_port, O(7) => OTMP_903_port, O(6) => 
                           OTMP_902_port, O(5) => OTMP_901_port, O(4) => 
                           OTMP_900_port, O(3) => OTMP_899_port, O(2) => 
                           OTMP_898_port, O(1) => OTMP_897_port, O(0) => n_1161
                           , A_so(63) => SHIFT_1023_port, A_so(62) => 
                           SHIFT_1022_port, A_so(61) => SHIFT_1021_port, 
                           A_so(60) => SHIFT_1020_port, A_so(59) => 
                           SHIFT_1019_port, A_so(58) => SHIFT_1018_port, 
                           A_so(57) => SHIFT_1017_port, A_so(56) => 
                           SHIFT_1016_port, A_so(55) => SHIFT_1015_port, 
                           A_so(54) => SHIFT_1014_port, A_so(53) => 
                           SHIFT_1013_port, A_so(52) => SHIFT_1012_port, 
                           A_so(51) => SHIFT_1011_port, A_so(50) => 
                           SHIFT_1010_port, A_so(49) => SHIFT_1009_port, 
                           A_so(48) => SHIFT_1008_port, A_so(47) => 
                           SHIFT_1007_port, A_so(46) => SHIFT_1006_port, 
                           A_so(45) => SHIFT_1005_port, A_so(44) => 
                           SHIFT_1004_port, A_so(43) => SHIFT_1003_port, 
                           A_so(42) => SHIFT_1002_port, A_so(41) => 
                           SHIFT_1001_port, A_so(40) => SHIFT_1000_port, 
                           A_so(39) => SHIFT_999_port, A_so(38) => 
                           SHIFT_998_port, A_so(37) => SHIFT_997_port, A_so(36)
                           => SHIFT_996_port, A_so(35) => SHIFT_995_port, 
                           A_so(34) => SHIFT_994_port, A_so(33) => 
                           SHIFT_993_port, A_so(32) => SHIFT_992_port, A_so(31)
                           => SHIFT_991_port, A_so(30) => SHIFT_990_port, 
                           A_so(29) => SHIFT_989_port, A_so(28) => 
                           SHIFT_988_port, A_so(27) => SHIFT_987_port, A_so(26)
                           => SHIFT_986_port, A_so(25) => SHIFT_985_port, 
                           A_so(24) => SHIFT_984_port, A_so(23) => 
                           SHIFT_983_port, A_so(22) => SHIFT_982_port, A_so(21)
                           => SHIFT_981_port, A_so(20) => SHIFT_980_port, 
                           A_so(19) => SHIFT_979_port, A_so(18) => 
                           SHIFT_978_port, A_so(17) => SHIFT_977_port, A_so(16)
                           => SHIFT_976_port, A_so(15) => SHIFT_975_port, 
                           A_so(14) => SHIFT_974_port, A_so(13) => 
                           SHIFT_973_port, A_so(12) => SHIFT_972_port, A_so(11)
                           => SHIFT_971_port, A_so(10) => SHIFT_970_port, 
                           A_so(9) => SHIFT_969_port, A_so(8) => SHIFT_968_port
                           , A_so(7) => SHIFT_967_port, A_so(6) => 
                           SHIFT_966_port, A_so(5) => SHIFT_965_port, A_so(4) 
                           => SHIFT_964_port, A_so(3) => SHIFT_963_port, 
                           A_so(2) => SHIFT_962_port, A_so(1) => n_1162, 
                           A_so(0) => n_1163, A_nso(63) => SHIFT_n_1023_port, 
                           A_nso(62) => SHIFT_n_1022_port, A_nso(61) => 
                           SHIFT_n_1021_port, A_nso(60) => SHIFT_n_1020_port, 
                           A_nso(59) => SHIFT_n_1019_port, A_nso(58) => 
                           SHIFT_n_1018_port, A_nso(57) => SHIFT_n_1017_port, 
                           A_nso(56) => SHIFT_n_1016_port, A_nso(55) => 
                           SHIFT_n_1015_port, A_nso(54) => SHIFT_n_1014_port, 
                           A_nso(53) => SHIFT_n_1013_port, A_nso(52) => 
                           SHIFT_n_1012_port, A_nso(51) => SHIFT_n_1011_port, 
                           A_nso(50) => SHIFT_n_1010_port, A_nso(49) => 
                           SHIFT_n_1009_port, A_nso(48) => SHIFT_n_1008_port, 
                           A_nso(47) => SHIFT_n_1007_port, A_nso(46) => 
                           SHIFT_n_1006_port, A_nso(45) => SHIFT_n_1005_port, 
                           A_nso(44) => SHIFT_n_1004_port, A_nso(43) => 
                           SHIFT_n_1003_port, A_nso(42) => SHIFT_n_1002_port, 
                           A_nso(41) => SHIFT_n_1001_port, A_nso(40) => 
                           SHIFT_n_1000_port, A_nso(39) => SHIFT_n_999_port, 
                           A_nso(38) => SHIFT_n_998_port, A_nso(37) => 
                           SHIFT_n_997_port, A_nso(36) => SHIFT_n_996_port, 
                           A_nso(35) => SHIFT_n_995_port, A_nso(34) => 
                           SHIFT_n_994_port, A_nso(33) => SHIFT_n_993_port, 
                           A_nso(32) => SHIFT_n_992_port, A_nso(31) => 
                           SHIFT_n_991_port, A_nso(30) => SHIFT_n_990_port, 
                           A_nso(29) => SHIFT_n_989_port, A_nso(28) => 
                           SHIFT_n_988_port, A_nso(27) => SHIFT_n_987_port, 
                           A_nso(26) => SHIFT_n_986_port, A_nso(25) => 
                           SHIFT_n_985_port, A_nso(24) => SHIFT_n_984_port, 
                           A_nso(23) => SHIFT_n_983_port, A_nso(22) => 
                           SHIFT_n_982_port, A_nso(21) => SHIFT_n_981_port, 
                           A_nso(20) => SHIFT_n_980_port, A_nso(19) => 
                           SHIFT_n_979_port, A_nso(18) => SHIFT_n_978_port, 
                           A_nso(17) => SHIFT_n_977_port, A_nso(16) => 
                           SHIFT_n_976_port, A_nso(15) => SHIFT_n_975_port, 
                           A_nso(14) => SHIFT_n_974_port, A_nso(13) => 
                           SHIFT_n_973_port, A_nso(12) => SHIFT_n_972_port, 
                           A_nso(11) => SHIFT_n_971_port, A_nso(10) => 
                           SHIFT_n_970_port, A_nso(9) => SHIFT_n_969_port, 
                           A_nso(8) => SHIFT_n_968_port, A_nso(7) => 
                           SHIFT_n_967_port, A_nso(6) => SHIFT_n_966_port, 
                           A_nso(5) => SHIFT_n_965_port, A_nso(4) => 
                           SHIFT_n_964_port, A_nso(3) => SHIFT_n_963_port, 
                           A_nso(2) => SHIFT_n_962_port, A_nso(1) => n_1164, 
                           A_nso(0) => n_1165);
   BOOTHENC_I_16 : BOOTHENC_NBIT64_i30 port map( A(63) => net46772, A(62) => 
                           net46773, A(61) => net46774, A(60) => net46775, 
                           A(59) => net46776, A(58) => net46777, A(57) => 
                           net46778, A(56) => net46779, A(55) => net46780, 
                           A(54) => net46781, A(53) => net46782, A(52) => 
                           net46783, A(51) => net46784, A(50) => net46785, 
                           A(49) => net46786, A(48) => net46787, A(47) => 
                           net46788, A(46) => net46789, A(45) => net46790, 
                           A(44) => net46791, A(43) => net46792, A(42) => 
                           net46793, A(41) => net46794, A(40) => net46795, 
                           A(39) => net46796, A(38) => net46797, A(37) => 
                           net46798, A(36) => net46799, A(35) => net46800, 
                           A(34) => net46801, A(33) => net46802, A(32) => 
                           net46803, A(31) => net46804, A(30) => net46805, 
                           A(29) => net46806, A(28) => net46807, A(27) => 
                           net46808, A(26) => net46809, A(25) => net46810, 
                           A(24) => net46811, A(23) => net46812, A(22) => 
                           net46813, A(21) => net46814, A(20) => net46815, 
                           A(19) => net46816, A(18) => net46817, A(17) => 
                           net46818, A(16) => net46819, A(15) => net46820, 
                           A(14) => net46821, A(13) => net46822, A(12) => 
                           net46823, A(11) => net46824, A(10) => net46825, A(9)
                           => net46826, A(8) => net46827, A(7) => net46828, 
                           A(6) => net46829, A(5) => net46830, A(4) => net46831
                           , A(3) => net46832, A(2) => net46833, A(1) => 
                           net46834, A(0) => net46835, A_n(63) => net46836, 
                           A_n(62) => net46837, A_n(61) => net46838, A_n(60) =>
                           net46839, A_n(59) => net46840, A_n(58) => net46841, 
                           A_n(57) => net46842, A_n(56) => net46843, A_n(55) =>
                           net46844, A_n(54) => net46845, A_n(53) => net46846, 
                           A_n(52) => net46847, A_n(51) => net46848, A_n(50) =>
                           net46849, A_n(49) => net46850, A_n(48) => net46851, 
                           A_n(47) => net46852, A_n(46) => net46853, A_n(45) =>
                           net46854, A_n(44) => net46855, A_n(43) => net46856, 
                           A_n(42) => net46857, A_n(41) => net46858, A_n(40) =>
                           net46859, A_n(39) => net46860, A_n(38) => net46861, 
                           A_n(37) => net46862, A_n(36) => net46863, A_n(35) =>
                           net46864, A_n(34) => net46865, A_n(33) => net46866, 
                           A_n(32) => net46867, A_n(31) => net46868, A_n(30) =>
                           net46869, A_n(29) => net46870, A_n(28) => net46871, 
                           A_n(27) => net46872, A_n(26) => net46873, A_n(25) =>
                           net46874, A_n(24) => net46875, A_n(23) => net46876, 
                           A_n(22) => net46877, A_n(21) => net46878, A_n(20) =>
                           net46879, A_n(19) => net46880, A_n(18) => net46881, 
                           A_n(17) => net46882, A_n(16) => net46883, A_n(15) =>
                           net46884, A_n(14) => net46885, A_n(13) => net46886, 
                           A_n(12) => net46887, A_n(11) => net46888, A_n(10) =>
                           net46889, A_n(9) => net46890, A_n(8) => net46891, 
                           A_n(7) => net46892, A_n(6) => net46893, A_n(5) => 
                           net46894, A_n(4) => net46895, A_n(3) => net46896, 
                           A_n(2) => net46897, A_n(1) => net46898, A_n(0) => 
                           net46899, A_ns(63) => SHIFT_n_1023_port, A_ns(62) =>
                           SHIFT_n_1022_port, A_ns(61) => SHIFT_n_1021_port, 
                           A_ns(60) => SHIFT_n_1020_port, A_ns(59) => 
                           SHIFT_n_1019_port, A_ns(58) => SHIFT_n_1018_port, 
                           A_ns(57) => SHIFT_n_1017_port, A_ns(56) => 
                           SHIFT_n_1016_port, A_ns(55) => SHIFT_n_1015_port, 
                           A_ns(54) => SHIFT_n_1014_port, A_ns(53) => 
                           SHIFT_n_1013_port, A_ns(52) => SHIFT_n_1012_port, 
                           A_ns(51) => SHIFT_n_1011_port, A_ns(50) => 
                           SHIFT_n_1010_port, A_ns(49) => SHIFT_n_1009_port, 
                           A_ns(48) => SHIFT_n_1008_port, A_ns(47) => 
                           SHIFT_n_1007_port, A_ns(46) => SHIFT_n_1006_port, 
                           A_ns(45) => SHIFT_n_1005_port, A_ns(44) => 
                           SHIFT_n_1004_port, A_ns(43) => SHIFT_n_1003_port, 
                           A_ns(42) => SHIFT_n_1002_port, A_ns(41) => 
                           SHIFT_n_1001_port, A_ns(40) => SHIFT_n_1000_port, 
                           A_ns(39) => SHIFT_n_999_port, A_ns(38) => 
                           SHIFT_n_998_port, A_ns(37) => SHIFT_n_997_port, 
                           A_ns(36) => SHIFT_n_996_port, A_ns(35) => 
                           SHIFT_n_995_port, A_ns(34) => SHIFT_n_994_port, 
                           A_ns(33) => SHIFT_n_993_port, A_ns(32) => 
                           SHIFT_n_992_port, A_ns(31) => SHIFT_n_991_port, 
                           A_ns(30) => SHIFT_n_990_port, A_ns(29) => 
                           SHIFT_n_989_port, A_ns(28) => SHIFT_n_988_port, 
                           A_ns(27) => SHIFT_n_987_port, A_ns(26) => 
                           SHIFT_n_986_port, A_ns(25) => SHIFT_n_985_port, 
                           A_ns(24) => SHIFT_n_984_port, A_ns(23) => 
                           SHIFT_n_983_port, A_ns(22) => SHIFT_n_982_port, 
                           A_ns(21) => SHIFT_n_981_port, A_ns(20) => 
                           SHIFT_n_980_port, A_ns(19) => SHIFT_n_979_port, 
                           A_ns(18) => SHIFT_n_978_port, A_ns(17) => 
                           SHIFT_n_977_port, A_ns(16) => SHIFT_n_976_port, 
                           A_ns(15) => SHIFT_n_975_port, A_ns(14) => 
                           SHIFT_n_974_port, A_ns(13) => SHIFT_n_973_port, 
                           A_ns(12) => SHIFT_n_972_port, A_ns(11) => 
                           SHIFT_n_971_port, A_ns(10) => SHIFT_n_970_port, 
                           A_ns(9) => SHIFT_n_969_port, A_ns(8) => 
                           SHIFT_n_968_port, A_ns(7) => SHIFT_n_967_port, 
                           A_ns(6) => SHIFT_n_966_port, A_ns(5) => 
                           SHIFT_n_965_port, A_ns(4) => SHIFT_n_964_port, 
                           A_ns(3) => SHIFT_n_963_port, A_ns(2) => 
                           SHIFT_n_962_port, A_ns(1) => SHIFT_n_961_port, 
                           A_ns(0) => SHIFT_n_960_port, A_s(63) => 
                           SHIFT_1023_port, A_s(62) => SHIFT_1022_port, A_s(61)
                           => SHIFT_1021_port, A_s(60) => SHIFT_1020_port, 
                           A_s(59) => SHIFT_1019_port, A_s(58) => 
                           SHIFT_1018_port, A_s(57) => SHIFT_1017_port, A_s(56)
                           => SHIFT_1016_port, A_s(55) => SHIFT_1015_port, 
                           A_s(54) => SHIFT_1014_port, A_s(53) => 
                           SHIFT_1013_port, A_s(52) => SHIFT_1012_port, A_s(51)
                           => SHIFT_1011_port, A_s(50) => SHIFT_1010_port, 
                           A_s(49) => SHIFT_1009_port, A_s(48) => 
                           SHIFT_1008_port, A_s(47) => SHIFT_1007_port, A_s(46)
                           => SHIFT_1006_port, A_s(45) => SHIFT_1005_port, 
                           A_s(44) => SHIFT_1004_port, A_s(43) => 
                           SHIFT_1003_port, A_s(42) => SHIFT_1002_port, A_s(41)
                           => SHIFT_1001_port, A_s(40) => SHIFT_1000_port, 
                           A_s(39) => SHIFT_999_port, A_s(38) => SHIFT_998_port
                           , A_s(37) => SHIFT_997_port, A_s(36) => 
                           SHIFT_996_port, A_s(35) => SHIFT_995_port, A_s(34) 
                           => SHIFT_994_port, A_s(33) => SHIFT_993_port, 
                           A_s(32) => SHIFT_992_port, A_s(31) => SHIFT_991_port
                           , A_s(30) => SHIFT_990_port, A_s(29) => 
                           SHIFT_989_port, A_s(28) => SHIFT_988_port, A_s(27) 
                           => SHIFT_987_port, A_s(26) => SHIFT_986_port, 
                           A_s(25) => SHIFT_985_port, A_s(24) => SHIFT_984_port
                           , A_s(23) => SHIFT_983_port, A_s(22) => 
                           SHIFT_982_port, A_s(21) => SHIFT_981_port, A_s(20) 
                           => SHIFT_980_port, A_s(19) => SHIFT_979_port, 
                           A_s(18) => SHIFT_978_port, A_s(17) => SHIFT_977_port
                           , A_s(16) => SHIFT_976_port, A_s(15) => 
                           SHIFT_975_port, A_s(14) => SHIFT_974_port, A_s(13) 
                           => SHIFT_973_port, A_s(12) => SHIFT_972_port, 
                           A_s(11) => SHIFT_971_port, A_s(10) => SHIFT_970_port
                           , A_s(9) => SHIFT_969_port, A_s(8) => SHIFT_968_port
                           , A_s(7) => SHIFT_967_port, A_s(6) => SHIFT_966_port
                           , A_s(5) => SHIFT_965_port, A_s(4) => SHIFT_964_port
                           , A_s(3) => SHIFT_963_port, A_s(2) => SHIFT_962_port
                           , A_s(1) => SHIFT_961_port, A_s(0) => SHIFT_960_port
                           , B(63) => B(31), B(62) => B(31), B(61) => B(31), 
                           B(60) => B(31), B(59) => B(31), B(58) => B(31), 
                           B(57) => B(31), B(56) => B(31), B(55) => B(31), 
                           B(54) => B(31), B(53) => B(31), B(52) => B(31), 
                           B(51) => B(31), B(50) => B(31), B(49) => B(31), 
                           B(48) => B(31), B(47) => B(31), B(46) => B(31), 
                           B(45) => B(31), B(44) => B(31), B(43) => B(31), 
                           B(42) => B(31), B(41) => B(31), B(40) => B(31), 
                           B(39) => B(31), B(38) => B(31), B(37) => B(31), 
                           B(36) => B(31), B(35) => B(31), B(34) => B(31), 
                           B(33) => B(31), B(32) => B(31), B(31) => B(31), 
                           B(30) => B(30), B(29) => B(29), B(28) => B(28), 
                           B(27) => B(27), B(26) => B(26), B(25) => B(25), 
                           B(24) => B(24), B(23) => B(23), B(22) => B(22), 
                           B(21) => B(21), B(20) => B(20), B(19) => B(19), 
                           B(18) => B(18), B(17) => B(17), B(16) => B(16), 
                           B(15) => B(15), B(14) => B(14), B(13) => B(13), 
                           B(12) => B(12), B(11) => B(11), B(10) => B(10), B(9)
                           => B(9), B(8) => B(8), B(7) => B(7), B(6) => B(6), 
                           B(5) => B(5), B(4) => B(4), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => B(0), O(63) => 
                           OTMP_1023_port, O(62) => OTMP_1022_port, O(61) => 
                           OTMP_1021_port, O(60) => OTMP_1020_port, O(59) => 
                           OTMP_1019_port, O(58) => OTMP_1018_port, O(57) => 
                           OTMP_1017_port, O(56) => OTMP_1016_port, O(55) => 
                           OTMP_1015_port, O(54) => OTMP_1014_port, O(53) => 
                           OTMP_1013_port, O(52) => OTMP_1012_port, O(51) => 
                           OTMP_1011_port, O(50) => OTMP_1010_port, O(49) => 
                           OTMP_1009_port, O(48) => OTMP_1008_port, O(47) => 
                           OTMP_1007_port, O(46) => OTMP_1006_port, O(45) => 
                           OTMP_1005_port, O(44) => OTMP_1004_port, O(43) => 
                           OTMP_1003_port, O(42) => OTMP_1002_port, O(41) => 
                           OTMP_1001_port, O(40) => OTMP_1000_port, O(39) => 
                           OTMP_999_port, O(38) => OTMP_998_port, O(37) => 
                           OTMP_997_port, O(36) => OTMP_996_port, O(35) => 
                           OTMP_995_port, O(34) => OTMP_994_port, O(33) => 
                           OTMP_993_port, O(32) => OTMP_992_port, O(31) => 
                           OTMP_991_port, O(30) => OTMP_990_port, O(29) => 
                           OTMP_989_port, O(28) => OTMP_988_port, O(27) => 
                           OTMP_987_port, O(26) => OTMP_986_port, O(25) => 
                           OTMP_985_port, O(24) => OTMP_984_port, O(23) => 
                           OTMP_983_port, O(22) => OTMP_982_port, O(21) => 
                           OTMP_981_port, O(20) => OTMP_980_port, O(19) => 
                           OTMP_979_port, O(18) => OTMP_978_port, O(17) => 
                           OTMP_977_port, O(16) => OTMP_976_port, O(15) => 
                           OTMP_975_port, O(14) => OTMP_974_port, O(13) => 
                           OTMP_973_port, O(12) => OTMP_972_port, O(11) => 
                           OTMP_971_port, O(10) => OTMP_970_port, O(9) => 
                           OTMP_969_port, O(8) => OTMP_968_port, O(7) => 
                           OTMP_967_port, O(6) => OTMP_966_port, O(5) => 
                           OTMP_965_port, O(4) => OTMP_964_port, O(3) => 
                           OTMP_963_port, O(2) => OTMP_962_port, O(1) => 
                           OTMP_961_port, O(0) => n_1166, A_so(63) => n_1167, 
                           A_so(62) => n_1168, A_so(61) => n_1169, A_so(60) => 
                           n_1170, A_so(59) => n_1171, A_so(58) => n_1172, 
                           A_so(57) => n_1173, A_so(56) => n_1174, A_so(55) => 
                           n_1175, A_so(54) => n_1176, A_so(53) => n_1177, 
                           A_so(52) => n_1178, A_so(51) => n_1179, A_so(50) => 
                           n_1180, A_so(49) => n_1181, A_so(48) => n_1182, 
                           A_so(47) => n_1183, A_so(46) => n_1184, A_so(45) => 
                           n_1185, A_so(44) => n_1186, A_so(43) => n_1187, 
                           A_so(42) => n_1188, A_so(41) => n_1189, A_so(40) => 
                           n_1190, A_so(39) => n_1191, A_so(38) => n_1192, 
                           A_so(37) => n_1193, A_so(36) => n_1194, A_so(35) => 
                           n_1195, A_so(34) => n_1196, A_so(33) => n_1197, 
                           A_so(32) => n_1198, A_so(31) => n_1199, A_so(30) => 
                           n_1200, A_so(29) => n_1201, A_so(28) => n_1202, 
                           A_so(27) => n_1203, A_so(26) => n_1204, A_so(25) => 
                           n_1205, A_so(24) => n_1206, A_so(23) => n_1207, 
                           A_so(22) => n_1208, A_so(21) => n_1209, A_so(20) => 
                           n_1210, A_so(19) => n_1211, A_so(18) => n_1212, 
                           A_so(17) => n_1213, A_so(16) => n_1214, A_so(15) => 
                           n_1215, A_so(14) => n_1216, A_so(13) => n_1217, 
                           A_so(12) => n_1218, A_so(11) => n_1219, A_so(10) => 
                           n_1220, A_so(9) => n_1221, A_so(8) => n_1222, 
                           A_so(7) => n_1223, A_so(6) => n_1224, A_so(5) => 
                           n_1225, A_so(4) => n_1226, A_so(3) => n_1227, 
                           A_so(2) => n_1228, A_so(1) => n_1229, A_so(0) => 
                           n_1230, A_nso(63) => n_1231, A_nso(62) => n_1232, 
                           A_nso(61) => n_1233, A_nso(60) => n_1234, A_nso(59) 
                           => n_1235, A_nso(58) => n_1236, A_nso(57) => n_1237,
                           A_nso(56) => n_1238, A_nso(55) => n_1239, A_nso(54) 
                           => n_1240, A_nso(53) => n_1241, A_nso(52) => n_1242,
                           A_nso(51) => n_1243, A_nso(50) => n_1244, A_nso(49) 
                           => n_1245, A_nso(48) => n_1246, A_nso(47) => n_1247,
                           A_nso(46) => n_1248, A_nso(45) => n_1249, A_nso(44) 
                           => n_1250, A_nso(43) => n_1251, A_nso(42) => n_1252,
                           A_nso(41) => n_1253, A_nso(40) => n_1254, A_nso(39) 
                           => n_1255, A_nso(38) => n_1256, A_nso(37) => n_1257,
                           A_nso(36) => n_1258, A_nso(35) => n_1259, A_nso(34) 
                           => n_1260, A_nso(33) => n_1261, A_nso(32) => n_1262,
                           A_nso(31) => n_1263, A_nso(30) => n_1264, A_nso(29) 
                           => n_1265, A_nso(28) => n_1266, A_nso(27) => n_1267,
                           A_nso(26) => n_1268, A_nso(25) => n_1269, A_nso(24) 
                           => n_1270, A_nso(23) => n_1271, A_nso(22) => n_1272,
                           A_nso(21) => n_1273, A_nso(20) => n_1274, A_nso(19) 
                           => n_1275, A_nso(18) => n_1276, A_nso(17) => n_1277,
                           A_nso(16) => n_1278, A_nso(15) => n_1279, A_nso(14) 
                           => n_1280, A_nso(13) => n_1281, A_nso(12) => n_1282,
                           A_nso(11) => n_1283, A_nso(10) => n_1284, A_nso(9) 
                           => n_1285, A_nso(8) => n_1286, A_nso(7) => n_1287, 
                           A_nso(6) => n_1288, A_nso(5) => n_1289, A_nso(4) => 
                           n_1290, A_nso(3) => n_1291, A_nso(2) => n_1292, 
                           A_nso(1) => n_1293, A_nso(0) => n_1294);
   ADDER2_2 : RCA_NBIT64_15 port map( A(63) => OTMP_63_port, A(62) => 
                           OTMP_62_port, A(61) => OTMP_61_port, A(60) => 
                           OTMP_60_port, A(59) => OTMP_59_port, A(58) => 
                           OTMP_58_port, A(57) => OTMP_57_port, A(56) => 
                           OTMP_56_port, A(55) => OTMP_55_port, A(54) => 
                           OTMP_54_port, A(53) => OTMP_53_port, A(52) => 
                           OTMP_52_port, A(51) => OTMP_51_port, A(50) => 
                           OTMP_50_port, A(49) => OTMP_49_port, A(48) => 
                           OTMP_48_port, A(47) => OTMP_47_port, A(46) => 
                           OTMP_46_port, A(45) => OTMP_45_port, A(44) => 
                           OTMP_44_port, A(43) => OTMP_43_port, A(42) => 
                           OTMP_42_port, A(41) => OTMP_41_port, A(40) => 
                           OTMP_40_port, A(39) => OTMP_39_port, A(38) => 
                           OTMP_38_port, A(37) => OTMP_37_port, A(36) => 
                           OTMP_36_port, A(35) => OTMP_35_port, A(34) => 
                           OTMP_34_port, A(33) => OTMP_33_port, A(32) => 
                           OTMP_32_port, A(31) => OTMP_31_port, A(30) => 
                           OTMP_30_port, A(29) => OTMP_29_port, A(28) => 
                           OTMP_28_port, A(27) => OTMP_27_port, A(26) => 
                           OTMP_26_port, A(25) => OTMP_25_port, A(24) => 
                           OTMP_24_port, A(23) => OTMP_23_port, A(22) => 
                           OTMP_22_port, A(21) => OTMP_21_port, A(20) => 
                           OTMP_20_port, A(19) => OTMP_19_port, A(18) => 
                           OTMP_18_port, A(17) => OTMP_17_port, A(16) => 
                           OTMP_16_port, A(15) => OTMP_15_port, A(14) => 
                           OTMP_14_port, A(13) => OTMP_13_port, A(12) => 
                           OTMP_12_port, A(11) => OTMP_11_port, A(10) => 
                           OTMP_10_port, A(9) => OTMP_9_port, A(8) => 
                           OTMP_8_port, A(7) => OTMP_7_port, A(6) => 
                           OTMP_6_port, A(5) => OTMP_5_port, A(4) => 
                           OTMP_4_port, A(3) => OTMP_3_port, A(2) => 
                           OTMP_2_port, A(1) => OTMP_1_port, A(0) => 
                           OTMP_0_port, B(63) => OTMP_127_port, B(62) => 
                           OTMP_126_port, B(61) => OTMP_125_port, B(60) => 
                           OTMP_124_port, B(59) => OTMP_123_port, B(58) => 
                           OTMP_122_port, B(57) => OTMP_121_port, B(56) => 
                           OTMP_120_port, B(55) => OTMP_119_port, B(54) => 
                           OTMP_118_port, B(53) => OTMP_117_port, B(52) => 
                           OTMP_116_port, B(51) => OTMP_115_port, B(50) => 
                           OTMP_114_port, B(49) => OTMP_113_port, B(48) => 
                           OTMP_112_port, B(47) => OTMP_111_port, B(46) => 
                           OTMP_110_port, B(45) => OTMP_109_port, B(44) => 
                           OTMP_108_port, B(43) => OTMP_107_port, B(42) => 
                           OTMP_106_port, B(41) => OTMP_105_port, B(40) => 
                           OTMP_104_port, B(39) => OTMP_103_port, B(38) => 
                           OTMP_102_port, B(37) => OTMP_101_port, B(36) => 
                           OTMP_100_port, B(35) => OTMP_99_port, B(34) => 
                           OTMP_98_port, B(33) => OTMP_97_port, B(32) => 
                           OTMP_96_port, B(31) => OTMP_95_port, B(30) => 
                           OTMP_94_port, B(29) => OTMP_93_port, B(28) => 
                           OTMP_92_port, B(27) => OTMP_91_port, B(26) => 
                           OTMP_90_port, B(25) => OTMP_89_port, B(24) => 
                           OTMP_88_port, B(23) => OTMP_87_port, B(22) => 
                           OTMP_86_port, B(21) => OTMP_85_port, B(20) => 
                           OTMP_84_port, B(19) => OTMP_83_port, B(18) => 
                           OTMP_82_port, B(17) => OTMP_81_port, B(16) => 
                           OTMP_80_port, B(15) => OTMP_79_port, B(14) => 
                           OTMP_78_port, B(13) => OTMP_77_port, B(12) => 
                           OTMP_76_port, B(11) => OTMP_75_port, B(10) => 
                           OTMP_74_port, B(9) => OTMP_73_port, B(8) => 
                           OTMP_72_port, B(7) => OTMP_71_port, B(6) => 
                           OTMP_70_port, B(5) => OTMP_69_port, B(4) => 
                           OTMP_68_port, B(3) => OTMP_67_port, B(2) => 
                           OTMP_66_port, B(1) => OTMP_65_port, B(0) => 
                           OTMP_64_port, Ci => X_Logic0_port, S(63) => 
                           PTMP_63_port, S(62) => PTMP_62_port, S(61) => 
                           PTMP_61_port, S(60) => PTMP_60_port, S(59) => 
                           PTMP_59_port, S(58) => PTMP_58_port, S(57) => 
                           PTMP_57_port, S(56) => PTMP_56_port, S(55) => 
                           PTMP_55_port, S(54) => PTMP_54_port, S(53) => 
                           PTMP_53_port, S(52) => PTMP_52_port, S(51) => 
                           PTMP_51_port, S(50) => PTMP_50_port, S(49) => 
                           PTMP_49_port, S(48) => PTMP_48_port, S(47) => 
                           PTMP_47_port, S(46) => PTMP_46_port, S(45) => 
                           PTMP_45_port, S(44) => PTMP_44_port, S(43) => 
                           PTMP_43_port, S(42) => PTMP_42_port, S(41) => 
                           PTMP_41_port, S(40) => PTMP_40_port, S(39) => 
                           PTMP_39_port, S(38) => PTMP_38_port, S(37) => 
                           PTMP_37_port, S(36) => PTMP_36_port, S(35) => 
                           PTMP_35_port, S(34) => PTMP_34_port, S(33) => 
                           PTMP_33_port, S(32) => PTMP_32_port, S(31) => 
                           PTMP_31_port, S(30) => PTMP_30_port, S(29) => 
                           PTMP_29_port, S(28) => PTMP_28_port, S(27) => 
                           PTMP_27_port, S(26) => PTMP_26_port, S(25) => 
                           PTMP_25_port, S(24) => PTMP_24_port, S(23) => 
                           PTMP_23_port, S(22) => PTMP_22_port, S(21) => 
                           PTMP_21_port, S(20) => PTMP_20_port, S(19) => 
                           PTMP_19_port, S(18) => PTMP_18_port, S(17) => 
                           PTMP_17_port, S(16) => PTMP_16_port, S(15) => 
                           PTMP_15_port, S(14) => PTMP_14_port, S(13) => 
                           PTMP_13_port, S(12) => PTMP_12_port, S(11) => 
                           PTMP_11_port, S(10) => PTMP_10_port, S(9) => 
                           PTMP_9_port, S(8) => PTMP_8_port, S(7) => 
                           PTMP_7_port, S(6) => PTMP_6_port, S(5) => 
                           PTMP_5_port, S(4) => PTMP_4_port, S(3) => 
                           PTMP_3_port, S(2) => PTMP_2_port, S(1) => 
                           PTMP_1_port, S(0) => PTMP_0_port, Co => n_1295);
   ADDERI_3 : RCA_NBIT64_29 port map( A(63) => PTMP_63_port, A(62) => 
                           PTMP_62_port, A(61) => PTMP_61_port, A(60) => 
                           PTMP_60_port, A(59) => PTMP_59_port, A(58) => 
                           PTMP_58_port, A(57) => PTMP_57_port, A(56) => 
                           PTMP_56_port, A(55) => PTMP_55_port, A(54) => 
                           PTMP_54_port, A(53) => PTMP_53_port, A(52) => 
                           PTMP_52_port, A(51) => PTMP_51_port, A(50) => 
                           PTMP_50_port, A(49) => PTMP_49_port, A(48) => 
                           PTMP_48_port, A(47) => PTMP_47_port, A(46) => 
                           PTMP_46_port, A(45) => PTMP_45_port, A(44) => 
                           PTMP_44_port, A(43) => PTMP_43_port, A(42) => 
                           PTMP_42_port, A(41) => PTMP_41_port, A(40) => 
                           PTMP_40_port, A(39) => PTMP_39_port, A(38) => 
                           PTMP_38_port, A(37) => PTMP_37_port, A(36) => 
                           PTMP_36_port, A(35) => PTMP_35_port, A(34) => 
                           PTMP_34_port, A(33) => PTMP_33_port, A(32) => 
                           PTMP_32_port, A(31) => PTMP_31_port, A(30) => 
                           PTMP_30_port, A(29) => PTMP_29_port, A(28) => 
                           PTMP_28_port, A(27) => PTMP_27_port, A(26) => 
                           PTMP_26_port, A(25) => PTMP_25_port, A(24) => 
                           PTMP_24_port, A(23) => PTMP_23_port, A(22) => 
                           PTMP_22_port, A(21) => PTMP_21_port, A(20) => 
                           PTMP_20_port, A(19) => PTMP_19_port, A(18) => 
                           PTMP_18_port, A(17) => PTMP_17_port, A(16) => 
                           PTMP_16_port, A(15) => PTMP_15_port, A(14) => 
                           PTMP_14_port, A(13) => PTMP_13_port, A(12) => 
                           PTMP_12_port, A(11) => PTMP_11_port, A(10) => 
                           PTMP_10_port, A(9) => PTMP_9_port, A(8) => 
                           PTMP_8_port, A(7) => PTMP_7_port, A(6) => 
                           PTMP_6_port, A(5) => PTMP_5_port, A(4) => 
                           PTMP_4_port, A(3) => PTMP_3_port, A(2) => 
                           PTMP_2_port, A(1) => PTMP_1_port, A(0) => 
                           PTMP_0_port, B(63) => OTMP_191_port, B(62) => 
                           OTMP_190_port, B(61) => OTMP_189_port, B(60) => 
                           OTMP_188_port, B(59) => OTMP_187_port, B(58) => 
                           OTMP_186_port, B(57) => OTMP_185_port, B(56) => 
                           OTMP_184_port, B(55) => OTMP_183_port, B(54) => 
                           OTMP_182_port, B(53) => OTMP_181_port, B(52) => 
                           OTMP_180_port, B(51) => OTMP_179_port, B(50) => 
                           OTMP_178_port, B(49) => OTMP_177_port, B(48) => 
                           OTMP_176_port, B(47) => OTMP_175_port, B(46) => 
                           OTMP_174_port, B(45) => OTMP_173_port, B(44) => 
                           OTMP_172_port, B(43) => OTMP_171_port, B(42) => 
                           OTMP_170_port, B(41) => OTMP_169_port, B(40) => 
                           OTMP_168_port, B(39) => OTMP_167_port, B(38) => 
                           OTMP_166_port, B(37) => OTMP_165_port, B(36) => 
                           OTMP_164_port, B(35) => OTMP_163_port, B(34) => 
                           OTMP_162_port, B(33) => OTMP_161_port, B(32) => 
                           OTMP_160_port, B(31) => OTMP_159_port, B(30) => 
                           OTMP_158_port, B(29) => OTMP_157_port, B(28) => 
                           OTMP_156_port, B(27) => OTMP_155_port, B(26) => 
                           OTMP_154_port, B(25) => OTMP_153_port, B(24) => 
                           OTMP_152_port, B(23) => OTMP_151_port, B(22) => 
                           OTMP_150_port, B(21) => OTMP_149_port, B(20) => 
                           OTMP_148_port, B(19) => OTMP_147_port, B(18) => 
                           OTMP_146_port, B(17) => OTMP_145_port, B(16) => 
                           OTMP_144_port, B(15) => OTMP_143_port, B(14) => 
                           OTMP_142_port, B(13) => OTMP_141_port, B(12) => 
                           OTMP_140_port, B(11) => OTMP_139_port, B(10) => 
                           OTMP_138_port, B(9) => OTMP_137_port, B(8) => 
                           OTMP_136_port, B(7) => OTMP_135_port, B(6) => 
                           OTMP_134_port, B(5) => OTMP_133_port, B(4) => 
                           OTMP_132_port, B(3) => OTMP_131_port, B(2) => 
                           OTMP_130_port, B(1) => OTMP_129_port, B(0) => 
                           OTMP_128_port, Ci => X_Logic0_port, S(63) => 
                           PTMP_127_port, S(62) => PTMP_126_port, S(61) => 
                           PTMP_125_port, S(60) => PTMP_124_port, S(59) => 
                           PTMP_123_port, S(58) => PTMP_122_port, S(57) => 
                           PTMP_121_port, S(56) => PTMP_120_port, S(55) => 
                           PTMP_119_port, S(54) => PTMP_118_port, S(53) => 
                           PTMP_117_port, S(52) => PTMP_116_port, S(51) => 
                           PTMP_115_port, S(50) => PTMP_114_port, S(49) => 
                           PTMP_113_port, S(48) => PTMP_112_port, S(47) => 
                           PTMP_111_port, S(46) => PTMP_110_port, S(45) => 
                           PTMP_109_port, S(44) => PTMP_108_port, S(43) => 
                           PTMP_107_port, S(42) => PTMP_106_port, S(41) => 
                           PTMP_105_port, S(40) => PTMP_104_port, S(39) => 
                           PTMP_103_port, S(38) => PTMP_102_port, S(37) => 
                           PTMP_101_port, S(36) => PTMP_100_port, S(35) => 
                           PTMP_99_port, S(34) => PTMP_98_port, S(33) => 
                           PTMP_97_port, S(32) => PTMP_96_port, S(31) => 
                           PTMP_95_port, S(30) => PTMP_94_port, S(29) => 
                           PTMP_93_port, S(28) => PTMP_92_port, S(27) => 
                           PTMP_91_port, S(26) => PTMP_90_port, S(25) => 
                           PTMP_89_port, S(24) => PTMP_88_port, S(23) => 
                           PTMP_87_port, S(22) => PTMP_86_port, S(21) => 
                           PTMP_85_port, S(20) => PTMP_84_port, S(19) => 
                           PTMP_83_port, S(18) => PTMP_82_port, S(17) => 
                           PTMP_81_port, S(16) => PTMP_80_port, S(15) => 
                           PTMP_79_port, S(14) => PTMP_78_port, S(13) => 
                           PTMP_77_port, S(12) => PTMP_76_port, S(11) => 
                           PTMP_75_port, S(10) => PTMP_74_port, S(9) => 
                           PTMP_73_port, S(8) => PTMP_72_port, S(7) => 
                           PTMP_71_port, S(6) => PTMP_70_port, S(5) => 
                           PTMP_69_port, S(4) => PTMP_68_port, S(3) => 
                           PTMP_67_port, S(2) => PTMP_66_port, S(1) => 
                           PTMP_65_port, S(0) => PTMP_64_port, Co => n_1296);
   ADDERI_4 : RCA_NBIT64_28 port map( A(63) => PTMP_127_port, A(62) => 
                           PTMP_126_port, A(61) => PTMP_125_port, A(60) => 
                           PTMP_124_port, A(59) => PTMP_123_port, A(58) => 
                           PTMP_122_port, A(57) => PTMP_121_port, A(56) => 
                           PTMP_120_port, A(55) => PTMP_119_port, A(54) => 
                           PTMP_118_port, A(53) => PTMP_117_port, A(52) => 
                           PTMP_116_port, A(51) => PTMP_115_port, A(50) => 
                           PTMP_114_port, A(49) => PTMP_113_port, A(48) => 
                           PTMP_112_port, A(47) => PTMP_111_port, A(46) => 
                           PTMP_110_port, A(45) => PTMP_109_port, A(44) => 
                           PTMP_108_port, A(43) => PTMP_107_port, A(42) => 
                           PTMP_106_port, A(41) => PTMP_105_port, A(40) => 
                           PTMP_104_port, A(39) => PTMP_103_port, A(38) => 
                           PTMP_102_port, A(37) => PTMP_101_port, A(36) => 
                           PTMP_100_port, A(35) => PTMP_99_port, A(34) => 
                           PTMP_98_port, A(33) => PTMP_97_port, A(32) => 
                           PTMP_96_port, A(31) => PTMP_95_port, A(30) => 
                           PTMP_94_port, A(29) => PTMP_93_port, A(28) => 
                           PTMP_92_port, A(27) => PTMP_91_port, A(26) => 
                           PTMP_90_port, A(25) => PTMP_89_port, A(24) => 
                           PTMP_88_port, A(23) => PTMP_87_port, A(22) => 
                           PTMP_86_port, A(21) => PTMP_85_port, A(20) => 
                           PTMP_84_port, A(19) => PTMP_83_port, A(18) => 
                           PTMP_82_port, A(17) => PTMP_81_port, A(16) => 
                           PTMP_80_port, A(15) => PTMP_79_port, A(14) => 
                           PTMP_78_port, A(13) => PTMP_77_port, A(12) => 
                           PTMP_76_port, A(11) => PTMP_75_port, A(10) => 
                           PTMP_74_port, A(9) => PTMP_73_port, A(8) => 
                           PTMP_72_port, A(7) => PTMP_71_port, A(6) => 
                           PTMP_70_port, A(5) => PTMP_69_port, A(4) => 
                           PTMP_68_port, A(3) => PTMP_67_port, A(2) => 
                           PTMP_66_port, A(1) => PTMP_65_port, A(0) => 
                           PTMP_64_port, B(63) => OTMP_255_port, B(62) => 
                           OTMP_254_port, B(61) => OTMP_253_port, B(60) => 
                           OTMP_252_port, B(59) => OTMP_251_port, B(58) => 
                           OTMP_250_port, B(57) => OTMP_249_port, B(56) => 
                           OTMP_248_port, B(55) => OTMP_247_port, B(54) => 
                           OTMP_246_port, B(53) => OTMP_245_port, B(52) => 
                           OTMP_244_port, B(51) => OTMP_243_port, B(50) => 
                           OTMP_242_port, B(49) => OTMP_241_port, B(48) => 
                           OTMP_240_port, B(47) => OTMP_239_port, B(46) => 
                           OTMP_238_port, B(45) => OTMP_237_port, B(44) => 
                           OTMP_236_port, B(43) => OTMP_235_port, B(42) => 
                           OTMP_234_port, B(41) => OTMP_233_port, B(40) => 
                           OTMP_232_port, B(39) => OTMP_231_port, B(38) => 
                           OTMP_230_port, B(37) => OTMP_229_port, B(36) => 
                           OTMP_228_port, B(35) => OTMP_227_port, B(34) => 
                           OTMP_226_port, B(33) => OTMP_225_port, B(32) => 
                           OTMP_224_port, B(31) => OTMP_223_port, B(30) => 
                           OTMP_222_port, B(29) => OTMP_221_port, B(28) => 
                           OTMP_220_port, B(27) => OTMP_219_port, B(26) => 
                           OTMP_218_port, B(25) => OTMP_217_port, B(24) => 
                           OTMP_216_port, B(23) => OTMP_215_port, B(22) => 
                           OTMP_214_port, B(21) => OTMP_213_port, B(20) => 
                           OTMP_212_port, B(19) => OTMP_211_port, B(18) => 
                           OTMP_210_port, B(17) => OTMP_209_port, B(16) => 
                           OTMP_208_port, B(15) => OTMP_207_port, B(14) => 
                           OTMP_206_port, B(13) => OTMP_205_port, B(12) => 
                           OTMP_204_port, B(11) => OTMP_203_port, B(10) => 
                           OTMP_202_port, B(9) => OTMP_201_port, B(8) => 
                           OTMP_200_port, B(7) => OTMP_199_port, B(6) => 
                           OTMP_198_port, B(5) => OTMP_197_port, B(4) => 
                           OTMP_196_port, B(3) => OTMP_195_port, B(2) => 
                           OTMP_194_port, B(1) => OTMP_193_port, B(0) => 
                           OTMP_192_port, Ci => X_Logic0_port, S(63) => 
                           PTMP_191_port, S(62) => PTMP_190_port, S(61) => 
                           PTMP_189_port, S(60) => PTMP_188_port, S(59) => 
                           PTMP_187_port, S(58) => PTMP_186_port, S(57) => 
                           PTMP_185_port, S(56) => PTMP_184_port, S(55) => 
                           PTMP_183_port, S(54) => PTMP_182_port, S(53) => 
                           PTMP_181_port, S(52) => PTMP_180_port, S(51) => 
                           PTMP_179_port, S(50) => PTMP_178_port, S(49) => 
                           PTMP_177_port, S(48) => PTMP_176_port, S(47) => 
                           PTMP_175_port, S(46) => PTMP_174_port, S(45) => 
                           PTMP_173_port, S(44) => PTMP_172_port, S(43) => 
                           PTMP_171_port, S(42) => PTMP_170_port, S(41) => 
                           PTMP_169_port, S(40) => PTMP_168_port, S(39) => 
                           PTMP_167_port, S(38) => PTMP_166_port, S(37) => 
                           PTMP_165_port, S(36) => PTMP_164_port, S(35) => 
                           PTMP_163_port, S(34) => PTMP_162_port, S(33) => 
                           PTMP_161_port, S(32) => PTMP_160_port, S(31) => 
                           PTMP_159_port, S(30) => PTMP_158_port, S(29) => 
                           PTMP_157_port, S(28) => PTMP_156_port, S(27) => 
                           PTMP_155_port, S(26) => PTMP_154_port, S(25) => 
                           PTMP_153_port, S(24) => PTMP_152_port, S(23) => 
                           PTMP_151_port, S(22) => PTMP_150_port, S(21) => 
                           PTMP_149_port, S(20) => PTMP_148_port, S(19) => 
                           PTMP_147_port, S(18) => PTMP_146_port, S(17) => 
                           PTMP_145_port, S(16) => PTMP_144_port, S(15) => 
                           PTMP_143_port, S(14) => PTMP_142_port, S(13) => 
                           PTMP_141_port, S(12) => PTMP_140_port, S(11) => 
                           PTMP_139_port, S(10) => PTMP_138_port, S(9) => 
                           PTMP_137_port, S(8) => PTMP_136_port, S(7) => 
                           PTMP_135_port, S(6) => PTMP_134_port, S(5) => 
                           PTMP_133_port, S(4) => PTMP_132_port, S(3) => 
                           PTMP_131_port, S(2) => PTMP_130_port, S(1) => 
                           PTMP_129_port, S(0) => PTMP_128_port, Co => n_1297);
   ADDERI_5 : RCA_NBIT64_27 port map( A(63) => PTMP_191_port, A(62) => 
                           PTMP_190_port, A(61) => PTMP_189_port, A(60) => 
                           PTMP_188_port, A(59) => PTMP_187_port, A(58) => 
                           PTMP_186_port, A(57) => PTMP_185_port, A(56) => 
                           PTMP_184_port, A(55) => PTMP_183_port, A(54) => 
                           PTMP_182_port, A(53) => PTMP_181_port, A(52) => 
                           PTMP_180_port, A(51) => PTMP_179_port, A(50) => 
                           PTMP_178_port, A(49) => PTMP_177_port, A(48) => 
                           PTMP_176_port, A(47) => PTMP_175_port, A(46) => 
                           PTMP_174_port, A(45) => PTMP_173_port, A(44) => 
                           PTMP_172_port, A(43) => PTMP_171_port, A(42) => 
                           PTMP_170_port, A(41) => PTMP_169_port, A(40) => 
                           PTMP_168_port, A(39) => PTMP_167_port, A(38) => 
                           PTMP_166_port, A(37) => PTMP_165_port, A(36) => 
                           PTMP_164_port, A(35) => PTMP_163_port, A(34) => 
                           PTMP_162_port, A(33) => PTMP_161_port, A(32) => 
                           PTMP_160_port, A(31) => PTMP_159_port, A(30) => 
                           PTMP_158_port, A(29) => PTMP_157_port, A(28) => 
                           PTMP_156_port, A(27) => PTMP_155_port, A(26) => 
                           PTMP_154_port, A(25) => PTMP_153_port, A(24) => 
                           PTMP_152_port, A(23) => PTMP_151_port, A(22) => 
                           PTMP_150_port, A(21) => PTMP_149_port, A(20) => 
                           PTMP_148_port, A(19) => PTMP_147_port, A(18) => 
                           PTMP_146_port, A(17) => PTMP_145_port, A(16) => 
                           PTMP_144_port, A(15) => PTMP_143_port, A(14) => 
                           PTMP_142_port, A(13) => PTMP_141_port, A(12) => 
                           PTMP_140_port, A(11) => PTMP_139_port, A(10) => 
                           PTMP_138_port, A(9) => PTMP_137_port, A(8) => 
                           PTMP_136_port, A(7) => PTMP_135_port, A(6) => 
                           PTMP_134_port, A(5) => PTMP_133_port, A(4) => 
                           PTMP_132_port, A(3) => PTMP_131_port, A(2) => 
                           PTMP_130_port, A(1) => PTMP_129_port, A(0) => 
                           PTMP_128_port, B(63) => OTMP_319_port, B(62) => 
                           OTMP_318_port, B(61) => OTMP_317_port, B(60) => 
                           OTMP_316_port, B(59) => OTMP_315_port, B(58) => 
                           OTMP_314_port, B(57) => OTMP_313_port, B(56) => 
                           OTMP_312_port, B(55) => OTMP_311_port, B(54) => 
                           OTMP_310_port, B(53) => OTMP_309_port, B(52) => 
                           OTMP_308_port, B(51) => OTMP_307_port, B(50) => 
                           OTMP_306_port, B(49) => OTMP_305_port, B(48) => 
                           OTMP_304_port, B(47) => OTMP_303_port, B(46) => 
                           OTMP_302_port, B(45) => OTMP_301_port, B(44) => 
                           OTMP_300_port, B(43) => OTMP_299_port, B(42) => 
                           OTMP_298_port, B(41) => OTMP_297_port, B(40) => 
                           OTMP_296_port, B(39) => OTMP_295_port, B(38) => 
                           OTMP_294_port, B(37) => OTMP_293_port, B(36) => 
                           OTMP_292_port, B(35) => OTMP_291_port, B(34) => 
                           OTMP_290_port, B(33) => OTMP_289_port, B(32) => 
                           OTMP_288_port, B(31) => OTMP_287_port, B(30) => 
                           OTMP_286_port, B(29) => OTMP_285_port, B(28) => 
                           OTMP_284_port, B(27) => OTMP_283_port, B(26) => 
                           OTMP_282_port, B(25) => OTMP_281_port, B(24) => 
                           OTMP_280_port, B(23) => OTMP_279_port, B(22) => 
                           OTMP_278_port, B(21) => OTMP_277_port, B(20) => 
                           OTMP_276_port, B(19) => OTMP_275_port, B(18) => 
                           OTMP_274_port, B(17) => OTMP_273_port, B(16) => 
                           OTMP_272_port, B(15) => OTMP_271_port, B(14) => 
                           OTMP_270_port, B(13) => OTMP_269_port, B(12) => 
                           OTMP_268_port, B(11) => OTMP_267_port, B(10) => 
                           OTMP_266_port, B(9) => OTMP_265_port, B(8) => 
                           OTMP_264_port, B(7) => OTMP_263_port, B(6) => 
                           OTMP_262_port, B(5) => OTMP_261_port, B(4) => 
                           OTMP_260_port, B(3) => OTMP_259_port, B(2) => 
                           OTMP_258_port, B(1) => OTMP_257_port, B(0) => 
                           OTMP_256_port, Ci => X_Logic0_port, S(63) => 
                           PTMP_255_port, S(62) => PTMP_254_port, S(61) => 
                           PTMP_253_port, S(60) => PTMP_252_port, S(59) => 
                           PTMP_251_port, S(58) => PTMP_250_port, S(57) => 
                           PTMP_249_port, S(56) => PTMP_248_port, S(55) => 
                           PTMP_247_port, S(54) => PTMP_246_port, S(53) => 
                           PTMP_245_port, S(52) => PTMP_244_port, S(51) => 
                           PTMP_243_port, S(50) => PTMP_242_port, S(49) => 
                           PTMP_241_port, S(48) => PTMP_240_port, S(47) => 
                           PTMP_239_port, S(46) => PTMP_238_port, S(45) => 
                           PTMP_237_port, S(44) => PTMP_236_port, S(43) => 
                           PTMP_235_port, S(42) => PTMP_234_port, S(41) => 
                           PTMP_233_port, S(40) => PTMP_232_port, S(39) => 
                           PTMP_231_port, S(38) => PTMP_230_port, S(37) => 
                           PTMP_229_port, S(36) => PTMP_228_port, S(35) => 
                           PTMP_227_port, S(34) => PTMP_226_port, S(33) => 
                           PTMP_225_port, S(32) => PTMP_224_port, S(31) => 
                           PTMP_223_port, S(30) => PTMP_222_port, S(29) => 
                           PTMP_221_port, S(28) => PTMP_220_port, S(27) => 
                           PTMP_219_port, S(26) => PTMP_218_port, S(25) => 
                           PTMP_217_port, S(24) => PTMP_216_port, S(23) => 
                           PTMP_215_port, S(22) => PTMP_214_port, S(21) => 
                           PTMP_213_port, S(20) => PTMP_212_port, S(19) => 
                           PTMP_211_port, S(18) => PTMP_210_port, S(17) => 
                           PTMP_209_port, S(16) => PTMP_208_port, S(15) => 
                           PTMP_207_port, S(14) => PTMP_206_port, S(13) => 
                           PTMP_205_port, S(12) => PTMP_204_port, S(11) => 
                           PTMP_203_port, S(10) => PTMP_202_port, S(9) => 
                           PTMP_201_port, S(8) => PTMP_200_port, S(7) => 
                           PTMP_199_port, S(6) => PTMP_198_port, S(5) => 
                           PTMP_197_port, S(4) => PTMP_196_port, S(3) => 
                           PTMP_195_port, S(2) => PTMP_194_port, S(1) => 
                           PTMP_193_port, S(0) => PTMP_192_port, Co => n_1298);
   ADDERI_6 : RCA_NBIT64_26 port map( A(63) => PTMP_255_port, A(62) => 
                           PTMP_254_port, A(61) => PTMP_253_port, A(60) => 
                           PTMP_252_port, A(59) => PTMP_251_port, A(58) => 
                           PTMP_250_port, A(57) => PTMP_249_port, A(56) => 
                           PTMP_248_port, A(55) => PTMP_247_port, A(54) => 
                           PTMP_246_port, A(53) => PTMP_245_port, A(52) => 
                           PTMP_244_port, A(51) => PTMP_243_port, A(50) => 
                           PTMP_242_port, A(49) => PTMP_241_port, A(48) => 
                           PTMP_240_port, A(47) => PTMP_239_port, A(46) => 
                           PTMP_238_port, A(45) => PTMP_237_port, A(44) => 
                           PTMP_236_port, A(43) => PTMP_235_port, A(42) => 
                           PTMP_234_port, A(41) => PTMP_233_port, A(40) => 
                           PTMP_232_port, A(39) => PTMP_231_port, A(38) => 
                           PTMP_230_port, A(37) => PTMP_229_port, A(36) => 
                           PTMP_228_port, A(35) => PTMP_227_port, A(34) => 
                           PTMP_226_port, A(33) => PTMP_225_port, A(32) => 
                           PTMP_224_port, A(31) => PTMP_223_port, A(30) => 
                           PTMP_222_port, A(29) => PTMP_221_port, A(28) => 
                           PTMP_220_port, A(27) => PTMP_219_port, A(26) => 
                           PTMP_218_port, A(25) => PTMP_217_port, A(24) => 
                           PTMP_216_port, A(23) => PTMP_215_port, A(22) => 
                           PTMP_214_port, A(21) => PTMP_213_port, A(20) => 
                           PTMP_212_port, A(19) => PTMP_211_port, A(18) => 
                           PTMP_210_port, A(17) => PTMP_209_port, A(16) => 
                           PTMP_208_port, A(15) => PTMP_207_port, A(14) => 
                           PTMP_206_port, A(13) => PTMP_205_port, A(12) => 
                           PTMP_204_port, A(11) => PTMP_203_port, A(10) => 
                           PTMP_202_port, A(9) => PTMP_201_port, A(8) => 
                           PTMP_200_port, A(7) => PTMP_199_port, A(6) => 
                           PTMP_198_port, A(5) => PTMP_197_port, A(4) => 
                           PTMP_196_port, A(3) => PTMP_195_port, A(2) => 
                           PTMP_194_port, A(1) => PTMP_193_port, A(0) => 
                           PTMP_192_port, B(63) => OTMP_383_port, B(62) => 
                           OTMP_382_port, B(61) => OTMP_381_port, B(60) => 
                           OTMP_380_port, B(59) => OTMP_379_port, B(58) => 
                           OTMP_378_port, B(57) => OTMP_377_port, B(56) => 
                           OTMP_376_port, B(55) => OTMP_375_port, B(54) => 
                           OTMP_374_port, B(53) => OTMP_373_port, B(52) => 
                           OTMP_372_port, B(51) => OTMP_371_port, B(50) => 
                           OTMP_370_port, B(49) => OTMP_369_port, B(48) => 
                           OTMP_368_port, B(47) => OTMP_367_port, B(46) => 
                           OTMP_366_port, B(45) => OTMP_365_port, B(44) => 
                           OTMP_364_port, B(43) => OTMP_363_port, B(42) => 
                           OTMP_362_port, B(41) => OTMP_361_port, B(40) => 
                           OTMP_360_port, B(39) => OTMP_359_port, B(38) => 
                           OTMP_358_port, B(37) => OTMP_357_port, B(36) => 
                           OTMP_356_port, B(35) => OTMP_355_port, B(34) => 
                           OTMP_354_port, B(33) => OTMP_353_port, B(32) => 
                           OTMP_352_port, B(31) => OTMP_351_port, B(30) => 
                           OTMP_350_port, B(29) => OTMP_349_port, B(28) => 
                           OTMP_348_port, B(27) => OTMP_347_port, B(26) => 
                           OTMP_346_port, B(25) => OTMP_345_port, B(24) => 
                           OTMP_344_port, B(23) => OTMP_343_port, B(22) => 
                           OTMP_342_port, B(21) => OTMP_341_port, B(20) => 
                           OTMP_340_port, B(19) => OTMP_339_port, B(18) => 
                           OTMP_338_port, B(17) => OTMP_337_port, B(16) => 
                           OTMP_336_port, B(15) => OTMP_335_port, B(14) => 
                           OTMP_334_port, B(13) => OTMP_333_port, B(12) => 
                           OTMP_332_port, B(11) => OTMP_331_port, B(10) => 
                           OTMP_330_port, B(9) => OTMP_329_port, B(8) => 
                           OTMP_328_port, B(7) => OTMP_327_port, B(6) => 
                           OTMP_326_port, B(5) => OTMP_325_port, B(4) => 
                           OTMP_324_port, B(3) => OTMP_323_port, B(2) => 
                           OTMP_322_port, B(1) => OTMP_321_port, B(0) => 
                           OTMP_320_port, Ci => X_Logic0_port, S(63) => 
                           PTMP_319_port, S(62) => PTMP_318_port, S(61) => 
                           PTMP_317_port, S(60) => PTMP_316_port, S(59) => 
                           PTMP_315_port, S(58) => PTMP_314_port, S(57) => 
                           PTMP_313_port, S(56) => PTMP_312_port, S(55) => 
                           PTMP_311_port, S(54) => PTMP_310_port, S(53) => 
                           PTMP_309_port, S(52) => PTMP_308_port, S(51) => 
                           PTMP_307_port, S(50) => PTMP_306_port, S(49) => 
                           PTMP_305_port, S(48) => PTMP_304_port, S(47) => 
                           PTMP_303_port, S(46) => PTMP_302_port, S(45) => 
                           PTMP_301_port, S(44) => PTMP_300_port, S(43) => 
                           PTMP_299_port, S(42) => PTMP_298_port, S(41) => 
                           PTMP_297_port, S(40) => PTMP_296_port, S(39) => 
                           PTMP_295_port, S(38) => PTMP_294_port, S(37) => 
                           PTMP_293_port, S(36) => PTMP_292_port, S(35) => 
                           PTMP_291_port, S(34) => PTMP_290_port, S(33) => 
                           PTMP_289_port, S(32) => PTMP_288_port, S(31) => 
                           PTMP_287_port, S(30) => PTMP_286_port, S(29) => 
                           PTMP_285_port, S(28) => PTMP_284_port, S(27) => 
                           PTMP_283_port, S(26) => PTMP_282_port, S(25) => 
                           PTMP_281_port, S(24) => PTMP_280_port, S(23) => 
                           PTMP_279_port, S(22) => PTMP_278_port, S(21) => 
                           PTMP_277_port, S(20) => PTMP_276_port, S(19) => 
                           PTMP_275_port, S(18) => PTMP_274_port, S(17) => 
                           PTMP_273_port, S(16) => PTMP_272_port, S(15) => 
                           PTMP_271_port, S(14) => PTMP_270_port, S(13) => 
                           PTMP_269_port, S(12) => PTMP_268_port, S(11) => 
                           PTMP_267_port, S(10) => PTMP_266_port, S(9) => 
                           PTMP_265_port, S(8) => PTMP_264_port, S(7) => 
                           PTMP_263_port, S(6) => PTMP_262_port, S(5) => 
                           PTMP_261_port, S(4) => PTMP_260_port, S(3) => 
                           PTMP_259_port, S(2) => PTMP_258_port, S(1) => 
                           PTMP_257_port, S(0) => PTMP_256_port, Co => n_1299);
   ADDERI_7 : RCA_NBIT64_25 port map( A(63) => PTMP_319_port, A(62) => 
                           PTMP_318_port, A(61) => PTMP_317_port, A(60) => 
                           PTMP_316_port, A(59) => PTMP_315_port, A(58) => 
                           PTMP_314_port, A(57) => PTMP_313_port, A(56) => 
                           PTMP_312_port, A(55) => PTMP_311_port, A(54) => 
                           PTMP_310_port, A(53) => PTMP_309_port, A(52) => 
                           PTMP_308_port, A(51) => PTMP_307_port, A(50) => 
                           PTMP_306_port, A(49) => PTMP_305_port, A(48) => 
                           PTMP_304_port, A(47) => PTMP_303_port, A(46) => 
                           PTMP_302_port, A(45) => PTMP_301_port, A(44) => 
                           PTMP_300_port, A(43) => PTMP_299_port, A(42) => 
                           PTMP_298_port, A(41) => PTMP_297_port, A(40) => 
                           PTMP_296_port, A(39) => PTMP_295_port, A(38) => 
                           PTMP_294_port, A(37) => PTMP_293_port, A(36) => 
                           PTMP_292_port, A(35) => PTMP_291_port, A(34) => 
                           PTMP_290_port, A(33) => PTMP_289_port, A(32) => 
                           PTMP_288_port, A(31) => PTMP_287_port, A(30) => 
                           PTMP_286_port, A(29) => PTMP_285_port, A(28) => 
                           PTMP_284_port, A(27) => PTMP_283_port, A(26) => 
                           PTMP_282_port, A(25) => PTMP_281_port, A(24) => 
                           PTMP_280_port, A(23) => PTMP_279_port, A(22) => 
                           PTMP_278_port, A(21) => PTMP_277_port, A(20) => 
                           PTMP_276_port, A(19) => PTMP_275_port, A(18) => 
                           PTMP_274_port, A(17) => PTMP_273_port, A(16) => 
                           PTMP_272_port, A(15) => PTMP_271_port, A(14) => 
                           PTMP_270_port, A(13) => PTMP_269_port, A(12) => 
                           PTMP_268_port, A(11) => PTMP_267_port, A(10) => 
                           PTMP_266_port, A(9) => PTMP_265_port, A(8) => 
                           PTMP_264_port, A(7) => PTMP_263_port, A(6) => 
                           PTMP_262_port, A(5) => PTMP_261_port, A(4) => 
                           PTMP_260_port, A(3) => PTMP_259_port, A(2) => 
                           PTMP_258_port, A(1) => PTMP_257_port, A(0) => 
                           PTMP_256_port, B(63) => OTMP_447_port, B(62) => 
                           OTMP_446_port, B(61) => OTMP_445_port, B(60) => 
                           OTMP_444_port, B(59) => OTMP_443_port, B(58) => 
                           OTMP_442_port, B(57) => OTMP_441_port, B(56) => 
                           OTMP_440_port, B(55) => OTMP_439_port, B(54) => 
                           OTMP_438_port, B(53) => OTMP_437_port, B(52) => 
                           OTMP_436_port, B(51) => OTMP_435_port, B(50) => 
                           OTMP_434_port, B(49) => OTMP_433_port, B(48) => 
                           OTMP_432_port, B(47) => OTMP_431_port, B(46) => 
                           OTMP_430_port, B(45) => OTMP_429_port, B(44) => 
                           OTMP_428_port, B(43) => OTMP_427_port, B(42) => 
                           OTMP_426_port, B(41) => OTMP_425_port, B(40) => 
                           OTMP_424_port, B(39) => OTMP_423_port, B(38) => 
                           OTMP_422_port, B(37) => OTMP_421_port, B(36) => 
                           OTMP_420_port, B(35) => OTMP_419_port, B(34) => 
                           OTMP_418_port, B(33) => OTMP_417_port, B(32) => 
                           OTMP_416_port, B(31) => OTMP_415_port, B(30) => 
                           OTMP_414_port, B(29) => OTMP_413_port, B(28) => 
                           OTMP_412_port, B(27) => OTMP_411_port, B(26) => 
                           OTMP_410_port, B(25) => OTMP_409_port, B(24) => 
                           OTMP_408_port, B(23) => OTMP_407_port, B(22) => 
                           OTMP_406_port, B(21) => OTMP_405_port, B(20) => 
                           OTMP_404_port, B(19) => OTMP_403_port, B(18) => 
                           OTMP_402_port, B(17) => OTMP_401_port, B(16) => 
                           OTMP_400_port, B(15) => OTMP_399_port, B(14) => 
                           OTMP_398_port, B(13) => OTMP_397_port, B(12) => 
                           OTMP_396_port, B(11) => OTMP_395_port, B(10) => 
                           OTMP_394_port, B(9) => OTMP_393_port, B(8) => 
                           OTMP_392_port, B(7) => OTMP_391_port, B(6) => 
                           OTMP_390_port, B(5) => OTMP_389_port, B(4) => 
                           OTMP_388_port, B(3) => OTMP_387_port, B(2) => 
                           OTMP_386_port, B(1) => OTMP_385_port, B(0) => 
                           OTMP_384_port, Ci => X_Logic0_port, S(63) => 
                           PTMP_383_port, S(62) => PTMP_382_port, S(61) => 
                           PTMP_381_port, S(60) => PTMP_380_port, S(59) => 
                           PTMP_379_port, S(58) => PTMP_378_port, S(57) => 
                           PTMP_377_port, S(56) => PTMP_376_port, S(55) => 
                           PTMP_375_port, S(54) => PTMP_374_port, S(53) => 
                           PTMP_373_port, S(52) => PTMP_372_port, S(51) => 
                           PTMP_371_port, S(50) => PTMP_370_port, S(49) => 
                           PTMP_369_port, S(48) => PTMP_368_port, S(47) => 
                           PTMP_367_port, S(46) => PTMP_366_port, S(45) => 
                           PTMP_365_port, S(44) => PTMP_364_port, S(43) => 
                           PTMP_363_port, S(42) => PTMP_362_port, S(41) => 
                           PTMP_361_port, S(40) => PTMP_360_port, S(39) => 
                           PTMP_359_port, S(38) => PTMP_358_port, S(37) => 
                           PTMP_357_port, S(36) => PTMP_356_port, S(35) => 
                           PTMP_355_port, S(34) => PTMP_354_port, S(33) => 
                           PTMP_353_port, S(32) => PTMP_352_port, S(31) => 
                           PTMP_351_port, S(30) => PTMP_350_port, S(29) => 
                           PTMP_349_port, S(28) => PTMP_348_port, S(27) => 
                           PTMP_347_port, S(26) => PTMP_346_port, S(25) => 
                           PTMP_345_port, S(24) => PTMP_344_port, S(23) => 
                           PTMP_343_port, S(22) => PTMP_342_port, S(21) => 
                           PTMP_341_port, S(20) => PTMP_340_port, S(19) => 
                           PTMP_339_port, S(18) => PTMP_338_port, S(17) => 
                           PTMP_337_port, S(16) => PTMP_336_port, S(15) => 
                           PTMP_335_port, S(14) => PTMP_334_port, S(13) => 
                           PTMP_333_port, S(12) => PTMP_332_port, S(11) => 
                           PTMP_331_port, S(10) => PTMP_330_port, S(9) => 
                           PTMP_329_port, S(8) => PTMP_328_port, S(7) => 
                           PTMP_327_port, S(6) => PTMP_326_port, S(5) => 
                           PTMP_325_port, S(4) => PTMP_324_port, S(3) => 
                           PTMP_323_port, S(2) => PTMP_322_port, S(1) => 
                           PTMP_321_port, S(0) => PTMP_320_port, Co => n_1300);
   ADDERI_8 : RCA_NBIT64_24 port map( A(63) => PTMP_383_port, A(62) => 
                           PTMP_382_port, A(61) => PTMP_381_port, A(60) => 
                           PTMP_380_port, A(59) => PTMP_379_port, A(58) => 
                           PTMP_378_port, A(57) => PTMP_377_port, A(56) => 
                           PTMP_376_port, A(55) => PTMP_375_port, A(54) => 
                           PTMP_374_port, A(53) => PTMP_373_port, A(52) => 
                           PTMP_372_port, A(51) => PTMP_371_port, A(50) => 
                           PTMP_370_port, A(49) => PTMP_369_port, A(48) => 
                           PTMP_368_port, A(47) => PTMP_367_port, A(46) => 
                           PTMP_366_port, A(45) => PTMP_365_port, A(44) => 
                           PTMP_364_port, A(43) => PTMP_363_port, A(42) => 
                           PTMP_362_port, A(41) => PTMP_361_port, A(40) => 
                           PTMP_360_port, A(39) => PTMP_359_port, A(38) => 
                           PTMP_358_port, A(37) => PTMP_357_port, A(36) => 
                           PTMP_356_port, A(35) => PTMP_355_port, A(34) => 
                           PTMP_354_port, A(33) => PTMP_353_port, A(32) => 
                           PTMP_352_port, A(31) => PTMP_351_port, A(30) => 
                           PTMP_350_port, A(29) => PTMP_349_port, A(28) => 
                           PTMP_348_port, A(27) => PTMP_347_port, A(26) => 
                           PTMP_346_port, A(25) => PTMP_345_port, A(24) => 
                           PTMP_344_port, A(23) => PTMP_343_port, A(22) => 
                           PTMP_342_port, A(21) => PTMP_341_port, A(20) => 
                           PTMP_340_port, A(19) => PTMP_339_port, A(18) => 
                           PTMP_338_port, A(17) => PTMP_337_port, A(16) => 
                           PTMP_336_port, A(15) => PTMP_335_port, A(14) => 
                           PTMP_334_port, A(13) => PTMP_333_port, A(12) => 
                           PTMP_332_port, A(11) => PTMP_331_port, A(10) => 
                           PTMP_330_port, A(9) => PTMP_329_port, A(8) => 
                           PTMP_328_port, A(7) => PTMP_327_port, A(6) => 
                           PTMP_326_port, A(5) => PTMP_325_port, A(4) => 
                           PTMP_324_port, A(3) => PTMP_323_port, A(2) => 
                           PTMP_322_port, A(1) => PTMP_321_port, A(0) => 
                           PTMP_320_port, B(63) => OTMP_511_port, B(62) => 
                           OTMP_510_port, B(61) => OTMP_509_port, B(60) => 
                           OTMP_508_port, B(59) => OTMP_507_port, B(58) => 
                           OTMP_506_port, B(57) => OTMP_505_port, B(56) => 
                           OTMP_504_port, B(55) => OTMP_503_port, B(54) => 
                           OTMP_502_port, B(53) => OTMP_501_port, B(52) => 
                           OTMP_500_port, B(51) => OTMP_499_port, B(50) => 
                           OTMP_498_port, B(49) => OTMP_497_port, B(48) => 
                           OTMP_496_port, B(47) => OTMP_495_port, B(46) => 
                           OTMP_494_port, B(45) => OTMP_493_port, B(44) => 
                           OTMP_492_port, B(43) => OTMP_491_port, B(42) => 
                           OTMP_490_port, B(41) => OTMP_489_port, B(40) => 
                           OTMP_488_port, B(39) => OTMP_487_port, B(38) => 
                           OTMP_486_port, B(37) => OTMP_485_port, B(36) => 
                           OTMP_484_port, B(35) => OTMP_483_port, B(34) => 
                           OTMP_482_port, B(33) => OTMP_481_port, B(32) => 
                           OTMP_480_port, B(31) => OTMP_479_port, B(30) => 
                           OTMP_478_port, B(29) => OTMP_477_port, B(28) => 
                           OTMP_476_port, B(27) => OTMP_475_port, B(26) => 
                           OTMP_474_port, B(25) => OTMP_473_port, B(24) => 
                           OTMP_472_port, B(23) => OTMP_471_port, B(22) => 
                           OTMP_470_port, B(21) => OTMP_469_port, B(20) => 
                           OTMP_468_port, B(19) => OTMP_467_port, B(18) => 
                           OTMP_466_port, B(17) => OTMP_465_port, B(16) => 
                           OTMP_464_port, B(15) => OTMP_463_port, B(14) => 
                           OTMP_462_port, B(13) => OTMP_461_port, B(12) => 
                           OTMP_460_port, B(11) => OTMP_459_port, B(10) => 
                           OTMP_458_port, B(9) => OTMP_457_port, B(8) => 
                           OTMP_456_port, B(7) => OTMP_455_port, B(6) => 
                           OTMP_454_port, B(5) => OTMP_453_port, B(4) => 
                           OTMP_452_port, B(3) => OTMP_451_port, B(2) => 
                           OTMP_450_port, B(1) => OTMP_449_port, B(0) => 
                           OTMP_448_port, Ci => X_Logic0_port, S(63) => 
                           PTMP_447_port, S(62) => PTMP_446_port, S(61) => 
                           PTMP_445_port, S(60) => PTMP_444_port, S(59) => 
                           PTMP_443_port, S(58) => PTMP_442_port, S(57) => 
                           PTMP_441_port, S(56) => PTMP_440_port, S(55) => 
                           PTMP_439_port, S(54) => PTMP_438_port, S(53) => 
                           PTMP_437_port, S(52) => PTMP_436_port, S(51) => 
                           PTMP_435_port, S(50) => PTMP_434_port, S(49) => 
                           PTMP_433_port, S(48) => PTMP_432_port, S(47) => 
                           PTMP_431_port, S(46) => PTMP_430_port, S(45) => 
                           PTMP_429_port, S(44) => PTMP_428_port, S(43) => 
                           PTMP_427_port, S(42) => PTMP_426_port, S(41) => 
                           PTMP_425_port, S(40) => PTMP_424_port, S(39) => 
                           PTMP_423_port, S(38) => PTMP_422_port, S(37) => 
                           PTMP_421_port, S(36) => PTMP_420_port, S(35) => 
                           PTMP_419_port, S(34) => PTMP_418_port, S(33) => 
                           PTMP_417_port, S(32) => PTMP_416_port, S(31) => 
                           PTMP_415_port, S(30) => PTMP_414_port, S(29) => 
                           PTMP_413_port, S(28) => PTMP_412_port, S(27) => 
                           PTMP_411_port, S(26) => PTMP_410_port, S(25) => 
                           PTMP_409_port, S(24) => PTMP_408_port, S(23) => 
                           PTMP_407_port, S(22) => PTMP_406_port, S(21) => 
                           PTMP_405_port, S(20) => PTMP_404_port, S(19) => 
                           PTMP_403_port, S(18) => PTMP_402_port, S(17) => 
                           PTMP_401_port, S(16) => PTMP_400_port, S(15) => 
                           PTMP_399_port, S(14) => PTMP_398_port, S(13) => 
                           PTMP_397_port, S(12) => PTMP_396_port, S(11) => 
                           PTMP_395_port, S(10) => PTMP_394_port, S(9) => 
                           PTMP_393_port, S(8) => PTMP_392_port, S(7) => 
                           PTMP_391_port, S(6) => PTMP_390_port, S(5) => 
                           PTMP_389_port, S(4) => PTMP_388_port, S(3) => 
                           PTMP_387_port, S(2) => PTMP_386_port, S(1) => 
                           PTMP_385_port, S(0) => PTMP_384_port, Co => n_1301);
   ADDERI_9 : RCA_NBIT64_23 port map( A(63) => PTMP_447_port, A(62) => 
                           PTMP_446_port, A(61) => PTMP_445_port, A(60) => 
                           PTMP_444_port, A(59) => PTMP_443_port, A(58) => 
                           PTMP_442_port, A(57) => PTMP_441_port, A(56) => 
                           PTMP_440_port, A(55) => PTMP_439_port, A(54) => 
                           PTMP_438_port, A(53) => PTMP_437_port, A(52) => 
                           PTMP_436_port, A(51) => PTMP_435_port, A(50) => 
                           PTMP_434_port, A(49) => PTMP_433_port, A(48) => 
                           PTMP_432_port, A(47) => PTMP_431_port, A(46) => 
                           PTMP_430_port, A(45) => PTMP_429_port, A(44) => 
                           PTMP_428_port, A(43) => PTMP_427_port, A(42) => 
                           PTMP_426_port, A(41) => PTMP_425_port, A(40) => 
                           PTMP_424_port, A(39) => PTMP_423_port, A(38) => 
                           PTMP_422_port, A(37) => PTMP_421_port, A(36) => 
                           PTMP_420_port, A(35) => PTMP_419_port, A(34) => 
                           PTMP_418_port, A(33) => PTMP_417_port, A(32) => 
                           PTMP_416_port, A(31) => PTMP_415_port, A(30) => 
                           PTMP_414_port, A(29) => PTMP_413_port, A(28) => 
                           PTMP_412_port, A(27) => PTMP_411_port, A(26) => 
                           PTMP_410_port, A(25) => PTMP_409_port, A(24) => 
                           PTMP_408_port, A(23) => PTMP_407_port, A(22) => 
                           PTMP_406_port, A(21) => PTMP_405_port, A(20) => 
                           PTMP_404_port, A(19) => PTMP_403_port, A(18) => 
                           PTMP_402_port, A(17) => PTMP_401_port, A(16) => 
                           PTMP_400_port, A(15) => PTMP_399_port, A(14) => 
                           PTMP_398_port, A(13) => PTMP_397_port, A(12) => 
                           PTMP_396_port, A(11) => PTMP_395_port, A(10) => 
                           PTMP_394_port, A(9) => PTMP_393_port, A(8) => 
                           PTMP_392_port, A(7) => PTMP_391_port, A(6) => 
                           PTMP_390_port, A(5) => PTMP_389_port, A(4) => 
                           PTMP_388_port, A(3) => PTMP_387_port, A(2) => 
                           PTMP_386_port, A(1) => PTMP_385_port, A(0) => 
                           PTMP_384_port, B(63) => OTMP_575_port, B(62) => 
                           OTMP_574_port, B(61) => OTMP_573_port, B(60) => 
                           OTMP_572_port, B(59) => OTMP_571_port, B(58) => 
                           OTMP_570_port, B(57) => OTMP_569_port, B(56) => 
                           OTMP_568_port, B(55) => OTMP_567_port, B(54) => 
                           OTMP_566_port, B(53) => OTMP_565_port, B(52) => 
                           OTMP_564_port, B(51) => OTMP_563_port, B(50) => 
                           OTMP_562_port, B(49) => OTMP_561_port, B(48) => 
                           OTMP_560_port, B(47) => OTMP_559_port, B(46) => 
                           OTMP_558_port, B(45) => OTMP_557_port, B(44) => 
                           OTMP_556_port, B(43) => OTMP_555_port, B(42) => 
                           OTMP_554_port, B(41) => OTMP_553_port, B(40) => 
                           OTMP_552_port, B(39) => OTMP_551_port, B(38) => 
                           OTMP_550_port, B(37) => OTMP_549_port, B(36) => 
                           OTMP_548_port, B(35) => OTMP_547_port, B(34) => 
                           OTMP_546_port, B(33) => OTMP_545_port, B(32) => 
                           OTMP_544_port, B(31) => OTMP_543_port, B(30) => 
                           OTMP_542_port, B(29) => OTMP_541_port, B(28) => 
                           OTMP_540_port, B(27) => OTMP_539_port, B(26) => 
                           OTMP_538_port, B(25) => OTMP_537_port, B(24) => 
                           OTMP_536_port, B(23) => OTMP_535_port, B(22) => 
                           OTMP_534_port, B(21) => OTMP_533_port, B(20) => 
                           OTMP_532_port, B(19) => OTMP_531_port, B(18) => 
                           OTMP_530_port, B(17) => OTMP_529_port, B(16) => 
                           OTMP_528_port, B(15) => OTMP_527_port, B(14) => 
                           OTMP_526_port, B(13) => OTMP_525_port, B(12) => 
                           OTMP_524_port, B(11) => OTMP_523_port, B(10) => 
                           OTMP_522_port, B(9) => OTMP_521_port, B(8) => 
                           OTMP_520_port, B(7) => OTMP_519_port, B(6) => 
                           OTMP_518_port, B(5) => OTMP_517_port, B(4) => 
                           OTMP_516_port, B(3) => OTMP_515_port, B(2) => 
                           OTMP_514_port, B(1) => OTMP_513_port, B(0) => 
                           OTMP_512_port, Ci => X_Logic0_port, S(63) => 
                           PTMP_511_port, S(62) => PTMP_510_port, S(61) => 
                           PTMP_509_port, S(60) => PTMP_508_port, S(59) => 
                           PTMP_507_port, S(58) => PTMP_506_port, S(57) => 
                           PTMP_505_port, S(56) => PTMP_504_port, S(55) => 
                           PTMP_503_port, S(54) => PTMP_502_port, S(53) => 
                           PTMP_501_port, S(52) => PTMP_500_port, S(51) => 
                           PTMP_499_port, S(50) => PTMP_498_port, S(49) => 
                           PTMP_497_port, S(48) => PTMP_496_port, S(47) => 
                           PTMP_495_port, S(46) => PTMP_494_port, S(45) => 
                           PTMP_493_port, S(44) => PTMP_492_port, S(43) => 
                           PTMP_491_port, S(42) => PTMP_490_port, S(41) => 
                           PTMP_489_port, S(40) => PTMP_488_port, S(39) => 
                           PTMP_487_port, S(38) => PTMP_486_port, S(37) => 
                           PTMP_485_port, S(36) => PTMP_484_port, S(35) => 
                           PTMP_483_port, S(34) => PTMP_482_port, S(33) => 
                           PTMP_481_port, S(32) => PTMP_480_port, S(31) => 
                           PTMP_479_port, S(30) => PTMP_478_port, S(29) => 
                           PTMP_477_port, S(28) => PTMP_476_port, S(27) => 
                           PTMP_475_port, S(26) => PTMP_474_port, S(25) => 
                           PTMP_473_port, S(24) => PTMP_472_port, S(23) => 
                           PTMP_471_port, S(22) => PTMP_470_port, S(21) => 
                           PTMP_469_port, S(20) => PTMP_468_port, S(19) => 
                           PTMP_467_port, S(18) => PTMP_466_port, S(17) => 
                           PTMP_465_port, S(16) => PTMP_464_port, S(15) => 
                           PTMP_463_port, S(14) => PTMP_462_port, S(13) => 
                           PTMP_461_port, S(12) => PTMP_460_port, S(11) => 
                           PTMP_459_port, S(10) => PTMP_458_port, S(9) => 
                           PTMP_457_port, S(8) => PTMP_456_port, S(7) => 
                           PTMP_455_port, S(6) => PTMP_454_port, S(5) => 
                           PTMP_453_port, S(4) => PTMP_452_port, S(3) => 
                           PTMP_451_port, S(2) => PTMP_450_port, S(1) => 
                           PTMP_449_port, S(0) => PTMP_448_port, Co => n_1302);
   ADDERI_10 : RCA_NBIT64_22 port map( A(63) => PTMP_511_port, A(62) => 
                           PTMP_510_port, A(61) => PTMP_509_port, A(60) => 
                           PTMP_508_port, A(59) => PTMP_507_port, A(58) => 
                           PTMP_506_port, A(57) => PTMP_505_port, A(56) => 
                           PTMP_504_port, A(55) => PTMP_503_port, A(54) => 
                           PTMP_502_port, A(53) => PTMP_501_port, A(52) => 
                           PTMP_500_port, A(51) => PTMP_499_port, A(50) => 
                           PTMP_498_port, A(49) => PTMP_497_port, A(48) => 
                           PTMP_496_port, A(47) => PTMP_495_port, A(46) => 
                           PTMP_494_port, A(45) => PTMP_493_port, A(44) => 
                           PTMP_492_port, A(43) => PTMP_491_port, A(42) => 
                           PTMP_490_port, A(41) => PTMP_489_port, A(40) => 
                           PTMP_488_port, A(39) => PTMP_487_port, A(38) => 
                           PTMP_486_port, A(37) => PTMP_485_port, A(36) => 
                           PTMP_484_port, A(35) => PTMP_483_port, A(34) => 
                           PTMP_482_port, A(33) => PTMP_481_port, A(32) => 
                           PTMP_480_port, A(31) => PTMP_479_port, A(30) => 
                           PTMP_478_port, A(29) => PTMP_477_port, A(28) => 
                           PTMP_476_port, A(27) => PTMP_475_port, A(26) => 
                           PTMP_474_port, A(25) => PTMP_473_port, A(24) => 
                           PTMP_472_port, A(23) => PTMP_471_port, A(22) => 
                           PTMP_470_port, A(21) => PTMP_469_port, A(20) => 
                           PTMP_468_port, A(19) => PTMP_467_port, A(18) => 
                           PTMP_466_port, A(17) => PTMP_465_port, A(16) => 
                           PTMP_464_port, A(15) => PTMP_463_port, A(14) => 
                           PTMP_462_port, A(13) => PTMP_461_port, A(12) => 
                           PTMP_460_port, A(11) => PTMP_459_port, A(10) => 
                           PTMP_458_port, A(9) => PTMP_457_port, A(8) => 
                           PTMP_456_port, A(7) => PTMP_455_port, A(6) => 
                           PTMP_454_port, A(5) => PTMP_453_port, A(4) => 
                           PTMP_452_port, A(3) => PTMP_451_port, A(2) => 
                           PTMP_450_port, A(1) => PTMP_449_port, A(0) => 
                           PTMP_448_port, B(63) => OTMP_639_port, B(62) => 
                           OTMP_638_port, B(61) => OTMP_637_port, B(60) => 
                           OTMP_636_port, B(59) => OTMP_635_port, B(58) => 
                           OTMP_634_port, B(57) => OTMP_633_port, B(56) => 
                           OTMP_632_port, B(55) => OTMP_631_port, B(54) => 
                           OTMP_630_port, B(53) => OTMP_629_port, B(52) => 
                           OTMP_628_port, B(51) => OTMP_627_port, B(50) => 
                           OTMP_626_port, B(49) => OTMP_625_port, B(48) => 
                           OTMP_624_port, B(47) => OTMP_623_port, B(46) => 
                           OTMP_622_port, B(45) => OTMP_621_port, B(44) => 
                           OTMP_620_port, B(43) => OTMP_619_port, B(42) => 
                           OTMP_618_port, B(41) => OTMP_617_port, B(40) => 
                           OTMP_616_port, B(39) => OTMP_615_port, B(38) => 
                           OTMP_614_port, B(37) => OTMP_613_port, B(36) => 
                           OTMP_612_port, B(35) => OTMP_611_port, B(34) => 
                           OTMP_610_port, B(33) => OTMP_609_port, B(32) => 
                           OTMP_608_port, B(31) => OTMP_607_port, B(30) => 
                           OTMP_606_port, B(29) => OTMP_605_port, B(28) => 
                           OTMP_604_port, B(27) => OTMP_603_port, B(26) => 
                           OTMP_602_port, B(25) => OTMP_601_port, B(24) => 
                           OTMP_600_port, B(23) => OTMP_599_port, B(22) => 
                           OTMP_598_port, B(21) => OTMP_597_port, B(20) => 
                           OTMP_596_port, B(19) => OTMP_595_port, B(18) => 
                           OTMP_594_port, B(17) => OTMP_593_port, B(16) => 
                           OTMP_592_port, B(15) => OTMP_591_port, B(14) => 
                           OTMP_590_port, B(13) => OTMP_589_port, B(12) => 
                           OTMP_588_port, B(11) => OTMP_587_port, B(10) => 
                           OTMP_586_port, B(9) => OTMP_585_port, B(8) => 
                           OTMP_584_port, B(7) => OTMP_583_port, B(6) => 
                           OTMP_582_port, B(5) => OTMP_581_port, B(4) => 
                           OTMP_580_port, B(3) => OTMP_579_port, B(2) => 
                           OTMP_578_port, B(1) => OTMP_577_port, B(0) => 
                           OTMP_576_port, Ci => X_Logic0_port, S(63) => 
                           PTMP_575_port, S(62) => PTMP_574_port, S(61) => 
                           PTMP_573_port, S(60) => PTMP_572_port, S(59) => 
                           PTMP_571_port, S(58) => PTMP_570_port, S(57) => 
                           PTMP_569_port, S(56) => PTMP_568_port, S(55) => 
                           PTMP_567_port, S(54) => PTMP_566_port, S(53) => 
                           PTMP_565_port, S(52) => PTMP_564_port, S(51) => 
                           PTMP_563_port, S(50) => PTMP_562_port, S(49) => 
                           PTMP_561_port, S(48) => PTMP_560_port, S(47) => 
                           PTMP_559_port, S(46) => PTMP_558_port, S(45) => 
                           PTMP_557_port, S(44) => PTMP_556_port, S(43) => 
                           PTMP_555_port, S(42) => PTMP_554_port, S(41) => 
                           PTMP_553_port, S(40) => PTMP_552_port, S(39) => 
                           PTMP_551_port, S(38) => PTMP_550_port, S(37) => 
                           PTMP_549_port, S(36) => PTMP_548_port, S(35) => 
                           PTMP_547_port, S(34) => PTMP_546_port, S(33) => 
                           PTMP_545_port, S(32) => PTMP_544_port, S(31) => 
                           PTMP_543_port, S(30) => PTMP_542_port, S(29) => 
                           PTMP_541_port, S(28) => PTMP_540_port, S(27) => 
                           PTMP_539_port, S(26) => PTMP_538_port, S(25) => 
                           PTMP_537_port, S(24) => PTMP_536_port, S(23) => 
                           PTMP_535_port, S(22) => PTMP_534_port, S(21) => 
                           PTMP_533_port, S(20) => PTMP_532_port, S(19) => 
                           PTMP_531_port, S(18) => PTMP_530_port, S(17) => 
                           PTMP_529_port, S(16) => PTMP_528_port, S(15) => 
                           PTMP_527_port, S(14) => PTMP_526_port, S(13) => 
                           PTMP_525_port, S(12) => PTMP_524_port, S(11) => 
                           PTMP_523_port, S(10) => PTMP_522_port, S(9) => 
                           PTMP_521_port, S(8) => PTMP_520_port, S(7) => 
                           PTMP_519_port, S(6) => PTMP_518_port, S(5) => 
                           PTMP_517_port, S(4) => PTMP_516_port, S(3) => 
                           PTMP_515_port, S(2) => PTMP_514_port, S(1) => 
                           PTMP_513_port, S(0) => PTMP_512_port, Co => n_1303);
   ADDERI_11 : RCA_NBIT64_21 port map( A(63) => PTMP_575_port, A(62) => 
                           PTMP_574_port, A(61) => PTMP_573_port, A(60) => 
                           PTMP_572_port, A(59) => PTMP_571_port, A(58) => 
                           PTMP_570_port, A(57) => PTMP_569_port, A(56) => 
                           PTMP_568_port, A(55) => PTMP_567_port, A(54) => 
                           PTMP_566_port, A(53) => PTMP_565_port, A(52) => 
                           PTMP_564_port, A(51) => PTMP_563_port, A(50) => 
                           PTMP_562_port, A(49) => PTMP_561_port, A(48) => 
                           PTMP_560_port, A(47) => PTMP_559_port, A(46) => 
                           PTMP_558_port, A(45) => PTMP_557_port, A(44) => 
                           PTMP_556_port, A(43) => PTMP_555_port, A(42) => 
                           PTMP_554_port, A(41) => PTMP_553_port, A(40) => 
                           PTMP_552_port, A(39) => PTMP_551_port, A(38) => 
                           PTMP_550_port, A(37) => PTMP_549_port, A(36) => 
                           PTMP_548_port, A(35) => PTMP_547_port, A(34) => 
                           PTMP_546_port, A(33) => PTMP_545_port, A(32) => 
                           PTMP_544_port, A(31) => PTMP_543_port, A(30) => 
                           PTMP_542_port, A(29) => PTMP_541_port, A(28) => 
                           PTMP_540_port, A(27) => PTMP_539_port, A(26) => 
                           PTMP_538_port, A(25) => PTMP_537_port, A(24) => 
                           PTMP_536_port, A(23) => PTMP_535_port, A(22) => 
                           PTMP_534_port, A(21) => PTMP_533_port, A(20) => 
                           PTMP_532_port, A(19) => PTMP_531_port, A(18) => 
                           PTMP_530_port, A(17) => PTMP_529_port, A(16) => 
                           PTMP_528_port, A(15) => PTMP_527_port, A(14) => 
                           PTMP_526_port, A(13) => PTMP_525_port, A(12) => 
                           PTMP_524_port, A(11) => PTMP_523_port, A(10) => 
                           PTMP_522_port, A(9) => PTMP_521_port, A(8) => 
                           PTMP_520_port, A(7) => PTMP_519_port, A(6) => 
                           PTMP_518_port, A(5) => PTMP_517_port, A(4) => 
                           PTMP_516_port, A(3) => PTMP_515_port, A(2) => 
                           PTMP_514_port, A(1) => PTMP_513_port, A(0) => 
                           PTMP_512_port, B(63) => OTMP_703_port, B(62) => 
                           OTMP_702_port, B(61) => OTMP_701_port, B(60) => 
                           OTMP_700_port, B(59) => OTMP_699_port, B(58) => 
                           OTMP_698_port, B(57) => OTMP_697_port, B(56) => 
                           OTMP_696_port, B(55) => OTMP_695_port, B(54) => 
                           OTMP_694_port, B(53) => OTMP_693_port, B(52) => 
                           OTMP_692_port, B(51) => OTMP_691_port, B(50) => 
                           OTMP_690_port, B(49) => OTMP_689_port, B(48) => 
                           OTMP_688_port, B(47) => OTMP_687_port, B(46) => 
                           OTMP_686_port, B(45) => OTMP_685_port, B(44) => 
                           OTMP_684_port, B(43) => OTMP_683_port, B(42) => 
                           OTMP_682_port, B(41) => OTMP_681_port, B(40) => 
                           OTMP_680_port, B(39) => OTMP_679_port, B(38) => 
                           OTMP_678_port, B(37) => OTMP_677_port, B(36) => 
                           OTMP_676_port, B(35) => OTMP_675_port, B(34) => 
                           OTMP_674_port, B(33) => OTMP_673_port, B(32) => 
                           OTMP_672_port, B(31) => OTMP_671_port, B(30) => 
                           OTMP_670_port, B(29) => OTMP_669_port, B(28) => 
                           OTMP_668_port, B(27) => OTMP_667_port, B(26) => 
                           OTMP_666_port, B(25) => OTMP_665_port, B(24) => 
                           OTMP_664_port, B(23) => OTMP_663_port, B(22) => 
                           OTMP_662_port, B(21) => OTMP_661_port, B(20) => 
                           OTMP_660_port, B(19) => OTMP_659_port, B(18) => 
                           OTMP_658_port, B(17) => OTMP_657_port, B(16) => 
                           OTMP_656_port, B(15) => OTMP_655_port, B(14) => 
                           OTMP_654_port, B(13) => OTMP_653_port, B(12) => 
                           OTMP_652_port, B(11) => OTMP_651_port, B(10) => 
                           OTMP_650_port, B(9) => OTMP_649_port, B(8) => 
                           OTMP_648_port, B(7) => OTMP_647_port, B(6) => 
                           OTMP_646_port, B(5) => OTMP_645_port, B(4) => 
                           OTMP_644_port, B(3) => OTMP_643_port, B(2) => 
                           OTMP_642_port, B(1) => OTMP_641_port, B(0) => 
                           OTMP_640_port, Ci => X_Logic0_port, S(63) => 
                           PTMP_639_port, S(62) => PTMP_638_port, S(61) => 
                           PTMP_637_port, S(60) => PTMP_636_port, S(59) => 
                           PTMP_635_port, S(58) => PTMP_634_port, S(57) => 
                           PTMP_633_port, S(56) => PTMP_632_port, S(55) => 
                           PTMP_631_port, S(54) => PTMP_630_port, S(53) => 
                           PTMP_629_port, S(52) => PTMP_628_port, S(51) => 
                           PTMP_627_port, S(50) => PTMP_626_port, S(49) => 
                           PTMP_625_port, S(48) => PTMP_624_port, S(47) => 
                           PTMP_623_port, S(46) => PTMP_622_port, S(45) => 
                           PTMP_621_port, S(44) => PTMP_620_port, S(43) => 
                           PTMP_619_port, S(42) => PTMP_618_port, S(41) => 
                           PTMP_617_port, S(40) => PTMP_616_port, S(39) => 
                           PTMP_615_port, S(38) => PTMP_614_port, S(37) => 
                           PTMP_613_port, S(36) => PTMP_612_port, S(35) => 
                           PTMP_611_port, S(34) => PTMP_610_port, S(33) => 
                           PTMP_609_port, S(32) => PTMP_608_port, S(31) => 
                           PTMP_607_port, S(30) => PTMP_606_port, S(29) => 
                           PTMP_605_port, S(28) => PTMP_604_port, S(27) => 
                           PTMP_603_port, S(26) => PTMP_602_port, S(25) => 
                           PTMP_601_port, S(24) => PTMP_600_port, S(23) => 
                           PTMP_599_port, S(22) => PTMP_598_port, S(21) => 
                           PTMP_597_port, S(20) => PTMP_596_port, S(19) => 
                           PTMP_595_port, S(18) => PTMP_594_port, S(17) => 
                           PTMP_593_port, S(16) => PTMP_592_port, S(15) => 
                           PTMP_591_port, S(14) => PTMP_590_port, S(13) => 
                           PTMP_589_port, S(12) => PTMP_588_port, S(11) => 
                           PTMP_587_port, S(10) => PTMP_586_port, S(9) => 
                           PTMP_585_port, S(8) => PTMP_584_port, S(7) => 
                           PTMP_583_port, S(6) => PTMP_582_port, S(5) => 
                           PTMP_581_port, S(4) => PTMP_580_port, S(3) => 
                           PTMP_579_port, S(2) => PTMP_578_port, S(1) => 
                           PTMP_577_port, S(0) => PTMP_576_port, Co => n_1304);
   ADDERI_12 : RCA_NBIT64_20 port map( A(63) => PTMP_639_port, A(62) => 
                           PTMP_638_port, A(61) => PTMP_637_port, A(60) => 
                           PTMP_636_port, A(59) => PTMP_635_port, A(58) => 
                           PTMP_634_port, A(57) => PTMP_633_port, A(56) => 
                           PTMP_632_port, A(55) => PTMP_631_port, A(54) => 
                           PTMP_630_port, A(53) => PTMP_629_port, A(52) => 
                           PTMP_628_port, A(51) => PTMP_627_port, A(50) => 
                           PTMP_626_port, A(49) => PTMP_625_port, A(48) => 
                           PTMP_624_port, A(47) => PTMP_623_port, A(46) => 
                           PTMP_622_port, A(45) => PTMP_621_port, A(44) => 
                           PTMP_620_port, A(43) => PTMP_619_port, A(42) => 
                           PTMP_618_port, A(41) => PTMP_617_port, A(40) => 
                           PTMP_616_port, A(39) => PTMP_615_port, A(38) => 
                           PTMP_614_port, A(37) => PTMP_613_port, A(36) => 
                           PTMP_612_port, A(35) => PTMP_611_port, A(34) => 
                           PTMP_610_port, A(33) => PTMP_609_port, A(32) => 
                           PTMP_608_port, A(31) => PTMP_607_port, A(30) => 
                           PTMP_606_port, A(29) => PTMP_605_port, A(28) => 
                           PTMP_604_port, A(27) => PTMP_603_port, A(26) => 
                           PTMP_602_port, A(25) => PTMP_601_port, A(24) => 
                           PTMP_600_port, A(23) => PTMP_599_port, A(22) => 
                           PTMP_598_port, A(21) => PTMP_597_port, A(20) => 
                           PTMP_596_port, A(19) => PTMP_595_port, A(18) => 
                           PTMP_594_port, A(17) => PTMP_593_port, A(16) => 
                           PTMP_592_port, A(15) => PTMP_591_port, A(14) => 
                           PTMP_590_port, A(13) => PTMP_589_port, A(12) => 
                           PTMP_588_port, A(11) => PTMP_587_port, A(10) => 
                           PTMP_586_port, A(9) => PTMP_585_port, A(8) => 
                           PTMP_584_port, A(7) => PTMP_583_port, A(6) => 
                           PTMP_582_port, A(5) => PTMP_581_port, A(4) => 
                           PTMP_580_port, A(3) => PTMP_579_port, A(2) => 
                           PTMP_578_port, A(1) => PTMP_577_port, A(0) => 
                           PTMP_576_port, B(63) => OTMP_767_port, B(62) => 
                           OTMP_766_port, B(61) => OTMP_765_port, B(60) => 
                           OTMP_764_port, B(59) => OTMP_763_port, B(58) => 
                           OTMP_762_port, B(57) => OTMP_761_port, B(56) => 
                           OTMP_760_port, B(55) => OTMP_759_port, B(54) => 
                           OTMP_758_port, B(53) => OTMP_757_port, B(52) => 
                           OTMP_756_port, B(51) => OTMP_755_port, B(50) => 
                           OTMP_754_port, B(49) => OTMP_753_port, B(48) => 
                           OTMP_752_port, B(47) => OTMP_751_port, B(46) => 
                           OTMP_750_port, B(45) => OTMP_749_port, B(44) => 
                           OTMP_748_port, B(43) => OTMP_747_port, B(42) => 
                           OTMP_746_port, B(41) => OTMP_745_port, B(40) => 
                           OTMP_744_port, B(39) => OTMP_743_port, B(38) => 
                           OTMP_742_port, B(37) => OTMP_741_port, B(36) => 
                           OTMP_740_port, B(35) => OTMP_739_port, B(34) => 
                           OTMP_738_port, B(33) => OTMP_737_port, B(32) => 
                           OTMP_736_port, B(31) => OTMP_735_port, B(30) => 
                           OTMP_734_port, B(29) => OTMP_733_port, B(28) => 
                           OTMP_732_port, B(27) => OTMP_731_port, B(26) => 
                           OTMP_730_port, B(25) => OTMP_729_port, B(24) => 
                           OTMP_728_port, B(23) => OTMP_727_port, B(22) => 
                           OTMP_726_port, B(21) => OTMP_725_port, B(20) => 
                           OTMP_724_port, B(19) => OTMP_723_port, B(18) => 
                           OTMP_722_port, B(17) => OTMP_721_port, B(16) => 
                           OTMP_720_port, B(15) => OTMP_719_port, B(14) => 
                           OTMP_718_port, B(13) => OTMP_717_port, B(12) => 
                           OTMP_716_port, B(11) => OTMP_715_port, B(10) => 
                           OTMP_714_port, B(9) => OTMP_713_port, B(8) => 
                           OTMP_712_port, B(7) => OTMP_711_port, B(6) => 
                           OTMP_710_port, B(5) => OTMP_709_port, B(4) => 
                           OTMP_708_port, B(3) => OTMP_707_port, B(2) => 
                           OTMP_706_port, B(1) => OTMP_705_port, B(0) => 
                           OTMP_704_port, Ci => X_Logic0_port, S(63) => 
                           PTMP_703_port, S(62) => PTMP_702_port, S(61) => 
                           PTMP_701_port, S(60) => PTMP_700_port, S(59) => 
                           PTMP_699_port, S(58) => PTMP_698_port, S(57) => 
                           PTMP_697_port, S(56) => PTMP_696_port, S(55) => 
                           PTMP_695_port, S(54) => PTMP_694_port, S(53) => 
                           PTMP_693_port, S(52) => PTMP_692_port, S(51) => 
                           PTMP_691_port, S(50) => PTMP_690_port, S(49) => 
                           PTMP_689_port, S(48) => PTMP_688_port, S(47) => 
                           PTMP_687_port, S(46) => PTMP_686_port, S(45) => 
                           PTMP_685_port, S(44) => PTMP_684_port, S(43) => 
                           PTMP_683_port, S(42) => PTMP_682_port, S(41) => 
                           PTMP_681_port, S(40) => PTMP_680_port, S(39) => 
                           PTMP_679_port, S(38) => PTMP_678_port, S(37) => 
                           PTMP_677_port, S(36) => PTMP_676_port, S(35) => 
                           PTMP_675_port, S(34) => PTMP_674_port, S(33) => 
                           PTMP_673_port, S(32) => PTMP_672_port, S(31) => 
                           PTMP_671_port, S(30) => PTMP_670_port, S(29) => 
                           PTMP_669_port, S(28) => PTMP_668_port, S(27) => 
                           PTMP_667_port, S(26) => PTMP_666_port, S(25) => 
                           PTMP_665_port, S(24) => PTMP_664_port, S(23) => 
                           PTMP_663_port, S(22) => PTMP_662_port, S(21) => 
                           PTMP_661_port, S(20) => PTMP_660_port, S(19) => 
                           PTMP_659_port, S(18) => PTMP_658_port, S(17) => 
                           PTMP_657_port, S(16) => PTMP_656_port, S(15) => 
                           PTMP_655_port, S(14) => PTMP_654_port, S(13) => 
                           PTMP_653_port, S(12) => PTMP_652_port, S(11) => 
                           PTMP_651_port, S(10) => PTMP_650_port, S(9) => 
                           PTMP_649_port, S(8) => PTMP_648_port, S(7) => 
                           PTMP_647_port, S(6) => PTMP_646_port, S(5) => 
                           PTMP_645_port, S(4) => PTMP_644_port, S(3) => 
                           PTMP_643_port, S(2) => PTMP_642_port, S(1) => 
                           PTMP_641_port, S(0) => PTMP_640_port, Co => n_1305);
   ADDERI_13 : RCA_NBIT64_19 port map( A(63) => PTMP_703_port, A(62) => 
                           PTMP_702_port, A(61) => PTMP_701_port, A(60) => 
                           PTMP_700_port, A(59) => PTMP_699_port, A(58) => 
                           PTMP_698_port, A(57) => PTMP_697_port, A(56) => 
                           PTMP_696_port, A(55) => PTMP_695_port, A(54) => 
                           PTMP_694_port, A(53) => PTMP_693_port, A(52) => 
                           PTMP_692_port, A(51) => PTMP_691_port, A(50) => 
                           PTMP_690_port, A(49) => PTMP_689_port, A(48) => 
                           PTMP_688_port, A(47) => PTMP_687_port, A(46) => 
                           PTMP_686_port, A(45) => PTMP_685_port, A(44) => 
                           PTMP_684_port, A(43) => PTMP_683_port, A(42) => 
                           PTMP_682_port, A(41) => PTMP_681_port, A(40) => 
                           PTMP_680_port, A(39) => PTMP_679_port, A(38) => 
                           PTMP_678_port, A(37) => PTMP_677_port, A(36) => 
                           PTMP_676_port, A(35) => PTMP_675_port, A(34) => 
                           PTMP_674_port, A(33) => PTMP_673_port, A(32) => 
                           PTMP_672_port, A(31) => PTMP_671_port, A(30) => 
                           PTMP_670_port, A(29) => PTMP_669_port, A(28) => 
                           PTMP_668_port, A(27) => PTMP_667_port, A(26) => 
                           PTMP_666_port, A(25) => PTMP_665_port, A(24) => 
                           PTMP_664_port, A(23) => PTMP_663_port, A(22) => 
                           PTMP_662_port, A(21) => PTMP_661_port, A(20) => 
                           PTMP_660_port, A(19) => PTMP_659_port, A(18) => 
                           PTMP_658_port, A(17) => PTMP_657_port, A(16) => 
                           PTMP_656_port, A(15) => PTMP_655_port, A(14) => 
                           PTMP_654_port, A(13) => PTMP_653_port, A(12) => 
                           PTMP_652_port, A(11) => PTMP_651_port, A(10) => 
                           PTMP_650_port, A(9) => PTMP_649_port, A(8) => 
                           PTMP_648_port, A(7) => PTMP_647_port, A(6) => 
                           PTMP_646_port, A(5) => PTMP_645_port, A(4) => 
                           PTMP_644_port, A(3) => PTMP_643_port, A(2) => 
                           PTMP_642_port, A(1) => PTMP_641_port, A(0) => 
                           PTMP_640_port, B(63) => OTMP_831_port, B(62) => 
                           OTMP_830_port, B(61) => OTMP_829_port, B(60) => 
                           OTMP_828_port, B(59) => OTMP_827_port, B(58) => 
                           OTMP_826_port, B(57) => OTMP_825_port, B(56) => 
                           OTMP_824_port, B(55) => OTMP_823_port, B(54) => 
                           OTMP_822_port, B(53) => OTMP_821_port, B(52) => 
                           OTMP_820_port, B(51) => OTMP_819_port, B(50) => 
                           OTMP_818_port, B(49) => OTMP_817_port, B(48) => 
                           OTMP_816_port, B(47) => OTMP_815_port, B(46) => 
                           OTMP_814_port, B(45) => OTMP_813_port, B(44) => 
                           OTMP_812_port, B(43) => OTMP_811_port, B(42) => 
                           OTMP_810_port, B(41) => OTMP_809_port, B(40) => 
                           OTMP_808_port, B(39) => OTMP_807_port, B(38) => 
                           OTMP_806_port, B(37) => OTMP_805_port, B(36) => 
                           OTMP_804_port, B(35) => OTMP_803_port, B(34) => 
                           OTMP_802_port, B(33) => OTMP_801_port, B(32) => 
                           OTMP_800_port, B(31) => OTMP_799_port, B(30) => 
                           OTMP_798_port, B(29) => OTMP_797_port, B(28) => 
                           OTMP_796_port, B(27) => OTMP_795_port, B(26) => 
                           OTMP_794_port, B(25) => OTMP_793_port, B(24) => 
                           OTMP_792_port, B(23) => OTMP_791_port, B(22) => 
                           OTMP_790_port, B(21) => OTMP_789_port, B(20) => 
                           OTMP_788_port, B(19) => OTMP_787_port, B(18) => 
                           OTMP_786_port, B(17) => OTMP_785_port, B(16) => 
                           OTMP_784_port, B(15) => OTMP_783_port, B(14) => 
                           OTMP_782_port, B(13) => OTMP_781_port, B(12) => 
                           OTMP_780_port, B(11) => OTMP_779_port, B(10) => 
                           OTMP_778_port, B(9) => OTMP_777_port, B(8) => 
                           OTMP_776_port, B(7) => OTMP_775_port, B(6) => 
                           OTMP_774_port, B(5) => OTMP_773_port, B(4) => 
                           OTMP_772_port, B(3) => OTMP_771_port, B(2) => 
                           OTMP_770_port, B(1) => OTMP_769_port, B(0) => 
                           OTMP_768_port, Ci => X_Logic0_port, S(63) => 
                           PTMP_767_port, S(62) => PTMP_766_port, S(61) => 
                           PTMP_765_port, S(60) => PTMP_764_port, S(59) => 
                           PTMP_763_port, S(58) => PTMP_762_port, S(57) => 
                           PTMP_761_port, S(56) => PTMP_760_port, S(55) => 
                           PTMP_759_port, S(54) => PTMP_758_port, S(53) => 
                           PTMP_757_port, S(52) => PTMP_756_port, S(51) => 
                           PTMP_755_port, S(50) => PTMP_754_port, S(49) => 
                           PTMP_753_port, S(48) => PTMP_752_port, S(47) => 
                           PTMP_751_port, S(46) => PTMP_750_port, S(45) => 
                           PTMP_749_port, S(44) => PTMP_748_port, S(43) => 
                           PTMP_747_port, S(42) => PTMP_746_port, S(41) => 
                           PTMP_745_port, S(40) => PTMP_744_port, S(39) => 
                           PTMP_743_port, S(38) => PTMP_742_port, S(37) => 
                           PTMP_741_port, S(36) => PTMP_740_port, S(35) => 
                           PTMP_739_port, S(34) => PTMP_738_port, S(33) => 
                           PTMP_737_port, S(32) => PTMP_736_port, S(31) => 
                           PTMP_735_port, S(30) => PTMP_734_port, S(29) => 
                           PTMP_733_port, S(28) => PTMP_732_port, S(27) => 
                           PTMP_731_port, S(26) => PTMP_730_port, S(25) => 
                           PTMP_729_port, S(24) => PTMP_728_port, S(23) => 
                           PTMP_727_port, S(22) => PTMP_726_port, S(21) => 
                           PTMP_725_port, S(20) => PTMP_724_port, S(19) => 
                           PTMP_723_port, S(18) => PTMP_722_port, S(17) => 
                           PTMP_721_port, S(16) => PTMP_720_port, S(15) => 
                           PTMP_719_port, S(14) => PTMP_718_port, S(13) => 
                           PTMP_717_port, S(12) => PTMP_716_port, S(11) => 
                           PTMP_715_port, S(10) => PTMP_714_port, S(9) => 
                           PTMP_713_port, S(8) => PTMP_712_port, S(7) => 
                           PTMP_711_port, S(6) => PTMP_710_port, S(5) => 
                           PTMP_709_port, S(4) => PTMP_708_port, S(3) => 
                           PTMP_707_port, S(2) => PTMP_706_port, S(1) => 
                           PTMP_705_port, S(0) => PTMP_704_port, Co => n_1306);
   ADDERI_14 : RCA_NBIT64_18 port map( A(63) => PTMP_767_port, A(62) => 
                           PTMP_766_port, A(61) => PTMP_765_port, A(60) => 
                           PTMP_764_port, A(59) => PTMP_763_port, A(58) => 
                           PTMP_762_port, A(57) => PTMP_761_port, A(56) => 
                           PTMP_760_port, A(55) => PTMP_759_port, A(54) => 
                           PTMP_758_port, A(53) => PTMP_757_port, A(52) => 
                           PTMP_756_port, A(51) => PTMP_755_port, A(50) => 
                           PTMP_754_port, A(49) => PTMP_753_port, A(48) => 
                           PTMP_752_port, A(47) => PTMP_751_port, A(46) => 
                           PTMP_750_port, A(45) => PTMP_749_port, A(44) => 
                           PTMP_748_port, A(43) => PTMP_747_port, A(42) => 
                           PTMP_746_port, A(41) => PTMP_745_port, A(40) => 
                           PTMP_744_port, A(39) => PTMP_743_port, A(38) => 
                           PTMP_742_port, A(37) => PTMP_741_port, A(36) => 
                           PTMP_740_port, A(35) => PTMP_739_port, A(34) => 
                           PTMP_738_port, A(33) => PTMP_737_port, A(32) => 
                           PTMP_736_port, A(31) => PTMP_735_port, A(30) => 
                           PTMP_734_port, A(29) => PTMP_733_port, A(28) => 
                           PTMP_732_port, A(27) => PTMP_731_port, A(26) => 
                           PTMP_730_port, A(25) => PTMP_729_port, A(24) => 
                           PTMP_728_port, A(23) => PTMP_727_port, A(22) => 
                           PTMP_726_port, A(21) => PTMP_725_port, A(20) => 
                           PTMP_724_port, A(19) => PTMP_723_port, A(18) => 
                           PTMP_722_port, A(17) => PTMP_721_port, A(16) => 
                           PTMP_720_port, A(15) => PTMP_719_port, A(14) => 
                           PTMP_718_port, A(13) => PTMP_717_port, A(12) => 
                           PTMP_716_port, A(11) => PTMP_715_port, A(10) => 
                           PTMP_714_port, A(9) => PTMP_713_port, A(8) => 
                           PTMP_712_port, A(7) => PTMP_711_port, A(6) => 
                           PTMP_710_port, A(5) => PTMP_709_port, A(4) => 
                           PTMP_708_port, A(3) => PTMP_707_port, A(2) => 
                           PTMP_706_port, A(1) => PTMP_705_port, A(0) => 
                           PTMP_704_port, B(63) => OTMP_895_port, B(62) => 
                           OTMP_894_port, B(61) => OTMP_893_port, B(60) => 
                           OTMP_892_port, B(59) => OTMP_891_port, B(58) => 
                           OTMP_890_port, B(57) => OTMP_889_port, B(56) => 
                           OTMP_888_port, B(55) => OTMP_887_port, B(54) => 
                           OTMP_886_port, B(53) => OTMP_885_port, B(52) => 
                           OTMP_884_port, B(51) => OTMP_883_port, B(50) => 
                           OTMP_882_port, B(49) => OTMP_881_port, B(48) => 
                           OTMP_880_port, B(47) => OTMP_879_port, B(46) => 
                           OTMP_878_port, B(45) => OTMP_877_port, B(44) => 
                           OTMP_876_port, B(43) => OTMP_875_port, B(42) => 
                           OTMP_874_port, B(41) => OTMP_873_port, B(40) => 
                           OTMP_872_port, B(39) => OTMP_871_port, B(38) => 
                           OTMP_870_port, B(37) => OTMP_869_port, B(36) => 
                           OTMP_868_port, B(35) => OTMP_867_port, B(34) => 
                           OTMP_866_port, B(33) => OTMP_865_port, B(32) => 
                           OTMP_864_port, B(31) => OTMP_863_port, B(30) => 
                           OTMP_862_port, B(29) => OTMP_861_port, B(28) => 
                           OTMP_860_port, B(27) => OTMP_859_port, B(26) => 
                           OTMP_858_port, B(25) => OTMP_857_port, B(24) => 
                           OTMP_856_port, B(23) => OTMP_855_port, B(22) => 
                           OTMP_854_port, B(21) => OTMP_853_port, B(20) => 
                           OTMP_852_port, B(19) => OTMP_851_port, B(18) => 
                           OTMP_850_port, B(17) => OTMP_849_port, B(16) => 
                           OTMP_848_port, B(15) => OTMP_847_port, B(14) => 
                           OTMP_846_port, B(13) => OTMP_845_port, B(12) => 
                           OTMP_844_port, B(11) => OTMP_843_port, B(10) => 
                           OTMP_842_port, B(9) => OTMP_841_port, B(8) => 
                           OTMP_840_port, B(7) => OTMP_839_port, B(6) => 
                           OTMP_838_port, B(5) => OTMP_837_port, B(4) => 
                           OTMP_836_port, B(3) => OTMP_835_port, B(2) => 
                           OTMP_834_port, B(1) => OTMP_833_port, B(0) => 
                           OTMP_832_port, Ci => X_Logic0_port, S(63) => 
                           PTMP_831_port, S(62) => PTMP_830_port, S(61) => 
                           PTMP_829_port, S(60) => PTMP_828_port, S(59) => 
                           PTMP_827_port, S(58) => PTMP_826_port, S(57) => 
                           PTMP_825_port, S(56) => PTMP_824_port, S(55) => 
                           PTMP_823_port, S(54) => PTMP_822_port, S(53) => 
                           PTMP_821_port, S(52) => PTMP_820_port, S(51) => 
                           PTMP_819_port, S(50) => PTMP_818_port, S(49) => 
                           PTMP_817_port, S(48) => PTMP_816_port, S(47) => 
                           PTMP_815_port, S(46) => PTMP_814_port, S(45) => 
                           PTMP_813_port, S(44) => PTMP_812_port, S(43) => 
                           PTMP_811_port, S(42) => PTMP_810_port, S(41) => 
                           PTMP_809_port, S(40) => PTMP_808_port, S(39) => 
                           PTMP_807_port, S(38) => PTMP_806_port, S(37) => 
                           PTMP_805_port, S(36) => PTMP_804_port, S(35) => 
                           PTMP_803_port, S(34) => PTMP_802_port, S(33) => 
                           PTMP_801_port, S(32) => PTMP_800_port, S(31) => 
                           PTMP_799_port, S(30) => PTMP_798_port, S(29) => 
                           PTMP_797_port, S(28) => PTMP_796_port, S(27) => 
                           PTMP_795_port, S(26) => PTMP_794_port, S(25) => 
                           PTMP_793_port, S(24) => PTMP_792_port, S(23) => 
                           PTMP_791_port, S(22) => PTMP_790_port, S(21) => 
                           PTMP_789_port, S(20) => PTMP_788_port, S(19) => 
                           PTMP_787_port, S(18) => PTMP_786_port, S(17) => 
                           PTMP_785_port, S(16) => PTMP_784_port, S(15) => 
                           PTMP_783_port, S(14) => PTMP_782_port, S(13) => 
                           PTMP_781_port, S(12) => PTMP_780_port, S(11) => 
                           PTMP_779_port, S(10) => PTMP_778_port, S(9) => 
                           PTMP_777_port, S(8) => PTMP_776_port, S(7) => 
                           PTMP_775_port, S(6) => PTMP_774_port, S(5) => 
                           PTMP_773_port, S(4) => PTMP_772_port, S(3) => 
                           PTMP_771_port, S(2) => PTMP_770_port, S(1) => 
                           PTMP_769_port, S(0) => PTMP_768_port, Co => n_1307);
   ADDERI_15 : RCA_NBIT64_17 port map( A(63) => PTMP_831_port, A(62) => 
                           PTMP_830_port, A(61) => PTMP_829_port, A(60) => 
                           PTMP_828_port, A(59) => PTMP_827_port, A(58) => 
                           PTMP_826_port, A(57) => PTMP_825_port, A(56) => 
                           PTMP_824_port, A(55) => PTMP_823_port, A(54) => 
                           PTMP_822_port, A(53) => PTMP_821_port, A(52) => 
                           PTMP_820_port, A(51) => PTMP_819_port, A(50) => 
                           PTMP_818_port, A(49) => PTMP_817_port, A(48) => 
                           PTMP_816_port, A(47) => PTMP_815_port, A(46) => 
                           PTMP_814_port, A(45) => PTMP_813_port, A(44) => 
                           PTMP_812_port, A(43) => PTMP_811_port, A(42) => 
                           PTMP_810_port, A(41) => PTMP_809_port, A(40) => 
                           PTMP_808_port, A(39) => PTMP_807_port, A(38) => 
                           PTMP_806_port, A(37) => PTMP_805_port, A(36) => 
                           PTMP_804_port, A(35) => PTMP_803_port, A(34) => 
                           PTMP_802_port, A(33) => PTMP_801_port, A(32) => 
                           PTMP_800_port, A(31) => PTMP_799_port, A(30) => 
                           PTMP_798_port, A(29) => PTMP_797_port, A(28) => 
                           PTMP_796_port, A(27) => PTMP_795_port, A(26) => 
                           PTMP_794_port, A(25) => PTMP_793_port, A(24) => 
                           PTMP_792_port, A(23) => PTMP_791_port, A(22) => 
                           PTMP_790_port, A(21) => PTMP_789_port, A(20) => 
                           PTMP_788_port, A(19) => PTMP_787_port, A(18) => 
                           PTMP_786_port, A(17) => PTMP_785_port, A(16) => 
                           PTMP_784_port, A(15) => PTMP_783_port, A(14) => 
                           PTMP_782_port, A(13) => PTMP_781_port, A(12) => 
                           PTMP_780_port, A(11) => PTMP_779_port, A(10) => 
                           PTMP_778_port, A(9) => PTMP_777_port, A(8) => 
                           PTMP_776_port, A(7) => PTMP_775_port, A(6) => 
                           PTMP_774_port, A(5) => PTMP_773_port, A(4) => 
                           PTMP_772_port, A(3) => PTMP_771_port, A(2) => 
                           PTMP_770_port, A(1) => PTMP_769_port, A(0) => 
                           PTMP_768_port, B(63) => OTMP_959_port, B(62) => 
                           OTMP_958_port, B(61) => OTMP_957_port, B(60) => 
                           OTMP_956_port, B(59) => OTMP_955_port, B(58) => 
                           OTMP_954_port, B(57) => OTMP_953_port, B(56) => 
                           OTMP_952_port, B(55) => OTMP_951_port, B(54) => 
                           OTMP_950_port, B(53) => OTMP_949_port, B(52) => 
                           OTMP_948_port, B(51) => OTMP_947_port, B(50) => 
                           OTMP_946_port, B(49) => OTMP_945_port, B(48) => 
                           OTMP_944_port, B(47) => OTMP_943_port, B(46) => 
                           OTMP_942_port, B(45) => OTMP_941_port, B(44) => 
                           OTMP_940_port, B(43) => OTMP_939_port, B(42) => 
                           OTMP_938_port, B(41) => OTMP_937_port, B(40) => 
                           OTMP_936_port, B(39) => OTMP_935_port, B(38) => 
                           OTMP_934_port, B(37) => OTMP_933_port, B(36) => 
                           OTMP_932_port, B(35) => OTMP_931_port, B(34) => 
                           OTMP_930_port, B(33) => OTMP_929_port, B(32) => 
                           OTMP_928_port, B(31) => OTMP_927_port, B(30) => 
                           OTMP_926_port, B(29) => OTMP_925_port, B(28) => 
                           OTMP_924_port, B(27) => OTMP_923_port, B(26) => 
                           OTMP_922_port, B(25) => OTMP_921_port, B(24) => 
                           OTMP_920_port, B(23) => OTMP_919_port, B(22) => 
                           OTMP_918_port, B(21) => OTMP_917_port, B(20) => 
                           OTMP_916_port, B(19) => OTMP_915_port, B(18) => 
                           OTMP_914_port, B(17) => OTMP_913_port, B(16) => 
                           OTMP_912_port, B(15) => OTMP_911_port, B(14) => 
                           OTMP_910_port, B(13) => OTMP_909_port, B(12) => 
                           OTMP_908_port, B(11) => OTMP_907_port, B(10) => 
                           OTMP_906_port, B(9) => OTMP_905_port, B(8) => 
                           OTMP_904_port, B(7) => OTMP_903_port, B(6) => 
                           OTMP_902_port, B(5) => OTMP_901_port, B(4) => 
                           OTMP_900_port, B(3) => OTMP_899_port, B(2) => 
                           OTMP_898_port, B(1) => OTMP_897_port, B(0) => 
                           OTMP_896_port, Ci => X_Logic0_port, S(63) => 
                           PTMP_895_port, S(62) => PTMP_894_port, S(61) => 
                           PTMP_893_port, S(60) => PTMP_892_port, S(59) => 
                           PTMP_891_port, S(58) => PTMP_890_port, S(57) => 
                           PTMP_889_port, S(56) => PTMP_888_port, S(55) => 
                           PTMP_887_port, S(54) => PTMP_886_port, S(53) => 
                           PTMP_885_port, S(52) => PTMP_884_port, S(51) => 
                           PTMP_883_port, S(50) => PTMP_882_port, S(49) => 
                           PTMP_881_port, S(48) => PTMP_880_port, S(47) => 
                           PTMP_879_port, S(46) => PTMP_878_port, S(45) => 
                           PTMP_877_port, S(44) => PTMP_876_port, S(43) => 
                           PTMP_875_port, S(42) => PTMP_874_port, S(41) => 
                           PTMP_873_port, S(40) => PTMP_872_port, S(39) => 
                           PTMP_871_port, S(38) => PTMP_870_port, S(37) => 
                           PTMP_869_port, S(36) => PTMP_868_port, S(35) => 
                           PTMP_867_port, S(34) => PTMP_866_port, S(33) => 
                           PTMP_865_port, S(32) => PTMP_864_port, S(31) => 
                           PTMP_863_port, S(30) => PTMP_862_port, S(29) => 
                           PTMP_861_port, S(28) => PTMP_860_port, S(27) => 
                           PTMP_859_port, S(26) => PTMP_858_port, S(25) => 
                           PTMP_857_port, S(24) => PTMP_856_port, S(23) => 
                           PTMP_855_port, S(22) => PTMP_854_port, S(21) => 
                           PTMP_853_port, S(20) => PTMP_852_port, S(19) => 
                           PTMP_851_port, S(18) => PTMP_850_port, S(17) => 
                           PTMP_849_port, S(16) => PTMP_848_port, S(15) => 
                           PTMP_847_port, S(14) => PTMP_846_port, S(13) => 
                           PTMP_845_port, S(12) => PTMP_844_port, S(11) => 
                           PTMP_843_port, S(10) => PTMP_842_port, S(9) => 
                           PTMP_841_port, S(8) => PTMP_840_port, S(7) => 
                           PTMP_839_port, S(6) => PTMP_838_port, S(5) => 
                           PTMP_837_port, S(4) => PTMP_836_port, S(3) => 
                           PTMP_835_port, S(2) => PTMP_834_port, S(1) => 
                           PTMP_833_port, S(0) => PTMP_832_port, Co => n_1308);
   ADDERI_16 : RCA_NBIT64_16 port map( A(63) => PTMP_895_port, A(62) => 
                           PTMP_894_port, A(61) => PTMP_893_port, A(60) => 
                           PTMP_892_port, A(59) => PTMP_891_port, A(58) => 
                           PTMP_890_port, A(57) => PTMP_889_port, A(56) => 
                           PTMP_888_port, A(55) => PTMP_887_port, A(54) => 
                           PTMP_886_port, A(53) => PTMP_885_port, A(52) => 
                           PTMP_884_port, A(51) => PTMP_883_port, A(50) => 
                           PTMP_882_port, A(49) => PTMP_881_port, A(48) => 
                           PTMP_880_port, A(47) => PTMP_879_port, A(46) => 
                           PTMP_878_port, A(45) => PTMP_877_port, A(44) => 
                           PTMP_876_port, A(43) => PTMP_875_port, A(42) => 
                           PTMP_874_port, A(41) => PTMP_873_port, A(40) => 
                           PTMP_872_port, A(39) => PTMP_871_port, A(38) => 
                           PTMP_870_port, A(37) => PTMP_869_port, A(36) => 
                           PTMP_868_port, A(35) => PTMP_867_port, A(34) => 
                           PTMP_866_port, A(33) => PTMP_865_port, A(32) => 
                           PTMP_864_port, A(31) => PTMP_863_port, A(30) => 
                           PTMP_862_port, A(29) => PTMP_861_port, A(28) => 
                           PTMP_860_port, A(27) => PTMP_859_port, A(26) => 
                           PTMP_858_port, A(25) => PTMP_857_port, A(24) => 
                           PTMP_856_port, A(23) => PTMP_855_port, A(22) => 
                           PTMP_854_port, A(21) => PTMP_853_port, A(20) => 
                           PTMP_852_port, A(19) => PTMP_851_port, A(18) => 
                           PTMP_850_port, A(17) => PTMP_849_port, A(16) => 
                           PTMP_848_port, A(15) => PTMP_847_port, A(14) => 
                           PTMP_846_port, A(13) => PTMP_845_port, A(12) => 
                           PTMP_844_port, A(11) => PTMP_843_port, A(10) => 
                           PTMP_842_port, A(9) => PTMP_841_port, A(8) => 
                           PTMP_840_port, A(7) => PTMP_839_port, A(6) => 
                           PTMP_838_port, A(5) => PTMP_837_port, A(4) => 
                           PTMP_836_port, A(3) => PTMP_835_port, A(2) => 
                           PTMP_834_port, A(1) => PTMP_833_port, A(0) => 
                           PTMP_832_port, B(63) => OTMP_1023_port, B(62) => 
                           OTMP_1022_port, B(61) => OTMP_1021_port, B(60) => 
                           OTMP_1020_port, B(59) => OTMP_1019_port, B(58) => 
                           OTMP_1018_port, B(57) => OTMP_1017_port, B(56) => 
                           OTMP_1016_port, B(55) => OTMP_1015_port, B(54) => 
                           OTMP_1014_port, B(53) => OTMP_1013_port, B(52) => 
                           OTMP_1012_port, B(51) => OTMP_1011_port, B(50) => 
                           OTMP_1010_port, B(49) => OTMP_1009_port, B(48) => 
                           OTMP_1008_port, B(47) => OTMP_1007_port, B(46) => 
                           OTMP_1006_port, B(45) => OTMP_1005_port, B(44) => 
                           OTMP_1004_port, B(43) => OTMP_1003_port, B(42) => 
                           OTMP_1002_port, B(41) => OTMP_1001_port, B(40) => 
                           OTMP_1000_port, B(39) => OTMP_999_port, B(38) => 
                           OTMP_998_port, B(37) => OTMP_997_port, B(36) => 
                           OTMP_996_port, B(35) => OTMP_995_port, B(34) => 
                           OTMP_994_port, B(33) => OTMP_993_port, B(32) => 
                           OTMP_992_port, B(31) => OTMP_991_port, B(30) => 
                           OTMP_990_port, B(29) => OTMP_989_port, B(28) => 
                           OTMP_988_port, B(27) => OTMP_987_port, B(26) => 
                           OTMP_986_port, B(25) => OTMP_985_port, B(24) => 
                           OTMP_984_port, B(23) => OTMP_983_port, B(22) => 
                           OTMP_982_port, B(21) => OTMP_981_port, B(20) => 
                           OTMP_980_port, B(19) => OTMP_979_port, B(18) => 
                           OTMP_978_port, B(17) => OTMP_977_port, B(16) => 
                           OTMP_976_port, B(15) => OTMP_975_port, B(14) => 
                           OTMP_974_port, B(13) => OTMP_973_port, B(12) => 
                           OTMP_972_port, B(11) => OTMP_971_port, B(10) => 
                           OTMP_970_port, B(9) => OTMP_969_port, B(8) => 
                           OTMP_968_port, B(7) => OTMP_967_port, B(6) => 
                           OTMP_966_port, B(5) => OTMP_965_port, B(4) => 
                           OTMP_964_port, B(3) => OTMP_963_port, B(2) => 
                           OTMP_962_port, B(1) => OTMP_961_port, B(0) => 
                           OTMP_960_port, Ci => X_Logic0_port, S(63) => S(63), 
                           S(62) => S(62), S(61) => S(61), S(60) => S(60), 
                           S(59) => S(59), S(58) => S(58), S(57) => S(57), 
                           S(56) => S(56), S(55) => S(55), S(54) => S(54), 
                           S(53) => S(53), S(52) => S(52), S(51) => S(51), 
                           S(50) => S(50), S(49) => S(49), S(48) => S(48), 
                           S(47) => S(47), S(46) => S(46), S(45) => S(45), 
                           S(44) => S(44), S(43) => S(43), S(42) => S(42), 
                           S(41) => S(41), S(40) => S(40), S(39) => S(39), 
                           S(38) => S(38), S(37) => S(37), S(36) => S(36), 
                           S(35) => S(35), S(34) => S(34), S(33) => S(33), 
                           S(32) => S(32), S(31) => S(31), S(30) => S(30), 
                           S(29) => S(29), S(28) => S(28), S(27) => S(27), 
                           S(26) => S(26), S(25) => S(25), S(24) => S(24), 
                           S(23) => S(23), S(22) => S(22), S(21) => S(21), 
                           S(20) => S(20), S(19) => S(19), S(18) => S(18), 
                           S(17) => S(17), S(16) => S(16), S(15) => S(15), 
                           S(14) => S(14), S(13) => S(13), S(12) => S(12), 
                           S(11) => S(11), S(10) => S(10), S(9) => S(9), S(8) 
                           => S(8), S(7) => S(7), S(6) => S(6), S(5) => S(5), 
                           S(4) => S(4), S(3) => S(3), S(2) => S(2), S(1) => 
                           S(1), S(0) => S(0), Co => n_1309);
   sub_82 : BOOTHMUL_NBIT32_1_DW01_sub_0 port map( A(31) => n4, A(30) => n4, 
                           A(29) => n4, A(28) => n4, A(27) => n4, A(26) => n4, 
                           A(25) => n4, A(24) => n4, A(23) => n4, A(22) => n4, 
                           A(21) => n4, A(20) => n4, A(19) => n4, A(18) => n4, 
                           A(17) => n4, A(16) => n4, A(15) => n4, A(14) => n4, 
                           A(13) => n4, A(12) => n4, A(11) => n4, A(10) => n4, 
                           A(9) => n4, A(8) => n4, A(7) => n4, A(6) => n4, A(5)
                           => n4, A(4) => n4, A(3) => n4, A(2) => n4, A(1) => 
                           n4, A(0) => n4, B(31) => A(31), B(30) => A(30), 
                           B(29) => A(29), B(28) => A(28), B(27) => A(27), 
                           B(26) => A(26), B(25) => A(25), B(24) => A(24), 
                           B(23) => A(23), B(22) => A(22), B(21) => A(21), 
                           B(20) => A(20), B(19) => A(19), B(18) => A(18), 
                           B(17) => A(17), B(16) => A(16), B(15) => A(15), 
                           B(14) => A(14), B(13) => A(13), B(12) => A(12), 
                           B(11) => A(11), B(10) => A(10), B(9) => A(9), B(8) 
                           => A(8), B(7) => A(7), B(6) => A(6), B(5) => A(5), 
                           B(4) => A(4), B(3) => A(3), B(2) => A(2), B(1) => 
                           A(1), B(0) => A(0), CI => n5, DIFF(31) => A_n_63, 
                           DIFF(30) => A_n_30_port, DIFF(29) => A_n_29_port, 
                           DIFF(28) => A_n_28_port, DIFF(27) => A_n_27_port, 
                           DIFF(26) => A_n_26_port, DIFF(25) => A_n_25_port, 
                           DIFF(24) => A_n_24_port, DIFF(23) => A_n_23_port, 
                           DIFF(22) => A_n_22_port, DIFF(21) => A_n_21_port, 
                           DIFF(20) => A_n_20_port, DIFF(19) => A_n_19_port, 
                           DIFF(18) => A_n_18_port, DIFF(17) => A_n_17_port, 
                           DIFF(16) => A_n_16_port, DIFF(15) => A_n_15_port, 
                           DIFF(14) => A_n_14_port, DIFF(13) => A_n_13_port, 
                           DIFF(12) => A_n_12_port, DIFF(11) => A_n_11_port, 
                           DIFF(10) => A_n_10_port, DIFF(9) => A_n_9_port, 
                           DIFF(8) => A_n_8_port, DIFF(7) => A_n_7_port, 
                           DIFF(6) => A_n_6_port, DIFF(5) => A_n_5_port, 
                           DIFF(4) => A_n_4_port, DIFF(3) => A_n_3_port, 
                           DIFF(2) => A_n_2_port, DIFF(1) => A_n_1_port, 
                           DIFF(0) => A_n_0_port, CO => n_1310);

end SYN_BEHAVIOURAL;
