PACKAGE CONSTANTS IS
   CONSTANT IVDELAY : TIME := 0.1 ns;
   CONSTANT NDDELAY : TIME := 0.2 ns;
   CONSTANT NDDELAYRISE : TIME := 0.6 ns;
   CONSTANT NDDELAYFALL : TIME := 0.4 ns;
   CONSTANT NRDELAY : TIME := 0.2 ns;
   CONSTANT DRCAS : TIME := 1 ns;
   CONSTANT DRCAC : TIME := 2 ns;
   CONSTANT NumBit : INTEGER := 32;
   CONSTANT TP_MUX : TIME := 0.5 ns;
END CONSTANTS;